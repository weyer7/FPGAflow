* NGSPICE file created from fpgacell.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_1 abstract view
.subckt sky130_fd_sc_hd__clkinv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

.subckt fpgacell CBeast_in[0] CBeast_in[10] CBeast_in[11] CBeast_in[12] CBeast_in[13]
+ CBeast_in[1] CBeast_in[2] CBeast_in[3] CBeast_in[4] CBeast_in[5] CBeast_in[6] CBeast_in[7]
+ CBeast_in[8] CBeast_in[9] CBeast_out[0] CBeast_out[10] CBeast_out[11] CBeast_out[12]
+ CBeast_out[13] CBeast_out[1] CBeast_out[2] CBeast_out[3] CBeast_out[4] CBeast_out[5]
+ CBeast_out[6] CBeast_out[7] CBeast_out[8] CBeast_out[9] CBnorth_in[0] CBnorth_in[10]
+ CBnorth_in[11] CBnorth_in[12] CBnorth_in[13] CBnorth_in[1] CBnorth_in[2] CBnorth_in[3]
+ CBnorth_in[4] CBnorth_in[5] CBnorth_in[6] CBnorth_in[7] CBnorth_in[8] CBnorth_in[9]
+ CBnorth_out[0] CBnorth_out[10] CBnorth_out[11] CBnorth_out[12] CBnorth_out[13] CBnorth_out[1]
+ CBnorth_out[2] CBnorth_out[3] CBnorth_out[4] CBnorth_out[5] CBnorth_out[6] CBnorth_out[7]
+ CBnorth_out[8] CBnorth_out[9] SBsouth_in[0] SBsouth_in[10] SBsouth_in[11] SBsouth_in[12]
+ SBsouth_in[13] SBsouth_in[1] SBsouth_in[2] SBsouth_in[3] SBsouth_in[4] SBsouth_in[5]
+ SBsouth_in[6] SBsouth_in[7] SBsouth_in[8] SBsouth_in[9] SBsouth_out[0] SBsouth_out[10]
+ SBsouth_out[11] SBsouth_out[12] SBsouth_out[13] SBsouth_out[1] SBsouth_out[2] SBsouth_out[3]
+ SBsouth_out[4] SBsouth_out[5] SBsouth_out[6] SBsouth_out[7] SBsouth_out[8] SBsouth_out[9]
+ SBwest_in[0] SBwest_in[10] SBwest_in[11] SBwest_in[12] SBwest_in[13] SBwest_in[1]
+ SBwest_in[2] SBwest_in[3] SBwest_in[4] SBwest_in[5] SBwest_in[6] SBwest_in[7] SBwest_in[8]
+ SBwest_in[9] SBwest_out[0] SBwest_out[10] SBwest_out[11] SBwest_out[12] SBwest_out[13]
+ SBwest_out[1] SBwest_out[2] SBwest_out[3] SBwest_out[4] SBwest_out[5] SBwest_out[6]
+ SBwest_out[7] SBwest_out[8] SBwest_out[9] clk config_data_in config_data_out config_en
+ le_clk le_en le_nrst nrst vccd1 vssd1
X_2037_ _1213_ SB0.route_sel\[105\] _0794_ vssd1 vssd1 vccd1 vccd1 _0795_ sky130_fd_sc_hd__a21bo_1
X_2106_ CB_1.config_dataA\[3\] _0851_ _0854_ _0861_ _0863_ vssd1 vssd1 vccd1 vccd1
+ _0864_ sky130_fd_sc_hd__o2111a_1
X_3086_ clknet_leaf_18_clk _0294_ net217 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[6\]
+ sky130_fd_sc_hd__dfstp_1
X_2939_ clknet_leaf_27_clk _0147_ net195 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[11\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_43_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3076__SET_B net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2724_ net169 CB_0.config_dataA\[11\] net253 vssd1 vssd1 vccd1 vccd1 _0260_ sky130_fd_sc_hd__mux2_1
X_1606_ net174 _0367_ CB_0.config_dataA\[2\] vssd1 vssd1 vccd1 vccd1 _0368_ sky130_fd_sc_hd__o21ai_1
X_2655_ SB0.route_sel\[55\] SB0.route_sel\[54\] net258 vssd1 vssd1 vccd1 vccd1 _0191_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_57_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout138 net140 vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout127 CB_0.le_outB vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__buf_2
X_2586_ CB_1.config_dataB\[6\] net184 net263 vssd1 vssd1 vccd1 vccd1 _0122_ sky130_fd_sc_hd__mux2_1
Xfanout149 CB_1.config_dataA\[8\] vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__clkbuf_2
X_1399_ SB0.route_sel\[71\] vssd1 vssd1 vccd1 vccd1 _1193_ sky130_fd_sc_hd__inv_2
X_1468_ net142 net143 vssd1 vssd1 vccd1 vccd1 _1262_ sky130_fd_sc_hd__nand2b_1
X_1537_ _1258_ _1329_ net9 vssd1 vssd1 vccd1 vccd1 _1331_ sky130_fd_sc_hd__a21o_1
X_3069_ clknet_leaf_9_clk _0277_ net209 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[9\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_19_Left_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1978__A2 _0359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2155__A2 _0816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1551__X _1345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_31_clk_A clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2091__A1 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2440_ SB0.route_sel\[106\] SB0.route_sel\[107\] vssd1 vssd1 vccd1 vccd1 _1137_ sky130_fd_sc_hd__nand2b_1
XFILLER_5_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2371_ _1281_ _0377_ _0822_ vssd1 vssd1 vccd1 vccd1 _1092_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_62_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2082__A1 net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2707_ SB0.route_sel\[107\] SB0.route_sel\[106\] net268 vssd1 vssd1 vccd1 vccd1 _0243_
+ sky130_fd_sc_hd__mux2_1
X_2569_ net392 LE_1A.config_data\[9\] net259 vssd1 vssd1 vccd1 vccd1 _0105_ sky130_fd_sc_hd__mux2_1
X_2638_ SB0.route_sel\[38\] SB0.route_sel\[37\] net241 vssd1 vssd1 vccd1 vccd1 _0174_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__1896__A1 net20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_4_Left_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1820__A1 _0447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1584__B1 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2128__A2 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input55_A SBwest_in[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input10_X net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1722__A net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1871_ LEI0.config_data\[38\] _0606_ _0620_ _1222_ _0632_ vssd1 vssd1 vccd1 vccd1
+ _0633_ sky130_fd_sc_hd__o221a_1
X_1940_ _0690_ _0698_ _0699_ CB_0.config_dataB\[2\] vssd1 vssd1 vccd1 vccd1 _0700_
+ sky130_fd_sc_hd__a2bb2o_2
X_2423_ SB0.route_sel\[19\] _1166_ _1168_ _1169_ vssd1 vssd1 vccd1 vccd1 _1126_ sky130_fd_sc_hd__a22o_1
X_2285_ CB_1.config_dataB\[15\] _1040_ vssd1 vssd1 vccd1 vccd1 _1041_ sky130_fd_sc_hd__nor2_1
X_2354_ _0500_ _1083_ _0501_ vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__a21o_1
XFILLER_52_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1566__B1 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1802__A1 net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout128_X net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input2_X net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input58_X net58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2070_ _0489_ _0826_ vssd1 vssd1 vccd1 vccd1 _0828_ sky130_fd_sc_hd__nand2_1
X_2972_ clknet_leaf_23_clk _0180_ net212 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[44\]
+ sky130_fd_sc_hd__dfstp_1
X_1785_ _0447_ _0391_ net172 vssd1 vssd1 vccd1 vccd1 _0547_ sky130_fd_sc_hd__mux2_1
X_1854_ _1321_ _1345_ _1221_ vssd1 vssd1 vccd1 vccd1 _0616_ sky130_fd_sc_hd__mux2_1
X_1923_ net27 net28 net16 net17 net167 net166 vssd1 vssd1 vccd1 vccd1 _0683_ sky130_fd_sc_hd__mux4_1
X_2406_ _1318_ _1114_ vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__nor2_1
X_2337_ _1321_ net125 _1301_ vssd1 vssd1 vccd1 vccd1 _1075_ sky130_fd_sc_hd__mux2_1
X_2199_ _0827_ _0831_ _0835_ _0838_ _1242_ CB_1.config_dataB\[1\] vssd1 vssd1 vccd1
+ vccd1 _0955_ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout192_A net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2268_ _1021_ _1022_ _1017_ vssd1 vssd1 vccd1 vccd1 _1024_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_35_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold63 LE_0A.config_data\[2\] vssd1 vssd1 vccd1 vccd1 net335 sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 LE_1B.config_data\[2\] vssd1 vssd1 vccd1 vccd1 net324 sky130_fd_sc_hd__dlygate4sd3_1
Xhold30 LE_1A.config_data\[14\] vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 LE_1A.config_data\[8\] vssd1 vssd1 vccd1 vccd1 net346 sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 LE_1A.config_data\[3\] vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 LEI0.config_data\[39\] vssd1 vssd1 vccd1 vccd1 net368 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_43_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold85 LE_0B.config_data\[5\] vssd1 vssd1 vccd1 vccd1 net357 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input18_A CBnorth_in[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_7_Left_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_5 net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1570_ _0328_ _0330_ _0331_ vssd1 vssd1 vccd1 vccd1 _0332_ sky130_fd_sc_hd__and3_1
XANTENNA__1950__A0 net23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2053_ SB0.route_sel\[28\] SB0.route_sel\[29\] vssd1 vssd1 vccd1 vccd1 _0811_ sky130_fd_sc_hd__nor2_1
X_2122_ net9 net10 net11 net12 net149 CB_1.config_dataA\[9\] vssd1 vssd1 vccd1 vccd1
+ _0880_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_32_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2955_ clknet_leaf_23_clk _0163_ net211 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[27\]
+ sky130_fd_sc_hd__dfstp_1
X_1837_ _1297_ _0578_ _0579_ _1273_ vssd1 vssd1 vccd1 vccd1 _0599_ sky130_fd_sc_hd__o22a_1
X_1906_ _1359_ _0335_ _0338_ _1228_ vssd1 vssd1 vccd1 vccd1 _0666_ sky130_fd_sc_hd__a31o_1
X_1768_ SB0.route_sel\[84\] SB0.route_sel\[85\] net44 vssd1 vssd1 vccd1 vccd1 _0530_
+ sky130_fd_sc_hd__and3_1
XANTENNA__2194__A0 net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2886_ LE_1B.sel_clk _0094_ net61 vssd1 vssd1 vccd1 vccd1 LE_1B.dff1_out sky130_fd_sc_hd__dfstp_1
XANTENNA__1941__A0 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1699_ net131 _1330_ _0457_ _0460_ _1333_ vssd1 vssd1 vccd1 vccd1 _0461_ sky130_fd_sc_hd__o32a_1
XFILLER_40_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1607__S0 LEI0.config_data\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_33_Left_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2185__A0 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput64 net64 vssd1 vssd1 vccd1 vccd1 CBeast_out[10] sky130_fd_sc_hd__buf_2
Xoutput75 net75 vssd1 vssd1 vccd1 vccd1 CBeast_out[8] sky130_fd_sc_hd__buf_2
Xoutput86 net86 vssd1 vssd1 vccd1 vccd1 CBnorth_out[5] sky130_fd_sc_hd__buf_2
XANTENNA__2385__X net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput97 net97 vssd1 vssd1 vccd1 vccd1 SBsouth_out[2] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2740_ net163 CB_0.config_dataB\[7\] net252 vssd1 vssd1 vccd1 vccd1 _0276_ sky130_fd_sc_hd__mux2_1
X_1622_ SB0.route_sel\[26\] SB0.route_sel\[27\] _0378_ _0381_ _0383_ vssd1 vssd1 vccd1
+ vccd1 _0384_ sky130_fd_sc_hd__a221o_1
X_2671_ SB0.route_sel\[71\] SB0.route_sel\[70\] net239 vssd1 vssd1 vccd1 vccd1 _0207_
+ sky130_fd_sc_hd__mux2_1
X_1553_ SB0.route_sel\[106\] SB0.route_sel\[107\] vssd1 vssd1 vccd1 vccd1 _1347_ sky130_fd_sc_hd__nand2_1
XANTENNA__1923__A0 net27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2191__A3 _0819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1484_ SB0.route_sel\[49\] SB0.route_sel\[48\] vssd1 vssd1 vccd1 vccd1 _1278_ sky130_fd_sc_hd__nand2_1
X_2036_ SB0.route_sel\[108\] SB0.route_sel\[109\] net119 _1212_ vssd1 vssd1 vccd1
+ vccd1 _0794_ sky130_fd_sc_hd__o22a_1
X_2105_ _0855_ _0862_ vssd1 vssd1 vccd1 vccd1 _0863_ sky130_fd_sc_hd__nand2b_1
X_3085_ clknet_leaf_19_clk _0293_ net217 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[5\]
+ sky130_fd_sc_hd__dfstp_2
XANTENNA__1786__S net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2938_ clknet_leaf_27_clk _0146_ net195 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[10\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_22_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2869_ clknet_leaf_3_clk net351 net201 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_43_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_51_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_5_clk_A clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1905__A0 _1345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2723_ CB_0.config_dataA\[11\] CB_0.config_dataA\[10\] net249 vssd1 vssd1 vccd1 vccd1
+ _0259_ sky130_fd_sc_hd__mux2_1
XFILLER_44_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1605_ CB_0.config_dataA\[1\] CB_0.config_dataA\[3\] vssd1 vssd1 vccd1 vccd1 _0367_
+ sky130_fd_sc_hd__nand2_1
X_2585_ net184 CB_1.config_dataB\[4\] net264 vssd1 vssd1 vccd1 vccd1 _0121_ sky130_fd_sc_hd__mux2_1
X_2654_ SB0.route_sel\[54\] SB0.route_sel\[53\] net260 vssd1 vssd1 vccd1 vccd1 _0190_
+ sky130_fd_sc_hd__mux2_1
X_1536_ net177 net178 vssd1 vssd1 vccd1 vccd1 _1330_ sky130_fd_sc_hd__or2_2
XANTENNA_fanout272_A net58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout139 net140 vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_57_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout128 net130 vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__buf_2
X_1467_ CB_1.config_dataA\[17\] net145 vssd1 vssd1 vccd1 vccd1 _1261_ sky130_fd_sc_hd__nand2_2
X_1398_ SB0.route_sel\[68\] vssd1 vssd1 vccd1 vccd1 _1192_ sky130_fd_sc_hd__inv_2
X_3068_ clknet_leaf_9_clk _0276_ net209 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[8\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2019_ CB_1.config_dataA\[5\] CB_1.config_dataA\[7\] vssd1 vssd1 vccd1 vccd1 _0777_
+ sky130_fd_sc_hd__nand2_1
XFILLER_50_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2155__A3 _0813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2095__B _0831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2091__A2 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1455__A net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2370_ _0381_ _1091_ _0383_ vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_20_Left_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2706_ SB0.route_sel\[106\] SB0.route_sel\[105\] net268 vssd1 vssd1 vccd1 vccd1 _0242_
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2499_ net387 LEI0.config_data\[36\] net270 vssd1 vssd1 vccd1 vccd1 _0038_ sky130_fd_sc_hd__mux2_1
XANTENNA__1896__A2 net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2568_ net403 net346 net259 vssd1 vssd1 vccd1 vccd1 _0104_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_12_Right_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2637_ SB0.route_sel\[37\] SB0.route_sel\[36\] net238 vssd1 vssd1 vccd1 vccd1 _0173_
+ sky130_fd_sc_hd__mux2_1
X_1519_ SB0.route_sel\[43\] SB0.route_sel\[42\] _1307_ _1310_ _1312_ vssd1 vssd1 vccd1
+ vccd1 _1313_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_21_Right_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_30_Right_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2128__A3 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1887__A2 _0645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input48_A SBwest_in[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1870_ _0630_ _0631_ _1222_ vssd1 vssd1 vccd1 vccd1 _0632_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_24_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2353_ net177 net178 _0456_ _0835_ vssd1 vssd1 vccd1 vccd1 _1083_ sky130_fd_sc_hd__a31o_1
X_2422_ SB0.route_sel\[17\] _1170_ vssd1 vssd1 vccd1 vccd1 _1125_ sky130_fd_sc_hd__nor2_1
XFILLER_37_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2284_ net1 net6 net7 net8 net180 net179 vssd1 vssd1 vccd1 vccd1 _1040_ sky130_fd_sc_hd__mux4_1
X_1999_ _0758_ vssd1 vssd1 vccd1 vccd1 _0759_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_30_clk_A clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1922_ _0513_ _0539_ _1225_ vssd1 vssd1 vccd1 vccd1 _0682_ sky130_fd_sc_hd__mux2_1
X_2971_ clknet_leaf_23_clk _0179_ net212 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[43\]
+ sky130_fd_sc_hd__dfstp_1
X_1784_ net171 net172 vssd1 vssd1 vccd1 vccd1 _0546_ sky130_fd_sc_hd__nand2_1
X_1853_ net169 _0359_ _0614_ vssd1 vssd1 vccd1 vccd1 _0615_ sky130_fd_sc_hd__o21a_1
X_2336_ net139 _1074_ _1275_ vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__mux2_1
X_2405_ SB0.route_sel\[47\] SB0.route_sel\[46\] SB0.route_sel\[41\] _1183_ _1113_
+ vssd1 vssd1 vccd1 vccd1 _1114_ sky130_fd_sc_hd__o221a_1
X_2198_ CB_1.config_dataB\[3\] _0949_ _0953_ vssd1 vssd1 vccd1 vccd1 _0954_ sky130_fd_sc_hd__o21ai_1
X_2267_ LE_1B.config_data\[0\] LE_1B.config_data\[1\] _0961_ vssd1 vssd1 vccd1 vccd1
+ _1023_ sky130_fd_sc_hd__mux2_1
XFILLER_1_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1787__B2 net22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1787__A1 net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold97 LEI0.config_data\[46\] vssd1 vssd1 vccd1 vccd1 net369 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 LE_0A.config_data\[12\] vssd1 vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_42_Left_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold64 LEI0.config_data\[26\] vssd1 vssd1 vccd1 vccd1 net336 sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 _0078_ vssd1 vssd1 vccd1 vccd1 net358 sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 LEI0.config_data\[22\] vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 LE_1B.config_data\[4\] vssd1 vssd1 vccd1 vccd1 net325 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 _0109_ vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 LE_1B.config_data\[7\] vssd1 vssd1 vccd1 vccd1 net347 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_51_Left_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_6 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_60_Left_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1950__A1 net24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_49_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1750__X _0512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2052_ _0778_ _0809_ CB_1.config_dataA\[6\] vssd1 vssd1 vccd1 vccd1 _0810_ sky130_fd_sc_hd__o21ai_1
X_2121_ net148 _0797_ _0877_ _0878_ vssd1 vssd1 vccd1 vccd1 _0879_ sky130_fd_sc_hd__a211o_1
XANTENNA__1466__B1 net12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1905_ _1345_ _1321_ _1297_ _1273_ net165 CB_0.config_dataB\[5\] vssd1 vssd1 vccd1
+ vccd1 _0665_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_32_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2885_ LE_1A.sel_clk _0093_ net61 vssd1 vssd1 vccd1 vccd1 LE_1A.dff0_out sky130_fd_sc_hd__dfrtp_1
X_2954_ clknet_leaf_24_clk _0162_ net211 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[26\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__1638__A net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1836_ CB_0.config_dataA\[11\] _0597_ _0595_ vssd1 vssd1 vccd1 vccd1 _0598_ sky130_fd_sc_hd__o21ai_1
XANTENNA__1941__A1 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2194__A1 net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1767_ _0525_ _0526_ _0527_ _0528_ vssd1 vssd1 vccd1 vccd1 _0529_ sky130_fd_sc_hd__a211oi_1
XPHY_EDGE_ROW_6_Right_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1698_ net143 net142 vssd1 vssd1 vccd1 vccd1 _0460_ sky130_fd_sc_hd__nand2b_1
X_2319_ net187 LE_1B.reset_mode vssd1 vssd1 vccd1 vccd1 _2319_/X sky130_fd_sc_hd__xor2_2
XFILLER_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput87 net87 vssd1 vssd1 vccd1 vccd1 CBnorth_out[6] sky130_fd_sc_hd__buf_2
XANTENNA__2185__A1 net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput65 net65 vssd1 vssd1 vccd1 vccd1 CBeast_out[11] sky130_fd_sc_hd__buf_2
Xoutput76 net76 vssd1 vssd1 vccd1 vccd1 CBeast_out[9] sky130_fd_sc_hd__buf_2
Xoutput98 net98 vssd1 vssd1 vccd1 vccd1 SBsouth_out[3] sky130_fd_sc_hd__buf_2
XFILLER_48_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output117_A net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input30_A SBsouth_in[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1696__B1 net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_59_Right_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_54_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1552_ _1273_ _1297_ _1321_ _1345_ _1165_ _1154_ vssd1 vssd1 vccd1 vccd1 _1346_ sky130_fd_sc_hd__mux4_1
XANTENNA__1923__A1 net28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2670_ SB0.route_sel\[70\] SB0.route_sel\[69\] net239 vssd1 vssd1 vccd1 vccd1 _0206_
+ sky130_fd_sc_hd__mux2_1
X_1621_ _1249_ _1261_ _0380_ vssd1 vssd1 vccd1 vccd1 _0383_ sky130_fd_sc_hd__nor3_1
X_1483_ net25 net125 _1276_ vssd1 vssd1 vccd1 vccd1 _1277_ sky130_fd_sc_hd__mux2_1
XANTENNA__1687__A0 _0391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2104_ _0838_ _0835_ net151 vssd1 vssd1 vccd1 vccd1 _0862_ sky130_fd_sc_hd__mux2_1
XFILLER_47_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3084_ clknet_leaf_19_clk _0292_ net217 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[4\]
+ sky130_fd_sc_hd__dfstp_1
X_2035_ _0784_ _0792_ _0781_ _0788_ _1237_ CB_1.config_dataA\[5\] vssd1 vssd1 vccd1
+ vccd1 _0793_ sky130_fd_sc_hd__mux4_1
XFILLER_22_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1611__A0 net22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2868_ clknet_leaf_3_clk _0076_ net201 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_2937_ clknet_leaf_28_clk _0145_ net188 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[9\]
+ sky130_fd_sc_hd__dfstp_1
X_1819_ _1217_ _0576_ _0580_ vssd1 vssd1 vccd1 vccd1 _0581_ sky130_fd_sc_hd__a21o_1
X_2799_ clknet_leaf_5_clk _0007_ net201 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_60_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1850__A0 net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1905__A1 _1321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input33_X net33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2722_ CB_0.config_dataA\[10\] CB_0.config_dataA\[9\] net249 vssd1 vssd1 vccd1 vccd1
+ _0258_ sky130_fd_sc_hd__mux2_1
X_1604_ _0364_ _0365_ vssd1 vssd1 vccd1 vccd1 _0366_ sky130_fd_sc_hd__nor2_1
Xfanout129 net130 vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__dlymetal6s2s_1
X_2584_ net185 CB_1.config_dataB\[3\] net257 vssd1 vssd1 vccd1 vccd1 _0120_ sky130_fd_sc_hd__mux2_1
X_2653_ SB0.route_sel\[53\] SB0.route_sel\[52\] net258 vssd1 vssd1 vccd1 vccd1 _0189_
+ sky130_fd_sc_hd__mux2_1
X_1535_ CB_1.config_dataB\[17\] CB_1.config_dataB\[16\] vssd1 vssd1 vccd1 vccd1 _1329_
+ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_57_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3067_ clknet_leaf_2_clk _0275_ net209 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[7\]
+ sky130_fd_sc_hd__dfstp_1
X_1397_ SB0.route_sel\[67\] vssd1 vssd1 vccd1 vccd1 _1191_ sky130_fd_sc_hd__inv_2
X_1466_ net177 net178 _1258_ net12 vssd1 vssd1 vccd1 vccd1 _1260_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout265_A net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2018_ LE_0B.config_data\[16\] _0775_ _0776_ _0646_ vssd1 vssd1 vccd1 vccd1 CB_0.le_outB
+ sky130_fd_sc_hd__o211a_1
XFILLER_6_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2560__A1 LE_1A.config_data\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2091__A3 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2171__S0 _0848_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2705_ SB0.route_sel\[105\] SB0.route_sel\[104\] net268 vssd1 vssd1 vccd1 vccd1 _0241_
+ sky130_fd_sc_hd__mux2_1
X_2636_ SB0.route_sel\[36\] SB0.route_sel\[35\] net239 vssd1 vssd1 vccd1 vccd1 _0172_
+ sky130_fd_sc_hd__mux2_1
X_2498_ net409 LEI0.config_data\[35\] net270 vssd1 vssd1 vccd1 vccd1 _0037_ sky130_fd_sc_hd__mux2_1
XANTENNA__1896__A3 net22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1449_ CB_1.config_dataB\[3\] vssd1 vssd1 vccd1 vccd1 _1243_ sky130_fd_sc_hd__inv_2
X_2567_ net346 net310 net259 vssd1 vssd1 vccd1 vccd1 _0103_ sky130_fd_sc_hd__mux2_1
X_1518_ _1249_ _1262_ _1309_ vssd1 vssd1 vccd1 vccd1 _1312_ sky130_fd_sc_hd__nor3_1
XANTENNA_clkbuf_leaf_4_clk_A clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3119_ clknet_leaf_30_clk _0327_ net187 vssd1 vssd1 vccd1 vccd1 LE_1B.reset_mode
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2297__B1 _1052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2144__S0 _0848_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2283_ _0819_ _0822_ _0816_ _0813_ net179 net180 vssd1 vssd1 vccd1 vccd1 _1039_ sky130_fd_sc_hd__mux4_1
X_2352_ _0348_ _1082_ _0350_ vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__a21o_1
X_2421_ _1123_ _1124_ _0444_ vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__a21boi_1
XFILLER_37_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout228_A net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1998_ CB_0.config_dataB\[14\] _0756_ _0757_ vssd1 vssd1 vccd1 vccd1 _0758_ sky130_fd_sc_hd__o21a_1
X_2619_ SB0.route_sel\[19\] SB0.route_sel\[18\] net232 vssd1 vssd1 vccd1 vccd1 _0155_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__2279__A0 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2294__A3 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input60_A le_en vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1852_ net169 _0339_ _0611_ vssd1 vssd1 vccd1 vccd1 _0614_ sky130_fd_sc_hd__a21oi_1
X_1921_ _0474_ _0493_ CB_0.config_dataB\[0\] vssd1 vssd1 vccd1 vccd1 _0681_ sky130_fd_sc_hd__mux2_1
X_2970_ clknet_leaf_22_clk _0178_ net212 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[42\]
+ sky130_fd_sc_hd__dfstp_1
X_1783_ net172 net171 vssd1 vssd1 vccd1 vccd1 _0545_ sky130_fd_sc_hd__nand2b_1
XANTENNA__1548__A2 _1328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2335_ _1297_ net125 _1276_ vssd1 vssd1 vccd1 vccd1 _1074_ sky130_fd_sc_hd__mux2_1
X_2266_ LE_1B.config_data\[2\] net120 net135 _0984_ _0986_ vssd1 vssd1 vccd1 vccd1
+ _1022_ sky130_fd_sc_hd__a32o_1
X_2404_ SB0.route_sel\[42\] SB0.route_sel\[43\] vssd1 vssd1 vccd1 vccd1 _1113_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_35_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2197_ CB_1.config_dataB\[1\] _1243_ _0950_ _0952_ vssd1 vssd1 vccd1 vccd1 _0953_
+ sky130_fd_sc_hd__o31a_1
XANTENNA_fanout133_X net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold87 LE_0A.config_data\[4\] vssd1 vssd1 vccd1 vccd1 net359 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 _0063_ vssd1 vssd1 vccd1 vccd1 net315 sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 _0047_ vssd1 vssd1 vccd1 vccd1 net370 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 LE_0B.config_data\[8\] vssd1 vssd1 vccd1 vccd1 net348 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 _0027_ vssd1 vssd1 vccd1 vccd1 net337 sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 LE_1A.config_data\[1\] vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 LE_1A.config_data\[6\] vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 LE_1B.config_data\[13\] vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 _0313_ vssd1 vssd1 vccd1 vccd1 net326 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_7 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1950__A2 net25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2120_ net148 _0803_ vssd1 vssd1 vccd1 vccd1 _0878_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_49_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2051_ _1238_ _0793_ _0808_ vssd1 vssd1 vccd1 vccd1 _0809_ sky130_fd_sc_hd__a21oi_1
X_1835_ CB_0.config_dataA\[8\] _1321_ _0596_ vssd1 vssd1 vccd1 vccd1 _0597_ sky130_fd_sc_hd__a21oi_1
X_1904_ _0650_ _0653_ _0663_ vssd1 vssd1 vccd1 vccd1 _0664_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_32_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2884_ clknet_leaf_29_clk _0092_ net186 vssd1 vssd1 vccd1 vccd1 LE_0B.reset_mode
+ sky130_fd_sc_hd__dfrtp_1
X_2953_ clknet_leaf_26_clk _0161_ net194 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[25\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__1654__A net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1941__A2 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2718__A1 net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1766_ net128 _1283_ _0459_ vssd1 vssd1 vccd1 vccd1 _0528_ sky130_fd_sc_hd__and3_1
X_1697_ net143 net142 vssd1 vssd1 vccd1 vccd1 _0459_ sky130_fd_sc_hd__and2b_1
X_2249_ CB_1.config_dataB\[10\] _0999_ _1002_ _1004_ vssd1 vssd1 vccd1 vccd1 _1005_
+ sky130_fd_sc_hd__a31o_1
X_2318_ net59 LE_1A.edge_mode vssd1 vssd1 vccd1 vccd1 LE_1A.sel_clk sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout250_X net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput77 net77 vssd1 vssd1 vccd1 vccd1 CBnorth_out[0] sky130_fd_sc_hd__buf_2
Xoutput88 net88 vssd1 vssd1 vccd1 vccd1 CBnorth_out[7] sky130_fd_sc_hd__buf_2
XANTENNA__1932__A2 _0359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput66 net66 vssd1 vssd1 vccd1 vccd1 CBeast_out[12] sky130_fd_sc_hd__buf_2
Xoutput99 net99 vssd1 vssd1 vccd1 vccd1 SBsouth_out[4] sky130_fd_sc_hd__buf_2
XANTENNA__1791__S1 net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input23_A CBnorth_in[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1482_ net160 net154 net156 net158 vssd1 vssd1 vccd1 vccd1 _1276_ sky130_fd_sc_hd__and4bb_1
X_1551_ _1342_ _1344_ vssd1 vssd1 vccd1 vccd1 _1345_ sky130_fd_sc_hd__and2_2
XANTENNA__1923__A2 net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1620_ SB0.route_sel\[26\] SB0.route_sel\[27\] vssd1 vssd1 vccd1 vccd1 _0382_ sky130_fd_sc_hd__nand2_1
X_3083_ clknet_leaf_15_clk _0291_ net223 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[3\]
+ sky130_fd_sc_hd__dfstp_2
X_2103_ _0858_ _0860_ CB_1.config_dataA\[2\] vssd1 vssd1 vccd1 vccd1 _0861_ sky130_fd_sc_hd__a21oi_1
X_2034_ _1342_ _0791_ vssd1 vssd1 vccd1 vccd1 _0792_ sky130_fd_sc_hd__and2_1
XFILLER_22_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1818_ CB_0.config_dataA\[9\] net170 _0391_ CB_0.config_dataA\[11\] vssd1 vssd1 vccd1
+ vccd1 _0580_ sky130_fd_sc_hd__a31o_1
X_2798_ clknet_leaf_5_clk net297 net205 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout210_A net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2867_ clknet_leaf_3_clk net317 net202 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_2936_ clknet_leaf_28_clk _0144_ net188 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[8\]
+ sky130_fd_sc_hd__dfstp_1
X_1749_ _1204_ SB0.route_sel\[93\] vssd1 vssd1 vccd1 vccd1 _0511_ sky130_fd_sc_hd__nor2_1
XANTENNA__1850__A1 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1905__A2 _1297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2158__A2 _0831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input26_X net26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2721_ CB_0.config_dataA\[9\] net170 net248 vssd1 vssd1 vccd1 vccd1 _0257_ sky130_fd_sc_hd__mux2_1
XFILLER_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2652_ SB0.route_sel\[52\] SB0.route_sel\[51\] net258 vssd1 vssd1 vccd1 vccd1 _0188_
+ sky130_fd_sc_hd__mux2_1
X_1534_ _1325_ _1326_ _1327_ vssd1 vssd1 vccd1 vccd1 _1328_ sky130_fd_sc_hd__a21o_1
X_1603_ _1214_ _1346_ _0340_ _0360_ vssd1 vssd1 vccd1 vccd1 _0365_ sky130_fd_sc_hd__a22o_1
X_2583_ CB_1.config_dataB\[3\] CB_1.config_dataB\[2\] net257 vssd1 vssd1 vccd1 vccd1
+ _0119_ sky130_fd_sc_hd__mux2_1
X_1465_ net175 net176 vssd1 vssd1 vccd1 vccd1 _1259_ sky130_fd_sc_hd__nand2b_1
X_3066_ clknet_leaf_2_clk _0274_ net209 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[6\]
+ sky130_fd_sc_hd__dfstp_1
X_2017_ _1234_ LE_0B.dff_out vssd1 vssd1 vccd1 vccd1 _0776_ sky130_fd_sc_hd__or2_1
X_1396_ SB0.route_sel\[57\] vssd1 vssd1 vccd1 vccd1 _1190_ sky130_fd_sc_hd__inv_2
X_2919_ clknet_leaf_15_clk _0127_ net222 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[11\]
+ sky130_fd_sc_hd__dfstp_2
XANTENNA_fanout258_A net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold140 LEI0.config_data\[15\] vssd1 vssd1 vccd1 vccd1 net412 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2171__S1 _0874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1814__A1 _0430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2704_ SB0.route_sel\[104\] SB0.route_sel\[103\] net265 vssd1 vssd1 vccd1 vccd1 _0240_
+ sky130_fd_sc_hd__mux2_1
X_2635_ SB0.route_sel\[35\] SB0.route_sel\[34\] net240 vssd1 vssd1 vccd1 vccd1 _0171_
+ sky130_fd_sc_hd__mux2_1
X_2497_ LEI0.config_data\[35\] net378 net270 vssd1 vssd1 vccd1 vccd1 _0036_ sky130_fd_sc_hd__mux2_1
X_1448_ CB_1.config_dataB\[0\] vssd1 vssd1 vccd1 vccd1 _1242_ sky130_fd_sc_hd__inv_2
XFILLER_4_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2566_ net310 net293 net259 vssd1 vssd1 vccd1 vccd1 _0102_ sky130_fd_sc_hd__mux2_1
X_1517_ SB0.route_sel\[43\] SB0.route_sel\[42\] vssd1 vssd1 vccd1 vccd1 _1311_ sky130_fd_sc_hd__nand2_1
X_3049_ clknet_leaf_7_clk _0257_ net205 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[9\]
+ sky130_fd_sc_hd__dfstp_2
X_1379_ SB0.route_sel\[31\] vssd1 vssd1 vccd1 vccd1 _1173_ sky130_fd_sc_hd__inv_2
X_3118_ clknet_leaf_30_clk _0326_ net187 vssd1 vssd1 vccd1 vccd1 LE_1B.reset_val sky130_fd_sc_hd__dfrtp_1
XFILLER_48_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2144__S1 _0874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1980__A0 net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2420_ SB0.route_sel\[19\] _1166_ SB0.route_sel\[20\] _1167_ vssd1 vssd1 vccd1 vccd1
+ _1124_ sky130_fd_sc_hd__o22a_1
X_2282_ _1031_ _1033_ _1036_ CB_1.config_dataB\[14\] vssd1 vssd1 vccd1 vccd1 _1038_
+ sky130_fd_sc_hd__o211a_1
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2351_ CB_1.config_dataB\[19\] net176 _1329_ _0803_ vssd1 vssd1 vccd1 vccd1 _1082_
+ sky130_fd_sc_hd__a31o_1
XFILLER_37_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1997_ _1231_ _0745_ _0744_ vssd1 vssd1 vccd1 vccd1 _0757_ sky130_fd_sc_hd__a21oi_1
XANTENNA__1799__A0 net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2549_ net331 net327 net242 vssd1 vssd1 vccd1 vccd1 _0086_ sky130_fd_sc_hd__mux2_1
X_2618_ SB0.route_sel\[18\] SB0.route_sel\[17\] net232 vssd1 vssd1 vccd1 vccd1 _0154_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__2279__A1 net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1962__A0 net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input53_A SBwest_in[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1851_ CB_0.config_dataA\[15\] _0610_ _0611_ _0612_ vssd1 vssd1 vccd1 vccd1 _0613_
+ sky130_fd_sc_hd__o22a_1
X_1920_ CB_0.config_dataB\[3\] _0679_ _0678_ vssd1 vssd1 vccd1 vccd1 _0680_ sky130_fd_sc_hd__o21ai_1
X_1782_ _0430_ net121 net172 vssd1 vssd1 vccd1 vccd1 _0544_ sky130_fd_sc_hd__mux2_1
X_2403_ _1318_ _1112_ vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_3_clk_A clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2334_ net138 _1073_ _1252_ vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__mux2_1
X_2196_ _0945_ _0951_ vssd1 vssd1 vccd1 vccd1 _0952_ sky130_fd_sc_hd__or2_1
X_2265_ net120 net135 LE_1B.config_data\[3\] vssd1 vssd1 vccd1 vccd1 _1021_ sky130_fd_sc_hd__a21boi_1
XANTENNA__2130__A0 _0819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold22 LE_0A.config_data\[1\] vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__dlygate4sd3_1
Xhold11 LE_1B.config_data\[1\] vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3088__SET_B net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold88 LEI0.config_data\[31\] vssd1 vssd1 vccd1 vccd1 net360 sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 LEI0.config_data\[33\] vssd1 vssd1 vccd1 vccd1 net371 sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 LE_0B.config_data\[2\] vssd1 vssd1 vccd1 vccd1 net316 sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 LE_0B.config_data\[12\] vssd1 vssd1 vccd1 vccd1 net327 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 _0081_ vssd1 vssd1 vccd1 vccd1 net349 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 LE_1A.config_data\[2\] vssd1 vssd1 vccd1 vccd1 net305 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 LE_1B.config_data\[11\] vssd1 vssd1 vccd1 vccd1 net338 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_8 CBeast_in[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1950__A3 net26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2050_ _0798_ _0799_ _0804_ _0807_ vssd1 vssd1 vccd1 vccd1 _0808_ sky130_fd_sc_hd__a31o_1
XFILLER_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2952_ clknet_leaf_28_clk _0160_ net195 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[24\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_19_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1834_ _1218_ _1342_ _1344_ CB_0.config_dataA\[9\] vssd1 vssd1 vccd1 vccd1 _0596_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__1926__A0 _0391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1903_ _0538_ _0655_ _0657_ _0512_ _0662_ vssd1 vssd1 vccd1 vccd1 _0663_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_32_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1765_ SB0.route_sel\[82\] SB0.route_sel\[83\] vssd1 vssd1 vccd1 vccd1 _0527_ sky130_fd_sc_hd__and2_1
X_2883_ clknet_leaf_29_clk _0091_ net186 vssd1 vssd1 vccd1 vccd1 LE_0B.reset_val sky130_fd_sc_hd__dfrtp_1
XANTENNA__1941__A3 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1696_ _1329_ _0456_ net13 vssd1 vssd1 vccd1 vccd1 _0458_ sky130_fd_sc_hd__a21o_1
X_2248_ _1003_ _1245_ CB_1.config_dataB\[10\] vssd1 vssd1 vccd1 vccd1 _1004_ sky130_fd_sc_hd__and3b_1
X_2317_ net186 LE_1A.reset_mode vssd1 vssd1 vccd1 vccd1 _2317_/X sky130_fd_sc_hd__xor2_2
X_2179_ LE_1A.config_data\[16\] _0934_ _0935_ _0646_ vssd1 vssd1 vccd1 vccd1 CB_1.le_outA
+ sky130_fd_sc_hd__o211a_1
XFILLER_25_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1917__A0 net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput78 net78 vssd1 vssd1 vccd1 vccd1 CBnorth_out[10] sky130_fd_sc_hd__buf_2
Xoutput89 net89 vssd1 vssd1 vccd1 vccd1 CBnorth_out[8] sky130_fd_sc_hd__buf_2
Xoutput67 net67 vssd1 vssd1 vccd1 vccd1 CBeast_out[13] sky130_fd_sc_hd__buf_2
XFILLER_63_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input16_A CBnorth_in[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_0__f_clk_X clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1908__A0 net23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1481_ _1251_ _1274_ vssd1 vssd1 vccd1 vccd1 _1275_ sky130_fd_sc_hd__nand2_1
XANTENNA__2333__A0 _1273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1923__A3 net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1550_ SB0.route_sel\[36\] _1176_ SB0.route_sel\[39\] _1178_ _1343_ vssd1 vssd1 vccd1
+ vccd1 _1344_ sky130_fd_sc_hd__a221o_1
XANTENNA__1687__A2 _0447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3082_ clknet_leaf_15_clk _0290_ net223 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[2\]
+ sky130_fd_sc_hd__dfstp_1
X_2102_ CB_1.config_dataA\[3\] _0856_ _0859_ _0855_ vssd1 vssd1 vccd1 vccd1 _0860_
+ sky130_fd_sc_hd__o22a_1
X_2033_ _1177_ SB0.route_sel\[38\] SB0.route_sel\[33\] _1179_ _0790_ vssd1 vssd1 vccd1
+ vccd1 _0791_ sky130_fd_sc_hd__a221o_1
XANTENNA__2822__Q LEI0.config_data\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2935_ clknet_leaf_28_clk _0143_ net188 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[7\]
+ sky130_fd_sc_hd__dfstp_1
X_1817_ CB_0.config_dataA\[9\] net170 vssd1 vssd1 vccd1 vccd1 _0579_ sky130_fd_sc_hd__nand2_1
X_2797_ clknet_leaf_5_clk _0005_ net203 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_1748_ SB0.route_sel\[94\] SB0.route_sel\[95\] vssd1 vssd1 vccd1 vccd1 _0510_ sky130_fd_sc_hd__and2b_1
X_2866_ clknet_leaf_3_clk net402 net201 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input8_A CBeast_in[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1679_ _1168_ _1169_ net49 SB0.route_sel\[21\] SB0.route_sel\[20\] vssd1 vssd1 vccd1
+ vccd1 _0441_ sky130_fd_sc_hd__o2111a_1
XANTENNA_fanout193_X net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1905__A3 _1273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_39_Left_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input19_X net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_48_Left_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1741__C net45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2720_ net170 CB_0.config_dataA\[7\] net249 vssd1 vssd1 vccd1 vccd1 _0256_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_57_Left_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1602_ CB_0.config_dataA\[1\] _1214_ _0363_ _0362_ vssd1 vssd1 vccd1 vccd1 _0364_
+ sky130_fd_sc_hd__o31a_1
X_2582_ CB_1.config_dataB\[2\] CB_1.config_dataB\[1\] net257 vssd1 vssd1 vccd1 vccd1
+ _0118_ sky130_fd_sc_hd__mux2_1
X_2651_ SB0.route_sel\[51\] SB0.route_sel\[50\] net258 vssd1 vssd1 vccd1 vccd1 _0187_
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1533_ net138 _1251_ _1324_ vssd1 vssd1 vccd1 vccd1 _1327_ sky130_fd_sc_hd__and3_1
X_1395_ SB0.route_sel\[60\] vssd1 vssd1 vccd1 vccd1 _1189_ sky130_fd_sc_hd__inv_2
X_1464_ net175 CB_1.config_dataB\[18\] vssd1 vssd1 vccd1 vccd1 _1258_ sky130_fd_sc_hd__and2b_2
XANTENNA__2306__B1 _1017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3065_ clknet_leaf_3_clk _0273_ net208 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[5\]
+ sky130_fd_sc_hd__dfstp_2
X_2016_ LE_0B.dff0_out LE_0B.dff1_out LE_0B.reset_val vssd1 vssd1 vccd1 vccd1 LE_0B.dff_out
+ sky130_fd_sc_hd__mux2_1
XANTENNA__1832__A2 _0339_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2918_ clknet_leaf_15_clk _0126_ net222 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[10\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_10_107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_30_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_clk
+ sky130_fd_sc_hd__clkbuf_8
Xhold141 LE_0A.config_data\[5\] vssd1 vssd1 vccd1 vccd1 net413 sky130_fd_sc_hd__dlygate4sd3_1
X_2849_ clknet_leaf_6_clk net377 net204 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold130 _0074_ vssd1 vssd1 vccd1 vccd1 net402 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_5_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_21_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_5_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wire121_A _0411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_12_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2703_ SB0.route_sel\[103\] SB0.route_sel\[102\] net264 vssd1 vssd1 vccd1 vccd1 _0239_
+ sky130_fd_sc_hd__mux2_1
X_2565_ net293 net291 net260 vssd1 vssd1 vccd1 vccd1 _0101_ sky130_fd_sc_hd__mux2_1
X_1516_ net132 _1259_ _1306_ _1309_ _1262_ vssd1 vssd1 vccd1 vccd1 _1310_ sky130_fd_sc_hd__o32a_1
X_2634_ SB0.route_sel\[34\] SB0.route_sel\[33\] net240 vssd1 vssd1 vccd1 vccd1 _0170_
+ sky130_fd_sc_hd__mux2_1
X_2496_ net378 net371 net269 vssd1 vssd1 vccd1 vccd1 _0035_ sky130_fd_sc_hd__mux2_1
X_1447_ CB_1.config_dataB\[1\] vssd1 vssd1 vccd1 vccd1 _1241_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_2_147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1378_ SB0.route_sel\[29\] vssd1 vssd1 vccd1 vccd1 _1172_ sky130_fd_sc_hd__inv_2
X_3117_ clknet_leaf_29_clk _0325_ net187 vssd1 vssd1 vccd1 vccd1 LE_1B.edge_mode sky130_fd_sc_hd__dfstp_1
X_3048_ clknet_leaf_7_clk _0256_ net206 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[8\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__2297__A2 _1017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1980__A1 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_24_Left_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2281_ net181 CB_1.config_dataB\[14\] CB_1.config_dataB\[15\] net179 vssd1 vssd1
+ vccd1 vccd1 _1037_ sky130_fd_sc_hd__and4b_1
Xclkbuf_leaf_1_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2350_ _1350_ _1351_ _1081_ _1352_ vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__a31o_1
XANTENNA__1799__A1 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1996_ CB_0.config_dataB\[15\] _0746_ _0748_ _0755_ vssd1 vssd1 vccd1 vccd1 _0756_
+ sky130_fd_sc_hd__o211a_1
XFILLER_20_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2548_ net327 LE_0B.config_data\[11\] net243 vssd1 vssd1 vccd1 vccd1 _0085_ sky130_fd_sc_hd__mux2_1
X_2617_ SB0.route_sel\[17\] SB0.route_sel\[16\] net231 vssd1 vssd1 vccd1 vccd1 _0153_
+ sky130_fd_sc_hd__mux2_1
X_2479_ net385 net374 net244 vssd1 vssd1 vccd1 vccd1 _0018_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_38_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1962__A1 net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload0 clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload0/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_7_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout270 net271 vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input46_A SBwest_in[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1850_ net18 net19 net169 vssd1 vssd1 vccd1 vccd1 _0612_ sky130_fd_sc_hd__mux2_1
X_1781_ _0366_ _0368_ _0370_ _0542_ vssd1 vssd1 vccd1 vccd1 _0543_ sky130_fd_sc_hd__o211a_2
X_2333_ _1273_ net124 _1253_ vssd1 vssd1 vccd1 vccd1 _1073_ sky130_fd_sc_hd__mux2_1
X_2402_ SB0.route_sel\[44\] _1181_ SB0.route_sel\[41\] SB0.route_sel\[40\] _1111_
+ vssd1 vssd1 vccd1 vccd1 _1112_ sky130_fd_sc_hd__o221a_1
XANTENNA__1800__S1 net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2195_ net2 net3 CB_1.config_dataB\[0\] vssd1 vssd1 vccd1 vccd1 _0951_ sky130_fd_sc_hd__mux2_1
X_2264_ LE_1B.config_data\[5\] _0961_ _0987_ _1019_ vssd1 vssd1 vccd1 vccd1 _1020_
+ sky130_fd_sc_hd__a211oi_1
XANTENNA__2130__A1 _0822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2116__X _0874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout233_A net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1979_ net23 net24 net25 net26 net162 CB_0.config_dataB\[13\] vssd1 vssd1 vccd1 vccd1
+ _0739_ sky130_fd_sc_hd__mux4_1
Xhold23 _0052_ vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 LE_0B.config_data\[9\] vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 _0085_ vssd1 vssd1 vccd1 vccd1 net328 sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 _0075_ vssd1 vssd1 vccd1 vccd1 net317 sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 _0309_ vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 _0032_ vssd1 vssd1 vccd1 vccd1 net361 sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 LE_0B.config_data\[3\] vssd1 vssd1 vccd1 vccd1 net350 sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 _0319_ vssd1 vssd1 vccd1 vccd1 net339 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_16_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_9 CBeast_in[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1902_ _0659_ _0661_ CB_0.config_dataB\[6\] vssd1 vssd1 vccd1 vccd1 _0662_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_32_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2951_ clknet_leaf_28_clk _0159_ net195 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[23\]
+ sky130_fd_sc_hd__dfstp_1
X_1833_ CB_0.config_dataA\[8\] _0359_ _0594_ vssd1 vssd1 vccd1 vccd1 _0595_ sky130_fd_sc_hd__o21ai_1
XANTENNA__1926__A1 _0447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_0_clk_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2882_ clknet_leaf_29_clk _0090_ net187 vssd1 vssd1 vccd1 vccd1 LE_0B.edge_mode sky130_fd_sc_hd__dfstp_1
X_1764_ net131 _1281_ _0457_ _0460_ _1284_ vssd1 vssd1 vccd1 vccd1 _0526_ sky130_fd_sc_hd__o32a_1
XPHY_EDGE_ROW_27_Left_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2351__A1 CB_1.config_dataB\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2316_ net59 LE_0B.edge_mode vssd1 vssd1 vccd1 vccd1 LE_0B.sel_clk sky130_fd_sc_hd__xnor2_1
X_1695_ net176 net175 vssd1 vssd1 vccd1 vccd1 _0457_ sky130_fd_sc_hd__nand2b_1
X_2247_ CB_1.config_dataB\[9\] CB_1.config_dataB\[11\] vssd1 vssd1 vccd1 vccd1 _1003_
+ sky130_fd_sc_hd__nand2_1
X_2178_ _1240_ LE_1A.dff_out vssd1 vssd1 vccd1 vccd1 _0935_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_11_Left_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1917__A1 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput79 net79 vssd1 vssd1 vccd1 vccd1 CBnorth_out[11] sky130_fd_sc_hd__buf_2
Xoutput68 net68 vssd1 vssd1 vccd1 vccd1 CBeast_out[1] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_46_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_2_clk_A clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_19_Right_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1908__A1 net24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1480_ CB_0.config_dataA\[16\] CB_0.config_dataA\[17\] vssd1 vssd1 vccd1 vccd1 _1274_
+ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_28_Right_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1687__A3 _0430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3081_ clknet_leaf_14_clk _0289_ net223 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[1\]
+ sky130_fd_sc_hd__dfstp_2
XPHY_EDGE_ROW_37_Right_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2101_ net2 net3 net151 vssd1 vssd1 vccd1 vccd1 _0859_ sky130_fd_sc_hd__mux2_1
X_2032_ SB0.route_sel\[36\] SB0.route_sel\[37\] vssd1 vssd1 vccd1 vccd1 _0790_ sky130_fd_sc_hd__nor2_1
X_2934_ clknet_leaf_27_clk _0142_ net195 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[6\]
+ sky130_fd_sc_hd__dfstp_1
X_2865_ clknet_leaf_30_clk _0073_ net190 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_1816_ _0577_ vssd1 vssd1 vccd1 vccd1 _0578_ sky130_fd_sc_hd__inv_2
X_2796_ clknet_leaf_5_clk _0004_ net203 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_46_Right_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1747_ SB0.route_sel\[90\] SB0.route_sel\[91\] vssd1 vssd1 vccd1 vccd1 _0509_ sky130_fd_sc_hd__nor2_1
X_1678_ SB0.route_sel\[19\] SB0.route_sel\[18\] _0436_ _0437_ _0439_ vssd1 vssd1 vccd1
+ vccd1 _0440_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_55_Right_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2023__Y _0781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output115_A net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2174__S0 _0848_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1532_ net124 net23 _1323_ vssd1 vssd1 vccd1 vccd1 _1326_ sky130_fd_sc_hd__mux2_1
X_1601_ net18 net19 net174 vssd1 vssd1 vccd1 vccd1 _0363_ sky130_fd_sc_hd__mux2_1
X_2581_ CB_1.config_dataB\[1\] CB_1.config_dataB\[0\] net257 vssd1 vssd1 vccd1 vccd1
+ _0117_ sky130_fd_sc_hd__mux2_1
XANTENNA__1766__A net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2650_ SB0.route_sel\[50\] SB0.route_sel\[49\] net258 vssd1 vssd1 vccd1 vccd1 _0186_
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1394_ SB0.route_sel\[59\] vssd1 vssd1 vccd1 vccd1 _1188_ sky130_fd_sc_hd__inv_2
X_1463_ net177 net178 vssd1 vssd1 vccd1 vccd1 _1257_ sky130_fd_sc_hd__nand2_1
X_3064_ clknet_leaf_3_clk _0272_ net208 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[4\]
+ sky130_fd_sc_hd__dfstp_1
X_2015_ _0734_ _0764_ _0768_ _0774_ vssd1 vssd1 vccd1 vccd1 _0775_ sky130_fd_sc_hd__o22a_1
X_2848_ clknet_leaf_6_clk _0056_ net204 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_2917_ clknet_leaf_15_clk _0125_ net222 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[9\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_12_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold142 LEI0.config_data\[18\] vssd1 vssd1 vccd1 vccd1 net414 sky130_fd_sc_hd__dlygate4sd3_1
Xhold120 LE_1A.config_data\[10\] vssd1 vssd1 vccd1 vccd1 net392 sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 LE_1A.config_data\[9\] vssd1 vssd1 vccd1 vccd1 net403 sky130_fd_sc_hd__dlygate4sd3_1
X_2779_ net347 net344 net235 vssd1 vssd1 vccd1 vccd1 _0315_ sky130_fd_sc_hd__mux2_1
XFILLER_58_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2233__B1 _0984_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input31_X net31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2702_ SB0.route_sel\[102\] SB0.route_sel\[101\] net264 vssd1 vssd1 vccd1 vccd1 _0238_
+ sky130_fd_sc_hd__mux2_1
X_2495_ net371 net354 net269 vssd1 vssd1 vccd1 vccd1 _0034_ sky130_fd_sc_hd__mux2_1
X_2633_ SB0.route_sel\[33\] SB0.route_sel\[32\] net238 vssd1 vssd1 vccd1 vccd1 _0169_
+ sky130_fd_sc_hd__mux2_1
X_2564_ net291 net278 net260 vssd1 vssd1 vccd1 vccd1 _0100_ sky130_fd_sc_hd__mux2_1
X_1515_ net144 net145 vssd1 vssd1 vccd1 vccd1 _1309_ sky130_fd_sc_hd__nand2b_1
XANTENNA__2828__Q LEI0.config_data\[35\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1446_ LE_1A.config_data\[16\] vssd1 vssd1 vccd1 vccd1 _1240_ sky130_fd_sc_hd__inv_2
X_1377_ SB0.route_sel\[27\] vssd1 vssd1 vccd1 vccd1 _1171_ sky130_fd_sc_hd__inv_2
X_3116_ clknet_leaf_30_clk _0324_ net187 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_3047_ clknet_leaf_7_clk _0255_ net206 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[7\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_fanout263_A net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2205__A _0957_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2280_ CB_1.config_dataB\[15\] _1034_ _1035_ _1028_ vssd1 vssd1 vccd1 vccd1 _1036_
+ sky130_fd_sc_hd__o22ai_1
X_1995_ net161 _0539_ _0743_ _0749_ _0754_ vssd1 vssd1 vccd1 vccd1 _0755_ sky130_fd_sc_hd__o311a_1
X_2616_ SB0.route_sel\[16\] SB0.route_sel\[15\] net231 vssd1 vssd1 vccd1 vccd1 _0152_
+ sky130_fd_sc_hd__mux2_1
X_2478_ net374 LEI0.config_data\[15\] net244 vssd1 vssd1 vccd1 vccd1 _0017_ sky130_fd_sc_hd__mux2_1
X_2547_ LE_0B.config_data\[11\] net300 net243 vssd1 vssd1 vccd1 vccd1 _0084_ sky130_fd_sc_hd__mux2_1
X_1429_ LE_0A.config_data\[16\] vssd1 vssd1 vccd1 vccd1 _1223_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_38_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload1 clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload1/X sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_21_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout271 net272 vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input39_A SBsouth_in[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout260 net261 vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__clkbuf_4
X_1780_ _0519_ _0541_ CB_0.config_dataA\[2\] vssd1 vssd1 vccd1 vccd1 _0542_ sky130_fd_sc_hd__a21o_1
XFILLER_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2332_ net137 _1072_ _0451_ vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__mux2_1
X_2401_ SB0.route_sel\[43\] SB0.route_sel\[42\] vssd1 vssd1 vccd1 vccd1 _1111_ sky130_fd_sc_hd__nand2b_1
XANTENNA__3054__SET_B net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2194_ net13 net14 CB_1.config_dataB\[0\] vssd1 vssd1 vccd1 vccd1 _0950_ sky130_fd_sc_hd__mux2_1
X_2263_ LE_1B.config_data\[4\] net120 net135 vssd1 vssd1 vccd1 vccd1 _1019_ sky130_fd_sc_hd__and3_1
XANTENNA__2130__A2 _0816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1978_ net161 _0359_ _0737_ vssd1 vssd1 vccd1 vccd1 _0738_ sky130_fd_sc_hd__o21a_1
Xhold68 LE_0A.config_data\[3\] vssd1 vssd1 vccd1 vccd1 net340 sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 LEI0.config_data\[3\] vssd1 vssd1 vccd1 vccd1 net329 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 LEI0.config_data\[5\] vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 _0082_ vssd1 vssd1 vccd1 vccd1 net307 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 _0077_ vssd1 vssd1 vccd1 vccd1 net351 sky130_fd_sc_hd__dlygate4sd3_1
Xhold13 LEI0.config_data\[23\] vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold46 LE_1B.config_data\[14\] vssd1 vssd1 vccd1 vccd1 net318 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_24_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2409__B1 _1342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1578__B _0339_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1832_ net170 _0339_ _0588_ vssd1 vssd1 vccd1 vccd1 _0594_ sky130_fd_sc_hd__a21oi_1
X_1901_ CB_0.config_dataB\[7\] _0656_ _0660_ _0654_ vssd1 vssd1 vccd1 vccd1 _0661_
+ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_32_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2881_ clknet_leaf_0_clk _0089_ net199 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[16\]
+ sky130_fd_sc_hd__dfrtp_2
X_2950_ clknet_leaf_28_clk _0158_ net189 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[22\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__1935__C _1297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1763_ _1280_ _0456_ net2 vssd1 vssd1 vccd1 vccd1 _0525_ sky130_fd_sc_hd__a21o_1
XANTENNA__2179__A2 _0934_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1694_ net176 net175 vssd1 vssd1 vccd1 vccd1 _0456_ sky130_fd_sc_hd__and2b_2
X_2246_ CB_1.config_dataB\[11\] _1000_ _1001_ _0991_ vssd1 vssd1 vccd1 vccd1 _1002_
+ sky130_fd_sc_hd__o22ai_1
X_2315_ net186 LE_0B.reset_mode vssd1 vssd1 vccd1 vccd1 _2315_/X sky130_fd_sc_hd__xor2_2
XANTENNA__1862__A1 _0430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2177_ LE_1A.dff0_out LE_1A.dff1_out LE_1A.reset_val vssd1 vssd1 vccd1 vccd1 LE_1A.dff_out
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout229_X net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1685__Y _0447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput69 net69 vssd1 vssd1 vccd1 vccd1 CBeast_out[2] sky130_fd_sc_hd__buf_2
XFILLER_0_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1908__A2 net25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3080_ clknet_leaf_14_clk _0288_ net225 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_2100_ _0852_ _0857_ vssd1 vssd1 vccd1 vccd1 _0858_ sky130_fd_sc_hd__or2_1
X_2031_ _0785_ _0786_ _0787_ _1294_ vssd1 vssd1 vccd1 vccd1 _0789_ sky130_fd_sc_hd__o31ai_2
X_1815_ _1217_ net170 vssd1 vssd1 vccd1 vccd1 _0577_ sky130_fd_sc_hd__nor2_1
X_2795_ clknet_leaf_5_clk net321 net199 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_2864_ LE_1A.sel_clk _0072_ net61 vssd1 vssd1 vccd1 vccd1 LE_1A.dff1_out sky130_fd_sc_hd__dfstp_1
X_2933_ clknet_leaf_28_clk _0141_ net195 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[5\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_15_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1746_ _0497_ _0498_ _0502_ _0507_ vssd1 vssd1 vccd1 vccd1 _0508_ sky130_fd_sc_hd__a22o_1
X_1677_ net128 _1283_ _0379_ vssd1 vssd1 vccd1 vccd1 _0439_ sky130_fd_sc_hd__and3_1
X_2229_ net136 net122 net130 net134 LEI0.config_data\[21\] LEI0.config_data\[22\]
+ vssd1 vssd1 vccd1 vccd1 _0985_ sky130_fd_sc_hd__mux4_1
XFILLER_53_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1599__A0 net23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input21_A CBnorth_in[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2174__S1 _0874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1462_ net138 _1254_ _1252_ vssd1 vssd1 vccd1 vccd1 _1256_ sky130_fd_sc_hd__mux2_1
X_1531_ _1251_ _1324_ vssd1 vssd1 vccd1 vccd1 _1325_ sky130_fd_sc_hd__nand2_1
XANTENNA__1762__A0 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1600_ CB_0.config_dataA\[3\] _0361_ vssd1 vssd1 vccd1 vccd1 _0362_ sky130_fd_sc_hd__or2_1
X_2580_ CB_1.config_dataB\[0\] CB_1.config_dataA\[19\] net257 vssd1 vssd1 vccd1 vccd1
+ _0116_ sky130_fd_sc_hd__mux2_1
X_3063_ clknet_leaf_3_clk _0271_ net208 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[3\]
+ sky130_fd_sc_hd__dfstp_1
X_1393_ SB0.route_sel\[49\] vssd1 vssd1 vccd1 vccd1 _1187_ sky130_fd_sc_hd__inv_2
X_2014_ _0730_ _0773_ _0758_ vssd1 vssd1 vccd1 vccd1 _0774_ sky130_fd_sc_hd__a21o_1
X_2847_ clknet_leaf_6_clk _0055_ net204 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_2916_ clknet_leaf_16_clk _0124_ net222 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[8\]
+ sky130_fd_sc_hd__dfstp_1
Xhold110 _0029_ vssd1 vssd1 vccd1 vccd1 net382 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_2_1__f_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2778_ net344 LE_1B.config_data\[5\] net235 vssd1 vssd1 vccd1 vccd1 _0314_ sky130_fd_sc_hd__mux2_1
Xhold132 LEI0.config_data\[43\] vssd1 vssd1 vccd1 vccd1 net404 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1753__A0 net27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1729_ SB0.route_sel\[76\] _1195_ SB0.route_sel\[79\] _1197_ _0490_ vssd1 vssd1 vccd1
+ vccd1 _0491_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_1_clk_A clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold121 _0105_ vssd1 vssd1 vccd1 vccd1 net393 sky130_fd_sc_hd__dlygate4sd3_1
Xhold143 LE_0A.reset_val vssd1 vssd1 vccd1 vccd1 net415 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_56_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1992__A0 net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input24_X net24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2701_ SB0.route_sel\[101\] SB0.route_sel\[100\] net264 vssd1 vssd1 vccd1 vccd1 _0237_
+ sky130_fd_sc_hd__mux2_1
X_2632_ SB0.route_sel\[32\] SB0.route_sel\[31\] net238 vssd1 vssd1 vccd1 vccd1 _0168_
+ sky130_fd_sc_hd__mux2_1
X_2494_ net354 LEI0.config_data\[31\] net269 vssd1 vssd1 vccd1 vccd1 _0033_ sky130_fd_sc_hd__mux2_1
X_1445_ LEI0.config_data\[44\] vssd1 vssd1 vccd1 vccd1 _1239_ sky130_fd_sc_hd__inv_2
X_2563_ net278 LE_1A.config_data\[3\] net260 vssd1 vssd1 vccd1 vccd1 _0099_ sky130_fd_sc_hd__mux2_1
X_1514_ net144 net145 vssd1 vssd1 vccd1 vccd1 _1308_ sky130_fd_sc_hd__and2b_1
X_3046_ clknet_leaf_7_clk _0254_ net206 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[6\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_2_149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1376_ SB0.route_sel\[16\] vssd1 vssd1 vccd1 vccd1 _1170_ sky130_fd_sc_hd__inv_2
X_3115_ clknet_leaf_30_clk _0323_ net189 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2463__A1 LEI0.config_data\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2151__A0 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2205__B _0960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1717__A0 net28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1994_ CB_0.config_dataB\[15\] _0750_ _0753_ vssd1 vssd1 vccd1 vccd1 _0754_ sky130_fd_sc_hd__o21ai_1
XANTENNA__1956__A0 _0430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload30 clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 clkload30/Y sky130_fd_sc_hd__inv_8
X_2615_ SB0.route_sel\[15\] SB0.route_sel\[14\] net231 vssd1 vssd1 vccd1 vccd1 _0151_
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1428_ CB_0.config_dataA\[14\] vssd1 vssd1 vccd1 vccd1 _1222_ sky130_fd_sc_hd__inv_2
X_2477_ net412 net386 net248 vssd1 vssd1 vccd1 vccd1 _0016_ sky130_fd_sc_hd__mux2_1
X_2546_ net300 net306 net243 vssd1 vssd1 vccd1 vccd1 _0083_ sky130_fd_sc_hd__mux2_1
XANTENNA__2133__A0 net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3029_ clknet_leaf_15_clk _0237_ net220 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[101\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_38_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload2 clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload2/X sky130_fd_sc_hd__clkbuf_8
XFILLER_11_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout272 net58 vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__buf_2
Xfanout250 net254 vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout261 net262 vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__clkbuf_4
XFILLER_42_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2400_ _1294_ _1110_ vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__and2_1
X_2331_ net123 _0473_ _0452_ vssd1 vssd1 vccd1 vccd1 _1072_ sky130_fd_sc_hd__mux2_1
X_2262_ _1017_ vssd1 vssd1 vccd1 vccd1 _1018_ sky130_fd_sc_hd__inv_2
X_2193_ net1 net6 net7 net8 CB_1.config_dataB\[0\] CB_1.config_dataB\[1\] vssd1 vssd1
+ vccd1 vccd1 _0949_ sky130_fd_sc_hd__mux4_1
XANTENNA__2130__A3 _0813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1977_ net161 _0339_ _0736_ vssd1 vssd1 vccd1 vccd1 _0737_ sky130_fd_sc_hd__a21oi_1
X_2529_ LE_0A.config_data\[16\] net343 net242 vssd1 vssd1 vccd1 vccd1 _0067_ sky130_fd_sc_hd__mux2_1
Xhold69 LE_0A.config_data\[11\] vssd1 vssd1 vccd1 vccd1 net341 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 LE_0A.config_data\[14\] vssd1 vssd1 vccd1 vccd1 net308 sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 _0006_ vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 LE_0A.config_data\[13\] vssd1 vssd1 vccd1 vccd1 net319 sky130_fd_sc_hd__dlygate4sd3_1
Xhold14 _0025_ vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold58 LE_1B.config_data\[3\] vssd1 vssd1 vccd1 vccd1 net330 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_43_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2345__A0 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input51_A SBwest_in[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1871__A2 _0606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1831_ CB_0.config_dataA\[11\] _0591_ _0592_ _0588_ vssd1 vssd1 vccd1 vccd1 _0593_
+ sky130_fd_sc_hd__o22a_1
X_1900_ net16 net17 net165 vssd1 vssd1 vccd1 vccd1 _0660_ sky130_fd_sc_hd__mux2_1
X_2880_ clknet_leaf_4_clk _0088_ net199 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_15_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1762_ net141 _0522_ _0520_ vssd1 vssd1 vccd1 vccd1 _0524_ sky130_fd_sc_hd__mux2_1
X_1693_ net137 _0453_ _0451_ vssd1 vssd1 vccd1 vccd1 _0455_ sky130_fd_sc_hd__mux2_1
X_2245_ net4 net5 net182 vssd1 vssd1 vccd1 vccd1 _1001_ sky130_fd_sc_hd__mux2_1
X_2314_ LE_0A.edge_mode net59 vssd1 vssd1 vccd1 vccd1 LE_0A.sel_clk sky130_fd_sc_hd__xnor2_1
X_2176_ _0930_ _0933_ _0928_ vssd1 vssd1 vccd1 vccd1 _0934_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_1_Right_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1853__A2 _0359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1908__A3 net26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input54_X net54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2030_ _0785_ _0786_ _0787_ _1294_ vssd1 vssd1 vccd1 vccd1 _0788_ sky130_fd_sc_hd__o31a_2
XTAP_TAPCELL_ROW_45_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2228__X _0984_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2932_ clknet_leaf_27_clk _0140_ net195 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[4\]
+ sky130_fd_sc_hd__dfstp_1
X_1814_ net121 _0430_ _1218_ vssd1 vssd1 vccd1 vccd1 _0576_ sky130_fd_sc_hd__mux2_1
X_2794_ clknet_leaf_5_clk _0002_ net199 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1745_ _0504_ _0506_ _0497_ vssd1 vssd1 vccd1 vccd1 _0507_ sky130_fd_sc_hd__a21oi_1
X_2863_ LE_0B.sel_clk _0071_ net61 vssd1 vssd1 vccd1 vccd1 LE_0B.dff0_out sky130_fd_sc_hd__dfrtp_1
XFILLER_15_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1676_ SB0.route_sel\[19\] SB0.route_sel\[18\] vssd1 vssd1 vccd1 vccd1 _0438_ sky130_fd_sc_hd__nand2_1
XANTENNA__1532__A1 net23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1835__A2 _1321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2228_ _0965_ _0971_ _0982_ _0983_ vssd1 vssd1 vccd1 vccd1 _0984_ sky130_fd_sc_hd__a211o_2
X_2159_ net1 net6 net7 net8 net147 CB_1.config_dataA\[13\] vssd1 vssd1 vccd1 vccd1
+ _0917_ sky130_fd_sc_hd__mux4_1
XFILLER_53_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1599__A1 net24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input14_A CBeast_in[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_24_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1530_ CB_0.config_dataA\[17\] CB_0.config_dataA\[16\] vssd1 vssd1 vccd1 vccd1 _1324_
+ sky130_fd_sc_hd__nor2_1
X_1461_ SB0.route_sel\[57\] SB0.route_sel\[56\] vssd1 vssd1 vccd1 vccd1 _1255_ sky130_fd_sc_hd__nand2_1
X_1392_ SB0.route_sel\[52\] vssd1 vssd1 vccd1 vccd1 _1186_ sky130_fd_sc_hd__inv_2
XANTENNA__2711__A0 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3062_ clknet_leaf_3_clk _0270_ net202 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[2\]
+ sky130_fd_sc_hd__dfstp_1
X_2013_ _0676_ _0771_ _0772_ _0769_ _0770_ vssd1 vssd1 vccd1 vccd1 _0773_ sky130_fd_sc_hd__o32a_1
Xclkbuf_leaf_15_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2915_ clknet_leaf_16_clk _0123_ net220 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[7\]
+ sky130_fd_sc_hd__dfstp_1
X_2846_ clknet_leaf_6_clk _0054_ net203 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold100 LE_0A.config_data\[10\] vssd1 vssd1 vccd1 vccd1 net372 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1753__A1 net28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold111 LEI0.config_data\[1\] vssd1 vssd1 vccd1 vccd1 net383 sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 LEI0.config_data\[25\] vssd1 vssd1 vccd1 vccd1 net394 sky130_fd_sc_hd__dlygate4sd3_1
X_1728_ SB0.route_sel\[74\] SB0.route_sel\[75\] vssd1 vssd1 vccd1 vccd1 _0490_ sky130_fd_sc_hd__nor2_1
X_2777_ LE_1B.config_data\[5\] net325 net235 vssd1 vssd1 vccd1 vccd1 _0313_ sky130_fd_sc_hd__mux2_1
Xhold133 LE_0B.reset_val vssd1 vssd1 vccd1 vccd1 net405 sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 LE_0B.config_data\[0\] vssd1 vssd1 vccd1 vccd1 net416 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input6_A CBeast_in[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1659_ net128 _1332_ _0379_ vssd1 vssd1 vccd1 vccd1 _0421_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_56_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1992__A1 net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input17_X net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2700_ SB0.route_sel\[100\] SB0.route_sel\[99\] net264 vssd1 vssd1 vccd1 vccd1 _0236_
+ sky130_fd_sc_hd__mux2_1
X_2631_ SB0.route_sel\[31\] SB0.route_sel\[30\] net237 vssd1 vssd1 vccd1 vccd1 _0167_
+ sky130_fd_sc_hd__mux2_1
X_2562_ net313 net305 net259 vssd1 vssd1 vccd1 vccd1 _0098_ sky130_fd_sc_hd__mux2_1
XANTENNA__1496__C net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2493_ net360 LEI0.config_data\[30\] net269 vssd1 vssd1 vccd1 vccd1 _0032_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_4_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1444_ CB_1.config_dataA\[7\] vssd1 vssd1 vccd1 vccd1 _1238_ sky130_fd_sc_hd__inv_2
X_1375_ SB0.route_sel\[22\] vssd1 vssd1 vccd1 vccd1 _1169_ sky130_fd_sc_hd__inv_2
X_1513_ _1258_ _1305_ net10 vssd1 vssd1 vccd1 vccd1 _1307_ sky130_fd_sc_hd__a21o_1
X_3045_ clknet_leaf_7_clk _0253_ net206 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[5\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_55_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3114_ clknet_leaf_30_clk _0322_ net191 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__1671__A0 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout249_A net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2829_ clknet_leaf_13_clk _0037_ net226 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[36\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input9_X net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2151__A1 net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1965__A1 _0512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1993_ _0736_ _0751_ _0752_ _0743_ vssd1 vssd1 vccd1 vccd1 _0753_ sky130_fd_sc_hd__o22a_1
XANTENNA__1788__A net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1956__A1 _0447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_0_clk_A clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2545_ net306 LE_0B.config_data\[8\] net243 vssd1 vssd1 vccd1 vccd1 _0082_ sky130_fd_sc_hd__mux2_1
XANTENNA__2131__B _0831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2614_ SB0.route_sel\[14\] SB0.route_sel\[13\] net231 vssd1 vssd1 vccd1 vccd1 _0150_
+ sky130_fd_sc_hd__mux2_1
Xclkload20 clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 clkload20/Y sky130_fd_sc_hd__inv_6
X_2476_ net386 net364 net248 vssd1 vssd1 vccd1 vccd1 _0015_ sky130_fd_sc_hd__mux2_1
X_1427_ net169 vssd1 vssd1 vccd1 vccd1 _1221_ sky130_fd_sc_hd__inv_2
XFILLER_28_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2133__A1 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3028_ clknet_leaf_10_clk _0236_ net220 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[100\]
+ sky130_fd_sc_hd__dfstp_1
Xclkload3 clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 clkload3/Y sky130_fd_sc_hd__clkinv_2
XFILLER_11_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout240 net241 vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__clkbuf_4
Xfanout251 net253 vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__clkbuf_4
Xfanout262 net58 vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__buf_2
XANTENNA__1635__A0 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_3__f_clk_X clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2330_ net138 _0477_ _0478_ _1071_ vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__a22o_1
X_2261_ _1005_ _1014_ _1016_ LEI0.config_data\[35\] vssd1 vssd1 vccd1 vccd1 _1017_
+ sky130_fd_sc_hd__o22a_2
X_2192_ CB_1.config_dataB\[3\] _0947_ vssd1 vssd1 vccd1 vccd1 _0948_ sky130_fd_sc_hd__or2_1
XFILLER_52_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1976_ CB_0.config_dataB\[13\] _1233_ vssd1 vssd1 vccd1 vccd1 _0736_ sky130_fd_sc_hd__or2_1
X_2528_ net343 net308 net246 vssd1 vssd1 vccd1 vccd1 _0066_ sky130_fd_sc_hd__mux2_1
Xhold26 LE_0A.config_data\[7\] vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 _0065_ vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 LEI0.config_data\[2\] vssd1 vssd1 vccd1 vccd1 net320 sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 LE_0B.config_data\[13\] vssd1 vssd1 vccd1 vccd1 net331 sky130_fd_sc_hd__dlygate4sd3_1
X_2459_ SB0.route_sel\[87\] SB0.route_sel\[86\] _1202_ SB0.route_sel\[80\] vssd1 vssd1
+ vccd1 vccd1 _1150_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_26_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold15 LE_1B.config_data\[8\] vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_10_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input44_A SBwest_in[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1830_ net18 net19 CB_0.config_dataA\[8\] vssd1 vssd1 vccd1 vccd1 _0592_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_40_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1761_ SB0.route_sel\[81\] SB0.route_sel\[80\] vssd1 vssd1 vccd1 vccd1 _0523_ sky130_fd_sc_hd__nand2_1
X_2313_ net190 LE_0A.reset_mode vssd1 vssd1 vccd1 vccd1 _2313_/X sky130_fd_sc_hd__xor2_2
X_1692_ SB0.route_sel\[65\] SB0.route_sel\[64\] vssd1 vssd1 vccd1 vccd1 _0454_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_48_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2244_ net9 net10 net11 net12 net182 CB_1.config_dataB\[9\] vssd1 vssd1 vccd1 vccd1
+ _1000_ sky130_fd_sc_hd__mux4_1
X_2175_ _0932_ _0931_ _0901_ vssd1 vssd1 vccd1 vccd1 _0933_ sky130_fd_sc_hd__mux2_1
X_1959_ net163 _0473_ _0718_ vssd1 vssd1 vccd1 vccd1 _0719_ sky130_fd_sc_hd__o21a_1
XANTENNA__2575__A1 LE_1A.config_data\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1829__A0 net23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input47_X net47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2254__A0 net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clknet_0_clk sky130_fd_sc_hd__clkbuf_16
X_2931_ clknet_leaf_27_clk _0139_ net194 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[3\]
+ sky130_fd_sc_hd__dfstp_1
X_1813_ LEI0.config_data\[26\] _0574_ vssd1 vssd1 vccd1 vccd1 _0575_ sky130_fd_sc_hd__and2b_1
X_1744_ SB0.route_sel\[90\] SB0.route_sel\[91\] _0505_ vssd1 vssd1 vccd1 vccd1 _0506_
+ sky130_fd_sc_hd__and3_1
X_2862_ clknet_leaf_0_clk _0070_ net192 vssd1 vssd1 vccd1 vccd1 LE_0A.reset_mode sky130_fd_sc_hd__dfrtp_1
X_2793_ clknet_leaf_29_clk _0001_ net186 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_15_Left_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1675_ net131 _1281_ _0377_ _0380_ _1284_ vssd1 vssd1 vccd1 vccd1 _0437_ sky130_fd_sc_hd__o32a_1
XPHY_EDGE_ROW_15_Right_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2227_ _0979_ _0980_ _0981_ _0975_ CB_1.config_dataB\[6\] vssd1 vssd1 vccd1 vccd1
+ _0983_ sky130_fd_sc_hd__o311a_1
X_2089_ net136 net122 net130 net134 LEI0.config_data\[18\] LEI0.config_data\[19\]
+ vssd1 vssd1 vccd1 vccd1 _0847_ sky130_fd_sc_hd__mux4_2
XPHY_EDGE_ROW_24_Right_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2158_ net147 _0831_ _0915_ vssd1 vssd1 vccd1 vccd1 _0916_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_51_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1599__A2 net25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2245__A0 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2154__X _0912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_33_Right_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_42_Right_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_51_Right_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1460_ net26 net123 _1253_ vssd1 vssd1 vccd1 vccd1 _1254_ sky130_fd_sc_hd__mux2_1
X_1391_ SB0.route_sel\[50\] vssd1 vssd1 vccd1 vccd1 _1185_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_60_Right_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2012_ _0700_ _0702_ LE_0B.config_data\[11\] vssd1 vssd1 vccd1 vccd1 _0772_ sky130_fd_sc_hd__a21boi_1
X_3061_ clknet_leaf_3_clk _0269_ net202 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[1\]
+ sky130_fd_sc_hd__dfstp_1
X_2845_ clknet_leaf_7_clk _0053_ net206 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_2914_ clknet_leaf_16_clk _0122_ net219 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[6\]
+ sky130_fd_sc_hd__dfstp_1
Xhold134 LEI0.config_data\[44\] vssd1 vssd1 vccd1 vccd1 net406 sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 LEI0.config_data\[27\] vssd1 vssd1 vccd1 vccd1 net384 sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 _0026_ vssd1 vssd1 vccd1 vccd1 net395 sky130_fd_sc_hd__dlygate4sd3_1
X_2776_ net325 net330 net236 vssd1 vssd1 vccd1 vccd1 _0312_ sky130_fd_sc_hd__mux2_1
X_1727_ _0475_ _0480_ _0485_ _0488_ vssd1 vssd1 vccd1 vccd1 _0489_ sky130_fd_sc_hd__a22o_2
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1658_ net131 _1330_ _0377_ _0380_ _1333_ vssd1 vssd1 vccd1 vccd1 _0420_ sky130_fd_sc_hd__o32a_1
XANTENNA__2421__Y net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold101 LE_1B.config_data\[10\] vssd1 vssd1 vccd1 vccd1 net373 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_56_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1589_ _0346_ _0348_ _0349_ _0350_ vssd1 vssd1 vccd1 vccd1 _0351_ sky130_fd_sc_hd__a211o_1
XANTENNA__2218__A0 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output113_A net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2492_ net398 LEI0.config_data\[29\] net269 vssd1 vssd1 vccd1 vccd1 _0031_ sky130_fd_sc_hd__mux2_1
X_2630_ SB0.route_sel\[30\] SB0.route_sel\[29\] net237 vssd1 vssd1 vccd1 vccd1 _0166_
+ sky130_fd_sc_hd__mux2_1
X_2561_ net305 net304 net259 vssd1 vssd1 vccd1 vccd1 _0097_ sky130_fd_sc_hd__mux2_1
X_1512_ net177 net178 vssd1 vssd1 vccd1 vccd1 _1306_ sky130_fd_sc_hd__nand2b_2
X_1443_ net150 vssd1 vssd1 vccd1 vccd1 _1237_ sky130_fd_sc_hd__inv_2
X_1374_ SB0.route_sel\[23\] vssd1 vssd1 vccd1 vccd1 _1168_ sky130_fd_sc_hd__inv_2
X_3113_ clknet_leaf_30_clk _0321_ net190 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__1671__A1 net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3044_ clknet_leaf_7_clk _0252_ net205 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[4\]
+ sky130_fd_sc_hd__dfstp_1
X_2828_ clknet_leaf_13_clk _0036_ net226 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[35\]
+ sky130_fd_sc_hd__dfrtp_1
X_2759_ CB_1.config_dataA\[7\] CB_1.config_dataA\[6\] net262 vssd1 vssd1 vccd1 vccd1
+ _0295_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_18_Left_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_45_Left_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_54_Left_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2061__Y _0819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_63_Left_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1992_ net16 net17 net161 vssd1 vssd1 vccd1 vccd1 _0752_ sky130_fd_sc_hd__mux2_1
Xclkload10 clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 clkload10/Y sky130_fd_sc_hd__inv_12
X_2475_ net364 LEI0.config_data\[12\] net248 vssd1 vssd1 vccd1 vccd1 _0014_ sky130_fd_sc_hd__mux2_1
X_2544_ net348 LE_0B.config_data\[7\] net243 vssd1 vssd1 vccd1 vccd1 _0081_ sky130_fd_sc_hd__mux2_1
X_2613_ SB0.route_sel\[13\] SB0.route_sel\[12\] net231 vssd1 vssd1 vccd1 vccd1 _0149_
+ sky130_fd_sc_hd__mux2_1
Xclkload21 clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 clkload21/Y sky130_fd_sc_hd__clkinvlp_4
X_1426_ net168 vssd1 vssd1 vccd1 vccd1 _1220_ sky130_fd_sc_hd__inv_2
XANTENNA__2133__A2 net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3027_ clknet_leaf_9_clk _0235_ net219 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[99\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout261_A net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2427__X net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload4 clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 clkload4/Y sky130_fd_sc_hd__bufinv_16
Xfanout263 net272 vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__clkbuf_4
Xfanout252 net253 vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__clkbuf_2
Xfanout241 net254 vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_3_Left_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout230 net233 vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__clkbuf_4
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2260_ _1015_ vssd1 vssd1 vccd1 vccd1 _1016_ sky130_fd_sc_hd__inv_2
X_2191_ _0813_ _0816_ _0822_ _0819_ _1241_ _1242_ vssd1 vssd1 vccd1 vccd1 _0947_ sky130_fd_sc_hd__mux4_1
XFILLER_60_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1975_ _1345_ _1321_ _1297_ _1273_ net161 CB_0.config_dataB\[13\] vssd1 vssd1 vccd1
+ vccd1 _0735_ sky130_fd_sc_hd__mux4_1
Xhold27 _0058_ vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__dlygate4sd3_1
X_2527_ net308 LE_0A.config_data\[13\] net246 vssd1 vssd1 vccd1 vccd1 _0065_ sky130_fd_sc_hd__mux2_1
X_2458_ SB0.route_sel\[82\] _1199_ vssd1 vssd1 vccd1 vccd1 _1149_ sky130_fd_sc_hd__nor2_1
X_1409_ SB0.route_sel\[91\] vssd1 vssd1 vccd1 vccd1 _1203_ sky130_fd_sc_hd__inv_2
Xhold38 LE_1A.config_data\[7\] vssd1 vssd1 vccd1 vccd1 net310 sky130_fd_sc_hd__dlygate4sd3_1
Xhold16 _0316_ vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 _0003_ vssd1 vssd1 vccd1 vccd1 net321 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2511__C1 net60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2389_ SB0.route_sel\[57\] SB0.route_sel\[56\] vssd1 vssd1 vccd1 vccd1 _1103_ sky130_fd_sc_hd__nor2_1
XFILLER_10_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1856__A1 _1297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1856__B2 _1273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input37_A SBsouth_in[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1760_ net16 net123 _0521_ vssd1 vssd1 vccd1 vccd1 _0522_ sky130_fd_sc_hd__mux2_1
X_1691_ net123 net27 _0452_ vssd1 vssd1 vccd1 vccd1 _0453_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_40_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2312_ LE_1B.config_data\[16\] _1065_ _1066_ _0646_ vssd1 vssd1 vccd1 vccd1 CB_1.le_outB
+ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_48_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2243_ CB_1.config_dataB\[9\] _0997_ _0998_ _0993_ _0996_ vssd1 vssd1 vccd1 vccd1
+ _0999_ sky130_fd_sc_hd__a32o_1
X_2174_ LE_1A.config_data\[13\] LE_1A.config_data\[15\] LE_1A.config_data\[12\] LE_1A.config_data\[14\]
+ _0848_ _0874_ vssd1 vssd1 vccd1 vccd1 _0932_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_31_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1958_ net163 _0493_ _0707_ vssd1 vssd1 vccd1 vccd1 _0718_ sky130_fd_sc_hd__a21oi_1
X_1889_ net121 _0430_ _0391_ _0447_ _1228_ CB_0.config_dataB\[5\] vssd1 vssd1 vccd1
+ vccd1 _0649_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_54_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1503__Y _1297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1407__A net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1829__A1 net24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload2_A clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_6_Left_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2254__A1 net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2861_ clknet_leaf_0_clk _0069_ net190 vssd1 vssd1 vccd1 vccd1 LE_0A.reset_val sky130_fd_sc_hd__dfrtp_1
X_2930_ clknet_leaf_27_clk _0138_ net194 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[2\]
+ sky130_fd_sc_hd__dfstp_1
X_1812_ net136 net122 net130 net134 LEI0.config_data\[24\] LEI0.config_data\[25\]
+ vssd1 vssd1 vccd1 vccd1 _0574_ sky130_fd_sc_hd__mux4_1
X_2792_ LE_0A.sel_clk _0000_ net61 vssd1 vssd1 vccd1 vccd1 LE_0A.dff1_out sky130_fd_sc_hd__dfstp_1
X_1743_ SB0.route_sel\[92\] SB0.route_sel\[93\] net31 vssd1 vssd1 vccd1 vccd1 _0505_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_7_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1674_ _1280_ _0376_ net7 vssd1 vssd1 vccd1 vccd1 _0436_ sky130_fd_sc_hd__a21o_1
X_2226_ net184 _1244_ CB_1.config_dataB\[6\] net183 vssd1 vssd1 vccd1 vccd1 _0982_
+ sky130_fd_sc_hd__and4_1
XFILLER_53_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout174_A CB_0.config_dataA\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3040__Q CB_0.config_dataA\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2245__A1 net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2088_ _0799_ _0832_ _0845_ _0824_ vssd1 vssd1 vccd1 vccd1 _0846_ sky130_fd_sc_hd__a211o_1
X_2157_ net147 _0828_ _0905_ vssd1 vssd1 vccd1 vccd1 _0915_ sky130_fd_sc_hd__a21oi_1
XANTENNA__1599__A3 net26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1508__A0 net24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2757__S net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_32_Left_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2064__Y _0822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3060_ clknet_leaf_10_clk _0268_ net221 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_1390_ SB0.route_sel\[51\] vssd1 vssd1 vccd1 vccd1 _1184_ sky130_fd_sc_hd__inv_2
X_2011_ LE_0B.config_data\[10\] _0700_ _0702_ vssd1 vssd1 vccd1 vccd1 _0771_ sky130_fd_sc_hd__and3_1
X_2844_ clknet_leaf_6_clk net295 net206 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_2913_ clknet_leaf_16_clk _0121_ net220 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[5\]
+ sky130_fd_sc_hd__dfstp_1
Xhold135 LEI0.config_data\[45\] vssd1 vssd1 vccd1 vccd1 net407 sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 LEI0.config_data\[17\] vssd1 vssd1 vccd1 vccd1 net385 sky130_fd_sc_hd__dlygate4sd3_1
Xhold102 LEI0.config_data\[16\] vssd1 vssd1 vccd1 vccd1 net374 sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 LEI0.config_data\[20\] vssd1 vssd1 vccd1 vccd1 net396 sky130_fd_sc_hd__dlygate4sd3_1
X_2775_ net330 net324 net236 vssd1 vssd1 vccd1 vccd1 _0311_ sky130_fd_sc_hd__mux2_1
X_1726_ _0483_ _0486_ _0487_ _0475_ vssd1 vssd1 vccd1 vccd1 _0488_ sky130_fd_sc_hd__a31oi_1
X_1657_ _1329_ _0376_ net1 vssd1 vssd1 vccd1 vccd1 _0419_ sky130_fd_sc_hd__a21o_1
X_1588_ _1249_ _0347_ vssd1 vssd1 vccd1 vccd1 _0350_ sky130_fd_sc_hd__nor2_1
XANTENNA__1910__A0 net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2209_ net183 _0964_ vssd1 vssd1 vccd1 vccd1 _0965_ sky130_fd_sc_hd__or2_1
XANTENNA__2218__A1 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_4_160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_2_0__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_2_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__1968__A0 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output106_A net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2491_ LEI0.config_data\[29\] net381 net251 vssd1 vssd1 vccd1 vccd1 _0030_ sky130_fd_sc_hd__mux2_1
X_1442_ LEI0.config_data\[20\] vssd1 vssd1 vccd1 vccd1 _1236_ sky130_fd_sc_hd__inv_2
X_2560_ net304 LE_1A.config_data\[0\] net259 vssd1 vssd1 vccd1 vccd1 _0096_ sky130_fd_sc_hd__mux2_1
X_1511_ CB_1.config_dataB\[17\] CB_1.config_dataB\[16\] vssd1 vssd1 vccd1 vccd1 _1305_
+ sky130_fd_sc_hd__and2b_1
X_3043_ clknet_leaf_5_clk _0251_ net205 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[3\]
+ sky130_fd_sc_hd__dfstp_2
X_1373_ SB0.route_sel\[21\] vssd1 vssd1 vccd1 vccd1 _1167_ sky130_fd_sc_hd__inv_2
X_3112_ clknet_leaf_30_clk net277 net190 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_18_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2827_ clknet_leaf_13_clk _0035_ net226 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[34\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2758_ CB_1.config_dataA\[6\] CB_1.config_dataA\[5\] net261 vssd1 vssd1 vccd1 vccd1
+ _0294_ sky130_fd_sc_hd__mux2_1
X_2689_ SB0.route_sel\[89\] SB0.route_sel\[88\] net240 vssd1 vssd1 vccd1 vccd1 _0225_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__2136__A0 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1709_ SB0.route_sel\[67\] SB0.route_sel\[66\] vssd1 vssd1 vccd1 vccd1 _0471_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_1_141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2375__B1 _0819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input22_X net22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1991_ net27 net28 net161 vssd1 vssd1 vccd1 vccd1 _0751_ sky130_fd_sc_hd__mux2_1
XANTENNA__1956__A3 _0391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload11 clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 clkload11/Y sky130_fd_sc_hd__clkinv_2
Xclkload22 clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 clkload22/Y sky130_fd_sc_hd__inv_4
X_2612_ SB0.route_sel\[12\] SB0.route_sel\[11\] net231 vssd1 vssd1 vccd1 vccd1 _0148_
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1425_ CB_0.config_dataA\[10\] vssd1 vssd1 vccd1 vccd1 _1219_ sky130_fd_sc_hd__inv_2
X_2474_ net408 LEI0.config_data\[11\] net248 vssd1 vssd1 vccd1 vccd1 _0013_ sky130_fd_sc_hd__mux2_1
X_2543_ net353 net311 net243 vssd1 vssd1 vccd1 vccd1 _0080_ sky130_fd_sc_hd__mux2_1
X_3026_ clknet_leaf_9_clk _0234_ net219 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[98\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__2133__A3 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout254_A net58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload5 clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 clkload5/Y sky130_fd_sc_hd__inv_6
XFILLER_50_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout253 net254 vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__clkbuf_2
Xfanout242 net245 vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__clkbuf_4
Xfanout220 net228 vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__clkbuf_4
Xfanout264 net272 vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__buf_2
XANTENNA__2765__S net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout231 net233 vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_29_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2190_ CB_1.config_dataB\[0\] _0945_ CB_1.config_dataB\[2\] vssd1 vssd1 vccd1 vccd1
+ _0946_ sky130_fd_sc_hd__o21ai_1
X_1974_ _0675_ _0704_ _0732_ _0733_ _0731_ vssd1 vssd1 vccd1 vccd1 _0734_ sky130_fd_sc_hd__o221a_1
XANTENNA__1626__A2 _0375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2526_ net319 net314 net246 vssd1 vssd1 vccd1 vccd1 _0064_ sky130_fd_sc_hd__mux2_1
Xhold28 LE_0B.config_data\[10\] vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 LE_0B.config_data\[6\] vssd1 vssd1 vccd1 vccd1 net311 sky130_fd_sc_hd__dlygate4sd3_1
X_2457_ _0534_ _1148_ vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__and2_1
X_1408_ SB0.route_sel\[81\] vssd1 vssd1 vccd1 vccd1 _1202_ sky130_fd_sc_hd__inv_2
X_2388_ _1101_ _1102_ _0469_ vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__a21boi_1
Xhold17 LE_1A.config_data\[12\] vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__dlygate4sd3_1
X_3009_ clknet_leaf_2_clk _0217_ net208 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[81\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_26_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1690_ net157 net159 net155 net153 vssd1 vssd1 vccd1 vccd1 _0452_ sky130_fd_sc_hd__or4b_1
XANTENNA__1792__B2 net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1792__A1 net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2242_ _1245_ _0788_ vssd1 vssd1 vccd1 vccd1 _0998_ sky130_fd_sc_hd__nand2_1
X_2311_ _1246_ LE_1B.dff_out vssd1 vssd1 vccd1 vccd1 _1066_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_48_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2173_ LE_1A.config_data\[9\] LE_1A.config_data\[11\] LE_1A.config_data\[8\] LE_1A.config_data\[10\]
+ _0848_ _0874_ vssd1 vssd1 vccd1 vccd1 _0931_ sky130_fd_sc_hd__mux4_1
X_1957_ CB_0.config_dataB\[11\] _0716_ vssd1 vssd1 vccd1 vccd1 _0717_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_31_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2732__A0 CB_0.config_dataB\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2509_ net397 net369 net269 vssd1 vssd1 vccd1 vccd1 _0048_ sky130_fd_sc_hd__mux2_1
X_1888_ net136 net122 net130 net134 LEI0.config_data\[15\] LEI0.config_data\[16\]
+ vssd1 vssd1 vccd1 vccd1 _0648_ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout217_A net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1560__B1_N net47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1829__A2 net25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2238__B _1318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_27_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1811_ LE_0A.config_data\[7\] LE_0A.config_data\[6\] _0543_ vssd1 vssd1 vccd1 vccd1
+ _0573_ sky130_fd_sc_hd__mux2_1
X_2860_ clknet_leaf_0_clk _0068_ net190 vssd1 vssd1 vccd1 vccd1 LE_0A.edge_mode sky130_fd_sc_hd__dfstp_1
X_2791_ LE_1B.reset_mode net400 net233 vssd1 vssd1 vccd1 vccd1 _0327_ sky130_fd_sc_hd__mux2_1
X_1673_ net136 _0433_ _0431_ vssd1 vssd1 vccd1 vccd1 _0435_ sky130_fd_sc_hd__mux2_1
X_1742_ SB0.route_sel\[95\] SB0.route_sel\[94\] _0503_ vssd1 vssd1 vccd1 vccd1 _0504_
+ sky130_fd_sc_hd__a21bo_1
X_2225_ net184 _0976_ _0977_ net183 vssd1 vssd1 vccd1 vccd1 _0981_ sky130_fd_sc_hd__o31a_1
XFILLER_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout167_A CB_0.config_dataB\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1987__B _0473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2087_ CB_1.config_dataA\[5\] net150 CB_1.config_dataA\[7\] _0835_ _0844_ vssd1 vssd1
+ vccd1 vccd1 _0845_ sky130_fd_sc_hd__a41o_1
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_18_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_clk
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_5_Right_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2156_ CB_1.config_dataA\[15\] _0913_ vssd1 vssd1 vccd1 vccd1 _0914_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_51_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout122_X net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2989_ clknet_leaf_23_clk _0197_ net211 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[61\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_8_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2080__Y _0838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input52_X net52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2010_ LE_0B.config_data\[8\] _0700_ _0702_ _0675_ vssd1 vssd1 vccd1 vccd1 _0770_
+ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_7_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2912_ clknet_leaf_16_clk _0120_ net219 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[4\]
+ sky130_fd_sc_hd__dfstp_1
X_2843_ clknet_leaf_6_clk _0051_ net203 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__1986__A1 _0430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2774_ net324 net283 net236 vssd1 vssd1 vccd1 vccd1 _0310_ sky130_fd_sc_hd__mux2_1
X_1725_ SB0.route_sel\[76\] SB0.route_sel\[77\] net42 vssd1 vssd1 vccd1 vccd1 _0487_
+ sky130_fd_sc_hd__a21bo_1
Xclkbuf_leaf_7_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_clk
+ sky130_fd_sc_hd__clkbuf_8
Xhold114 LEI0.config_data\[14\] vssd1 vssd1 vccd1 vccd1 net386 sky130_fd_sc_hd__dlygate4sd3_1
Xhold136 LEI0.config_data\[12\] vssd1 vssd1 vccd1 vccd1 net408 sky130_fd_sc_hd__dlygate4sd3_1
Xhold125 CB_0.config_data_inA vssd1 vssd1 vccd1 vccd1 net397 sky130_fd_sc_hd__dlygate4sd3_1
X_1656_ net141 _0417_ _0415_ vssd1 vssd1 vccd1 vccd1 _0418_ sky130_fd_sc_hd__mux2_1
Xhold103 _0017_ vssd1 vssd1 vccd1 vccd1 net375 sky130_fd_sc_hd__dlygate4sd3_1
X_1587_ SB0.route_sel\[98\] SB0.route_sel\[99\] vssd1 vssd1 vccd1 vccd1 _0349_ sky130_fd_sc_hd__and2_1
XANTENNA__1910__A1 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2208_ _0816_ _0819_ _0813_ _0822_ _1244_ net184 vssd1 vssd1 vccd1 vccd1 _0964_ sky130_fd_sc_hd__mux4_1
X_2139_ _0835_ net148 vssd1 vssd1 vccd1 vccd1 _0897_ sky130_fd_sc_hd__nand2b_1
XANTENNA__1674__B1 net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2218__A2 net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2768__S net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input12_A CBeast_in[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1701__A net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1968__A1 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2090__B1 _0847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1510_ net139 _1302_ _1299_ vssd1 vssd1 vccd1 vccd1 _1304_ sky130_fd_sc_hd__mux2_2
X_1441_ CB_1.config_dataA\[3\] vssd1 vssd1 vccd1 vccd1 _1235_ sky130_fd_sc_hd__inv_2
X_2490_ net381 LEI0.config_data\[27\] net251 vssd1 vssd1 vccd1 vccd1 _0029_ sky130_fd_sc_hd__mux2_1
XANTENNA__1656__A0 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3042_ clknet_leaf_5_clk _0250_ net205 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[2\]
+ sky130_fd_sc_hd__dfstp_1
X_1372_ SB0.route_sel\[18\] vssd1 vssd1 vccd1 vccd1 _1166_ sky130_fd_sc_hd__inv_2
X_3111_ clknet_leaf_31_clk net339 net190 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_61_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2081__A0 net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2826_ clknet_leaf_13_clk _0034_ net226 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[33\]
+ sky130_fd_sc_hd__dfrtp_1
X_2688_ SB0.route_sel\[88\] SB0.route_sel\[87\] net252 vssd1 vssd1 vccd1 vccd1 _0224_
+ sky130_fd_sc_hd__mux2_1
X_2757_ CB_1.config_dataA\[5\] CB_1.config_dataA\[4\] net261 vssd1 vssd1 vccd1 vccd1
+ _0293_ sky130_fd_sc_hd__mux2_1
X_1708_ _1193_ SB0.route_sel\[70\] vssd1 vssd1 vccd1 vccd1 _0470_ sky130_fd_sc_hd__nor2_1
XANTENNA_input4_A CBeast_in[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2136__A1 net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1639_ SB0.route_sel\[11\] SB0.route_sel\[10\] _0398_ _0399_ _0400_ vssd1 vssd1 vccd1
+ vccd1 _0401_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_1_142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2176__X _0934_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input15_X net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1990_ net15 net20 net21 net22 net161 CB_0.config_dataB\[13\] vssd1 vssd1 vccd1 vccd1
+ _0750_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_15_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload12 clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 clkload12/X sky130_fd_sc_hd__clkbuf_4
X_2542_ net311 LE_0B.config_data\[5\] net242 vssd1 vssd1 vccd1 vccd1 _0079_ sky130_fd_sc_hd__mux2_1
XANTENNA__2262__A _1017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2611_ SB0.route_sel\[11\] SB0.route_sel\[10\] net238 vssd1 vssd1 vccd1 vccd1 _0147_
+ sky130_fd_sc_hd__mux2_1
Xclkload23 clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 clkload23/Y sky130_fd_sc_hd__clkinv_8
X_1424_ net170 vssd1 vssd1 vccd1 vccd1 _1218_ sky130_fd_sc_hd__inv_2
X_2473_ LEI0.config_data\[11\] net380 net264 vssd1 vssd1 vccd1 vccd1 _0012_ sky130_fd_sc_hd__mux2_1
X_3025_ clknet_leaf_9_clk _0233_ net219 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[97\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_36_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout247_A net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload6 clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 clkload6/Y sky130_fd_sc_hd__clkinvlp_4
X_2809_ clknet_leaf_5_clk net375 net201 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[16\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout221 net228 vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__clkbuf_4
Xfanout265 net272 vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__clkbuf_4
Xfanout210 net229 vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__clkbuf_2
Xfanout254 net58 vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__buf_2
Xfanout243 net245 vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input7_X net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout232 net233 vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_37_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2284__A0 net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2036__B1 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1973_ LE_0B.config_data\[7\] _0703_ _0676_ vssd1 vssd1 vccd1 vccd1 _0733_ sky130_fd_sc_hd__a21o_1
XANTENNA__2339__A1 _1345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2525_ net314 LE_0A.config_data\[11\] net246 vssd1 vssd1 vccd1 vccd1 _0063_ sky130_fd_sc_hd__mux2_1
Xhold29 _0084_ vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__dlygate4sd3_1
X_1407_ net2 vssd1 vssd1 vccd1 vccd1 _1201_ sky130_fd_sc_hd__inv_2
X_2456_ SB0.route_sel\[82\] _1199_ _1200_ SB0.route_sel\[85\] _1147_ vssd1 vssd1 vccd1
+ vccd1 _1148_ sky130_fd_sc_hd__a221o_1
X_2387_ _1191_ SB0.route_sel\[66\] SB0.route_sel\[65\] _1194_ vssd1 vssd1 vccd1 vccd1
+ _1102_ sky130_fd_sc_hd__o22a_1
Xhold18 _0107_ vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__dlygate4sd3_1
X_3008_ clknet_leaf_1_clk _0216_ net196 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[80\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_26_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2266__B1 _0984_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2241_ net182 _0781_ vssd1 vssd1 vccd1 vccd1 _0997_ sky130_fd_sc_hd__nand2_1
X_2172_ _0902_ _0929_ _0901_ vssd1 vssd1 vccd1 vccd1 _0930_ sky130_fd_sc_hd__mux2_1
X_2310_ LE_1B.dff0_out LE_1B.dff1_out LE_1B.reset_val vssd1 vssd1 vccd1 vccd1 LE_1B.dff_out
+ sky130_fd_sc_hd__mux2_1
X_1956_ _0430_ _0447_ net121 _0391_ CB_0.config_dataB\[9\] net163 vssd1 vssd1 vccd1
+ vccd1 _0716_ sky130_fd_sc_hd__mux4_1
X_1887_ LE_0A.config_data\[16\] _0645_ _0646_ _0647_ vssd1 vssd1 vccd1 vccd1 CB_0.le_outA
+ sky130_fd_sc_hd__o211a_1
XANTENNA__1743__B1_N net31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2508_ net369 LEI0.config_data\[45\] net269 vssd1 vssd1 vccd1 vccd1 _0047_ sky130_fd_sc_hd__mux2_1
XANTENNA__2596__S net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2439_ _1136_ _0336_ vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_54_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1829__A3 net26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input42_A SBsouth_in[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1810_ _1215_ _0560_ _0571_ _0559_ vssd1 vssd1 vccd1 vccd1 _0572_ sky130_fd_sc_hd__a211o_1
X_1741_ SB0.route_sel\[92\] SB0.route_sel\[93\] net45 vssd1 vssd1 vccd1 vccd1 _0503_
+ sky130_fd_sc_hd__and3_1
XFILLER_7_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2790_ net400 LE_1B.edge_mode net233 vssd1 vssd1 vccd1 vccd1 _0326_ sky130_fd_sc_hd__mux2_1
XFILLER_7_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1672_ SB0.route_sel\[17\] SB0.route_sel\[16\] vssd1 vssd1 vccd1 vccd1 _0434_ sky130_fd_sc_hd__nand2_1
X_2224_ _0781_ _0962_ _0963_ _0789_ vssd1 vssd1 vccd1 vccd1 _0980_ sky130_fd_sc_hd__a2bb2o_1
X_2155_ _0819_ _0822_ _0816_ _0813_ CB_1.config_dataA\[13\] net146 vssd1 vssd1 vccd1
+ vccd1 _0913_ sky130_fd_sc_hd__mux4_1
X_2086_ _0778_ _0838_ _0843_ CB_1.config_dataA\[6\] vssd1 vssd1 vccd1 vccd1 _0844_
+ sky130_fd_sc_hd__a211o_1
X_1939_ net166 _1225_ CB_0.config_dataB\[3\] vssd1 vssd1 vccd1 vccd1 _0699_ sky130_fd_sc_hd__and3_1
X_2988_ clknet_leaf_23_clk _0196_ net211 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[60\]
+ sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_11_Right_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_20_Right_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2089__X _0847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input45_X net45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1986__A2 _0391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2911_ clknet_leaf_16_clk _0119_ net213 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[3\]
+ sky130_fd_sc_hd__dfstp_2
Xhold115 LEI0.config_data\[37\] vssd1 vssd1 vccd1 vccd1 net387 sky130_fd_sc_hd__dlygate4sd3_1
Xhold104 LE_0A.config_data\[6\] vssd1 vssd1 vccd1 vccd1 net376 sky130_fd_sc_hd__dlygate4sd3_1
Xhold126 LEI0.config_data\[30\] vssd1 vssd1 vccd1 vccd1 net398 sky130_fd_sc_hd__dlygate4sd3_1
X_1724_ _1196_ _1197_ net56 SB0.route_sel\[77\] SB0.route_sel\[76\] vssd1 vssd1 vccd1
+ vccd1 _0486_ sky130_fd_sc_hd__o2111ai_1
X_2773_ net283 LE_1B.config_data\[0\] net236 vssd1 vssd1 vccd1 vccd1 _0309_ sky130_fd_sc_hd__mux2_1
X_2842_ LE_0B.sel_clk _0050_ net61 vssd1 vssd1 vccd1 vccd1 LE_0B.dff1_out sky130_fd_sc_hd__dfstp_1
Xhold137 LEI0.config_data\[36\] vssd1 vssd1 vccd1 vccd1 net409 sky130_fd_sc_hd__dlygate4sd3_1
X_1655_ net127 net15 _0414_ vssd1 vssd1 vccd1 vccd1 _0417_ sky130_fd_sc_hd__mux2_1
X_1586_ net131 _1330_ _1348_ _0347_ vssd1 vssd1 vccd1 vccd1 _0348_ sky130_fd_sc_hd__o31a_1
X_2207_ CB_1.config_dataB\[5\] _1244_ vssd1 vssd1 vccd1 vccd1 _0963_ sky130_fd_sc_hd__and2_1
X_2069_ _0489_ _0826_ vssd1 vssd1 vccd1 vccd1 _0827_ sky130_fd_sc_hd__and2_1
X_2138_ _0877_ _0893_ _0895_ _0892_ vssd1 vssd1 vccd1 vccd1 _0896_ sky130_fd_sc_hd__o211a_1
XANTENNA__1977__A2 _0339_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2218__A3 net12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1968__A2 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2090__B2 _1236_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2372__X net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1371_ net174 vssd1 vssd1 vccd1 vccd1 _1165_ sky130_fd_sc_hd__inv_2
X_1440_ LE_0B.config_data\[16\] vssd1 vssd1 vccd1 vccd1 _1234_ sky130_fd_sc_hd__inv_2
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3110_ clknet_leaf_31_clk _0318_ net190 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_3041_ clknet_leaf_5_clk _0249_ net205 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[1\]
+ sky130_fd_sc_hd__dfstp_2
XTAP_TAPCELL_ROW_61_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2825_ clknet_leaf_13_clk net355 net225 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[32\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__1959__A2 _0473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2081__A1 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2687_ SB0.route_sel\[87\] SB0.route_sel\[86\] net251 vssd1 vssd1 vccd1 vccd1 _0223_
+ sky130_fd_sc_hd__mux2_1
X_2756_ net150 CB_1.config_dataA\[3\] net261 vssd1 vssd1 vccd1 vccd1 _0292_ sky130_fd_sc_hd__mux2_1
X_1707_ _0468_ _0464_ _0455_ _0454_ vssd1 vssd1 vccd1 vccd1 _0469_ sky130_fd_sc_hd__a2bb2o_1
X_1638_ net128 _1308_ _0379_ vssd1 vssd1 vccd1 vccd1 _0400_ sky130_fd_sc_hd__and3_1
X_1569_ net154 net156 _1248_ _1300_ vssd1 vssd1 vccd1 vccd1 _0331_ sky130_fd_sc_hd__nand4_1
XANTENNA__2457__X net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output111_A net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2472_ net380 LEI0.config_data\[9\] net263 vssd1 vssd1 vccd1 vccd1 _0011_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_41_Left_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload24 clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 clkload24/Y sky130_fd_sc_hd__bufinv_16
Xclkload13 clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 clkload13/Y sky130_fd_sc_hd__bufinv_16
X_2541_ net357 LE_0B.config_data\[4\] net242 vssd1 vssd1 vccd1 vccd1 _0078_ sky130_fd_sc_hd__mux2_1
X_2610_ SB0.route_sel\[10\] SB0.route_sel\[9\] net238 vssd1 vssd1 vccd1 vccd1 _0146_
+ sky130_fd_sc_hd__mux2_1
X_1423_ CB_0.config_dataA\[9\] vssd1 vssd1 vccd1 vccd1 _1217_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_50_Left_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3024_ clknet_leaf_9_clk _0232_ net219 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[96\]
+ sky130_fd_sc_hd__dfstp_1
X_2808_ clknet_leaf_5_clk _0016_ net205 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload7 clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 clkload7/Y sky130_fd_sc_hd__bufinv_16
Xfanout200 net202 vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__clkbuf_2
Xfanout222 net228 vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__clkbuf_4
X_2739_ CB_0.config_dataB\[7\] CB_0.config_dataB\[6\] net252 vssd1 vssd1 vccd1 vccd1
+ _0275_ sky130_fd_sc_hd__mux2_1
Xfanout211 net213 vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__clkbuf_4
Xfanout266 net272 vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__clkbuf_4
Xfanout244 net245 vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_29_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout233 net254 vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__clkbuf_2
Xfanout255 net257 vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_12_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2284__A1 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1972_ LE_0B.config_data\[6\] _0700_ _0702_ vssd1 vssd1 vccd1 vccd1 _0732_ sky130_fd_sc_hd__and3_1
X_2524_ net341 LE_0A.config_data\[10\] net246 vssd1 vssd1 vccd1 vccd1 _0062_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_49_Right_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2455_ SB0.route_sel\[81\] SB0.route_sel\[80\] vssd1 vssd1 vccd1 vccd1 _1147_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_58_Right_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1406_ SB0.route_sel\[84\] vssd1 vssd1 vccd1 vccd1 _1200_ sky130_fd_sc_hd__inv_2
Xhold19 LE_1A.config_data\[5\] vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__dlygate4sd3_1
X_2386_ SB0.route_sel\[71\] SB0.route_sel\[70\] vssd1 vssd1 vccd1 vccd1 _1101_ sky130_fd_sc_hd__or2_1
XFILLER_51_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3007_ clknet_leaf_1_clk _0215_ net196 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[79\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_24_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1527__A _1318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2240_ _0994_ _0995_ CB_1.config_dataB\[11\] vssd1 vssd1 vccd1 vccd1 _0996_ sky130_fd_sc_hd__a21o_1
X_2171_ LE_1A.config_data\[1\] LE_1A.config_data\[3\] LE_1A.config_data\[0\] LE_1A.config_data\[2\]
+ _0848_ _0874_ vssd1 vssd1 vccd1 vccd1 _0929_ sky130_fd_sc_hd__mux4_1
XANTENNA__2257__A1 _0831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1955_ CB_0.config_dataB\[10\] _0714_ vssd1 vssd1 vccd1 vccd1 _0715_ sky130_fd_sc_hd__nand2_1
X_1886_ _1223_ LE_0A.dff_out vssd1 vssd1 vccd1 vccd1 _0647_ sky130_fd_sc_hd__or2_1
X_2507_ net407 net406 net269 vssd1 vssd1 vccd1 vccd1 _0046_ sky130_fd_sc_hd__mux2_1
X_2438_ SB0.route_sel\[108\] _1211_ SB0.route_sel\[104\] SB0.route_sel\[105\] _1135_
+ vssd1 vssd1 vccd1 vccd1 _1136_ sky130_fd_sc_hd__o221a_1
XANTENNA__2193__A0 net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout262_X net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2369_ _1257_ _0377_ _0813_ vssd1 vssd1 vccd1 vccd1 _1091_ sky130_fd_sc_hd__o21ai_1
XFILLER_24_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input35_A SBsouth_in[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1671_ net127 net21 _0432_ vssd1 vssd1 vccd1 vccd1 _0433_ sky130_fd_sc_hd__mux2_1
XFILLER_30_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1740_ SB0.route_sel\[90\] SB0.route_sel\[91\] _0499_ _0500_ _0501_ vssd1 vssd1 vccd1
+ vccd1 _0502_ sky130_fd_sc_hd__a221o_1
XANTENNA__1630__A _0391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2154_ net139 net126 net129 net133 LEI0.config_data\[42\] LEI0.config_data\[43\]
+ vssd1 vssd1 vccd1 vccd1 _0912_ sky130_fd_sc_hd__mux4_2
X_2223_ net185 _0784_ _0978_ vssd1 vssd1 vccd1 vccd1 _0979_ sky130_fd_sc_hd__a21oi_1
X_2085_ _0800_ _0840_ _0842_ vssd1 vssd1 vccd1 vccd1 _0843_ sky130_fd_sc_hd__o21a_1
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2987_ clknet_leaf_22_clk _0195_ net212 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[59\]
+ sky130_fd_sc_hd__dfstp_1
X_1869_ _0622_ _0623_ _0625_ _0627_ vssd1 vssd1 vccd1 vccd1 _0631_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout222_A net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1938_ _0692_ _0697_ CB_0.config_dataB\[2\] vssd1 vssd1 vccd1 vccd1 _0698_ sky130_fd_sc_hd__o21a_1
XANTENNA__2469__A1 LEI0.config_data\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload0_A clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1986__A3 _0447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2910_ clknet_leaf_17_clk _0118_ net213 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[2\]
+ sky130_fd_sc_hd__dfstp_1
X_2841_ LE_0A.sel_clk _0049_ net61 vssd1 vssd1 vccd1 vccd1 LE_0A.dff0_out sky130_fd_sc_hd__dfrtp_1
Xhold116 _0038_ vssd1 vssd1 vccd1 vccd1 net388 sky130_fd_sc_hd__dlygate4sd3_1
Xhold105 _0057_ vssd1 vssd1 vccd1 vccd1 net377 sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 LEI0.config_data\[41\] vssd1 vssd1 vccd1 vccd1 net410 sky130_fd_sc_hd__dlygate4sd3_1
X_1654_ net122 _0414_ vssd1 vssd1 vccd1 vccd1 _0416_ sky130_fd_sc_hd__nor2_1
Xhold127 LEI0.config_data\[8\] vssd1 vssd1 vccd1 vccd1 net399 sky130_fd_sc_hd__dlygate4sd3_1
X_2772_ net356 LE_0A.reset_mode net236 vssd1 vssd1 vccd1 vccd1 _0308_ sky130_fd_sc_hd__mux2_1
X_1723_ _0481_ _0482_ _0483_ _0484_ vssd1 vssd1 vccd1 vccd1 _0485_ sky130_fd_sc_hd__a211o_1
XFILLER_7_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2206_ net184 net185 vssd1 vssd1 vccd1 vccd1 _0962_ sky130_fd_sc_hd__nand2_1
X_1585_ net144 net145 net142 net143 vssd1 vssd1 vccd1 vccd1 _0347_ sky130_fd_sc_hd__or4bb_1
X_2068_ _1196_ SB0.route_sel\[78\] SB0.route_sel\[73\] _1198_ _0825_ vssd1 vssd1 vccd1
+ vccd1 _0826_ sky130_fd_sc_hd__a221o_1
X_2137_ _0883_ _0894_ vssd1 vssd1 vccd1 vccd1 _0895_ sky130_fd_sc_hd__or2_1
XFILLER_5_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2154__A3 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1665__A2 _0418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1968__A3 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1370_ SB0.route_sel\[8\] vssd1 vssd1 vccd1 vccd1 _1164_ sky130_fd_sc_hd__inv_2
XFILLER_4_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2145__A3 _0781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3040_ clknet_leaf_13_clk _0248_ net225 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[0\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_18_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2824_ clknet_leaf_13_clk net361 net225 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2369__B1 _0813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2081__A2 net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2755_ CB_1.config_dataA\[3\] CB_1.config_dataA\[2\] net267 vssd1 vssd1 vccd1 vccd1
+ _0291_ sky130_fd_sc_hd__mux2_1
X_2686_ SB0.route_sel\[86\] SB0.route_sel\[85\] net251 vssd1 vssd1 vccd1 vccd1 _0222_
+ sky130_fd_sc_hd__mux2_1
X_1637_ net131 _1306_ _0377_ _0380_ _1309_ vssd1 vssd1 vccd1 vccd1 _0399_ sky130_fd_sc_hd__o32a_1
X_1706_ _0462_ _0466_ _0467_ _0454_ vssd1 vssd1 vccd1 vccd1 _0468_ sky130_fd_sc_hd__a31o_1
XFILLER_58_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1568_ _0329_ CB_0.config_dataA\[17\] CB_0.config_dataA\[16\] vssd1 vssd1 vccd1 vccd1
+ _0330_ sky130_fd_sc_hd__or3b_1
X_1499_ _1287_ _1291_ _1292_ _1278_ vssd1 vssd1 vccd1 vccd1 _1293_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_1_144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1422_ CB_0.config_dataA\[7\] vssd1 vssd1 vccd1 vccd1 _1216_ sky130_fd_sc_hd__inv_2
Xclkload14 clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 clkload14/Y sky130_fd_sc_hd__clkinv_2
X_2471_ LEI0.config_data\[9\] net399 net266 vssd1 vssd1 vccd1 vccd1 _0010_ sky130_fd_sc_hd__mux2_1
Xclkload25 clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 clkload25/Y sky130_fd_sc_hd__clkinvlp_4
X_2540_ LE_0B.config_data\[4\] net350 net244 vssd1 vssd1 vccd1 vccd1 _0077_ sky130_fd_sc_hd__mux2_1
XANTENNA__1462__X _1256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3023_ clknet_leaf_9_clk _0231_ net219 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[95\]
+ sky130_fd_sc_hd__dfstp_1
X_2807_ clknet_leaf_6_clk _0015_ net205 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_2738_ CB_0.config_dataB\[6\] CB_0.config_dataB\[5\] net252 vssd1 vssd1 vccd1 vccd1
+ _0274_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout135_A _0960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload8 clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 clkload8/Y sky130_fd_sc_hd__inv_6
XFILLER_59_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout245 net250 vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__clkbuf_2
Xfanout201 net202 vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__clkbuf_4
Xfanout223 net228 vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__clkbuf_2
Xfanout234 net236 vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__clkbuf_4
Xfanout212 net213 vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__buf_2
Xfanout256 net257 vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__buf_2
X_2669_ SB0.route_sel\[69\] SB0.route_sel\[68\] net239 vssd1 vssd1 vccd1 vccd1 _0205_
+ sky130_fd_sc_hd__mux2_1
Xfanout267 net272 vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_29_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input20_X net20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2284__A2 net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_23_Left_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1971_ _0730_ vssd1 vssd1 vccd1 vccd1 _0731_ sky130_fd_sc_hd__inv_2
X_2523_ net372 net332 net246 vssd1 vssd1 vccd1 vccd1 _0061_ sky130_fd_sc_hd__mux2_1
X_1405_ SB0.route_sel\[83\] vssd1 vssd1 vccd1 vccd1 _1199_ sky130_fd_sc_hd__inv_2
X_2454_ _1145_ _1146_ _0508_ vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__o21a_1
X_2385_ _0469_ _1100_ vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__and2_1
Xinput1 CBeast_in[0] vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_26_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3006_ clknet_leaf_1_clk _0214_ net192 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[78\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__1483__A0 net25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1527__B _1320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1453__A net60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2170_ _0925_ _0926_ _0927_ _0912_ _1239_ vssd1 vssd1 vccd1 vccd1 _0928_ sky130_fd_sc_hd__a32o_1
X_1954_ net163 _0705_ _0709_ _0713_ vssd1 vssd1 vccd1 vccd1 _0714_ sky130_fd_sc_hd__a2bb2o_1
X_1885_ LE_0A.dff0_out LE_0A.dff1_out LE_0A.reset_val vssd1 vssd1 vccd1 vccd1 LE_0A.dff_out
+ sky130_fd_sc_hd__mux2_1
XANTENNA__2717__A0 net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2193__A1 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2506_ net406 net404 net269 vssd1 vssd1 vccd1 vccd1 _0045_ sky130_fd_sc_hd__mux2_1
X_2437_ SB0.route_sel\[107\] SB0.route_sel\[106\] vssd1 vssd1 vccd1 vccd1 _1135_ sky130_fd_sc_hd__nand2b_1
X_2368_ _1335_ _1090_ _1337_ vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__a21o_1
X_2299_ LE_1B.config_data\[14\] net120 net135 _0984_ _0986_ vssd1 vssd1 vccd1 vccd1
+ _1055_ sky130_fd_sc_hd__a32o_1
XFILLER_21_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input28_A CBnorth_in[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2239__A2 _1342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2391__X net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1670_ net159 net153 net155 net157 vssd1 vssd1 vccd1 vccd1 _0432_ sky130_fd_sc_hd__or4b_1
XFILLER_7_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2222_ _1244_ _1342_ _0791_ CB_1.config_dataB\[7\] CB_1.config_dataB\[5\] vssd1 vssd1
+ vccd1 vccd1 _0978_ sky130_fd_sc_hd__a311o_1
X_2084_ CB_1.config_dataA\[7\] _0839_ _0841_ _0777_ vssd1 vssd1 vccd1 vccd1 _0842_
+ sky130_fd_sc_hd__o22a_1
X_2153_ CB_1.config_dataA\[13\] CB_1.config_dataA\[15\] vssd1 vssd1 vccd1 vccd1 _0911_
+ sky130_fd_sc_hd__nand2_1
X_1937_ _0694_ _0695_ _0696_ _1226_ vssd1 vssd1 vccd1 vccd1 _0697_ sky130_fd_sc_hd__o31a_1
XPHY_EDGE_ROW_26_Left_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2986_ clknet_leaf_23_clk _0194_ net212 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[58\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__1629__Y _0391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1799_ net18 net19 net172 vssd1 vssd1 vccd1 vccd1 _0561_ sky130_fd_sc_hd__mux2_1
X_1868_ _0628_ _0629_ CB_0.config_dataA\[15\] vssd1 vssd1 vccd1 vccd1 _0630_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout215_A net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_10_Left_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1601__A0 net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_19_clk_A clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2840_ clknet_leaf_14_clk _0048_ net225 vssd1 vssd1 vccd1 vccd1 CB_0.config_data_inA
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2093__A0 _0819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2771_ net142 net143 net262 vssd1 vssd1 vccd1 vccd1 _0307_ sky130_fd_sc_hd__mux2_1
Xhold106 LEI0.config_data\[34\] vssd1 vssd1 vccd1 vccd1 net378 sky130_fd_sc_hd__dlygate4sd3_1
X_1653_ CB_0.config_dataA\[17\] CB_0.config_dataA\[16\] CB_0.config_dataA\[19\] CB_0.config_dataA\[18\]
+ vssd1 vssd1 vccd1 vccd1 _0415_ sky130_fd_sc_hd__or4_1
Xhold117 LEI0.config_data\[7\] vssd1 vssd1 vccd1 vccd1 net389 sky130_fd_sc_hd__dlygate4sd3_1
X_1584_ net175 CB_1.config_dataB\[18\] _1329_ net4 vssd1 vssd1 vccd1 vccd1 _0346_
+ sky130_fd_sc_hd__a31o_1
Xhold139 LE_1A.reset_val vssd1 vssd1 vccd1 vccd1 net411 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_194 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_Right_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold128 LE_1B.reset_val vssd1 vssd1 vccd1 vccd1 net400 sky130_fd_sc_hd__dlygate4sd3_1
X_1722_ net128 _1308_ _0459_ vssd1 vssd1 vccd1 vccd1 _0484_ sky130_fd_sc_hd__and3_1
XANTENNA__2296__X _1052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2205_ _0957_ _0960_ vssd1 vssd1 vccd1 vccd1 _0961_ sky130_fd_sc_hd__nand2_1
X_2067_ SB0.route_sel\[76\] SB0.route_sel\[77\] vssd1 vssd1 vccd1 vccd1 _0825_ sky130_fd_sc_hd__nor2_1
X_2136_ net2 net3 net148 vssd1 vssd1 vccd1 vccd1 _0894_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout218_X net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2969_ clknet_leaf_24_clk _0177_ net212 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[41\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__1898__A0 net27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1551__A _1342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2557__A net60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2276__B _0781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2823_ clknet_leaf_14_clk _0031_ net225 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_2754_ CB_1.config_dataA\[2\] CB_1.config_dataA\[1\] net267 vssd1 vssd1 vccd1 vccd1
+ _0290_ sky130_fd_sc_hd__mux2_1
XANTENNA__2081__A3 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1705_ SB0.route_sel\[68\] SB0.route_sel\[69\] net41 vssd1 vssd1 vccd1 vccd1 _0467_
+ sky130_fd_sc_hd__a21bo_1
X_1567_ CB_0.config_dataA\[19\] CB_0.config_dataA\[18\] vssd1 vssd1 vccd1 vccd1 _0329_
+ sky130_fd_sc_hd__nand2_1
X_2685_ SB0.route_sel\[85\] SB0.route_sel\[84\] net240 vssd1 vssd1 vccd1 vccd1 _0221_
+ sky130_fd_sc_hd__mux2_1
X_1636_ _1305_ _0376_ net6 vssd1 vssd1 vccd1 vccd1 _0398_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_1_145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1498_ SB0.route_sel\[52\] SB0.route_sel\[53\] net39 vssd1 vssd1 vccd1 vccd1 _1292_
+ sky130_fd_sc_hd__a21bo_1
X_2119_ CB_1.config_dataA\[9\] CB_1.config_dataA\[11\] vssd1 vssd1 vccd1 vccd1 _0877_
+ sky130_fd_sc_hd__nand2b_1
X_3099_ clknet_leaf_25_clk _0307_ net213 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[19\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_22_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input10_A CBeast_in[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2048__A0 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload26 clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 clkload26/Y sky130_fd_sc_hd__clkinv_8
Xclkload15 clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 clkload15/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_15_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1421_ LEI0.config_data\[14\] vssd1 vssd1 vccd1 vccd1 _1215_ sky130_fd_sc_hd__inv_2
X_2470_ net399 net389 net266 vssd1 vssd1 vccd1 vccd1 _0009_ sky130_fd_sc_hd__mux2_1
X_3022_ clknet_leaf_9_clk _0230_ net219 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[94\]
+ sky130_fd_sc_hd__dfstp_1
X_2806_ clknet_leaf_6_clk net365 net205 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_2737_ CB_0.config_dataB\[5\] net165 net251 vssd1 vssd1 vccd1 vccd1 _0273_ sky130_fd_sc_hd__mux2_1
XANTENNA__2211__A0 net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2668_ SB0.route_sel\[68\] SB0.route_sel\[67\] net240 vssd1 vssd1 vccd1 vccd1 _0204_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout128_A net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload9 clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 clkload9/Y sky130_fd_sc_hd__clkinv_1
Xfanout246 net250 vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__clkbuf_4
Xfanout224 net227 vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__clkbuf_4
Xfanout268 net271 vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout202 net207 vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input2_A CBeast_in[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout235 net236 vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__clkbuf_4
Xfanout257 net262 vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__clkbuf_4
Xfanout213 net218 vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__clkbuf_4
X_1619_ net131 _1257_ _0377_ _0380_ _1261_ vssd1 vssd1 vccd1 vccd1 _0381_ sky130_fd_sc_hd__o32a_1
X_2599_ net175 net176 net255 vssd1 vssd1 vccd1 vccd1 _0135_ sky130_fd_sc_hd__mux2_1
XANTENNA__2278__A0 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1680__B1_N net35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input58_A config_en vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input13_X net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1970_ _0715_ _0727_ _0729_ LEI0.config_data\[29\] vssd1 vssd1 vccd1 vccd1 _0730_
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__2284__A3 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2522_ net332 net322 net247 vssd1 vssd1 vccd1 vccd1 _0060_ sky130_fd_sc_hd__mux2_1
X_2453_ SB0.route_sel\[95\] SB0.route_sel\[94\] SB0.route_sel\[88\] _1205_ vssd1 vssd1
+ vccd1 vccd1 _1146_ sky130_fd_sc_hd__a2bb2o_1
X_2384_ _1191_ SB0.route_sel\[66\] _1192_ SB0.route_sel\[69\] _1099_ vssd1 vssd1 vccd1
+ vccd1 _1100_ sky130_fd_sc_hd__a221o_1
X_1404_ SB0.route_sel\[72\] vssd1 vssd1 vccd1 vccd1 _1198_ sky130_fd_sc_hd__inv_2
Xinput2 CBeast_in[10] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_4
XFILLER_36_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3005_ clknet_leaf_1_clk _0213_ net192 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[77\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_fanout245_A net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input5_X net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_38_Left_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2257__A3 _0838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1953_ _1230_ _0706_ _0712_ vssd1 vssd1 vccd1 vccd1 _0713_ sky130_fd_sc_hd__a21oi_1
X_1884_ net230 net186 vssd1 vssd1 vccd1 vccd1 _0646_ sky130_fd_sc_hd__and2b_1
X_2505_ net404 LEI0.config_data\[42\] net270 vssd1 vssd1 vccd1 vccd1 _0044_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_47_Left_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2193__A2 net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2436_ _1133_ _1134_ _0427_ vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__o21a_1
X_2367_ _1258_ _1329_ _0792_ vssd1 vssd1 vccd1 vccd1 _1090_ sky130_fd_sc_hd__a21o_1
X_2298_ net120 net135 LE_1B.config_data\[15\] vssd1 vssd1 vccd1 vccd1 _1054_ sky130_fd_sc_hd__a21boi_1
XPHY_EDGE_ROW_56_Left_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2239__A3 _0791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2221_ _0356_ _0802_ net185 vssd1 vssd1 vccd1 vccd1 _0977_ sky130_fd_sc_hd__a21oi_1
X_2152_ CB_1.config_dataA\[15\] _0908_ _0909_ _0905_ vssd1 vssd1 vccd1 vccd1 _0910_
+ sky130_fd_sc_hd__o22a_1
XANTENNA__3084__SET_B net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2083_ net2 net3 net150 vssd1 vssd1 vccd1 vccd1 _0841_ sky130_fd_sc_hd__mux2_1
X_1867_ net27 net28 net16 net17 net169 net168 vssd1 vssd1 vccd1 vccd1 _0629_ sky130_fd_sc_hd__mux4_1
X_1936_ CB_0.config_dataB\[1\] net167 _1273_ vssd1 vssd1 vccd1 vccd1 _0696_ sky130_fd_sc_hd__and3_1
X_2985_ clknet_leaf_23_clk _0193_ net211 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[57\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_21_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1798_ net136 net127 net130 net134 LEI0.config_data\[12\] LEI0.config_data\[13\]
+ vssd1 vssd1 vccd1 vccd1 _0560_ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout208_A net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput60 le_en vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_59_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2419_ SB0.route_sel\[17\] SB0.route_sel\[16\] vssd1 vssd1 vccd1 vccd1 _1123_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_42_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1601__A1 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2157__A2 _0828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input40_A SBsouth_in[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2093__A1 _0822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2770_ net143 net144 net257 vssd1 vssd1 vccd1 vccd1 _0306_ sky130_fd_sc_hd__mux2_1
X_1721_ SB0.route_sel\[74\] SB0.route_sel\[75\] vssd1 vssd1 vccd1 vccd1 _0483_ sky130_fd_sc_hd__and2_1
X_1583_ net138 _0343_ _0341_ vssd1 vssd1 vccd1 vccd1 _0345_ sky130_fd_sc_hd__mux2_1
X_1652_ net157 net159 net153 net155 vssd1 vssd1 vccd1 vccd1 _0414_ sky130_fd_sc_hd__or4_1
Xhold107 LEI0.config_data\[4\] vssd1 vssd1 vccd1 vccd1 net379 sky130_fd_sc_hd__dlygate4sd3_1
Xhold118 LEI0.config_data\[19\] vssd1 vssd1 vccd1 vccd1 net390 sky130_fd_sc_hd__dlygate4sd3_1
Xhold129 LE_0B.config_data\[1\] vssd1 vssd1 vccd1 vccd1 net401 sky130_fd_sc_hd__dlygate4sd3_1
X_2204_ _0944_ _0946_ _0959_ LEI0.config_data\[11\] vssd1 vssd1 vccd1 vccd1 _0960_
+ sky130_fd_sc_hd__o22a_1
X_2135_ net13 net14 net148 vssd1 vssd1 vccd1 vccd1 _0893_ sky130_fd_sc_hd__mux2_1
X_2066_ CB_1.config_dataA\[7\] _0823_ vssd1 vssd1 vccd1 vccd1 _0824_ sky130_fd_sc_hd__nor2_1
XANTENNA__1656__X _0418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1919_ net23 net24 net25 net26 net167 net166 vssd1 vssd1 vccd1 vccd1 _0679_ sky130_fd_sc_hd__mux4_1
X_2899_ clknet_leaf_21_clk net290 net215 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_2968_ clknet_leaf_26_clk _0176_ net211 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[40\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__1898__A1 net28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1551__B _1344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1822__B2 _0512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1889__A1 _0430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2397__X net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2753_ CB_1.config_dataA\[1\] net152 net267 vssd1 vssd1 vccd1 vccd1 _0289_ sky130_fd_sc_hd__mux2_1
X_2822_ clknet_leaf_2_clk _0030_ net208 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[29\]
+ sky130_fd_sc_hd__dfrtp_2
X_2684_ SB0.route_sel\[84\] SB0.route_sel\[83\] net240 vssd1 vssd1 vccd1 vccd1 _0220_
+ sky130_fd_sc_hd__mux2_1
X_1704_ SB0.route_sel\[71\] SB0.route_sel\[70\] _0465_ vssd1 vssd1 vccd1 vccd1 _0466_
+ sky130_fd_sc_hd__a21bo_1
X_1566_ net154 net156 _1300_ net19 vssd1 vssd1 vccd1 vccd1 _0328_ sky130_fd_sc_hd__a31o_1
X_1635_ net136 _0395_ _0393_ vssd1 vssd1 vccd1 vccd1 _0397_ sky130_fd_sc_hd__mux2_1
X_1497_ SB0.route_sel\[55\] SB0.route_sel\[54\] _1290_ vssd1 vssd1 vccd1 vccd1 _1291_
+ sky130_fd_sc_hd__a21bo_1
X_2049_ CB_1.config_dataA\[7\] _0805_ _0806_ _0800_ vssd1 vssd1 vccd1 vccd1 _0807_
+ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_1_146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3098_ clknet_leaf_24_clk _0306_ net213 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[18\]
+ sky130_fd_sc_hd__dfstp_1
X_2118_ CB_1.config_dataA\[11\] _0875_ vssd1 vssd1 vccd1 vccd1 _0876_ sky130_fd_sc_hd__nand2b_1
XANTENNA_clkbuf_leaf_18_clk_A clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2048__A1 net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload16 clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 clkload16/Y sky130_fd_sc_hd__inv_12
Xclkload27 clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 clkload27/Y sky130_fd_sc_hd__inv_4
X_1420_ CB_0.config_dataA\[3\] vssd1 vssd1 vccd1 vccd1 _1214_ sky130_fd_sc_hd__inv_2
X_3021_ clknet_leaf_25_clk _0229_ net198 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[93\]
+ sky130_fd_sc_hd__dfstp_1
X_2805_ clknet_leaf_5_clk _0013_ net205 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2804__Q LEI0.config_data\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1798__A0 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2736_ net165 CB_0.config_dataB\[3\] net251 vssd1 vssd1 vccd1 vccd1 _0272_ sky130_fd_sc_hd__mux2_1
XANTENNA__2211__A1 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2667_ SB0.route_sel\[67\] SB0.route_sel\[66\] net240 vssd1 vssd1 vccd1 vccd1 _0203_
+ sky130_fd_sc_hd__mux2_1
X_1618_ net142 net143 vssd1 vssd1 vccd1 vccd1 _0380_ sky130_fd_sc_hd__or2_1
Xfanout269 net271 vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__clkbuf_4
Xfanout203 net207 vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__clkbuf_4
Xfanout247 net250 vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__clkbuf_2
Xfanout225 net227 vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__clkbuf_4
XANTENNA__2278__A1 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout236 net254 vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__buf_2
Xfanout214 net217 vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__clkbuf_4
Xfanout258 net261 vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__clkbuf_4
X_1549_ SB0.route_sel\[35\] SB0.route_sel\[34\] vssd1 vssd1 vccd1 vccd1 _1343_ sky130_fd_sc_hd__nor2_1
X_2598_ net176 CB_1.config_dataB\[17\] net261 vssd1 vssd1 vccd1 vccd1 _0134_ sky130_fd_sc_hd__mux2_1
XANTENNA__1789__A0 net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1961__A0 net27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2441__A1 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2521_ net322 net298 net247 vssd1 vssd1 vccd1 vccd1 _0059_ sky130_fd_sc_hd__mux2_1
X_2452_ SB0.route_sel\[90\] _1203_ vssd1 vssd1 vccd1 vccd1 _1145_ sky130_fd_sc_hd__nor2_1
X_1403_ SB0.route_sel\[78\] vssd1 vssd1 vccd1 vccd1 _1197_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_18_Right_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2383_ SB0.route_sel\[65\] SB0.route_sel\[64\] vssd1 vssd1 vccd1 vccd1 _1099_ sky130_fd_sc_hd__nor2_1
Xinput3 CBeast_in[11] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_27_Right_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3004_ clknet_leaf_1_clk _0212_ net191 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[76\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_fanout140_A net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2719_ CB_0.config_dataA\[7\] CB_0.config_dataA\[6\] net249 vssd1 vssd1 vccd1 vccd1
+ _0255_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_36_Right_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_45_Right_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_54_Right_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_63_Right_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2111__A0 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1883_ _0644_ _0637_ _0633_ vssd1 vssd1 vccd1 vccd1 _0645_ sky130_fd_sc_hd__mux2_1
X_1952_ CB_0.config_dataB\[11\] _0710_ _0711_ _0707_ vssd1 vssd1 vccd1 vccd1 _0712_
+ sky130_fd_sc_hd__o22a_1
X_2504_ LEI0.config_data\[42\] net410 net270 vssd1 vssd1 vccd1 vccd1 _0043_ sky130_fd_sc_hd__mux2_1
XANTENNA__1925__A0 net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2193__A3 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2435_ _1160_ SB0.route_sel\[1\] _1157_ _1158_ vssd1 vssd1 vccd1 vccd1 _1134_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_fanout188_A net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2366_ _1310_ _1089_ _1312_ vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__a21o_1
X_2297_ _0990_ _1017_ _1020_ _1052_ vssd1 vssd1 vccd1 vccd1 _1053_ sky130_fd_sc_hd__o31a_1
XFILLER_20_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2902__Q LE_1A.config_data\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2220_ _1358_ _0334_ _0796_ net185 vssd1 vssd1 vccd1 vccd1 _0976_ sky130_fd_sc_hd__o31a_1
X_2082_ net13 net14 net150 vssd1 vssd1 vccd1 vccd1 _0840_ sky130_fd_sc_hd__mux2_1
X_2151_ net4 net5 net146 vssd1 vssd1 vccd1 vccd1 _0909_ sky130_fd_sc_hd__mux2_1
XFILLER_53_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2984_ clknet_leaf_22_clk _0192_ net214 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[56\]
+ sky130_fd_sc_hd__dfstp_1
X_1866_ net15 net20 net21 net22 net169 net168 vssd1 vssd1 vccd1 vccd1 _0628_ sky130_fd_sc_hd__mux4_1
X_1797_ CB_0.config_dataA\[6\] _0558_ vssd1 vssd1 vccd1 vccd1 _0559_ sky130_fd_sc_hd__and2b_1
X_1935_ net166 _1225_ _1297_ vssd1 vssd1 vccd1 vccd1 _0695_ sky130_fd_sc_hd__and3_1
Xinput61 le_nrst vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__buf_2
Xinput50 SBwest_in[3] vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_59_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2323__A0 _0359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2418_ _1121_ _1122_ _0388_ vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__o21a_1
X_2349_ _1306_ _1348_ _0797_ vssd1 vssd1 vccd1 vccd1 _1081_ sky130_fd_sc_hd__o21ai_1
XFILLER_52_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Right_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input33_A SBsouth_in[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2093__A2 _0816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold108 LEI0.config_data\[10\] vssd1 vssd1 vccd1 vccd1 net380 sky130_fd_sc_hd__dlygate4sd3_1
X_1651_ SB0.route_sel\[0\] SB0.route_sel\[1\] vssd1 vssd1 vccd1 vccd1 _0413_ sky130_fd_sc_hd__nand2_1
X_1720_ net131 _1306_ _0457_ _0460_ _1309_ vssd1 vssd1 vccd1 vccd1 _0482_ sky130_fd_sc_hd__o32a_1
XANTENNA__1762__X _0524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1582_ SB0.route_sel\[96\] SB0.route_sel\[97\] vssd1 vssd1 vccd1 vccd1 _0344_ sky130_fd_sc_hd__nand2_1
Xhold119 _0020_ vssd1 vssd1 vccd1 vccd1 net391 sky130_fd_sc_hd__dlygate4sd3_1
X_2203_ _0958_ vssd1 vssd1 vccd1 vccd1 _0959_ sky130_fd_sc_hd__inv_2
X_2065_ _0816_ _0819_ _0813_ _0822_ _1237_ CB_1.config_dataA\[5\] vssd1 vssd1 vccd1
+ vccd1 _0823_ sky130_fd_sc_hd__mux4_1
XFILLER_26_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2134_ CB_1.config_dataA\[11\] _0891_ vssd1 vssd1 vccd1 vccd1 _0892_ sky130_fd_sc_hd__or2_1
X_2967_ clknet_leaf_26_clk _0175_ net198 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[39\]
+ sky130_fd_sc_hd__dfstp_1
X_1849_ _1220_ CB_0.config_dataA\[15\] vssd1 vssd1 vccd1 vccd1 _0611_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout220_A net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1918_ net166 _1226_ _0677_ vssd1 vssd1 vccd1 vccd1 _0678_ sky130_fd_sc_hd__or3_1
X_2898_ clknet_leaf_21_clk net334 net215 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_4_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_20_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__1889__A2 _0391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2821_ clknet_leaf_3_clk net382 net208 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_11_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2752_ net152 net154 net268 vssd1 vssd1 vccd1 vccd1 _0288_ sky130_fd_sc_hd__mux2_1
X_2683_ SB0.route_sel\[83\] SB0.route_sel\[82\] net239 vssd1 vssd1 vccd1 vccd1 _0219_
+ sky130_fd_sc_hd__mux2_1
X_1634_ SB0.route_sel\[9\] SB0.route_sel\[8\] vssd1 vssd1 vccd1 vccd1 _0396_ sky130_fd_sc_hd__nand2_1
X_1703_ SB0.route_sel\[68\] SB0.route_sel\[69\] net55 vssd1 vssd1 vccd1 vccd1 _0465_
+ sky130_fd_sc_hd__and3_1
X_1565_ _1347_ _1353_ _1357_ vssd1 vssd1 vccd1 vccd1 _1359_ sky130_fd_sc_hd__a21o_1
X_1496_ SB0.route_sel\[52\] SB0.route_sel\[53\] net53 vssd1 vssd1 vccd1 vccd1 _1290_
+ sky130_fd_sc_hd__and3_1
X_2048_ net4 net5 net150 vssd1 vssd1 vccd1 vccd1 _0806_ sky130_fd_sc_hd__mux2_1
X_3097_ clknet_leaf_24_clk _0305_ net211 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[17\]
+ sky130_fd_sc_hd__dfstp_1
X_2117_ _0792_ _0788_ _0784_ _0781_ CB_1.config_dataA\[9\] net149 vssd1 vssd1 vccd1
+ vccd1 _0875_ sky130_fd_sc_hd__mux4_1
XANTENNA__1804__A2 _0359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload28 clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 clkload28/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__1577__X _0339_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload17 clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 clkload17/Y sky130_fd_sc_hd__clkinv_8
XFILLER_48_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2201__X _0957_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_0_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_clk
+ sky130_fd_sc_hd__clkbuf_8
X_3020_ clknet_leaf_25_clk _0228_ net213 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[92\]
+ sky130_fd_sc_hd__dfstp_1
X_2804_ clknet_leaf_10_clk _0012_ net220 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[11\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__1798__A1 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout204 net207 vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__clkbuf_2
X_2735_ CB_0.config_dataB\[3\] CB_0.config_dataB\[2\] net251 vssd1 vssd1 vccd1 vccd1
+ _0271_ sky130_fd_sc_hd__mux2_1
XANTENNA__1970__B2 LEI0.config_data\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2211__A2 net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1617_ net142 net143 vssd1 vssd1 vccd1 vccd1 _0379_ sky130_fd_sc_hd__nor2_1
X_2666_ SB0.route_sel\[66\] SB0.route_sel\[65\] net240 vssd1 vssd1 vccd1 vccd1 _0202_
+ sky130_fd_sc_hd__mux2_1
X_2597_ CB_1.config_dataB\[17\] net178 net261 vssd1 vssd1 vccd1 vccd1 _0133_ sky130_fd_sc_hd__mux2_1
Xfanout248 net250 vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__clkbuf_4
Xfanout226 net227 vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__buf_2
XANTENNA__2278__A2 net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout215 net217 vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__clkbuf_4
X_1479_ _1271_ _1272_ _1270_ vssd1 vssd1 vccd1 vccd1 _1273_ sky130_fd_sc_hd__a21boi_4
Xfanout237 net241 vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__clkbuf_4
Xfanout259 net261 vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__clkbuf_4
X_1548_ _1322_ _1328_ _1338_ _1341_ vssd1 vssd1 vccd1 vccd1 _1342_ sky130_fd_sc_hd__a22o_2
XANTENNA__1789__A1 net20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1961__A1 net28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1844__Y _0606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2520_ net298 LE_0A.config_data\[6\] net247 vssd1 vssd1 vccd1 vccd1 _0058_ sky130_fd_sc_hd__mux2_1
X_2451_ _0508_ _1144_ vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__and2_1
X_1402_ SB0.route_sel\[79\] vssd1 vssd1 vccd1 vccd1 _1196_ sky130_fd_sc_hd__inv_2
Xinput4 CBeast_in[12] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__buf_2
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_17_clk_A clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2382_ _1097_ _1098_ _0489_ vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__o21a_1
X_3003_ clknet_leaf_1_clk _0211_ net191 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[75\]
+ sky130_fd_sc_hd__dfstp_1
Xclkbuf_2_1__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_2_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_34_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2718_ CB_0.config_dataA\[6\] net171 net249 vssd1 vssd1 vccd1 vccd1 _0254_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout133_A net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2649_ SB0.route_sel\[49\] SB0.route_sel\[48\] net258 vssd1 vssd1 vccd1 vccd1 _0185_
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2111__A1 net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1882_ _0643_ _0640_ _0602_ vssd1 vssd1 vccd1 vccd1 _0644_ sky130_fd_sc_hd__mux2_1
X_1951_ net18 net19 net164 vssd1 vssd1 vccd1 vccd1 _0711_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_31_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2503_ LEI0.config_data\[41\] net362 net268 vssd1 vssd1 vccd1 vccd1 _0042_ sky130_fd_sc_hd__mux2_1
XANTENNA__1925__A1 net20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2434_ _1155_ SB0.route_sel\[2\] vssd1 vssd1 vccd1 vccd1 _1133_ sky130_fd_sc_hd__nor2_1
X_2365_ _1258_ _1305_ _0784_ vssd1 vssd1 vccd1 vccd1 _1089_ sky130_fd_sc_hd__a21o_1
X_2296_ _1037_ _1038_ _1049_ _1051_ CB_0.config_data_inA vssd1 vssd1 vccd1 vccd1 _1052_
+ sky130_fd_sc_hd__o32a_2
XANTENNA_fanout136_X net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout250_A net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2081_ net1 net6 net7 net8 net150 CB_1.config_dataA\[5\] vssd1 vssd1 vccd1 vccd1
+ _0839_ sky130_fd_sc_hd__mux4_1
X_2150_ net9 net10 net11 net12 net146 CB_1.config_dataA\[13\] vssd1 vssd1 vccd1 vccd1
+ _0908_ sky130_fd_sc_hd__mux4_1
X_1934_ net167 _1345_ _0693_ _1224_ vssd1 vssd1 vccd1 vccd1 _0694_ sky130_fd_sc_hd__o211a_1
X_2983_ clknet_leaf_22_clk _0191_ net214 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[55\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__1479__Y _1273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1796_ _0548_ _0552_ _0553_ _0557_ vssd1 vssd1 vccd1 vccd1 _0558_ sky130_fd_sc_hd__o2bb2a_1
Xinput62 nrst vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__clkbuf_1
X_1865_ _1220_ _0624_ _0626_ vssd1 vssd1 vccd1 vccd1 _0627_ sky130_fd_sc_hd__a21oi_1
Xinput40 SBsouth_in[7] vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__clkbuf_1
Xinput51 SBwest_in[4] vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__buf_1
X_2348_ net137 _1080_ _0415_ vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__mux2_1
X_2417_ SB0.route_sel\[25\] _1175_ _1173_ _1174_ vssd1 vssd1 vccd1 vccd1 _1122_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_42_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2279_ net4 net5 net181 vssd1 vssd1 vccd1 vccd1 _1035_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_50_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input26_A CBnorth_in[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2093__A3 _0813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2173__S0 _0848_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1581_ net18 net125 _0342_ vssd1 vssd1 vccd1 vccd1 _0343_ sky130_fd_sc_hd__mux2_1
X_1650_ net121 vssd1 vssd1 vccd1 vccd1 _0412_ sky130_fd_sc_hd__inv_2
Xhold109 LEI0.config_data\[28\] vssd1 vssd1 vccd1 vccd1 net381 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2250__A0 _0816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2204__X _0960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output94_A net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2202_ net140 net124 net129 net133 LEI0.config_data\[9\] LEI0.config_data\[10\] vssd1
+ vssd1 vccd1 vccd1 _0958_ sky130_fd_sc_hd__mux4_1
XFILLER_26_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2064_ _0444_ _0821_ vssd1 vssd1 vccd1 vccd1 _0822_ sky130_fd_sc_hd__nand2_4
X_2133_ net1 net6 net7 net8 net149 CB_1.config_dataA\[9\] vssd1 vssd1 vccd1 vccd1
+ _0891_ sky130_fd_sc_hd__mux4_1
X_1917_ net18 net19 net167 vssd1 vssd1 vccd1 vccd1 _0677_ sky130_fd_sc_hd__mux2_1
X_2897_ clknet_leaf_21_clk net393 net215 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_2966_ clknet_leaf_26_clk _0174_ net198 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[38\]
+ sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_14_Left_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1848_ net23 net24 net25 net26 CB_0.config_dataA\[12\] CB_0.config_dataA\[13\] vssd1
+ vssd1 vccd1 vccd1 _0610_ sky130_fd_sc_hd__mux4_1
X_1779_ _0449_ _0540_ CB_0.config_dataA\[3\] vssd1 vssd1 vccd1 vccd1 _0541_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout213_A net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1889__A3 _0447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2299__B1 _0984_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2751_ net154 net156 net271 vssd1 vssd1 vccd1 vccd1 _0287_ sky130_fd_sc_hd__mux2_1
X_2820_ clknet_leaf_2_clk _0028_ net208 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_1633_ net122 net20 _0394_ vssd1 vssd1 vccd1 vccd1 _0395_ sky130_fd_sc_hd__mux2_1
X_1564_ _1347_ _1353_ _1357_ vssd1 vssd1 vccd1 vccd1 _1358_ sky130_fd_sc_hd__a21oi_2
X_2682_ SB0.route_sel\[82\] SB0.route_sel\[81\] net251 vssd1 vssd1 vccd1 vccd1 _0218_
+ sky130_fd_sc_hd__mux2_1
X_1702_ _0458_ _0461_ _0462_ _0463_ vssd1 vssd1 vccd1 vccd1 _0464_ sky130_fd_sc_hd__a211oi_1
X_1495_ _1282_ _1286_ _1287_ _1288_ vssd1 vssd1 vccd1 vccd1 _1289_ sky130_fd_sc_hd__a211oi_1
X_2116_ _0864_ _0872_ _0873_ _0850_ LEI0.config_data\[8\] vssd1 vssd1 vccd1 vccd1
+ _0874_ sky130_fd_sc_hd__o32a_2
X_2047_ net9 net10 net11 net12 net150 CB_1.config_dataA\[5\] vssd1 vssd1 vccd1 vccd1
+ _0805_ sky130_fd_sc_hd__mux4_1
XANTENNA__2462__A0 LEI0.config_data\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3096_ clknet_leaf_20_clk _0304_ net218 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[16\]
+ sky130_fd_sc_hd__dfstp_1
X_2949_ clknet_leaf_30_clk _0157_ net189 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[21\]
+ sky130_fd_sc_hd__dfstp_1
Xclkload29 clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 clkload29/Y sky130_fd_sc_hd__inv_6
Xclkload18 clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 clkload18/Y sky130_fd_sc_hd__clkinv_8
XANTENNA__1472__C net54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2803_ clknet_leaf_10_clk _0011_ net220 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_2734_ CB_0.config_dataB\[2\] net166 net245 vssd1 vssd1 vccd1 vccd1 _0270_ sky130_fd_sc_hd__mux2_1
XANTENNA__1798__A2 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2211__A3 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout227 net228 vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout205 net207 vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__clkbuf_4
X_2596_ CB_1.config_dataB\[16\] CB_1.config_dataB\[15\] net261 vssd1 vssd1 vccd1 vccd1
+ _0132_ sky130_fd_sc_hd__mux2_1
Xfanout238 net241 vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__clkbuf_4
X_1547_ _1336_ _1339_ _1340_ SB0.route_sel\[32\] SB0.route_sel\[33\] vssd1 vssd1 vccd1
+ vccd1 _1341_ sky130_fd_sc_hd__o311a_1
Xfanout216 net217 vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__clkbuf_4
X_2665_ SB0.route_sel\[65\] SB0.route_sel\[64\] net240 vssd1 vssd1 vccd1 vccd1 _0201_
+ sky130_fd_sc_hd__mux2_1
X_1616_ net177 net178 _0376_ net8 vssd1 vssd1 vccd1 vccd1 _0378_ sky130_fd_sc_hd__a31o_1
Xfanout249 net250 vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__buf_2
XANTENNA__2278__A3 net12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1478_ SB0.route_sel\[58\] SB0.route_sel\[59\] _1189_ SB0.route_sel\[61\] vssd1 vssd1
+ vccd1 vccd1 _1272_ sky130_fd_sc_hd__o22a_1
X_3079_ clknet_leaf_12_clk _0287_ net227 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[19\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_37_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2202__A3 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_17_Left_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2450_ SB0.route_sel\[90\] _1203_ _1204_ SB0.route_sel\[93\] _1143_ vssd1 vssd1 vccd1
+ vccd1 _1144_ sky130_fd_sc_hd__a221o_1
X_2381_ SB0.route_sel\[73\] _1198_ _1196_ _1197_ vssd1 vssd1 vccd1 vccd1 _1098_ sky130_fd_sc_hd__a2bb2o_1
X_1401_ SB0.route_sel\[77\] vssd1 vssd1 vccd1 vccd1 _1195_ sky130_fd_sc_hd__inv_2
XFILLER_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput5 CBeast_in[13] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__buf_2
X_3002_ clknet_leaf_1_clk _0210_ net196 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[74\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_34_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2717_ net171 net173 net249 vssd1 vssd1 vccd1 vccd1 _0253_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout126_A net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2648_ SB0.route_sel\[48\] SB0.route_sel\[47\] net258 vssd1 vssd1 vccd1 vccd1 _0184_
+ sky130_fd_sc_hd__mux2_1
X_2579_ LE_1B.dff0_out _1247_ _1153_ vssd1 vssd1 vccd1 vccd1 _0115_ sky130_fd_sc_hd__a21bo_1
XFILLER_27_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1934__A2 _1345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_2_Left_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input56_A SBwest_in[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input11_X net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1950_ net23 net24 net25 net26 net163 CB_0.config_dataB\[9\] vssd1 vssd1 vccd1 vccd1
+ _0710_ sky130_fd_sc_hd__mux4_1
XFILLER_18_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2502_ net362 net368 net268 vssd1 vssd1 vccd1 vccd1 _0041_ sky130_fd_sc_hd__mux2_1
X_1881_ _0642_ _0641_ _0572_ vssd1 vssd1 vccd1 vccd1 _0643_ sky130_fd_sc_hd__mux2_1
XANTENNA__1925__A2 net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2433_ _1131_ _1132_ _0427_ vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__o21a_1
X_2364_ _1286_ _1088_ _1288_ vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__a21o_1
XFILLER_56_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2295_ _1050_ vssd1 vssd1 vccd1 vccd1 _1051_ sky130_fd_sc_hd__inv_2
XANTENNA_10 CBnorth_in[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1861__B2 _0512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input3_X net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_2_0__f_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_16_clk_A clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2080_ _0836_ _0837_ _0534_ vssd1 vssd1 vccd1 vccd1 _0838_ sky130_fd_sc_hd__a21boi_4
X_1933_ _1318_ _1320_ CB_0.config_dataB\[0\] vssd1 vssd1 vccd1 vccd1 _0693_ sky130_fd_sc_hd__o21ai_1
X_2982_ clknet_leaf_20_clk _0190_ net216 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[54\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_21_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1795_ _1216_ _0554_ _0556_ vssd1 vssd1 vccd1 vccd1 _0557_ sky130_fd_sc_hd__o21a_1
X_1864_ net168 net169 _0391_ CB_0.config_dataA\[15\] vssd1 vssd1 vccd1 vccd1 _0626_
+ sky130_fd_sc_hd__a31o_1
Xinput30 SBsouth_in[10] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__buf_1
Xinput41 SBsouth_in[8] vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__buf_1
Xinput52 SBwest_in[5] vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__buf_1
X_2347_ _0414_ _0430_ _0416_ vssd1 vssd1 vccd1 vccd1 _1080_ sky130_fd_sc_hd__a21oi_1
X_2278_ net9 net10 net11 net12 net181 net179 vssd1 vssd1 vccd1 vccd1 _1034_ sky130_fd_sc_hd__mux4_1
XANTENNA__2400__X net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2416_ SB0.route_sel\[26\] _1171_ vssd1 vssd1 vccd1 vccd1 _1121_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout193_A net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2924__SET_B net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input19_A CBnorth_in[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2173__S1 _0874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1580_ net158 net160 net154 net156 vssd1 vssd1 vccd1 vccd1 _0342_ sky130_fd_sc_hd__and4bb_1
XANTENNA__2250__A1 _0819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2201_ _0948_ _0954_ _0956_ CB_1.config_dataB\[2\] vssd1 vssd1 vccd1 vccd1 _0957_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__1513__B1 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2132_ net148 _0828_ _0877_ _0889_ vssd1 vssd1 vccd1 vccd1 _0890_ sky130_fd_sc_hd__a211o_1
X_2063_ _1168_ SB0.route_sel\[22\] SB0.route_sel\[17\] _1170_ _0820_ vssd1 vssd1 vccd1
+ vccd1 _0821_ sky130_fd_sc_hd__a221o_1
X_1847_ net168 net169 vssd1 vssd1 vccd1 vccd1 _0609_ sky130_fd_sc_hd__nand2_1
X_1916_ _0675_ vssd1 vssd1 vccd1 vccd1 _0676_ sky130_fd_sc_hd__inv_2
X_2896_ clknet_leaf_21_clk _0104_ net215 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_2965_ clknet_leaf_26_clk _0173_ net195 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[37\]
+ sky130_fd_sc_hd__dfstp_1
X_1778_ _0474_ _0493_ _0539_ _0513_ CB_0.config_dataA\[0\] CB_0.config_dataA\[1\]
+ vssd1 vssd1 vccd1 vccd1 _0540_ sky130_fd_sc_hd__mux4_1
XANTENNA__1752__A0 net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1807__A1 _1297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1807__B2 _1273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1991__A0 net27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2091__S0 LEI0.config_data\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_31_Left_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2750_ net156 net158 net271 vssd1 vssd1 vccd1 vccd1 _0286_ sky130_fd_sc_hd__mux2_1
X_2681_ SB0.route_sel\[81\] SB0.route_sel\[80\] net251 vssd1 vssd1 vccd1 vccd1 _0217_
+ sky130_fd_sc_hd__mux2_1
X_1701_ net128 _1332_ _0459_ vssd1 vssd1 vccd1 vccd1 _0463_ sky130_fd_sc_hd__and3_1
XANTENNA__1734__A0 net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1632_ net157 net153 net155 net159 vssd1 vssd1 vccd1 vccd1 _0394_ sky130_fd_sc_hd__or4b_1
X_1563_ SB0.route_sel\[104\] SB0.route_sel\[105\] _1356_ vssd1 vssd1 vccd1 vccd1 _1357_
+ sky130_fd_sc_hd__nand3_1
X_1494_ _1249_ _1285_ vssd1 vssd1 vccd1 vccd1 _1288_ sky130_fd_sc_hd__nor2_1
X_2115_ CB_1.config_dataA\[2\] _0867_ _0871_ vssd1 vssd1 vccd1 vccd1 _0873_ sky130_fd_sc_hd__and3_1
X_3095_ clknet_leaf_20_clk _0303_ net216 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[15\]
+ sky130_fd_sc_hd__dfstp_2
X_2046_ _0356_ _0802_ net150 vssd1 vssd1 vccd1 vccd1 _0804_ sky130_fd_sc_hd__a21o_1
XANTENNA__1677__A net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2879_ clknet_leaf_4_clk net274 net199 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_2948_ clknet_leaf_30_clk _0156_ net189 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[20\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_13_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2150__A0 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload19 clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 clkload19/Y sky130_fd_sc_hd__clkinv_8
XANTENNA_input41_X net41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1798__A3 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2802_ clknet_leaf_14_clk _0010_ net225 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_2733_ net166 net167 net245 vssd1 vssd1 vccd1 vccd1 _0269_ sky130_fd_sc_hd__mux2_1
X_2664_ SB0.route_sel\[64\] SB0.route_sel\[63\] net237 vssd1 vssd1 vccd1 vccd1 _0200_
+ sky130_fd_sc_hd__mux2_1
Xfanout228 net229 vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__buf_2
Xfanout206 net207 vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__buf_2
X_2595_ CB_1.config_dataB\[15\] CB_1.config_dataB\[14\] net267 vssd1 vssd1 vccd1 vccd1
+ _0131_ sky130_fd_sc_hd__mux2_1
Xfanout239 net240 vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__clkbuf_4
Xfanout217 net218 vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__clkbuf_4
X_1477_ SB0.route_sel\[62\] SB0.route_sel\[63\] vssd1 vssd1 vccd1 vccd1 _1271_ sky130_fd_sc_hd__nand2b_1
X_1546_ SB0.route_sel\[36\] SB0.route_sel\[37\] net37 vssd1 vssd1 vccd1 vccd1 _1340_
+ sky130_fd_sc_hd__a21boi_1
X_1615_ net175 net176 vssd1 vssd1 vccd1 vccd1 _0377_ sky130_fd_sc_hd__or2_2
X_3078_ clknet_leaf_12_clk _0286_ net227 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[18\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_54_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2029_ _1187_ SB0.route_sel\[48\] vssd1 vssd1 vccd1 vccd1 _0787_ sky130_fd_sc_hd__nor2_1
XANTENNA__1946__A0 _1345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2371__B1 _0822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2123__A0 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3096__SET_B net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1400_ SB0.route_sel\[64\] vssd1 vssd1 vccd1 vccd1 _1194_ sky130_fd_sc_hd__inv_2
X_2380_ SB0.route_sel\[74\] SB0.route_sel\[75\] vssd1 vssd1 vccd1 vccd1 _1097_ sky130_fd_sc_hd__and2b_1
Xinput6 CBeast_in[1] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__buf_2
X_3001_ clknet_leaf_1_clk _0209_ net196 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[73\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_34_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2716_ net173 CB_0.config_dataA\[3\] net248 vssd1 vssd1 vccd1 vccd1 _0252_ sky130_fd_sc_hd__mux2_1
X_2647_ SB0.route_sel\[47\] SB0.route_sel\[46\] net256 vssd1 vssd1 vccd1 vccd1 _0183_
+ sky130_fd_sc_hd__mux2_1
X_1529_ net157 net159 net153 net155 vssd1 vssd1 vccd1 vccd1 _1323_ sky130_fd_sc_hd__or4b_1
X_2578_ LE_1A.reset_mode net411 net230 vssd1 vssd1 vccd1 vccd1 _0114_ sky130_fd_sc_hd__mux2_1
XFILLER_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1919__A0 net23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_14_Right_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2026__A _1318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_23_Right_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input49_A SBwest_in[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1880_ LE_0A.config_data\[9\] LE_0A.config_data\[8\] _0543_ vssd1 vssd1 vccd1 vccd1
+ _0642_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_32_Right_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2501_ net368 LEI0.config_data\[38\] net268 vssd1 vssd1 vccd1 vccd1 _0040_ sky130_fd_sc_hd__mux2_1
XANTENNA__1925__A3 net22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2294_ net139 net126 net129 net133 LEI0.config_data\[45\] LEI0.config_data\[46\]
+ vssd1 vssd1 vccd1 vccd1 _1050_ sky130_fd_sc_hd__mux4_1
XANTENNA__2335__A0 _1297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_41_Right_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2432_ SB0.route_sel\[0\] SB0.route_sel\[1\] _1155_ SB0.route_sel\[2\] vssd1 vssd1
+ vccd1 vccd1 _1132_ sky130_fd_sc_hd__a2bb2o_1
X_2363_ _1258_ _1280_ _0788_ vssd1 vssd1 vccd1 vccd1 _1088_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_50_Right_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_11 net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout236_A net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2574__A0 LE_1A.config_data\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1852__A2 _0339_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2927__Q CB_1.config_dataB\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2096__A2 _0828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput20 CBnorth_in[1] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__buf_2
X_1863_ _0447_ _0607_ vssd1 vssd1 vccd1 vccd1 _0625_ sky130_fd_sc_hd__nand2_1
XANTENNA__1936__C _1273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1932_ net167 _0359_ _0691_ CB_0.config_dataB\[3\] _1224_ vssd1 vssd1 vccd1 vccd1
+ _0692_ sky130_fd_sc_hd__o2111a_1
Xinput31 SBsouth_in[11] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__buf_1
X_2981_ clknet_leaf_22_clk _0189_ net214 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[53\]
+ sky130_fd_sc_hd__dfstp_1
X_1794_ net171 _1216_ _0555_ vssd1 vssd1 vccd1 vccd1 _0556_ sky130_fd_sc_hd__or3_1
Xinput42 SBsouth_in[9] vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__buf_1
X_2415_ _1119_ _1120_ _0388_ vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__o21a_1
Xinput53 SBwest_in[6] vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__buf_1
XANTENNA__2308__B1 _1052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2346_ net137 _1079_ _0393_ vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__mux2_1
XFILLER_37_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2277_ net180 _0789_ _1032_ net179 vssd1 vssd1 vccd1 vccd1 _1033_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout186_A net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1834__A2 _1342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout141_X net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2250__A2 _0813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_23_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_clk
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_44_Left_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_53_Left_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2200_ CB_1.config_dataB\[3\] _0955_ vssd1 vssd1 vccd1 vccd1 _0956_ sky130_fd_sc_hd__nand2_1
X_2131_ net148 _0831_ vssd1 vssd1 vccd1 vccd1 _0889_ sky130_fd_sc_hd__nor2_1
X_2062_ SB0.route_sel\[20\] SB0.route_sel\[21\] vssd1 vssd1 vccd1 vccd1 _0820_ sky130_fd_sc_hd__nor2_1
X_2964_ clknet_leaf_26_clk _0172_ net196 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[36\]
+ sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_62_Left_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1846_ net168 _1221_ vssd1 vssd1 vccd1 vccd1 _0608_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_14_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1915_ _1227_ _0648_ _0664_ _0674_ vssd1 vssd1 vccd1 vccd1 _0675_ sky130_fd_sc_hd__a22o_1
X_1777_ _0535_ _0536_ _0537_ _0534_ vssd1 vssd1 vccd1 vccd1 _0539_ sky130_fd_sc_hd__o31ai_2
X_2895_ clknet_leaf_21_clk _0103_ net215 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_15_clk_A clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1752__A1 net20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_4_Right_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2329_ _0476_ _0492_ vssd1 vssd1 vccd1 vccd1 _1071_ sky130_fd_sc_hd__or2_1
XFILLER_40_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1991__A1 net28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2034__A _1342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input31_A SBsouth_in[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output118_A net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1631_ CB_0.config_dataA\[19\] CB_0.config_dataA\[18\] _1298_ vssd1 vssd1 vccd1 vccd1
+ _0393_ sky130_fd_sc_hd__or3b_1
X_2680_ SB0.route_sel\[80\] SB0.route_sel\[79\] net239 vssd1 vssd1 vccd1 vccd1 _0216_
+ sky130_fd_sc_hd__mux2_1
X_1700_ SB0.route_sel\[67\] SB0.route_sel\[66\] vssd1 vssd1 vccd1 vccd1 _0462_ sky130_fd_sc_hd__and2_1
X_1562_ SB0.route_sel\[108\] SB0.route_sel\[109\] _1354_ _1355_ _1347_ vssd1 vssd1
+ vccd1 vccd1 _1356_ sky130_fd_sc_hd__a311o_1
Xclkbuf_leaf_3_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1493_ _1184_ _1185_ vssd1 vssd1 vccd1 vccd1 _1287_ sky130_fd_sc_hd__nor2_1
XFILLER_39_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2114_ net152 CB_1.config_dataA\[2\] CB_1.config_dataA\[3\] CB_1.config_dataA\[1\]
+ vssd1 vssd1 vccd1 vccd1 _0872_ sky130_fd_sc_hd__and4b_1
X_2045_ _0356_ _0802_ vssd1 vssd1 vccd1 vccd1 _0803_ sky130_fd_sc_hd__and2_2
X_3094_ clknet_leaf_20_clk _0302_ net216 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[14\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_clkbuf_2_2__f_clk_X clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2947_ clknet_leaf_30_clk _0155_ net189 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[19\]
+ sky130_fd_sc_hd__dfstp_1
X_1829_ net23 net24 net25 net26 net170 CB_0.config_dataA\[9\] vssd1 vssd1 vccd1 vccd1
+ _0591_ sky130_fd_sc_hd__mux4_1
X_2878_ clknet_leaf_4_clk _0086_ net199 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2150__A1 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2801_ clknet_leaf_14_clk _0009_ net222 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2732_ CB_0.config_dataB\[0\] CB_0.config_dataA\[19\] net265 vssd1 vssd1 vccd1 vccd1
+ _0268_ sky130_fd_sc_hd__mux2_1
X_2594_ CB_1.config_dataB\[14\] CB_1.config_dataB\[13\] net267 vssd1 vssd1 vccd1 vccd1
+ _0130_ sky130_fd_sc_hd__mux2_1
X_2663_ SB0.route_sel\[63\] SB0.route_sel\[62\] net255 vssd1 vssd1 vccd1 vccd1 _0199_
+ sky130_fd_sc_hd__mux2_1
X_1614_ net175 net176 vssd1 vssd1 vccd1 vccd1 _0376_ sky130_fd_sc_hd__nor2_1
Xfanout207 net229 vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout229 net62 vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__buf_2
Xfanout218 net229 vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__clkbuf_2
X_1476_ _1269_ _1265_ _1256_ _1255_ vssd1 vssd1 vccd1 vccd1 _1270_ sky130_fd_sc_hd__a2bb2o_1
X_1545_ _1177_ _1178_ net51 SB0.route_sel\[37\] SB0.route_sel\[36\] vssd1 vssd1 vccd1
+ vccd1 _1339_ sky130_fd_sc_hd__o2111a_1
X_3077_ clknet_leaf_12_clk _0285_ net224 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[17\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_fanout266_A net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2028_ SB0.route_sel\[52\] SB0.route_sel\[53\] vssd1 vssd1 vccd1 vccd1 _0786_ sky130_fd_sc_hd__nor2_1
XANTENNA__1946__A1 _1321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2199__A1 _0831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1705__B1_N net41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2123__A1 net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput7 CBeast_in[2] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__buf_2
X_3000_ clknet_leaf_1_clk _0208_ net196 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[72\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_34_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2715_ CB_0.config_dataA\[3\] CB_0.config_dataA\[2\] net248 vssd1 vssd1 vccd1 vccd1
+ _0251_ sky130_fd_sc_hd__mux2_1
XANTENNA__2403__Y net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2577_ net411 LE_1A.edge_mode net230 vssd1 vssd1 vccd1 vccd1 _0113_ sky130_fd_sc_hd__mux2_1
X_2646_ SB0.route_sel\[46\] SB0.route_sel\[45\] net256 vssd1 vssd1 vccd1 vccd1 _0182_
+ sky130_fd_sc_hd__mux2_1
X_1459_ net153 net155 net157 net159 vssd1 vssd1 vccd1 vccd1 _1253_ sky130_fd_sc_hd__and4b_1
X_1528_ SB0.route_sel\[33\] SB0.route_sel\[32\] vssd1 vssd1 vccd1 vccd1 _1322_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout171_X net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1616__B1 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1919__A1 net24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1778__S0 CB_0.config_dataA\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1607__A0 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output100_A net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2500_ LEI0.config_data\[38\] net387 net268 vssd1 vssd1 vccd1 vccd1 _0039_ sky130_fd_sc_hd__mux2_1
X_2431_ SB0.route_sel\[4\] _1156_ vssd1 vssd1 vccd1 vccd1 _1131_ sky130_fd_sc_hd__nor2_1
X_2293_ CB_1.config_dataB\[14\] _1046_ _1048_ vssd1 vssd1 vccd1 vccd1 _1049_ sky130_fd_sc_hd__and3b_1
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2099__A0 net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2362_ _1263_ _1087_ _1264_ vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__a21o_1
XFILLER_24_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2629_ SB0.route_sel\[29\] SB0.route_sel\[28\] net237 vssd1 vssd1 vccd1 vccd1 _0165_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__2014__B1 _0758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input61_A le_nrst vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1843__A3 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2980_ clknet_leaf_22_clk _0188_ net214 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[52\]
+ sky130_fd_sc_hd__dfstp_1
X_1793_ net27 net28 net172 vssd1 vssd1 vccd1 vccd1 _0555_ sky130_fd_sc_hd__mux2_1
Xinput21 CBnorth_in[2] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__buf_2
X_1862_ net121 _0430_ _1221_ vssd1 vssd1 vccd1 vccd1 _0624_ sky130_fd_sc_hd__mux2_1
Xinput10 CBeast_in[5] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__buf_2
X_1931_ net167 _0339_ vssd1 vssd1 vccd1 vccd1 _0691_ sky130_fd_sc_hd__nand2_1
XANTENNA__2253__A0 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput43 SBwest_in[0] vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__clkbuf_1
Xinput32 SBsouth_in[12] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__buf_1
Xinput54 SBwest_in[7] vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__buf_1
X_2414_ SB0.route_sel\[25\] SB0.route_sel\[24\] SB0.route_sel\[26\] _1171_ vssd1 vssd1
+ vccd1 vccd1 _1120_ sky130_fd_sc_hd__a2bb2o_1
X_2345_ net122 _0412_ _0394_ vssd1 vssd1 vccd1 vccd1 _1079_ sky130_fd_sc_hd__mux2_1
X_2276_ net180 _0781_ vssd1 vssd1 vccd1 vccd1 _1032_ sky130_fd_sc_hd__nand2_1
XANTENNA__2409__X net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1598__A2 _0359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1834__A3 _1344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2244__A0 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout134_X net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2250__A3 _0822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2061_ _0427_ _0818_ vssd1 vssd1 vccd1 vccd1 _0819_ sky130_fd_sc_hd__nand2_4
X_2130_ _0819_ _0822_ _0816_ _0813_ CB_1.config_dataA\[9\] net149 vssd1 vssd1 vccd1
+ vccd1 _0888_ sky130_fd_sc_hd__mux4_1
XFILLER_19_241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1914_ _0655_ _0673_ CB_0.config_dataB\[6\] vssd1 vssd1 vccd1 vccd1 _0674_ sky130_fd_sc_hd__o21ai_1
XFILLER_34_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2963_ clknet_leaf_25_clk _0171_ net197 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[35\]
+ sky130_fd_sc_hd__dfstp_1
X_1845_ _1220_ net169 vssd1 vssd1 vccd1 vccd1 _0607_ sky130_fd_sc_hd__nor2_1
X_1776_ _0535_ _0536_ _0537_ _0534_ vssd1 vssd1 vccd1 vccd1 _0538_ sky130_fd_sc_hd__o31a_2
X_2894_ clknet_leaf_21_clk _0102_ net215 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2328_ net137 _1070_ _0520_ vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__mux2_1
XANTENNA__1752__A2 net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2259_ net139 net126 net129 net133 LEI0.config_data\[33\] LEI0.config_data\[34\]
+ vssd1 vssd1 vccd1 vccd1 _1015_ sky130_fd_sc_hd__mux4_1
XANTENNA__2034__B _0791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input24_A CBnorth_in[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2208__A0 _0816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1630_ _0391_ vssd1 vssd1 vccd1 vccd1 _0392_ sky130_fd_sc_hd__inv_2
XANTENNA__1783__B net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output92_A net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1561_ SB0.route_sel\[108\] SB0.route_sel\[109\] net33 vssd1 vssd1 vccd1 vccd1 _1355_
+ sky130_fd_sc_hd__a21oi_1
X_1492_ net131 _1259_ _1281_ _1285_ vssd1 vssd1 vccd1 vccd1 _1286_ sky130_fd_sc_hd__o31a_1
X_2044_ _1208_ SB0.route_sel\[102\] _1210_ SB0.route_sel\[97\] _0801_ vssd1 vssd1
+ vccd1 vccd1 _0802_ sky130_fd_sc_hd__a221o_1
X_2113_ _1235_ _0865_ _0870_ vssd1 vssd1 vccd1 vccd1 _0871_ sky130_fd_sc_hd__a21oi_1
X_3093_ clknet_leaf_20_clk _0301_ net217 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[13\]
+ sky130_fd_sc_hd__dfstp_2
X_2877_ clknet_leaf_4_clk net328 net200 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2406__Y net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2946_ clknet_leaf_30_clk _0154_ net189 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[18\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_17_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1759_ net159 net155 net153 net157 vssd1 vssd1 vccd1 vccd1 _0521_ sky130_fd_sc_hd__and4bb_1
X_1828_ _0586_ _0589_ CB_0.config_dataA\[11\] vssd1 vssd1 vccd1 vccd1 _0590_ sky130_fd_sc_hd__mux2_1
XANTENNA__2150__A2 net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input27_X net27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2731_ CB_0.config_dataA\[19\] CB_0.config_dataA\[18\] net265 vssd1 vssd1 vccd1 vccd1
+ _0267_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_14_clk_A clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2800_ clknet_leaf_14_clk _0008_ net222 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1613_ net137 _0373_ _0371_ vssd1 vssd1 vccd1 vccd1 _0375_ sky130_fd_sc_hd__mux2_1
XANTENNA__1794__A net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2593_ net179 net181 net267 vssd1 vssd1 vccd1 vccd1 _0129_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_29_clk_A clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2662_ SB0.route_sel\[62\] SB0.route_sel\[61\] net255 vssd1 vssd1 vccd1 vccd1 _0198_
+ sky130_fd_sc_hd__mux2_1
X_1544_ SB0.route_sel\[35\] SB0.route_sel\[34\] _1331_ _1335_ _1337_ vssd1 vssd1 vccd1
+ vccd1 _1338_ sky130_fd_sc_hd__a221o_1
Xfanout208 net210 vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__clkbuf_4
Xfanout219 net220 vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__clkbuf_4
X_1475_ SB0.route_sel\[58\] SB0.route_sel\[59\] _1267_ _1268_ _1255_ vssd1 vssd1 vccd1
+ vccd1 _1269_ sky130_fd_sc_hd__a41o_1
XANTENNA__2132__A2 _0828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3076_ clknet_leaf_12_clk _0284_ net228 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[16\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_39_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout259_A net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2027_ SB0.route_sel\[55\] SB0.route_sel\[54\] vssd1 vssd1 vccd1 vccd1 _0785_ sky130_fd_sc_hd__and2b_1
XANTENNA__1946__A2 _1297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2929_ clknet_leaf_27_clk _0137_ net194 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[1\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_20_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput8 CBeast_in[3] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__buf_2
X_2714_ CB_0.config_dataA\[2\] CB_0.config_dataA\[1\] net248 vssd1 vssd1 vccd1 vccd1
+ _0250_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_34_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1561__B1 net33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1527_ _1318_ _1320_ vssd1 vssd1 vccd1 vccd1 _1321_ sky130_fd_sc_hd__nor2_2
X_2645_ SB0.route_sel\[45\] SB0.route_sel\[44\] net256 vssd1 vssd1 vccd1 vccd1 _0181_
+ sky130_fd_sc_hd__mux2_1
X_2576_ LE_1A.edge_mode LE_1A.config_data\[16\] net230 vssd1 vssd1 vccd1 vccd1 _0112_
+ sky130_fd_sc_hd__mux2_1
X_1458_ _1250_ _1251_ vssd1 vssd1 vccd1 vccd1 _1252_ sky130_fd_sc_hd__nand2b_1
X_1389_ SB0.route_sel\[40\] vssd1 vssd1 vccd1 vccd1 _1183_ sky130_fd_sc_hd__inv_2
X_3059_ clknet_leaf_11_clk _0267_ net221 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[19\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1919__A2 net25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2224__A1_N _0781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1552__A0 _1273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1607__A1 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1791__A0 _0473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2430_ _1129_ _1130_ _0407_ vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__a21boi_1
X_2361_ net177 net178 _1258_ _0781_ vssd1 vssd1 vccd1 vccd1 _1087_ sky130_fd_sc_hd__a31o_1
XFILLER_49_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2292_ CB_1.config_dataB\[15\] _1047_ vssd1 vssd1 vccd1 vccd1 _1048_ sky130_fd_sc_hd__nand2_1
XANTENNA__2099__A1 net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1782__A0 _0430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2559_ LE_1A.config_data\[0\] LE_0B.reset_mode net230 vssd1 vssd1 vccd1 vccd1 _0095_
+ sky130_fd_sc_hd__mux2_1
X_2628_ SB0.route_sel\[28\] SB0.route_sel\[27\] net237 vssd1 vssd1 vccd1 vccd1 _0164_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__1837__A1 _1297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1837__B2 _1273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1921__S CB_0.config_dataB\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input54_A SBwest_in[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1930_ CB_0.config_dataB\[2\] _0680_ _0688_ _0689_ vssd1 vssd1 vccd1 vccd1 _0690_
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__2253__A1 net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1792_ net16 _0545_ _0546_ net17 vssd1 vssd1 vccd1 vccd1 _0554_ sky130_fd_sc_hd__o22a_1
Xinput22 CBnorth_in[3] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__buf_2
X_1861_ _0538_ _0608_ _0609_ _0512_ CB_0.config_dataA\[15\] vssd1 vssd1 vccd1 vccd1
+ _0623_ sky130_fd_sc_hd__o221a_1
Xinput11 CBeast_in[6] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__buf_2
Xinput55 SBwest_in[8] vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__buf_1
Xinput44 SBwest_in[10] vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__buf_1
Xinput33 SBsouth_in[13] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__buf_1
X_2344_ net137 _1078_ _0431_ vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__mux2_1
X_2413_ SB0.route_sel\[28\] _1172_ vssd1 vssd1 vccd1 vccd1 _1119_ sky130_fd_sc_hd__nor2_1
X_2275_ _1029_ _1030_ CB_1.config_dataB\[15\] _1027_ vssd1 vssd1 vccd1 vccd1 _1031_
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__2492__A1 LEI0.config_data\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2244__A1 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout241_A net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1755__A0 net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout127_X net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input1_X net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2180__A0 _0781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1522__A3 net52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2474__A1 LEI0.config_data\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2060_ _1157_ SB0.route_sel\[6\] _1160_ SB0.route_sel\[1\] _0817_ vssd1 vssd1 vccd1
+ vccd1 _0818_ sky130_fd_sc_hd__a221o_1
XFILLER_19_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1913_ _1229_ _0665_ _0672_ vssd1 vssd1 vccd1 vccd1 _0673_ sky130_fd_sc_hd__a21oi_1
X_2893_ clknet_leaf_21_clk _0101_ net216 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_2962_ clknet_leaf_25_clk _0170_ net197 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[34\]
+ sky130_fd_sc_hd__dfstp_1
X_1844_ _0605_ vssd1 vssd1 vccd1 vccd1 _0606_ sky130_fd_sc_hd__inv_2
XANTENNA__1752__A3 net22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1775_ _1200_ SB0.route_sel\[85\] vssd1 vssd1 vccd1 vccd1 _0537_ sky130_fd_sc_hd__nor2_1
XANTENNA__1737__B1 net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2327_ _0538_ net123 _0521_ vssd1 vssd1 vccd1 vccd1 _1070_ sky130_fd_sc_hd__mux2_1
X_2258_ CB_1.config_dataB\[11\] _1013_ _1007_ CB_1.config_dataB\[10\] _1012_ vssd1
+ vssd1 vccd1 vccd1 _1014_ sky130_fd_sc_hd__a2111oi_1
XANTENNA__2162__A0 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2189_ CB_1.config_dataB\[1\] CB_1.config_dataB\[3\] vssd1 vssd1 vccd1 vccd1 _0945_
+ sky130_fd_sc_hd__nand2_1
XANTENNA_input17_A CBnorth_in[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1900__A0 net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2208__A1 _0819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_9_Left_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1560_ net119 SB0.route_sel\[110\] net47 vssd1 vssd1 vccd1 vccd1 _1354_ sky130_fd_sc_hd__a21bo_1
XANTENNA__1719__B1 net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2112_ CB_1.config_dataA\[3\] _0868_ _0869_ _0852_ vssd1 vssd1 vccd1 vccd1 _0870_
+ sky130_fd_sc_hd__o22a_1
X_1491_ CB_1.config_dataA\[16\] net142 net143 net144 vssd1 vssd1 vccd1 vccd1 _1285_
+ sky130_fd_sc_hd__or4bb_1
X_2043_ SB0.route_sel\[100\] SB0.route_sel\[101\] vssd1 vssd1 vccd1 vccd1 _0801_ sky130_fd_sc_hd__nor2_1
X_3092_ clknet_leaf_20_clk _0300_ net216 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[12\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_60_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1827_ net27 net28 net16 net17 net170 CB_0.config_dataA\[9\] vssd1 vssd1 vccd1 vccd1
+ _0589_ sky130_fd_sc_hd__mux4_1
X_2876_ clknet_leaf_4_clk net301 net200 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_2945_ clknet_leaf_30_clk _0153_ net188 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[17\]
+ sky130_fd_sc_hd__dfstp_1
X_1758_ _1274_ _0450_ vssd1 vssd1 vccd1 vccd1 _0520_ sky130_fd_sc_hd__nand2_1
X_1689_ _1324_ _0450_ vssd1 vssd1 vccd1 vccd1 _0451_ sky130_fd_sc_hd__nand2_1
XANTENNA__2135__A0 net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input9_A CBeast_in[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3085__SET_B net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2150__A3 net12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_35_Left_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2760__S net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2730_ CB_0.config_dataA\[18\] CB_0.config_dataA\[17\] net265 vssd1 vssd1 vccd1 vccd1
+ _0266_ sky130_fd_sc_hd__mux2_1
X_2661_ SB0.route_sel\[61\] SB0.route_sel\[60\] net255 vssd1 vssd1 vccd1 vccd1 _0197_
+ sky130_fd_sc_hd__mux2_1
X_2592_ net181 CB_1.config_dataB\[11\] net266 vssd1 vssd1 vccd1 vccd1 _0128_ sky130_fd_sc_hd__mux2_1
Xfanout209 net210 vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__clkbuf_2
X_1474_ SB0.route_sel\[60\] SB0.route_sel\[61\] net40 vssd1 vssd1 vccd1 vccd1 _1268_
+ sky130_fd_sc_hd__a21bo_1
X_1612_ SB0.route_sel\[25\] SB0.route_sel\[24\] vssd1 vssd1 vccd1 vccd1 _0374_ sky130_fd_sc_hd__nand2_1
X_1543_ _1249_ _1334_ vssd1 vssd1 vccd1 vccd1 _1337_ sky130_fd_sc_hd__nor2_1
X_3075_ clknet_leaf_10_clk _0283_ net221 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[15\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_59_Left_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2026_ _1318_ _0783_ vssd1 vssd1 vccd1 vccd1 _0784_ sky130_fd_sc_hd__nor2_2
XANTENNA__1946__A3 _1273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2859_ clknet_leaf_4_clk _0067_ net199 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2199__A3 _0838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2433__X net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2928_ clknet_leaf_23_clk _0136_ net194 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[0\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_20_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_2_3__f_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput9 CBeast_in[4] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__buf_2
X_2713_ CB_0.config_dataA\[1\] net174 net248 vssd1 vssd1 vccd1 vccd1 _0249_ sky130_fd_sc_hd__mux2_1
X_2644_ SB0.route_sel\[44\] SB0.route_sel\[43\] net256 vssd1 vssd1 vccd1 vccd1 _0180_
+ sky130_fd_sc_hd__mux2_1
X_1457_ CB_0.config_dataA\[19\] CB_0.config_dataA\[18\] vssd1 vssd1 vccd1 vccd1 _1251_
+ sky130_fd_sc_hd__and2b_1
X_2575_ LE_1A.config_data\[16\] LE_1A.config_data\[15\] net231 vssd1 vssd1 vccd1 vccd1
+ _0111_ sky130_fd_sc_hd__mux2_1
X_1526_ _1180_ SB0.route_sel\[45\] _1182_ SB0.route_sel\[46\] _1319_ vssd1 vssd1 vccd1
+ vccd1 _1320_ sky130_fd_sc_hd__o221a_1
X_3058_ clknet_leaf_12_clk _0266_ net221 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[18\]
+ sky130_fd_sc_hd__dfstp_2
XANTENNA_fanout271_A net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1388_ SB0.route_sel\[47\] vssd1 vssd1 vccd1 vccd1 _1182_ sky130_fd_sc_hd__inv_2
XFILLER_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2009_ _0700_ _0702_ LE_0B.config_data\[9\] vssd1 vssd1 vccd1 vccd1 _0769_ sky130_fd_sc_hd__a21boi_1
XANTENNA__1919__A3 net26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1552__A1 _1297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_13_clk_A clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1607__A2 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_28_clk_A clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2073__X _0831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1791__A1 _0492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2291_ _0831_ _0838_ _0827_ _0835_ net179 net180 vssd1 vssd1 vccd1 vccd1 _1047_ sky130_fd_sc_hd__mux4_1
X_2360_ _0461_ _1086_ _0463_ vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__a21o_1
XFILLER_49_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_10_Right_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_22_Left_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2559__A0 LE_1A.config_data\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput110 net110 vssd1 vssd1 vccd1 vccd1 SBwest_out[1] sky130_fd_sc_hd__buf_2
X_2627_ SB0.route_sel\[27\] SB0.route_sel\[26\] net255 vssd1 vssd1 vccd1 vccd1 _0163_
+ sky130_fd_sc_hd__mux2_1
X_2489_ net384 net336 net251 vssd1 vssd1 vccd1 vccd1 _0028_ sky130_fd_sc_hd__mux2_1
X_2558_ LE_1B.dff1_out _1247_ _1153_ vssd1 vssd1 vccd1 vccd1 _0094_ sky130_fd_sc_hd__a21bo_1
X_1509_ SB0.route_sel\[41\] SB0.route_sel\[40\] vssd1 vssd1 vccd1 vccd1 _1303_ sky130_fd_sc_hd__nand2_1
XFILLER_23_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input47_A SBwest_in[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1860_ _1221_ _0473_ _0621_ net168 vssd1 vssd1 vccd1 vccd1 _0622_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_44_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_26_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_14_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput23 CBnorth_in[4] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__buf_2
X_1791_ _0473_ _0492_ _0538_ _0512_ net172 net171 vssd1 vssd1 vccd1 vccd1 _0553_ sky130_fd_sc_hd__mux4_1
Xinput12 CBeast_in[7] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__buf_2
Xinput56 SBwest_in[9] vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__buf_1
Xinput45 SBwest_in[11] vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__buf_1
Xinput34 SBsouth_in[1] vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__buf_1
X_2343_ net122 _0448_ _0432_ vssd1 vssd1 vccd1 vccd1 _1078_ sky130_fd_sc_hd__mux2_1
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2274_ net180 _0797_ _1028_ vssd1 vssd1 vccd1 vccd1 _1030_ sky130_fd_sc_hd__a21oi_1
X_2412_ _1117_ _1118_ _1342_ vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__o21a_1
XFILLER_37_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_17_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1989_ _1232_ _0513_ _0743_ vssd1 vssd1 vccd1 vccd1 _0749_ sky130_fd_sc_hd__or3_1
XANTENNA__2244__A2 net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1755__A1 net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2070__Y _0828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1843_ net139 net125 net129 net133 LEI0.config_data\[36\] LEI0.config_data\[37\]
+ vssd1 vssd1 vccd1 vccd1 _0605_ sky130_fd_sc_hd__mux4_1
X_1912_ _0651_ _0666_ _0667_ _0671_ vssd1 vssd1 vccd1 vccd1 _0672_ sky130_fd_sc_hd__a31o_1
XANTENNA__2261__X _1017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2892_ clknet_leaf_21_clk _0100_ net216 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_2961_ clknet_leaf_26_clk _0169_ net195 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[33\]
+ sky130_fd_sc_hd__dfstp_1
Xclkbuf_leaf_6_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1774_ SB0.route_sel\[86\] SB0.route_sel\[87\] vssd1 vssd1 vccd1 vccd1 _0536_ sky130_fd_sc_hd__and2b_1
X_2326_ net137 _1069_ _0494_ vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__mux2_1
X_2257_ _0827_ _0831_ _0835_ _0838_ _1245_ CB_1.config_dataB\[9\] vssd1 vssd1 vccd1
+ vccd1 _1013_ sky130_fd_sc_hd__mux4_1
XANTENNA__2162__A1 net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1673__A0 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_40_Left_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2188_ _1243_ _0936_ _0943_ vssd1 vssd1 vccd1 vccd1 _0944_ sky130_fd_sc_hd__a21oi_1
XANTENNA__2758__S net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1900__A1 net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2208__A2 _0813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2241__B _0781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1490_ net145 net144 vssd1 vssd1 vccd1 vccd1 _1284_ sky130_fd_sc_hd__nand2b_1
Xhold1 LE_0B.config_data\[14\] vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__dlygate4sd3_1
X_2111_ net4 net5 net152 vssd1 vssd1 vccd1 vccd1 _0869_ sky130_fd_sc_hd__mux2_1
X_2042_ CB_1.config_dataA\[5\] _1238_ vssd1 vssd1 vccd1 vccd1 _0800_ sky130_fd_sc_hd__or2_1
X_3091_ clknet_leaf_21_clk _0299_ net216 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[11\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1655__A0 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_8_Right_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1826_ _1217_ CB_0.config_dataA\[11\] vssd1 vssd1 vccd1 vccd1 _0588_ sky130_fd_sc_hd__nand2_1
X_2875_ clknet_leaf_4_clk _0083_ net200 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_2944_ clknet_leaf_30_clk _0152_ net188 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[16\]
+ sky130_fd_sc_hd__dfstp_1
X_1688_ CB_0.config_dataA\[18\] CB_0.config_dataA\[19\] vssd1 vssd1 vccd1 vccd1 _0450_
+ sky130_fd_sc_hd__and2b_1
X_1757_ _0516_ _0518_ vssd1 vssd1 vccd1 vccd1 _0519_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_39_Right_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2135__A1 net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2309_ _1025_ _1053_ _1063_ _1064_ vssd1 vssd1 vccd1 vccd1 _1065_ sky130_fd_sc_hd__a22oi_2
XPHY_EDGE_ROW_48_Right_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_57_Right_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output116_A net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1611_ net22 net123 _0372_ vssd1 vssd1 vccd1 vccd1 _0373_ sky130_fd_sc_hd__mux2_1
X_2660_ SB0.route_sel\[60\] SB0.route_sel\[59\] net255 vssd1 vssd1 vccd1 vccd1 _0196_
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2591_ CB_1.config_dataB\[11\] CB_1.config_dataB\[10\] net266 vssd1 vssd1 vccd1 vccd1
+ _0127_ sky130_fd_sc_hd__mux2_1
X_1473_ SB0.route_sel\[63\] SB0.route_sel\[62\] _1266_ vssd1 vssd1 vccd1 vccd1 _1267_
+ sky130_fd_sc_hd__a21bo_1
X_1542_ SB0.route_sel\[35\] SB0.route_sel\[34\] vssd1 vssd1 vccd1 vccd1 _1336_ sky130_fd_sc_hd__nand2_1
X_3074_ clknet_leaf_10_clk _0282_ net221 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[14\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_35_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2025_ _1180_ _1181_ _0782_ vssd1 vssd1 vccd1 vccd1 _0783_ sky130_fd_sc_hd__a21oi_1
XFILLER_62_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2927_ clknet_leaf_24_clk _0135_ net211 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[19\]
+ sky130_fd_sc_hd__dfstp_1
X_1809_ _1216_ _0567_ _0570_ _0564_ CB_0.config_dataA\[6\] vssd1 vssd1 vccd1 vccd1
+ _0571_ sky130_fd_sc_hd__o221a_1
X_2858_ clknet_leaf_5_clk _0066_ net203 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__1800__A0 net23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2789_ LE_1B.edge_mode LE_1B.config_data\[16\] net233 vssd1 vssd1 vccd1 vccd1 _0325_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_20_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1867__A0 net27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2771__S net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input32_X net32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2283__A0 _0819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2712_ CB_0.config_dataA\[0\] net397 net269 vssd1 vssd1 vccd1 vccd1 _0248_ sky130_fd_sc_hd__mux2_1
X_2574_ LE_1A.config_data\[15\] net302 net258 vssd1 vssd1 vccd1 vccd1 _0110_ sky130_fd_sc_hd__mux2_1
X_2643_ SB0.route_sel\[43\] SB0.route_sel\[42\] net256 vssd1 vssd1 vccd1 vccd1 _0179_
+ sky130_fd_sc_hd__mux2_1
X_1456_ CB_0.config_dataA\[17\] CB_0.config_dataA\[16\] vssd1 vssd1 vccd1 vccd1 _1250_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__1613__X _0375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1525_ SB0.route_sel\[43\] SB0.route_sel\[42\] vssd1 vssd1 vccd1 vccd1 _1319_ sky130_fd_sc_hd__or2_1
X_1387_ SB0.route_sel\[45\] vssd1 vssd1 vccd1 vccd1 _1181_ sky130_fd_sc_hd__inv_2
X_3057_ clknet_leaf_11_clk _0265_ net221 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[17\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__1864__A3 _0391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout264_A net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2008_ _0675_ _0765_ _0766_ _0767_ _0731_ vssd1 vssd1 vccd1 vccd1 _0768_ sky130_fd_sc_hd__o221a_1
XANTENNA__2510__A1 _0645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1552__A2 _1321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1607__A3 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2290_ _1041_ _1043_ _1045_ _1039_ CB_1.config_dataB\[15\] vssd1 vssd1 vccd1 vccd1
+ _1046_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_47_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput111 net111 vssd1 vssd1 vccd1 vccd1 SBwest_out[2] sky130_fd_sc_hd__buf_2
Xoutput100 net100 vssd1 vssd1 vccd1 vccd1 SBsouth_out[5] sky130_fd_sc_hd__buf_2
X_2626_ SB0.route_sel\[26\] SB0.route_sel\[25\] net255 vssd1 vssd1 vccd1 vccd1 _0162_
+ sky130_fd_sc_hd__mux2_1
X_2557_ net60 _1065_ vssd1 vssd1 vccd1 vccd1 _1153_ sky130_fd_sc_hd__nand2_1
X_1508_ net24 net125 _1301_ vssd1 vssd1 vccd1 vccd1 _1302_ sky130_fd_sc_hd__mux2_1
X_1439_ CB_0.config_dataB\[15\] vssd1 vssd1 vccd1 vccd1 _1233_ sky130_fd_sc_hd__inv_2
X_2488_ net336 LEI0.config_data\[25\] net244 vssd1 vssd1 vccd1 vccd1 _0027_ sky130_fd_sc_hd__mux2_1
X_3109_ clknet_leaf_0_clk net281 net190 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_23_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2793__Q LEI0.config_data\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1790_ CB_0.config_dataA\[7\] _0549_ _0550_ _0551_ vssd1 vssd1 vccd1 vccd1 _0552_
+ sky130_fd_sc_hd__o22ai_1
Xinput13 CBeast_in[8] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__buf_2
Xinput57 config_data_in vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__clkbuf_1
Xinput24 CBnorth_in[5] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__buf_2
Xinput46 SBwest_in[12] vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__buf_1
Xinput35 SBsouth_in[2] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__buf_1
X_2411_ SB0.route_sel\[33\] _1179_ _1177_ _1178_ vssd1 vssd1 vccd1 vccd1 _1118_ sky130_fd_sc_hd__a2bb2o_1
X_2342_ net137 _1077_ _0371_ vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__mux2_1
X_2273_ net180 _0803_ vssd1 vssd1 vccd1 vccd1 _1029_ sky130_fd_sc_hd__or2_1
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2244__A3 net12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2229__A0 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1988_ net161 _0493_ _0736_ _0747_ vssd1 vssd1 vccd1 vccd1 _0748_ sky130_fd_sc_hd__a211o_1
XANTENNA__3039__Q net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_12_clk_A clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout227_A net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_27_clk_A clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2609_ SB0.route_sel\[9\] SB0.route_sel\[8\] net231 vssd1 vssd1 vccd1 vccd1 _0145_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_58_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2329__B _0492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1691__A1 net27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2468__A0 LEI0.config_data\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_2_2__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_2_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_41_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout190 net192 vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__clkbuf_4
XANTENNA__2171__A2 LE_1A.config_data\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1711__X _0473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2960_ clknet_leaf_27_clk _0168_ net195 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[32\]
+ sky130_fd_sc_hd__dfstp_1
X_1842_ _0603_ _0573_ _0572_ vssd1 vssd1 vccd1 vccd1 _0604_ sky130_fd_sc_hd__mux2_1
X_1911_ CB_0.config_dataB\[5\] _1229_ _0670_ _0669_ vssd1 vssd1 vccd1 vccd1 _0671_
+ sky130_fd_sc_hd__o31a_1
X_1773_ SB0.route_sel\[82\] SB0.route_sel\[83\] vssd1 vssd1 vccd1 vccd1 _0535_ sky130_fd_sc_hd__nor2_1
X_2891_ clknet_leaf_20_clk net279 net216 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_2325_ _0512_ net123 _0495_ vssd1 vssd1 vccd1 vccd1 _1069_ sky130_fd_sc_hd__mux2_1
X_2256_ _1003_ _1009_ _1011_ vssd1 vssd1 vccd1 vccd1 _1012_ sky130_fd_sc_hd__o21a_1
X_2187_ _1241_ CB_1.config_dataB\[3\] _0937_ _0938_ _0942_ vssd1 vssd1 vccd1 vccd1
+ _0943_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_63_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2208__A3 _0822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2 _0087_ vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__dlygate4sd3_1
X_2110_ net9 net10 net11 net12 net152 CB_1.config_dataA\[1\] vssd1 vssd1 vccd1 vccd1
+ _0868_ sky130_fd_sc_hd__mux4_1
X_2041_ CB_1.config_dataA\[5\] _1238_ vssd1 vssd1 vccd1 vccd1 _0799_ sky130_fd_sc_hd__nor2_1
X_3090_ clknet_leaf_20_clk _0298_ net216 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[10\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__1655__A1 net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2943_ clknet_leaf_28_clk _0151_ net188 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[15\]
+ sky130_fd_sc_hd__dfstp_1
X_1825_ CB_0.config_dataA\[11\] _0577_ vssd1 vssd1 vccd1 vccd1 _0587_ sky130_fd_sc_hd__nand2_1
X_1756_ CB_0.config_dataA\[3\] _0514_ _0517_ _0367_ vssd1 vssd1 vccd1 vccd1 _0518_
+ sky130_fd_sc_hd__o22a_1
X_2874_ clknet_leaf_4_clk net307 net200 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_1687_ _0391_ net121 _0447_ _0430_ _1154_ _1165_ vssd1 vssd1 vccd1 vccd1 _0449_ sky130_fd_sc_hd__mux4_1
X_2308_ _1018_ _1058_ _1052_ vssd1 vssd1 vccd1 vccd1 _1064_ sky130_fd_sc_hd__a21oi_1
XANTENNA__1999__A _0758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2239_ _1245_ _1342_ _0791_ CB_1.config_dataB\[9\] vssd1 vssd1 vccd1 vccd1 _0995_
+ sky130_fd_sc_hd__a31oi_1
XTAP_TAPCELL_ROW_0_132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1949__A2 _0339_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1526__X _1320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input22_A CBnorth_in[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1610_ net153 net155 net157 net159 vssd1 vssd1 vccd1 vccd1 _0372_ sky130_fd_sc_hd__and4bb_1
X_2590_ CB_1.config_dataB\[10\] CB_1.config_dataB\[9\] net266 vssd1 vssd1 vccd1 vccd1
+ _0126_ sky130_fd_sc_hd__mux2_1
XFILLER_12_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1472_ SB0.route_sel\[60\] SB0.route_sel\[61\] net54 vssd1 vssd1 vccd1 vccd1 _1266_
+ sky130_fd_sc_hd__and3_1
X_1541_ net132 _1259_ _1330_ _1334_ vssd1 vssd1 vccd1 vccd1 _1335_ sky130_fd_sc_hd__o31a_1
X_3073_ clknet_leaf_10_clk _0281_ net221 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[13\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2024_ _1182_ SB0.route_sel\[46\] SB0.route_sel\[41\] _1183_ vssd1 vssd1 vccd1 vccd1
+ _0782_ sky130_fd_sc_hd__a22o_1
X_2857_ clknet_leaf_5_clk net309 net203 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__1800__A1 net24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2926_ clknet_leaf_18_clk _0134_ net217 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[18\]
+ sky130_fd_sc_hd__dfstp_1
X_1808_ _0550_ _0568_ _0569_ vssd1 vssd1 vccd1 vccd1 _0570_ sky130_fd_sc_hd__o21a_1
X_2788_ LE_1B.config_data\[16\] net366 net233 vssd1 vssd1 vccd1 vccd1 _0324_ sky130_fd_sc_hd__mux2_1
X_1739_ _1249_ _1261_ _0460_ vssd1 vssd1 vccd1 vccd1 _0501_ sky130_fd_sc_hd__nor3_1
XANTENNA__1867__A1 net28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2347__A2 _0430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1555__B1 net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input25_X net25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2711_ net119 SB0.route_sel\[110\] net266 vssd1 vssd1 vccd1 vccd1 _0247_ sky130_fd_sc_hd__mux2_1
XANTENNA__2283__A1 _0822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2573_ net302 LE_1A.config_data\[13\] net258 vssd1 vssd1 vccd1 vccd1 _0109_ sky130_fd_sc_hd__mux2_1
X_2642_ SB0.route_sel\[42\] SB0.route_sel\[41\] net256 vssd1 vssd1 vccd1 vccd1 _0178_
+ sky130_fd_sc_hd__mux2_1
X_1524_ _1303_ _1304_ _1313_ _1317_ vssd1 vssd1 vccd1 vccd1 _1318_ sky130_fd_sc_hd__a22oi_4
X_1386_ SB0.route_sel\[44\] vssd1 vssd1 vccd1 vccd1 _1180_ sky130_fd_sc_hd__inv_2
X_1455_ net128 vssd1 vssd1 vccd1 vccd1 _1249_ sky130_fd_sc_hd__inv_2
X_3056_ clknet_leaf_11_clk _0264_ net221 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[16\]
+ sky130_fd_sc_hd__dfstp_1
X_2007_ LE_0B.config_data\[15\] _0703_ _0676_ vssd1 vssd1 vccd1 vccd1 _0767_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout257_A net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1785__A0 _0447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2460__X net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2909_ clknet_leaf_17_clk _0117_ net213 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[1\]
+ sky130_fd_sc_hd__dfstp_2
XANTENNA__1552__A3 _1345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1537__B1 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1791__A3 _0512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1507_ net158 net154 net156 net160 vssd1 vssd1 vccd1 vccd1 _1301_ sky130_fd_sc_hd__and4bb_1
Xoutput112 net112 vssd1 vssd1 vccd1 vccd1 SBwest_out[3] sky130_fd_sc_hd__buf_2
X_2487_ net394 LEI0.config_data\[24\] net244 vssd1 vssd1 vccd1 vccd1 _0026_ sky130_fd_sc_hd__mux2_1
X_2556_ LE_1A.dff0_out _1247_ _1152_ vssd1 vssd1 vccd1 vccd1 _0093_ sky130_fd_sc_hd__a21o_1
Xoutput101 net101 vssd1 vssd1 vccd1 vccd1 SBsouth_out[6] sky130_fd_sc_hd__buf_2
X_2625_ SB0.route_sel\[25\] SB0.route_sel\[24\] net237 vssd1 vssd1 vccd1 vccd1 _0161_
+ sky130_fd_sc_hd__mux2_1
X_1438_ net161 vssd1 vssd1 vccd1 vccd1 _1232_ sky130_fd_sc_hd__inv_2
X_1369_ SB0.route_sel\[15\] vssd1 vssd1 vccd1 vccd1 _1163_ sky130_fd_sc_hd__inv_2
X_3108_ clknet_leaf_0_clk net288 net190 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_53_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3060__Q CB_0.config_dataB\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3039_ clknet_leaf_14_clk _0247_ net222 vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__dfstp_2
XFILLER_11_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1534__X _1328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2183__A0 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput25 CBnorth_in[6] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__buf_2
Xinput14 CBeast_in[9] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_4
Xinput36 SBsouth_in[3] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__clkbuf_1
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2341_ _0392_ net123 _0372_ vssd1 vssd1 vccd1 vccd1 _1077_ sky130_fd_sc_hd__mux2_1
Xinput58 config_en vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__clkbuf_2
Xinput47 SBwest_in[13] vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2410_ SB0.route_sel\[34\] SB0.route_sel\[35\] vssd1 vssd1 vccd1 vccd1 _1117_ sky130_fd_sc_hd__and2b_1
X_2272_ net179 CB_1.config_dataB\[15\] vssd1 vssd1 vccd1 vccd1 _1028_ sky130_fd_sc_hd__nand2b_1
XFILLER_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2229__A1 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1987_ net161 _0473_ vssd1 vssd1 vccd1 vccd1 _0747_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout122_A net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2539_ net350 net316 net244 vssd1 vssd1 vccd1 vccd1 _0076_ sky130_fd_sc_hd__mux2_1
XANTENNA__2165__A0 _0838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2608_ SB0.route_sel\[8\] SB0.route_sel\[7\] net231 vssd1 vssd1 vccd1 vccd1 _0144_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__2597__S net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1979__A0 net23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input52_A SBwest_in[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout180 CB_1.config_dataB\[12\] vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__buf_2
Xfanout191 net192 vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__clkbuf_4
X_1910_ net18 net19 net165 vssd1 vssd1 vccd1 vccd1 _0670_ sky130_fd_sc_hd__mux2_1
X_2890_ clknet_leaf_22_clk _0098_ net215 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__1682__A2 _0435_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1841_ LE_0A.config_data\[5\] LE_0A.config_data\[4\] _0543_ vssd1 vssd1 vccd1 vccd1
+ _0603_ sky130_fd_sc_hd__mux2_1
XANTENNA__1985__A3 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1772_ _0533_ _0529_ _0524_ _0523_ vssd1 vssd1 vccd1 vccd1 _0534_ sky130_fd_sc_hd__a2bb2o_1
X_2324_ net140 _1068_ _0341_ vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__mux2_1
X_2255_ CB_1.config_dataB\[11\] _1008_ _1010_ _0991_ vssd1 vssd1 vccd1 vccd1 _1011_
+ sky130_fd_sc_hd__o22a_1
X_2186_ CB_1.config_dataB\[1\] _1243_ _0941_ _0940_ vssd1 vssd1 vccd1 vccd1 _0942_
+ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_63_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2799__Q LEI0.config_data\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_11_clk_A clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold3 LE_0B.config_data\[15\] vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__dlygate4sd3_1
X_2040_ _1359_ _0335_ _0795_ _1237_ vssd1 vssd1 vccd1 vccd1 _0798_ sky130_fd_sc_hd__a31o_1
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2873_ clknet_leaf_4_clk net349 net200 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_2942_ clknet_leaf_28_clk _0150_ net188 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[14\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_clkbuf_leaf_26_clk_A clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1686_ _0447_ vssd1 vssd1 vccd1 vccd1 _0448_ sky130_fd_sc_hd__inv_2
X_1824_ net15 net20 net21 net22 net170 CB_0.config_dataA\[9\] vssd1 vssd1 vccd1 vccd1
+ _0586_ sky130_fd_sc_hd__mux4_1
X_1755_ net16 net17 net174 vssd1 vssd1 vccd1 vccd1 _0517_ sky130_fd_sc_hd__mux2_1
X_2238_ _1245_ _1318_ _0783_ vssd1 vssd1 vccd1 vccd1 _0994_ sky130_fd_sc_hd__or3_1
X_2307_ _0988_ _1059_ _1062_ vssd1 vssd1 vccd1 vccd1 _1063_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_0_133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2169_ _0904_ _0907_ _0910_ CB_1.config_dataA\[14\] vssd1 vssd1 vccd1 vccd1 _0927_
+ sky130_fd_sc_hd__or4b_1
XANTENNA__2359__B1 _0831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input15_A CBnorth_in[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2925__SET_B net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1540_ CB_1.config_dataA\[17\] CB_1.config_dataA\[16\] net142 CB_1.config_dataA\[18\]
+ vssd1 vssd1 vccd1 vccd1 _1334_ sky130_fd_sc_hd__or4b_1
X_1471_ SB0.route_sel\[58\] SB0.route_sel\[59\] _1260_ _1263_ _1264_ vssd1 vssd1 vccd1
+ vccd1 _1265_ sky130_fd_sc_hd__a221oi_1
XANTENNA__2117__A3 _0781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3072_ clknet_leaf_9_clk _0280_ net220 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[12\]
+ sky130_fd_sc_hd__dfstp_1
X_2023_ _0779_ _0780_ _1270_ vssd1 vssd1 vccd1 vccd1 _0781_ sky130_fd_sc_hd__a21boi_4
X_1807_ _1297_ _0545_ _0546_ _1273_ vssd1 vssd1 vccd1 vccd1 _0569_ sky130_fd_sc_hd__o22a_1
X_2856_ clknet_leaf_5_clk _0064_ net203 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__1800__A2 net25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2925_ clknet_leaf_18_clk _0133_ net217 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[17\]
+ sky130_fd_sc_hd__dfstp_1
X_1669_ CB_0.config_dataA\[19\] CB_0.config_dataA\[18\] _1274_ vssd1 vssd1 vccd1 vccd1
+ _0431_ sky130_fd_sc_hd__or3b_1
XPHY_EDGE_ROW_37_Left_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2787_ net366 net318 net230 vssd1 vssd1 vccd1 vccd1 _0323_ sky130_fd_sc_hd__mux2_1
X_1738_ net131 _1257_ _0457_ _0460_ _1261_ vssd1 vssd1 vccd1 vccd1 _0500_ sky130_fd_sc_hd__o32a_1
XANTENNA__1867__A2 net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input7_A CBeast_in[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_46_Left_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input18_X net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2283__A2 _0816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2710_ SB0.route_sel\[110\] SB0.route_sel\[109\] net266 vssd1 vssd1 vccd1 vccd1 _0246_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__2035__A2 _0781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1454_ net125 vssd1 vssd1 vccd1 vccd1 _1248_ sky130_fd_sc_hd__inv_2
X_2572_ net323 net289 net259 vssd1 vssd1 vccd1 vccd1 _0108_ sky130_fd_sc_hd__mux2_1
X_2641_ SB0.route_sel\[41\] SB0.route_sel\[40\] net256 vssd1 vssd1 vccd1 vccd1 _0177_
+ sky130_fd_sc_hd__mux2_1
X_1523_ _1315_ _1316_ _1303_ vssd1 vssd1 vccd1 vccd1 _1317_ sky130_fd_sc_hd__o21ba_1
X_3055_ clknet_leaf_11_clk _0263_ net221 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[15\]
+ sky130_fd_sc_hd__dfstp_2
X_1385_ SB0.route_sel\[32\] vssd1 vssd1 vccd1 vccd1 _1179_ sky130_fd_sc_hd__inv_2
X_2006_ LE_0B.config_data\[14\] _0700_ _0702_ vssd1 vssd1 vccd1 vccd1 _0766_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_33_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1785__A1 _0391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2839_ clknet_leaf_13_clk net370 net225 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[46\]
+ sky130_fd_sc_hd__dfrtp_1
X_2908_ clknet_leaf_17_clk _0116_ net213 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[0\]
+ sky130_fd_sc_hd__dfstp_2
XTAP_TAPCELL_ROW_56_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1730__X _0492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_29_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_30_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2624_ SB0.route_sel\[24\] SB0.route_sel\[23\] net238 vssd1 vssd1 vccd1 vccd1 _0160_
+ sky130_fd_sc_hd__mux2_1
X_1506_ net158 net160 vssd1 vssd1 vccd1 vccd1 _1300_ sky130_fd_sc_hd__and2b_1
X_1437_ LEI0.config_data\[41\] vssd1 vssd1 vccd1 vccd1 _1231_ sky130_fd_sc_hd__inv_2
Xoutput113 net113 vssd1 vssd1 vccd1 vccd1 SBwest_out[4] sky130_fd_sc_hd__buf_2
X_2486_ LEI0.config_data\[24\] net285 net244 vssd1 vssd1 vccd1 vccd1 _0025_ sky130_fd_sc_hd__mux2_1
X_2555_ LE_0B.reset_mode net405 net230 vssd1 vssd1 vccd1 vccd1 _0092_ sky130_fd_sc_hd__mux2_1
Xoutput102 net102 vssd1 vssd1 vccd1 vccd1 SBsouth_out[7] sky130_fd_sc_hd__buf_2
XFILLER_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3038_ clknet_leaf_14_clk _0246_ net222 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[110\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1368_ SB0.route_sel\[12\] vssd1 vssd1 vccd1 vccd1 _1162_ sky130_fd_sc_hd__inv_2
X_3107_ clknet_leaf_1_clk _0315_ net191 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2183__A1 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_44_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1550__X _1344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput26 CBnorth_in[7] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__buf_2
Xinput15 CBnorth_in[0] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__buf_2
Xinput48 SBwest_in[1] vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__clkbuf_1
Xinput37 SBsouth_in[4] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__buf_1
Xinput59 le_clk vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__clkbuf_2
X_2340_ _1325_ _1076_ _1327_ vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__a21o_1
X_2271_ net179 _1026_ vssd1 vssd1 vccd1 vccd1 _1027_ sky130_fd_sc_hd__nor2_1
XANTENNA__2174__A1 LE_1A.config_data\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2229__A2 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1986_ net121 _0430_ _0391_ _0447_ _1232_ CB_0.config_dataB\[13\] vssd1 vssd1 vccd1
+ vccd1 _0746_ sky130_fd_sc_hd__mux4_1
XANTENNA__1635__X _0397_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_9_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2607_ SB0.route_sel\[7\] SB0.route_sel\[6\] net231 vssd1 vssd1 vccd1 vccd1 _0143_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_58_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2469_ net389 LEI0.config_data\[6\] net266 vssd1 vssd1 vccd1 vccd1 _0008_ sky130_fd_sc_hd__mux2_1
X_2538_ net316 LE_0B.config_data\[1\] net245 vssd1 vssd1 vccd1 vccd1 _0075_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout272_X net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1979__A1 net24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1903__B2 _0512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input45_A SBwest_in[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout170 CB_0.config_dataA\[8\] vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__buf_2
Xfanout181 CB_1.config_dataB\[12\] vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout192 net193 vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__clkbuf_4
XFILLER_19_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1840_ CB_0.config_dataA\[10\] _0587_ _0600_ _0601_ _0575_ vssd1 vssd1 vccd1 vccd1
+ _0602_ sky130_fd_sc_hd__a311o_1
X_1771_ _0527_ _0531_ _0532_ _0523_ vssd1 vssd1 vccd1 vccd1 _0533_ sky130_fd_sc_hd__a31o_1
XFILLER_6_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2323_ _0359_ net125 _0342_ vssd1 vssd1 vccd1 vccd1 _1068_ sky130_fd_sc_hd__mux2_1
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2254_ net13 net14 net182 vssd1 vssd1 vccd1 vccd1 _1010_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_63_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2185_ net4 net5 CB_1.config_dataB\[0\] vssd1 vssd1 vccd1 vccd1 _0941_ sky130_fd_sc_hd__mux2_1
XANTENNA__1830__A0 net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1969_ _0728_ vssd1 vssd1 vccd1 vccd1 _0729_ sky130_fd_sc_hd__inv_2
XANTENNA__2083__A0 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1821__A0 _0473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1888__A0 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4 LE_1B.config_data\[12\] vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__dlygate4sd3_1
X_1823_ CB_0.config_dataA\[9\] _0583_ _0584_ vssd1 vssd1 vccd1 vccd1 _0585_ sky130_fd_sc_hd__o21a_1
X_2872_ clknet_leaf_4_clk _0080_ net199 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__1812__A0 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2065__A0 _0816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2941_ clknet_leaf_28_clk _0149_ net188 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[13\]
+ sky130_fd_sc_hd__dfstp_1
X_1754_ CB_0.config_dataA\[1\] _1214_ _0515_ vssd1 vssd1 vccd1 vccd1 _0516_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_29_Left_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1685_ _0444_ _0446_ vssd1 vssd1 vccd1 vccd1 _0447_ sky130_fd_sc_hd__nand2_4
XFILLER_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2237_ net182 _0797_ _0991_ _0992_ vssd1 vssd1 vccd1 vccd1 _0993_ sky130_fd_sc_hd__a211o_1
X_2306_ _0987_ _1060_ _1061_ _1017_ vssd1 vssd1 vccd1 vccd1 _1062_ sky130_fd_sc_hd__o31a_1
XPHY_EDGE_ROW_13_Left_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2099_ net13 net14 net151 vssd1 vssd1 vccd1 vccd1 _0857_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2168_ _0911_ net146 CB_1.config_dataA\[14\] vssd1 vssd1 vccd1 vccd1 _0926_ sky130_fd_sc_hd__or3b_1
XPHY_EDGE_ROW_17_Right_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Right_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_35_Right_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2047__A0 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1470_ _1249_ _1261_ _1262_ vssd1 vssd1 vccd1 vccd1 _1264_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_22_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_44_Right_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3071_ clknet_leaf_9_clk _0279_ net219 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[11\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_53_Right_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2286__A0 net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2022_ SB0.route_sel\[60\] SB0.route_sel\[61\] _1190_ SB0.route_sel\[56\] vssd1 vssd1
+ vccd1 vccd1 _0780_ sky130_fd_sc_hd__o22a_1
X_1806_ _1345_ _1321_ net172 vssd1 vssd1 vccd1 vccd1 _0568_ sky130_fd_sc_hd__mux2_1
X_2855_ clknet_leaf_5_clk net315 net203 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__1800__A3 net26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2924_ clknet_leaf_18_clk _0132_ net217 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[16\]
+ sky130_fd_sc_hd__dfstp_1
X_2786_ net318 net282 net234 vssd1 vssd1 vccd1 vccd1 _0322_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_62_Right_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1599_ net23 net24 net25 net26 net174 CB_0.config_dataA\[1\] vssd1 vssd1 vccd1 vccd1
+ _0361_ sky130_fd_sc_hd__mux4_1
X_1737_ net177 net178 _0456_ net3 vssd1 vssd1 vccd1 vccd1 _0499_ sky130_fd_sc_hd__a31o_1
X_1668_ _0427_ _0429_ vssd1 vssd1 vccd1 vccd1 _0430_ sky130_fd_sc_hd__nand2_4
XANTENNA__1867__A3 net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_10_clk_A clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_25_clk_A clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output114_A net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2283__A3 _0813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2268__B1 _1017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2640_ SB0.route_sel\[40\] SB0.route_sel\[39\] net255 vssd1 vssd1 vccd1 vccd1 _0176_
+ sky130_fd_sc_hd__mux2_1
X_1453_ net60 vssd1 vssd1 vccd1 vccd1 _1247_ sky130_fd_sc_hd__inv_2
X_2571_ net289 LE_1A.config_data\[11\] net259 vssd1 vssd1 vccd1 vccd1 _0107_ sky130_fd_sc_hd__mux2_1
X_1522_ SB0.route_sel\[44\] SB0.route_sel\[45\] net52 _1314_ _1311_ vssd1 vssd1 vccd1
+ vccd1 _1316_ sky130_fd_sc_hd__a41o_1
X_3054_ clknet_leaf_8_clk _0262_ net210 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[14\]
+ sky130_fd_sc_hd__dfstp_1
X_2005_ LE_0B.config_data\[12\] LE_0B.config_data\[13\] _0703_ vssd1 vssd1 vccd1 vccd1
+ _0765_ sky130_fd_sc_hd__mux2_1
X_1384_ SB0.route_sel\[38\] vssd1 vssd1 vccd1 vccd1 _1178_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_33_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2907_ LE_1B.sel_clk _0115_ net61 vssd1 vssd1 vccd1 vccd1 LE_1B.dff0_out sky130_fd_sc_hd__dfrtp_1
X_2838_ clknet_leaf_13_clk _0046_ net225 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[45\]
+ sky130_fd_sc_hd__dfrtp_1
X_2769_ net144 net145 net255 vssd1 vssd1 vccd1 vccd1 _0305_ sky130_fd_sc_hd__mux2_1
XFILLER_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_16_Left_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1548__X _1342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2379__X net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input30_X net30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput114 net114 vssd1 vssd1 vccd1 vccd1 SBwest_out[5] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_30_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2554_ net405 LE_0B.edge_mode net230 vssd1 vssd1 vccd1 vccd1 _0091_ sky130_fd_sc_hd__mux2_1
Xoutput103 net103 vssd1 vssd1 vccd1 vccd1 SBsouth_out[8] sky130_fd_sc_hd__buf_2
X_2623_ SB0.route_sel\[23\] SB0.route_sel\[22\] net238 vssd1 vssd1 vccd1 vccd1 _0159_
+ sky130_fd_sc_hd__mux2_1
X_1505_ _1251_ _1298_ vssd1 vssd1 vccd1 vccd1 _1299_ sky130_fd_sc_hd__nand2_1
X_1436_ CB_0.config_dataB\[11\] vssd1 vssd1 vccd1 vccd1 _1230_ sky130_fd_sc_hd__inv_2
X_2485_ net285 net292 net235 vssd1 vssd1 vccd1 vccd1 _0024_ sky130_fd_sc_hd__mux2_1
X_1367_ SB0.route_sel\[11\] vssd1 vssd1 vccd1 vccd1 _1161_ sky130_fd_sc_hd__inv_2
X_3037_ clknet_leaf_14_clk _0245_ net224 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[109\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_fanout262_A net58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3106_ clknet_leaf_1_clk net345 net191 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2183__A2 net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_1_Left_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput16 CBnorth_in[10] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__buf_2
Xinput27 CBnorth_in[8] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__buf_2
Xinput38 SBsouth_in[5] vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput49 SBwest_in[2] vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__buf_1
X_2270_ _0792_ _0784_ net180 vssd1 vssd1 vccd1 vccd1 _1026_ sky130_fd_sc_hd__mux2_1
XANTENNA__2229__A3 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1985_ net139 net125 net129 net133 LEI0.config_data\[39\] LEI0.config_data\[40\]
+ vssd1 vssd1 vccd1 vccd1 _0745_ sky130_fd_sc_hd__mux4_1
X_2537_ net401 LE_0B.config_data\[0\] net242 vssd1 vssd1 vccd1 vccd1 _0074_ sky130_fd_sc_hd__mux2_1
X_2606_ SB0.route_sel\[6\] SB0.route_sel\[5\] net238 vssd1 vssd1 vccd1 vccd1 _0142_
+ sky130_fd_sc_hd__mux2_1
X_2468_ LEI0.config_data\[6\] net296 net244 vssd1 vssd1 vccd1 vccd1 _0007_ sky130_fd_sc_hd__mux2_1
X_1419_ SB0.route_sel\[104\] vssd1 vssd1 vccd1 vccd1 _1213_ sky130_fd_sc_hd__inv_2
X_2399_ SB0.route_sel\[51\] _1185_ _1187_ SB0.route_sel\[48\] _1109_ vssd1 vssd1 vccd1
+ vccd1 _1110_ sky130_fd_sc_hd__a221o_1
XANTENNA__1979__A2 net25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input38_A SBsouth_in[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout171 CB_0.config_dataA\[5\] vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__buf_2
Xfanout160 CB_0.config_dataB\[16\] vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__buf_1
XFILLER_47_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout182 CB_1.config_dataB\[8\] vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__buf_2
Xfanout193 net229 vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_6_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1770_ SB0.route_sel\[84\] SB0.route_sel\[85\] net30 vssd1 vssd1 vccd1 vccd1 _0532_
+ sky130_fd_sc_hd__a21bo_1
X_2322_ _0330_ _0331_ _1067_ _0333_ vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__a31o_1
X_2253_ net2 net3 net182 vssd1 vssd1 vccd1 vccd1 _1009_ sky130_fd_sc_hd__mux2_1
X_2184_ CB_1.config_dataB\[3\] _0939_ vssd1 vssd1 vccd1 vccd1 _0940_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_63_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2083__A1 net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1830__A1 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1899_ CB_0.config_dataB\[5\] _1229_ _0658_ vssd1 vssd1 vccd1 vccd1 _0659_ sky130_fd_sc_hd__or3_1
X_1968_ net136 net122 net130 net134 LEI0.config_data\[27\] LEI0.config_data\[28\]
+ vssd1 vssd1 vccd1 vccd1 _0728_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_3_154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1821__A1 _0492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2074__A1 _0831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1888__A1 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold5 _0320_ vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2065__A1 _0819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2940_ clknet_leaf_28_clk _0148_ net188 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[12\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_17_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1822_ _0538_ _0578_ _0579_ _0512_ CB_0.config_dataA\[11\] vssd1 vssd1 vccd1 vccd1
+ _0584_ sky130_fd_sc_hd__o221a_1
XANTENNA__1576__B1 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1753_ net27 net28 net174 vssd1 vssd1 vccd1 vccd1 _0515_ sky130_fd_sc_hd__mux2_1
XANTENNA__1812__A1 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2871_ clknet_leaf_4_clk net312 net199 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1684_ SB0.route_sel\[20\] _1167_ SB0.route_sel\[23\] _1169_ _0445_ vssd1 vssd1 vccd1
+ vccd1 _0446_ sky130_fd_sc_hd__a221o_1
XFILLER_38_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2236_ _0356_ _0802_ net182 vssd1 vssd1 vccd1 vccd1 _0992_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_0_135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout175_A CB_1.config_dataB\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1500__B1 _1279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2167_ CB_1.config_dataA\[14\] _0914_ _0916_ _0924_ vssd1 vssd1 vccd1 vccd1 _0925_
+ sky130_fd_sc_hd__or4_1
X_2305_ LE_1B.config_data\[8\] net120 net135 vssd1 vssd1 vccd1 vccd1 _1061_ sky130_fd_sc_hd__and3_1
X_2098_ net1 net6 net7 net8 net151 CB_1.config_dataA\[1\] vssd1 vssd1 vccd1 vccd1
+ _0856_ sky130_fd_sc_hd__mux4_1
XFILLER_21_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout228_X net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout130_X net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2047__A1 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_30_Left_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input60_X net60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2286__A1 net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3070_ clknet_leaf_9_clk _0278_ net209 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[10\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_35_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2021_ SB0.route_sel\[63\] SB0.route_sel\[62\] vssd1 vssd1 vccd1 vccd1 _0779_ sky130_fd_sc_hd__nand2b_1
XANTENNA_output69_A net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2923_ clknet_leaf_14_clk _0131_ net223 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[15\]
+ sky130_fd_sc_hd__dfstp_2
X_1805_ _0564_ _0566_ _0545_ vssd1 vssd1 vccd1 vccd1 _0567_ sky130_fd_sc_hd__o21a_1
X_1736_ net137 _0496_ _0494_ vssd1 vssd1 vccd1 vccd1 _0498_ sky130_fd_sc_hd__mux2_1
X_2854_ clknet_leaf_6_clk net342 net203 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2210__A1 _0831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2785_ net282 net276 net234 vssd1 vssd1 vccd1 vccd1 _0321_ sky130_fd_sc_hd__mux2_1
X_1598_ net174 _0359_ CB_0.config_dataA\[3\] _1154_ vssd1 vssd1 vccd1 vccd1 _0360_
+ sky130_fd_sc_hd__o211a_1
X_1667_ SB0.route_sel\[4\] _1156_ SB0.route_sel\[7\] _1158_ _0428_ vssd1 vssd1 vccd1
+ vccd1 _0429_ sky130_fd_sc_hd__a221o_1
X_2219_ net183 _0974_ _0973_ vssd1 vssd1 vccd1 vccd1 _0975_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_28_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1960__A0 net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input20_A CBnorth_in[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2570_ net333 LE_1A.config_data\[10\] net259 vssd1 vssd1 vccd1 vccd1 _0106_ sky130_fd_sc_hd__mux2_1
XANTENNA__1951__A0 net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2288__A net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1521_ _1180_ _1181_ net38 vssd1 vssd1 vccd1 vccd1 _1315_ sky130_fd_sc_hd__o21a_1
X_1452_ LE_1B.config_data\[16\] vssd1 vssd1 vccd1 vccd1 _1246_ sky130_fd_sc_hd__inv_2
X_1383_ SB0.route_sel\[39\] vssd1 vssd1 vccd1 vccd1 _1177_ sky130_fd_sc_hd__inv_2
X_3053_ clknet_leaf_8_clk _0261_ net210 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[13\]
+ sky130_fd_sc_hd__dfstp_1
X_2004_ _0730_ _0761_ _0763_ _0759_ vssd1 vssd1 vccd1 vccd1 _0764_ sky130_fd_sc_hd__a31o_1
XFILLER_35_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2906_ clknet_leaf_29_clk _0114_ net186 vssd1 vssd1 vccd1 vccd1 LE_1A.reset_mode
+ sky130_fd_sc_hd__dfrtp_1
X_2837_ clknet_leaf_13_clk _0045_ net225 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[44\]
+ sky130_fd_sc_hd__dfrtp_1
X_2699_ SB0.route_sel\[99\] SB0.route_sel\[98\] net263 vssd1 vssd1 vccd1 vccd1 _0235_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__2195__A0 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1719_ _1305_ _0456_ net14 vssd1 vssd1 vccd1 vccd1 _0481_ sky130_fd_sc_hd__a21o_1
X_2768_ net145 CB_1.config_dataA\[15\] net262 vssd1 vssd1 vccd1 vccd1 _0304_ sky130_fd_sc_hd__mux2_1
XANTENNA__2498__A1 LEI0.config_data\[35\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1933__B1 CB_0.config_dataB\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2110__A0 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input23_X net23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_30_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1504_ CB_0.config_dataA\[17\] CB_0.config_dataA\[16\] vssd1 vssd1 vccd1 vccd1 _1298_
+ sky130_fd_sc_hd__and2b_1
Xoutput115 net115 vssd1 vssd1 vccd1 vccd1 SBwest_out[6] sky130_fd_sc_hd__buf_2
Xoutput104 net104 vssd1 vssd1 vccd1 vccd1 SBsouth_out[9] sky130_fd_sc_hd__buf_2
X_2553_ LE_0B.edge_mode LE_0B.config_data\[16\] net230 vssd1 vssd1 vccd1 vccd1 _0090_
+ sky130_fd_sc_hd__mux2_1
X_2622_ SB0.route_sel\[22\] SB0.route_sel\[21\] net232 vssd1 vssd1 vccd1 vccd1 _0158_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__2510__S net60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1435_ CB_0.config_dataB\[7\] vssd1 vssd1 vccd1 vccd1 _1229_ sky130_fd_sc_hd__inv_2
X_2484_ net292 net367 net235 vssd1 vssd1 vccd1 vccd1 _0023_ sky130_fd_sc_hd__mux2_1
X_3105_ clknet_leaf_1_clk net326 net191 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_1366_ SB0.route_sel\[0\] vssd1 vssd1 vccd1 vccd1 _1160_ sky130_fd_sc_hd__inv_2
X_3036_ clknet_leaf_14_clk _0244_ net224 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[108\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__2101__A0 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout210_X net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_24_clk_A clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2183__A3 net12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput28 CBnorth_in[9] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__buf_2
Xinput17 CBnorth_in[11] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__buf_2
Xinput39 SBsouth_in[6] vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__clkbuf_1
XANTENNA__2159__A0 net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1984_ _0738_ _0742_ _0743_ net162 CB_0.config_dataB\[14\] vssd1 vssd1 vccd1 vccd1
+ _0744_ sky130_fd_sc_hd__o221a_1
X_2467_ net296 LEI0.config_data\[4\] net248 vssd1 vssd1 vccd1 vccd1 _0006_ sky130_fd_sc_hd__mux2_1
X_2605_ SB0.route_sel\[5\] SB0.route_sel\[4\] net238 vssd1 vssd1 vccd1 vccd1 _0141_
+ sky130_fd_sc_hd__mux2_1
X_2536_ net416 LE_1B.reset_mode net234 vssd1 vssd1 vccd1 vccd1 _0073_ sky130_fd_sc_hd__mux2_1
X_1418_ SB0.route_sel\[110\] vssd1 vssd1 vccd1 vccd1 _1212_ sky130_fd_sc_hd__inv_2
X_2398_ SB0.route_sel\[55\] SB0.route_sel\[54\] vssd1 vssd1 vccd1 vccd1 _1109_ sky130_fd_sc_hd__nor2_1
XANTENNA__1979__A3 net26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3019_ clknet_leaf_25_clk _0227_ net213 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[91\]
+ sky130_fd_sc_hd__dfstp_1
Xfanout172 net173 vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__buf_2
Xfanout161 CB_0.config_dataB\[12\] vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__buf_2
Xfanout183 CB_1.config_dataB\[7\] vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__clkbuf_2
Xfanout150 CB_1.config_dataA\[4\] vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout194 net198 vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__clkbuf_4
XFILLER_19_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2321_ net154 net156 _1300_ _0336_ _0338_ vssd1 vssd1 vccd1 vccd1 _1067_ sky130_fd_sc_hd__a32o_1
X_2252_ net1 net6 net7 net8 net182 CB_1.config_dataB\[9\] vssd1 vssd1 vccd1 vccd1
+ _1008_ sky130_fd_sc_hd__mux4_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2183_ net9 net10 net11 net12 CB_1.config_dataB\[0\] CB_1.config_dataB\[1\] vssd1
+ vssd1 vccd1 vccd1 _0939_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_63_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1898_ net27 net28 net165 vssd1 vssd1 vccd1 vccd1 _0658_ sky130_fd_sc_hd__mux2_1
X_1967_ CB_0.config_dataB\[10\] _0717_ _0719_ _0726_ vssd1 vssd1 vccd1 vccd1 _0727_
+ sky130_fd_sc_hd__or4_1
XANTENNA_fanout218_A net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout120_A _0957_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2519_ net376 LE_0A.config_data\[5\] net247 vssd1 vssd1 vccd1 vccd1 _0057_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_3_155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input50_A SBwest_in[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1888__A2 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold6 LE_1A.config_data\[4\] vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_60_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1812__A2 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2870_ clknet_leaf_4_clk net358 net199 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2065__A2 _0813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1821_ _0473_ _0492_ CB_0.config_dataA\[8\] vssd1 vssd1 vccd1 vccd1 _0583_ sky130_fd_sc_hd__mux2_1
X_1752_ net15 net20 net21 net22 net174 CB_0.config_dataA\[1\] vssd1 vssd1 vccd1 vccd1
+ _0514_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_10_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1683_ SB0.route_sel\[19\] SB0.route_sel\[18\] vssd1 vssd1 vccd1 vccd1 _0445_ sky130_fd_sc_hd__nor2_1
X_2304_ net120 net135 LE_1B.config_data\[9\] vssd1 vssd1 vccd1 vccd1 _1060_ sky130_fd_sc_hd__a21boi_1
X_2235_ CB_1.config_dataB\[9\] CB_1.config_dataB\[11\] vssd1 vssd1 vccd1 vccd1 _0991_
+ sky130_fd_sc_hd__nand2b_1
X_2097_ CB_1.config_dataA\[1\] CB_1.config_dataA\[3\] vssd1 vssd1 vccd1 vccd1 _0855_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_0_136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2166_ CB_1.config_dataA\[13\] CB_1.config_dataA\[15\] _0923_ _0922_ vssd1 vssd1
+ vccd1 vccd1 _0924_ sky130_fd_sc_hd__a31o_1
XANTENNA__1803__A2 _0339_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_3_Right_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2999_ clknet_leaf_25_clk _0207_ net196 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[71\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_39_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2047__A2 net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input53_X net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2020_ net150 _0777_ vssd1 vssd1 vccd1 vccd1 _0778_ sky130_fd_sc_hd__nor2_1
XFILLER_62_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2853_ clknet_leaf_6_clk _0061_ net203 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_2922_ clknet_leaf_14_clk _0130_ net223 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[14\]
+ sky130_fd_sc_hd__dfstp_1
X_1804_ net172 _0359_ _0565_ vssd1 vssd1 vccd1 vccd1 _0566_ sky130_fd_sc_hd__o21a_1
X_1735_ SB0.route_sel\[88\] SB0.route_sel\[89\] vssd1 vssd1 vccd1 vccd1 _0497_ sky130_fd_sc_hd__nand2_1
X_1666_ SB0.route_sel\[3\] SB0.route_sel\[2\] vssd1 vssd1 vccd1 vccd1 _0428_ sky130_fd_sc_hd__nor2_1
X_2784_ net276 LE_1B.config_data\[11\] net234 vssd1 vssd1 vccd1 vccd1 _0320_ sky130_fd_sc_hd__mux2_1
X_1597_ _0356_ _0358_ vssd1 vssd1 vccd1 vccd1 _0359_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_36_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2218_ net9 net10 net11 net12 net185 net184 vssd1 vssd1 vccd1 vccd1 _0974_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_28_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2149_ net146 _0803_ _0906_ vssd1 vssd1 vccd1 vccd1 _0907_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_11_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1960__A1 net20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input13_A CBeast_in[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1476__B1 _1256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1951__A1 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1520_ SB0.route_sel\[47\] SB0.route_sel\[46\] vssd1 vssd1 vccd1 vccd1 _1314_ sky130_fd_sc_hd__nand2_1
X_1451_ net182 vssd1 vssd1 vccd1 vccd1 _1245_ sky130_fd_sc_hd__inv_2
X_1382_ SB0.route_sel\[37\] vssd1 vssd1 vccd1 vccd1 _1176_ sky130_fd_sc_hd__inv_2
X_3052_ clknet_leaf_8_clk _0260_ net210 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[12\]
+ sky130_fd_sc_hd__dfstp_1
X_2003_ LE_0B.config_data\[1\] _0703_ _0762_ _0675_ vssd1 vssd1 vccd1 vccd1 _0763_
+ sky130_fd_sc_hd__a211o_1
X_2836_ clknet_leaf_13_clk _0044_ net226 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[43\]
+ sky130_fd_sc_hd__dfrtp_1
X_2905_ clknet_leaf_29_clk _0113_ net186 vssd1 vssd1 vccd1 vccd1 LE_1A.reset_val sky130_fd_sc_hd__dfrtp_1
X_1718_ _0479_ net138 _0477_ vssd1 vssd1 vccd1 vccd1 _0480_ sky130_fd_sc_hd__mux2_1
X_2698_ SB0.route_sel\[98\] SB0.route_sel\[97\] net263 vssd1 vssd1 vccd1 vccd1 _0234_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__2195__A1 net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1649_ _0408_ _0409_ _0410_ _0407_ vssd1 vssd1 vccd1 vccd1 _0411_ sky130_fd_sc_hd__o31ai_2
X_2767_ CB_1.config_dataA\[15\] CB_1.config_dataA\[14\] net260 vssd1 vssd1 vccd1 vccd1
+ _0303_ sky130_fd_sc_hd__mux2_1
XANTENNA_input5_A CBeast_in[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1933__A1 _1318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2110__A1 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input16_X net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3086__SET_B net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput116 net116 vssd1 vssd1 vccd1 vccd1 SBwest_out[7] sky130_fd_sc_hd__buf_2
XANTENNA__1924__A1 _0430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput105 net105 vssd1 vssd1 vccd1 vccd1 SBwest_out[0] sky130_fd_sc_hd__buf_2
X_2552_ LE_0B.config_data\[16\] net275 net242 vssd1 vssd1 vccd1 vccd1 _0089_ sky130_fd_sc_hd__mux2_1
X_2483_ net367 net396 net235 vssd1 vssd1 vccd1 vccd1 _0022_ sky130_fd_sc_hd__mux2_1
X_2621_ SB0.route_sel\[21\] SB0.route_sel\[20\] net232 vssd1 vssd1 vccd1 vccd1 _0157_
+ sky130_fd_sc_hd__mux2_1
X_1503_ _1295_ _1296_ _1294_ vssd1 vssd1 vccd1 vccd1 _1297_ sky130_fd_sc_hd__a21boi_4
X_3035_ clknet_leaf_14_clk _0243_ net224 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[107\]
+ sky130_fd_sc_hd__dfstp_1
X_1434_ net165 vssd1 vssd1 vccd1 vccd1 _1228_ sky130_fd_sc_hd__inv_2
X_3104_ clknet_leaf_0_clk _0312_ net192 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_1365_ net29 vssd1 vssd1 vccd1 vccd1 _1159_ sky130_fd_sc_hd__inv_2
XANTENNA__2101__A1 net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout248_A net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1649__Y _0411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2819_ clknet_leaf_3_clk net337 net201 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input8_X net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput18 CBnorth_in[12] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_52_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput29 SBsouth_in[0] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_1
XANTENNA__2159__A1 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2331__A1 _0473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1983_ CB_0.config_dataB\[13\] CB_0.config_dataB\[15\] vssd1 vssd1 vccd1 vccd1 _0743_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__1485__X _1279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2604_ SB0.route_sel\[4\] SB0.route_sel\[3\] net238 vssd1 vssd1 vccd1 vccd1 _0140_
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2466_ net379 net329 net246 vssd1 vssd1 vccd1 vccd1 _0005_ sky130_fd_sc_hd__mux2_1
X_1417_ SB0.route_sel\[109\] vssd1 vssd1 vccd1 vccd1 _1211_ sky130_fd_sc_hd__inv_2
X_2535_ LE_1A.dff1_out _1247_ _1152_ vssd1 vssd1 vccd1 vccd1 _0072_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout198_A net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3018_ clknet_leaf_2_clk _0226_ net198 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[90\]
+ sky130_fd_sc_hd__dfstp_1
X_2397_ _1294_ _1108_ vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__and2_2
Xfanout140 net141 vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout173 CB_0.config_dataA\[4\] vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__clkbuf_2
Xfanout162 CB_0.config_dataB\[12\] vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout184 CB_1.config_dataB\[5\] vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__buf_2
Xfanout151 net152 vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout195 net198 vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__clkbuf_4
XFILLER_63_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1824__A0 net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2251_ CB_1.config_dataB\[11\] _1006_ vssd1 vssd1 vccd1 vccd1 _1007_ sky130_fd_sc_hd__nor2_1
X_2320_ net59 LE_1B.edge_mode vssd1 vssd1 vccd1 vccd1 LE_1B.sel_clk sky130_fd_sc_hd__xnor2_1
X_2182_ _0356_ _0802_ CB_1.config_dataB\[0\] vssd1 vssd1 vccd1 vccd1 _0938_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_23_clk_A clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1966_ CB_0.config_dataB\[9\] CB_0.config_dataB\[11\] _0725_ _0724_ vssd1 vssd1 vccd1
+ vccd1 _0726_ sky130_fd_sc_hd__a31o_1
X_1897_ _1228_ _0654_ vssd1 vssd1 vccd1 vccd1 _0657_ sky130_fd_sc_hd__nor2_1
X_2518_ net413 net359 net247 vssd1 vssd1 vccd1 vccd1 _0056_ sky130_fd_sc_hd__mux2_1
X_2449_ SB0.route_sel\[88\] SB0.route_sel\[89\] vssd1 vssd1 vccd1 vccd1 _1143_ sky130_fd_sc_hd__nor2_1
XANTENNA__1806__A0 _1345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1888__A3 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input43_A SBwest_in[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold7 _0099_ vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_60_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1820_ _0447_ _0577_ _0581_ vssd1 vssd1 vccd1 vccd1 _0582_ sky130_fd_sc_hd__a21oi_1
XANTENNA__1812__A3 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2065__A3 _0822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1751_ _0509_ _0510_ _0511_ _0508_ vssd1 vssd1 vccd1 vccd1 _0513_ sky130_fd_sc_hd__o31ai_2
X_1682_ _0434_ _0435_ _0440_ _0443_ vssd1 vssd1 vccd1 vccd1 _0444_ sky130_fd_sc_hd__a22o_2
X_2234_ LE_1B.config_data\[7\] _0961_ _0989_ vssd1 vssd1 vccd1 vccd1 _0990_ sky130_fd_sc_hd__a21oi_1
X_2303_ LE_1B.config_data\[10\] LE_1B.config_data\[11\] _0961_ vssd1 vssd1 vccd1 vccd1
+ _1059_ sky130_fd_sc_hd__mux2_1
X_2096_ net151 _0828_ _0852_ _0853_ vssd1 vssd1 vccd1 vccd1 _0854_ sky130_fd_sc_hd__a211o_1
X_2165_ _0838_ _0835_ net147 vssd1 vssd1 vccd1 vccd1 _0923_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1949_ net164 _0339_ _0707_ _0708_ vssd1 vssd1 vccd1 vccd1 _0709_ sky130_fd_sc_hd__a211o_1
XANTENNA__2213__A0 net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2998_ clknet_leaf_1_clk _0206_ net196 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[70\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__1673__X _0435_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2047__A3 net12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input46_X net46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_13_Right_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1803_ net172 _0339_ CB_0.config_dataA\[5\] vssd1 vssd1 vccd1 vccd1 _0565_ sky130_fd_sc_hd__a21oi_1
X_2852_ clknet_leaf_6_clk _0060_ net204 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_2921_ clknet_leaf_14_clk _0129_ net222 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[13\]
+ sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_22_Right_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2783_ net338 LE_1B.config_data\[10\] net234 vssd1 vssd1 vccd1 vccd1 _0319_ sky130_fd_sc_hd__mux2_1
X_1734_ net17 net123 _0495_ vssd1 vssd1 vccd1 vccd1 _0496_ sky130_fd_sc_hd__mux2_1
X_1596_ SB0.route_sel\[100\] _1207_ SB0.route_sel\[103\] _1209_ _0357_ vssd1 vssd1
+ vccd1 vccd1 _0358_ sky130_fd_sc_hd__a221o_1
XANTENNA__2210__A3 _0838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1665_ _0413_ _0418_ _0422_ _0426_ vssd1 vssd1 vccd1 vccd1 _0427_ sky130_fd_sc_hd__a22o_2
X_2217_ _0972_ net184 net183 vssd1 vssd1 vccd1 vccd1 _0973_ sky130_fd_sc_hd__or3b_1
XPHY_EDGE_ROW_31_Right_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2079_ SB0.route_sel\[84\] SB0.route_sel\[85\] _1202_ SB0.route_sel\[80\] vssd1 vssd1
+ vccd1 vccd1 _0837_ sky130_fd_sc_hd__o22a_1
X_2148_ net146 _0797_ _0905_ vssd1 vssd1 vccd1 vccd1 _0906_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_40_Right_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1960__A2 net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1450_ net185 vssd1 vssd1 vccd1 vccd1 _1244_ sky130_fd_sc_hd__inv_2
X_3051_ clknet_leaf_7_clk _0259_ net206 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[11\]
+ sky130_fd_sc_hd__dfstp_2
XANTENNA__2259__A3 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1381_ SB0.route_sel\[24\] vssd1 vssd1 vccd1 vccd1 _1175_ sky130_fd_sc_hd__inv_2
X_2002_ LE_0B.config_data\[0\] _0700_ _0702_ vssd1 vssd1 vccd1 vccd1 _0762_ sky130_fd_sc_hd__and3_1
XFILLER_35_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2835_ clknet_leaf_13_clk _0043_ net226 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[42\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_0_clk_X clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2904_ clknet_leaf_29_clk _0112_ net186 vssd1 vssd1 vccd1 vccd1 LE_1A.edge_mode sky130_fd_sc_hd__dfstp_1
X_2766_ CB_1.config_dataA\[14\] CB_1.config_dataA\[13\] net260 vssd1 vssd1 vccd1 vccd1
+ _0302_ sky130_fd_sc_hd__mux2_1
X_1579_ CB_0.config_dataA\[17\] CB_0.config_dataA\[16\] _0329_ vssd1 vssd1 vccd1 vccd1
+ _0341_ sky130_fd_sc_hd__or3_1
X_1717_ net28 net123 _0476_ vssd1 vssd1 vccd1 vccd1 _0479_ sky130_fd_sc_hd__mux2_1
X_2697_ SB0.route_sel\[97\] SB0.route_sel\[96\] net263 vssd1 vssd1 vccd1 vccd1 _0233_
+ sky130_fd_sc_hd__mux2_1
X_1648_ _1162_ SB0.route_sel\[13\] vssd1 vssd1 vccd1 vccd1 _0410_ sky130_fd_sc_hd__nor2_1
XFILLER_25_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1933__A2 _1320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2110__A2 net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output112_A net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2620_ SB0.route_sel\[20\] SB0.route_sel\[19\] net232 vssd1 vssd1 vccd1 vccd1 _0156_
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput106 net106 vssd1 vssd1 vccd1 vccd1 SBwest_out[10] sky130_fd_sc_hd__buf_2
Xoutput117 net117 vssd1 vssd1 vccd1 vccd1 SBwest_out[8] sky130_fd_sc_hd__buf_2
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1433_ LEI0.config_data\[17\] vssd1 vssd1 vccd1 vccd1 _1227_ sky130_fd_sc_hd__inv_2
X_2551_ net275 net273 net242 vssd1 vssd1 vccd1 vccd1 _0088_ sky130_fd_sc_hd__mux2_1
X_2482_ net396 net390 net235 vssd1 vssd1 vccd1 vccd1 _0021_ sky130_fd_sc_hd__mux2_1
X_1502_ SB0.route_sel\[51\] SB0.route_sel\[50\] _1186_ SB0.route_sel\[53\] vssd1 vssd1
+ vccd1 vccd1 _1296_ sky130_fd_sc_hd__o22a_1
X_3034_ clknet_leaf_12_clk _0242_ net224 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[106\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__1931__B _0339_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3103_ clknet_leaf_0_clk _0311_ net192 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_1364_ SB0.route_sel\[6\] vssd1 vssd1 vccd1 vccd1 _1158_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_43_Left_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1659__A net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2749_ net158 net160 net271 vssd1 vssd1 vccd1 vccd1 _0285_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_52_Left_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1591__B1_N net32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2818_ clknet_leaf_3_clk net395 net201 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_61_Left_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput19 CBnorth_in[13] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_52_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2159__A2 net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1982_ _1233_ _0735_ _0741_ vssd1 vssd1 vccd1 vccd1 _0742_ sky130_fd_sc_hd__a21o_1
X_2534_ net60 _0934_ vssd1 vssd1 vccd1 vccd1 _1152_ sky130_fd_sc_hd__and2_1
X_2603_ SB0.route_sel\[3\] SB0.route_sel\[2\] net237 vssd1 vssd1 vccd1 vccd1 _0139_
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2465_ net329 net320 net246 vssd1 vssd1 vccd1 vccd1 _0004_ sky130_fd_sc_hd__mux2_1
X_1416_ SB0.route_sel\[96\] vssd1 vssd1 vccd1 vccd1 _1210_ sky130_fd_sc_hd__inv_2
X_2396_ _1184_ SB0.route_sel\[50\] _1186_ SB0.route_sel\[53\] _1107_ vssd1 vssd1 vccd1
+ vccd1 _1108_ sky130_fd_sc_hd__a221o_1
X_3017_ clknet_leaf_2_clk _0225_ net197 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[89\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_fanout260_A net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_5_Left_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout152 CB_1.config_dataA\[0\] vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__clkbuf_2
Xfanout174 CB_0.config_dataA\[0\] vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__buf_2
Xfanout163 CB_0.config_dataB\[8\] vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__buf_2
Xfanout185 CB_1.config_dataB\[4\] vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__clkbuf_4
Xfanout141 CB_0.le_outA vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__buf_2
Xfanout130 CB_1.le_outA vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__clkbuf_4
Xfanout196 net197 vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1824__A1 net20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1760__A0 net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2250_ _0816_ _0819_ _0813_ _0822_ _1245_ CB_1.config_dataB\[9\] vssd1 vssd1 vccd1
+ vccd1 _1006_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_63_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2181_ _1359_ _0335_ _0795_ _1242_ vssd1 vssd1 vccd1 vccd1 _0937_ sky130_fd_sc_hd__a31o_1
XFILLER_18_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1965_ _0538_ _0512_ net163 vssd1 vssd1 vccd1 vccd1 _0725_ sky130_fd_sc_hd__mux2_1
X_2517_ net359 net340 net247 vssd1 vssd1 vccd1 vccd1 _0055_ sky130_fd_sc_hd__mux2_1
X_1896_ net15 net20 net21 net22 net165 CB_0.config_dataB\[5\] vssd1 vssd1 vccd1 vccd1
+ _0656_ sky130_fd_sc_hd__mux4_1
X_2448_ _1141_ _1142_ _0356_ vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__o21a_1
X_2379_ _1095_ _1096_ _0489_ vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_3_157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1806__A1 _1321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1990__A0 net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input36_A SBsouth_in[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold8 LE_1B.config_data\[9\] vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_60_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1750_ _0509_ _0510_ _0511_ _0508_ vssd1 vssd1 vccd1 vccd1 _0512_ sky130_fd_sc_hd__o31a_2
XFILLER_15_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1681_ _0438_ _0441_ _0442_ SB0.route_sel\[16\] SB0.route_sel\[17\] vssd1 vssd1 vccd1
+ vccd1 _0443_ sky130_fd_sc_hd__o311a_1
X_2233_ LE_1B.config_data\[6\] net120 net135 _0984_ _0986_ vssd1 vssd1 vccd1 vccd1
+ _0989_ sky130_fd_sc_hd__a32o_1
X_2302_ _0987_ _1056_ _1057_ _1054_ _1055_ vssd1 vssd1 vccd1 vccd1 _1058_ sky130_fd_sc_hd__o32a_1
X_2164_ _0905_ _0919_ _0921_ _0918_ vssd1 vssd1 vccd1 vccd1 _0922_ sky130_fd_sc_hd__o211a_1
X_2095_ net151 _0831_ vssd1 vssd1 vccd1 vccd1 _0853_ sky130_fd_sc_hd__nor2_1
XANTENNA__2461__A1 _0645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout223_A net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1879_ LE_0A.config_data\[11\] LE_0A.config_data\[10\] _0543_ vssd1 vssd1 vccd1 vccd1
+ _0641_ sky130_fd_sc_hd__mux2_1
X_1948_ net164 _0359_ vssd1 vssd1 vccd1 vccd1 _0708_ sky130_fd_sc_hd__nor2_1
XANTENNA__2213__A1 net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2997_ clknet_leaf_25_clk _0205_ net196 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[69\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_44_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_22_clk_A clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2204__B2 LEI0.config_data\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_8_Left_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2920_ clknet_leaf_15_clk _0128_ net222 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[12\]
+ sky130_fd_sc_hd__dfstp_1
Xclkbuf_2_3__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_2_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA_clkload1_A clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1802_ net171 _1216_ _0561_ _0563_ vssd1 vssd1 vccd1 vccd1 _0564_ sky130_fd_sc_hd__o31a_1
X_1733_ net155 net153 net159 net157 vssd1 vssd1 vccd1 vccd1 _0495_ sky130_fd_sc_hd__and4b_1
X_2851_ clknet_leaf_6_clk _0059_ net204 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_2782_ net373 net280 net234 vssd1 vssd1 vccd1 vccd1 _0318_ sky130_fd_sc_hd__mux2_1
X_1595_ SB0.route_sel\[98\] SB0.route_sel\[99\] vssd1 vssd1 vccd1 vccd1 _0357_ sky130_fd_sc_hd__nor2_1
X_1664_ SB0.route_sel\[3\] SB0.route_sel\[2\] _0425_ _0413_ vssd1 vssd1 vccd1 vccd1
+ _0426_ sky130_fd_sc_hd__a31oi_1
X_2216_ net4 net5 net185 vssd1 vssd1 vccd1 vccd1 _0972_ sky130_fd_sc_hd__mux2_1
X_2147_ CB_1.config_dataA\[13\] CB_1.config_dataA\[15\] vssd1 vssd1 vccd1 vccd1 _0905_
+ sky130_fd_sc_hd__nand2b_1
X_2078_ SB0.route_sel\[87\] SB0.route_sel\[86\] vssd1 vssd1 vccd1 vccd1 _0836_ sky130_fd_sc_hd__nand2b_1
XANTENNA__1668__Y _0430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1960__A3 net22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_34_Left_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2122__A0 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1380_ SB0.route_sel\[30\] vssd1 vssd1 vccd1 vccd1 _1174_ sky130_fd_sc_hd__inv_2
X_3050_ clknet_leaf_7_clk _0258_ net206 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[10\]
+ sky130_fd_sc_hd__dfstp_1
X_2001_ LE_0B.config_data\[3\] _0703_ _0760_ _0676_ vssd1 vssd1 vccd1 vccd1 _0761_
+ sky130_fd_sc_hd__a211o_1
XANTENNA__2361__B1 _0781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2903_ clknet_leaf_28_clk _0111_ net188 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_2834_ clknet_leaf_12_clk net363 net224 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[41\]
+ sky130_fd_sc_hd__dfrtp_1
X_1716_ _1248_ _0476_ _0477_ vssd1 vssd1 vccd1 vccd1 _0478_ sky130_fd_sc_hd__a21oi_1
X_2696_ SB0.route_sel\[96\] SB0.route_sel\[95\] net263 vssd1 vssd1 vccd1 vccd1 _0232_
+ sky130_fd_sc_hd__mux2_1
X_2765_ CB_1.config_dataA\[13\] net146 net261 vssd1 vssd1 vccd1 vccd1 _0301_ sky130_fd_sc_hd__mux2_1
X_1578_ net174 _0339_ vssd1 vssd1 vccd1 vccd1 _0340_ sky130_fd_sc_hd__nand2_1
X_1647_ SB0.route_sel\[11\] SB0.route_sel\[10\] vssd1 vssd1 vccd1 vccd1 _0409_ sky130_fd_sc_hd__nor2_1
XANTENNA__3052__SET_B net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2104__A0 _0838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1558__C net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2343__A0 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2110__A3 net12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output105_A net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput107 net107 vssd1 vssd1 vccd1 vccd1 SBwest_out[11] sky130_fd_sc_hd__buf_2
X_2550_ net273 LE_0B.config_data\[13\] net242 vssd1 vssd1 vccd1 vccd1 _0087_ sky130_fd_sc_hd__mux2_1
Xoutput118 net118 vssd1 vssd1 vccd1 vccd1 SBwest_out[9] sky130_fd_sc_hd__buf_2
X_1432_ CB_0.config_dataB\[3\] vssd1 vssd1 vccd1 vccd1 _1226_ sky130_fd_sc_hd__inv_2
X_2481_ net390 LEI0.config_data\[18\] net244 vssd1 vssd1 vccd1 vccd1 _0020_ sky130_fd_sc_hd__mux2_1
X_1363_ SB0.route_sel\[7\] vssd1 vssd1 vccd1 vccd1 _1157_ sky130_fd_sc_hd__inv_2
X_1501_ SB0.route_sel\[54\] SB0.route_sel\[55\] vssd1 vssd1 vccd1 vccd1 _1295_ sky130_fd_sc_hd__nand2b_1
X_3033_ clknet_leaf_12_clk _0241_ net224 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[105\]
+ sky130_fd_sc_hd__dfstp_2
X_3102_ clknet_leaf_0_clk _0310_ net192 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__1860__A2 _0473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout136_A net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2748_ net159 CB_0.config_dataB\[15\] net272 vssd1 vssd1 vccd1 vccd1 _0284_ sky130_fd_sc_hd__mux2_1
X_2817_ clknet_leaf_3_clk net286 net201 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_2679_ SB0.route_sel\[79\] SB0.route_sel\[78\] net239 vssd1 vssd1 vccd1 vccd1 _0215_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__2325__A0 _0512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2159__A3 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2033__X _0791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input21_X net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1981_ CB_0.config_dataB\[15\] _0739_ _0740_ _0736_ vssd1 vssd1 vccd1 vccd1 _0741_
+ sky130_fd_sc_hd__o22a_1
X_2602_ SB0.route_sel\[2\] SB0.route_sel\[1\] net237 vssd1 vssd1 vccd1 vccd1 _0138_
+ sky130_fd_sc_hd__mux2_1
X_2533_ LE_0B.dff0_out _1247_ _1151_ vssd1 vssd1 vccd1 vccd1 _0071_ sky130_fd_sc_hd__a21o_1
XFILLER_9_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_21_Left_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2464_ net320 LEI0.config_data\[1\] net242 vssd1 vssd1 vccd1 vccd1 _0003_ sky130_fd_sc_hd__mux2_1
X_1415_ SB0.route_sel\[102\] vssd1 vssd1 vccd1 vccd1 _1209_ sky130_fd_sc_hd__inv_2
XFILLER_28_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2395_ SB0.route_sel\[49\] SB0.route_sel\[48\] vssd1 vssd1 vccd1 vccd1 _1107_ sky130_fd_sc_hd__nor2_1
XANTENNA__1833__A2 _0359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3016_ clknet_leaf_2_clk _0224_ net209 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[88\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__2086__A2 _0838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout253_A net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_31_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_2_1__f_clk_X clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout120 _0957_ vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__buf_2
Xfanout131 net132 vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__buf_2
Xfanout153 CB_0.config_dataB\[19\] vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__clkbuf_2
XFILLER_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout164 CB_0.config_dataB\[8\] vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout197 net198 vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__clkbuf_4
Xfanout186 net193 vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_6_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout175 CB_1.config_dataB\[19\] vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__buf_2
Xfanout142 CB_1.config_dataA\[19\] vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__clkbuf_2
XFILLER_63_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1824__A2 net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_22_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_33_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2180_ _0781_ _0784_ _0788_ _0792_ _1241_ _1242_ vssd1 vssd1 vccd1 vccd1 _0936_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_63_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_13_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1964_ _0707_ _0721_ _0723_ vssd1 vssd1 vccd1 vccd1 _0724_ sky130_fd_sc_hd__o21a_1
X_1895_ net165 _0654_ vssd1 vssd1 vccd1 vccd1 _0655_ sky130_fd_sc_hd__nor2_1
X_2516_ net340 net335 net246 vssd1 vssd1 vccd1 vccd1 _0054_ sky130_fd_sc_hd__mux2_1
X_2447_ _1206_ SB0.route_sel\[99\] _1208_ _1209_ vssd1 vssd1 vccd1 vccd1 _1142_ sky130_fd_sc_hd__a22o_1
X_2378_ SB0.route_sel\[76\] _1195_ SB0.route_sel\[73\] SB0.route_sel\[72\] vssd1 vssd1
+ vccd1 vccd1 _1096_ sky130_fd_sc_hd__o22ai_1
XTAP_TAPCELL_ROW_3_158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1863__A _0447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1990__A1 net20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold9 _0317_ vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input29_A SBsouth_in[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1597__X _0359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2222__A2 _1342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1680_ SB0.route_sel\[20\] SB0.route_sel\[21\] net35 vssd1 vssd1 vccd1 vccd1 _0442_
+ sky130_fd_sc_hd__a21boi_1
X_2301_ LE_1B.config_data\[12\] net120 net135 vssd1 vssd1 vccd1 vccd1 _1057_ sky130_fd_sc_hd__and3_1
XFILLER_38_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_2_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2163_ _0911_ _0920_ vssd1 vssd1 vccd1 vccd1 _0921_ sky130_fd_sc_hd__or2_1
X_2232_ _0987_ vssd1 vssd1 vccd1 vccd1 _0988_ sky130_fd_sc_hd__inv_2
X_2094_ CB_1.config_dataA\[1\] _1235_ vssd1 vssd1 vccd1 vccd1 _0852_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_0_139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1878_ _0639_ _0638_ _0572_ vssd1 vssd1 vccd1 vccd1 _0640_ sky130_fd_sc_hd__mux2_1
X_1947_ CB_0.config_dataB\[9\] _1230_ vssd1 vssd1 vccd1 vccd1 _0707_ sky130_fd_sc_hd__or2_1
XANTENNA__2213__A2 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout216_A net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2996_ clknet_leaf_25_clk _0204_ net197 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[68\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1488__B1 net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2850_ clknet_leaf_6_clk net299 net204 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_1801_ CB_0.config_dataA\[7\] _0562_ vssd1 vssd1 vccd1 vccd1 _0563_ sky130_fd_sc_hd__or2_1
X_1732_ _1250_ _0450_ vssd1 vssd1 vccd1 vccd1 _0494_ sky130_fd_sc_hd__nand2b_1
X_1663_ _0424_ _1159_ _0423_ vssd1 vssd1 vccd1 vccd1 _0425_ sky130_fd_sc_hd__mux2_1
X_2781_ net280 LE_1B.config_data\[8\] net234 vssd1 vssd1 vccd1 vccd1 _0317_ sky130_fd_sc_hd__mux2_1
X_1594_ _0344_ _0345_ _0351_ _0355_ vssd1 vssd1 vccd1 vccd1 _0356_ sky130_fd_sc_hd__a22o_2
XPHY_EDGE_ROW_7_Right_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2215_ net183 _0966_ _0970_ vssd1 vssd1 vccd1 vccd1 _0971_ sky130_fd_sc_hd__a21oi_1
X_2077_ _0833_ _0834_ _0508_ vssd1 vssd1 vccd1 vccd1 _0835_ sky130_fd_sc_hd__a21boi_4
X_2146_ CB_1.config_dataA\[15\] _0903_ vssd1 vssd1 vccd1 vccd1 _0904_ sky130_fd_sc_hd__and2b_1
X_2979_ clknet_leaf_22_clk _0187_ net214 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[51\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__2122__A1 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1633__A0 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2000_ LE_0B.config_data\[2\] _0700_ _0702_ vssd1 vssd1 vccd1 vccd1 _0760_ sky130_fd_sc_hd__and3_1
X_2833_ clknet_leaf_12_clk _0041_ net224 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[40\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_23_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2902_ clknet_leaf_22_clk _0110_ net214 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_1715_ _1298_ _0450_ vssd1 vssd1 vccd1 vccd1 _0477_ sky130_fd_sc_hd__and2_1
X_2695_ SB0.route_sel\[95\] SB0.route_sel\[94\] net263 vssd1 vssd1 vccd1 vccd1 _0231_
+ sky130_fd_sc_hd__mux2_1
X_1646_ _1163_ SB0.route_sel\[14\] vssd1 vssd1 vccd1 vccd1 _0408_ sky130_fd_sc_hd__nor2_1
X_2764_ net146 CB_1.config_dataA\[11\] net260 vssd1 vssd1 vccd1 vccd1 _0300_ sky130_fd_sc_hd__mux2_1
X_1577_ _1358_ _0334_ _0338_ vssd1 vssd1 vccd1 vccd1 _0339_ sky130_fd_sc_hd__or3b_4
XANTENNA_clkbuf_leaf_21_clk_A clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2129_ LEI0.config_data\[32\] _0886_ vssd1 vssd1 vccd1 vccd1 _0887_ sky130_fd_sc_hd__nand2b_1
XANTENNA__1854__A0 _1321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input11_A CBeast_in[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput108 net108 vssd1 vssd1 vccd1 vccd1 SBwest_out[12] sky130_fd_sc_hd__buf_2
X_2480_ net414 net385 net244 vssd1 vssd1 vccd1 vccd1 _0019_ sky130_fd_sc_hd__mux2_1
Xoutput119 net119 vssd1 vssd1 vccd1 vccd1 config_data_out sky130_fd_sc_hd__buf_2
X_1500_ _1293_ _1289_ _1279_ _1278_ vssd1 vssd1 vccd1 vccd1 _1294_ sky130_fd_sc_hd__a2bb2o_1
Xoutput90 net90 vssd1 vssd1 vccd1 vccd1 CBnorth_out[9] sky130_fd_sc_hd__buf_2
X_1431_ net167 vssd1 vssd1 vccd1 vccd1 _1225_ sky130_fd_sc_hd__inv_2
X_3101_ clknet_leaf_0_clk net284 net192 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_1362_ SB0.route_sel\[5\] vssd1 vssd1 vccd1 vccd1 _1156_ sky130_fd_sc_hd__inv_2
X_3032_ clknet_leaf_10_clk _0240_ net221 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[104\]
+ sky130_fd_sc_hd__dfstp_2
XANTENNA__2098__A0 net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2926__SET_B net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout129_A net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2816_ clknet_leaf_0_clk _0024_ net191 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_2747_ CB_0.config_dataB\[15\] CB_0.config_dataB\[14\] net265 vssd1 vssd1 vccd1 vccd1
+ _0283_ sky130_fd_sc_hd__mux2_1
X_2678_ SB0.route_sel\[78\] SB0.route_sel\[77\] net236 vssd1 vssd1 vccd1 vccd1 _0214_
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1629_ _0388_ _0390_ vssd1 vssd1 vccd1 vccd1 _0391_ sky130_fd_sc_hd__nand2_4
XANTENNA_input3_A CBeast_in[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2089__A0 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2461__S net60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input59_A le_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1827__A0 net27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input14_X net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1980_ net18 net19 net162 vssd1 vssd1 vccd1 vccd1 _0740_ sky130_fd_sc_hd__mux2_1
XANTENNA__2252__A0 net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2463_ net383 LEI0.config_data\[0\] net242 vssd1 vssd1 vccd1 vccd1 _0002_ sky130_fd_sc_hd__mux2_1
X_2532_ LE_0A.reset_mode net415 net236 vssd1 vssd1 vccd1 vccd1 _0070_ sky130_fd_sc_hd__mux2_1
X_2601_ SB0.route_sel\[1\] SB0.route_sel\[0\] net237 vssd1 vssd1 vccd1 vccd1 _0137_
+ sky130_fd_sc_hd__mux2_1
X_1414_ SB0.route_sel\[103\] vssd1 vssd1 vccd1 vccd1 _1208_ sky130_fd_sc_hd__inv_2
X_3015_ clknet_leaf_2_clk _0223_ net208 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[87\]
+ sky130_fd_sc_hd__dfstp_1
X_2394_ _1105_ _1106_ _1270_ vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__o21a_1
XANTENNA__2491__A0 LEI0.config_data\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout246_A net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1686__A _0447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout154 CB_0.config_dataB\[19\] vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__clkbuf_2
Xfanout165 CB_0.config_dataB\[4\] vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input6_X net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout132 net133 vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__buf_1
Xfanout143 CB_1.config_dataA\[18\] vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__clkbuf_2
XFILLER_63_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout198 net229 vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout187 net193 vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__buf_2
Xfanout176 CB_1.config_dataB\[18\] vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__buf_2
XANTENNA__1824__A3 net22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1883__X _0645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2473__A0 LEI0.config_data\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1963_ CB_0.config_dataB\[11\] _0720_ _0722_ _0705_ vssd1 vssd1 vccd1 vccd1 _0723_
+ sky130_fd_sc_hd__o22a_1
X_1894_ CB_0.config_dataB\[5\] CB_0.config_dataB\[7\] vssd1 vssd1 vccd1 vccd1 _0654_
+ sky130_fd_sc_hd__nand2_1
X_2515_ net335 net294 net249 vssd1 vssd1 vccd1 vccd1 _0053_ sky130_fd_sc_hd__mux2_1
X_2446_ _1210_ SB0.route_sel\[97\] vssd1 vssd1 vccd1 vccd1 _1141_ sky130_fd_sc_hd__nor2_1
X_2377_ SB0.route_sel\[75\] SB0.route_sel\[74\] vssd1 vssd1 vccd1 vccd1 _1095_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_3_159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_49_Left_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2216__A0 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1990__A2 net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_58_Left_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2222__A3 _0791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2231_ _0984_ _0986_ vssd1 vssd1 vccd1 vccd1 _0987_ sky130_fd_sc_hd__nand2_2
X_2300_ net120 net135 LE_1B.config_data\[13\] vssd1 vssd1 vccd1 vccd1 _1056_ sky130_fd_sc_hd__a21boi_1
X_2093_ _0819_ _0822_ _0816_ _0813_ CB_1.config_dataA\[1\] net151 vssd1 vssd1 vccd1
+ vccd1 _0851_ sky130_fd_sc_hd__mux4_1
X_2162_ net2 net3 net147 vssd1 vssd1 vccd1 vccd1 _0920_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1948__B _0359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2995_ clknet_leaf_25_clk _0203_ net197 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[67\]
+ sky130_fd_sc_hd__dfstp_1
X_1877_ LE_0A.config_data\[13\] LE_0A.config_data\[12\] _0543_ vssd1 vssd1 vccd1 vccd1
+ _0639_ sky130_fd_sc_hd__mux2_1
X_1946_ _1345_ _1321_ _1297_ _1273_ net163 CB_0.config_dataB\[9\] vssd1 vssd1 vccd1
+ vccd1 _0706_ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout209_A net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2213__A3 net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2429_ _1161_ SB0.route_sel\[10\] SB0.route_sel\[9\] _1164_ vssd1 vssd1 vccd1 vccd1
+ _1130_ sky130_fd_sc_hd__o22a_1
XANTENNA_input41_A SBsouth_in[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2140__A2 _0838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1800_ net23 net24 net25 net26 net173 net171 vssd1 vssd1 vccd1 vccd1 _0562_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_13_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1784__A net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1731_ _0489_ _0491_ vssd1 vssd1 vccd1 vccd1 _0493_ sky130_fd_sc_hd__nand2_2
X_1662_ SB0.route_sel\[7\] SB0.route_sel\[6\] net43 vssd1 vssd1 vccd1 vccd1 _0424_
+ sky130_fd_sc_hd__a21bo_1
X_2780_ net287 LE_1B.config_data\[7\] net234 vssd1 vssd1 vccd1 vccd1 _0316_ sky130_fd_sc_hd__mux2_1
X_1593_ _0352_ _0354_ _0344_ vssd1 vssd1 vccd1 vccd1 _0355_ sky130_fd_sc_hd__o21ba_1
X_2214_ net183 _0969_ _0968_ CB_1.config_dataB\[6\] vssd1 vssd1 vccd1 vccd1 _0970_
+ sky130_fd_sc_hd__a211o_1
XFILLER_53_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2076_ SB0.route_sel\[92\] SB0.route_sel\[93\] SB0.route_sel\[88\] _1205_ vssd1 vssd1
+ vccd1 vccd1 _0834_ sky130_fd_sc_hd__o22a_1
X_2145_ _0792_ _0788_ _0784_ _0781_ CB_1.config_dataA\[13\] net146 vssd1 vssd1 vccd1
+ vccd1 _0903_ sky130_fd_sc_hd__mux4_1
XFILLER_61_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1929_ _0681_ _0682_ _0684_ _0686_ net166 _1226_ vssd1 vssd1 vccd1 vccd1 _0689_ sky130_fd_sc_hd__mux4_1
X_2978_ clknet_leaf_22_clk _0186_ net214 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[50\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_55_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2122__A2 net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1633__A1 net20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold90 LEI0.config_data\[40\] vssd1 vssd1 vccd1 vccd1 net362 sky130_fd_sc_hd__dlygate4sd3_1
X_2832_ clknet_leaf_12_clk _0040_ net224 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[39\]
+ sky130_fd_sc_hd__dfrtp_1
X_2901_ clknet_leaf_22_clk net303 net214 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_2763_ CB_1.config_dataA\[11\] CB_1.config_dataA\[10\] net260 vssd1 vssd1 vccd1 vccd1
+ _0299_ sky130_fd_sc_hd__mux2_1
X_1714_ net157 net155 net153 net160 vssd1 vssd1 vccd1 vccd1 _0476_ sky130_fd_sc_hd__and4bb_1
X_1576_ SB0.route_sel\[108\] _1211_ net119 _1212_ _0337_ vssd1 vssd1 vccd1 vccd1 _0338_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__2403__A _1318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2694_ SB0.route_sel\[94\] SB0.route_sel\[93\] net263 vssd1 vssd1 vccd1 vccd1 _0230_
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1645_ _0396_ _0397_ _0401_ _0406_ vssd1 vssd1 vccd1 vccd1 _0407_ sky130_fd_sc_hd__a22o_1
X_2128_ net139 net125 net128 net133 LEI0.config_data\[30\] LEI0.config_data\[31\]
+ vssd1 vssd1 vccd1 vccd1 _0886_ sky130_fd_sc_hd__mux4_1
XFILLER_26_147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2059_ SB0.route_sel\[4\] SB0.route_sel\[5\] vssd1 vssd1 vccd1 vccd1 _0817_ sky130_fd_sc_hd__nor2_1
XFILLER_41_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1854__A1 _1345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_55_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput109 net109 vssd1 vssd1 vccd1 vccd1 SBwest_out[13] sky130_fd_sc_hd__buf_2
X_1430_ net166 vssd1 vssd1 vccd1 vccd1 _1224_ sky130_fd_sc_hd__inv_2
Xoutput80 net80 vssd1 vssd1 vccd1 vccd1 CBnorth_out[12] sky130_fd_sc_hd__buf_2
X_3031_ clknet_leaf_10_clk _0239_ net220 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[103\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__2098__A1 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3100_ clknet_leaf_0_clk _0308_ net192 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_1361_ SB0.route_sel\[3\] vssd1 vssd1 vccd1 vccd1 _1155_ sky130_fd_sc_hd__inv_2
Xoutput91 net91 vssd1 vssd1 vccd1 vccd1 SBsouth_out[0] sky130_fd_sc_hd__buf_2
X_2746_ CB_0.config_dataB\[14\] CB_0.config_dataB\[13\] net265 vssd1 vssd1 vccd1 vccd1
+ _0282_ sky130_fd_sc_hd__mux2_1
X_2815_ clknet_leaf_0_clk _0023_ net191 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_2677_ SB0.route_sel\[77\] SB0.route_sel\[76\] net235 vssd1 vssd1 vccd1 vccd1 _0213_
+ sky130_fd_sc_hd__mux2_1
X_1559_ _1349_ _1350_ _1351_ _1352_ vssd1 vssd1 vccd1 vccd1 _1353_ sky130_fd_sc_hd__a31o_1
X_1628_ SB0.route_sel\[28\] _1172_ SB0.route_sel\[31\] _1174_ _0389_ vssd1 vssd1 vccd1
+ vccd1 _0390_ sky130_fd_sc_hd__a221o_1
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2089__A1 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2261__B2 LEI0.config_data\[35\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1772__B1 _0524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1827__A1 net28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output110_A net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2252__A1 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2600_ SB0.route_sel\[0\] CB_1.config_dataB\[19\] net237 vssd1 vssd1 vccd1 vccd1
+ _0136_ sky130_fd_sc_hd__mux2_1
XFILLER_9_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_20_clk_A clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1413_ SB0.route_sel\[101\] vssd1 vssd1 vccd1 vccd1 _1207_ sky130_fd_sc_hd__inv_2
XANTENNA__1763__B1 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2531_ net415 LE_0A.edge_mode net234 vssd1 vssd1 vccd1 vccd1 _0069_ sky130_fd_sc_hd__mux2_1
X_2462_ LEI0.config_data\[0\] LE_1A.reset_mode net230 vssd1 vssd1 vccd1 vccd1 _0001_
+ sky130_fd_sc_hd__mux2_1
X_2393_ SB0.route_sel\[63\] SB0.route_sel\[62\] _1190_ SB0.route_sel\[56\] vssd1 vssd1
+ vccd1 vccd1 _1106_ sky130_fd_sc_hd__a2bb2o_1
X_3014_ clknet_leaf_2_clk _0222_ net208 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[86\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_3_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2415__X net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2729_ CB_0.config_dataA\[17\] CB_0.config_dataA\[16\] net265 vssd1 vssd1 vccd1 vccd1
+ _0265_ sky130_fd_sc_hd__mux2_1
Xfanout155 CB_0.config_dataB\[18\] vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__clkbuf_2
Xfanout199 net202 vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__clkbuf_4
Xfanout166 CB_0.config_dataB\[1\] vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__buf_2
Xfanout122 net127 vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__buf_2
Xfanout177 CB_1.config_dataB\[17\] vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout188 net193 vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__clkbuf_4
Xfanout133 net134 vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__buf_2
Xfanout144 CB_1.config_dataA\[17\] vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_29_Right_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Right_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_47_Right_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2170__B1 _0912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_56_Right_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1962_ net16 net17 net164 vssd1 vssd1 vccd1 vccd1 _0722_ sky130_fd_sc_hd__mux2_1
XFILLER_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1893_ _1228_ _0492_ _0651_ _0652_ vssd1 vssd1 vccd1 vccd1 _0653_ sky130_fd_sc_hd__o211a_1
X_2514_ net294 LE_0A.config_data\[0\] net249 vssd1 vssd1 vccd1 vccd1 _0052_ sky130_fd_sc_hd__mux2_1
X_2445_ _1139_ _1140_ _0356_ vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__a21boi_2
X_2376_ _0420_ _1094_ _0421_ vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__a21o_1
XANTENNA__2161__A0 net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2129__Y _0887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout189_A net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1975__A0 _1345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2216__A1 net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1990__A3 net22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2230_ LEI0.config_data\[23\] _0985_ vssd1 vssd1 vccd1 vccd1 _0986_ sky130_fd_sc_hd__nand2b_1
XANTENNA__2143__B1 _0887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2231__A _0984_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2092_ _0849_ vssd1 vssd1 vccd1 vccd1 _0850_ sky130_fd_sc_hd__inv_2
X_2161_ net13 net14 net146 vssd1 vssd1 vccd1 vccd1 _0919_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_2_2__f_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1945_ CB_0.config_dataB\[9\] CB_0.config_dataB\[11\] vssd1 vssd1 vccd1 vccd1 _0705_
+ sky130_fd_sc_hd__nand2_1
XFILLER_9_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2406__A _1318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2994_ clknet_leaf_25_clk _0202_ net197 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[66\]
+ sky130_fd_sc_hd__dfstp_1
X_1876_ LE_0A.config_data\[15\] LE_0A.config_data\[14\] _0543_ vssd1 vssd1 vccd1 vccd1
+ _0638_ sky130_fd_sc_hd__mux2_1
XANTENNA__1725__B1_N net42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2428_ SB0.route_sel\[15\] SB0.route_sel\[14\] vssd1 vssd1 vccd1 vccd1 _1129_ sky130_fd_sc_hd__or2_1
X_2359_ _1329_ _0456_ _0831_ vssd1 vssd1 vccd1 vccd1 _1086_ sky130_fd_sc_hd__a21o_1
XFILLER_56_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout261_X net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2373__B1 _0816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input34_A SBsouth_in[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1592_ _0349_ _0353_ vssd1 vssd1 vccd1 vccd1 _0354_ sky130_fd_sc_hd__nand2_1
X_1730_ _0489_ _0491_ vssd1 vssd1 vccd1 vccd1 _0492_ sky130_fd_sc_hd__and2_1
XANTENNA__2600__A1 CB_1.config_dataB\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1661_ SB0.route_sel\[4\] SB0.route_sel\[5\] vssd1 vssd1 vccd1 vccd1 _0423_ sky130_fd_sc_hd__nand2_1
XFILLER_38_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2213_ net13 net14 net2 net3 net185 net184 vssd1 vssd1 vccd1 vccd1 _0969_ sky130_fd_sc_hd__mux4_1
X_2144_ LE_1A.config_data\[5\] LE_1A.config_data\[7\] LE_1A.config_data\[4\] LE_1A.config_data\[6\]
+ _0848_ _0874_ vssd1 vssd1 vccd1 vccd1 _0902_ sky130_fd_sc_hd__mux4_1
XFILLER_53_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2075_ SB0.route_sel\[95\] SB0.route_sel\[94\] vssd1 vssd1 vccd1 vccd1 _0833_ sky130_fd_sc_hd__nand2b_1
X_1859_ _1221_ _0493_ vssd1 vssd1 vccd1 vccd1 _0621_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout221_A net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1928_ CB_0.config_dataB\[3\] _0683_ _0687_ vssd1 vssd1 vccd1 vccd1 _0688_ sky130_fd_sc_hd__a21oi_1
X_2977_ clknet_leaf_22_clk _0185_ net214 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[49\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__2355__B1 _0838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2122__A3 net12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold80 LE_0A.config_data\[0\] vssd1 vssd1 vccd1 vccd1 net352 sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 _0042_ vssd1 vssd1 vccd1 vccd1 net363 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_50_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2900_ clknet_leaf_21_clk _0108_ net215 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_2831_ clknet_leaf_13_clk _0039_ net224 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[38\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_33_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1713_ SB0.route_sel\[73\] SB0.route_sel\[72\] vssd1 vssd1 vccd1 vccd1 _0475_ sky130_fd_sc_hd__nand2_1
X_2762_ CB_1.config_dataA\[10\] CB_1.config_dataA\[9\] net260 vssd1 vssd1 vccd1 vccd1
+ _0298_ sky130_fd_sc_hd__mux2_1
X_1575_ SB0.route_sel\[106\] SB0.route_sel\[107\] vssd1 vssd1 vccd1 vccd1 _0337_ sky130_fd_sc_hd__nor2_1
XANTENNA__2337__A0 _1321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2693_ SB0.route_sel\[93\] SB0.route_sel\[92\] net241 vssd1 vssd1 vccd1 vccd1 _0229_
+ sky130_fd_sc_hd__mux2_1
X_1644_ _0403_ _0405_ _0396_ vssd1 vssd1 vccd1 vccd1 _0406_ sky130_fd_sc_hd__a21oi_1
XFILLER_58_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1560__A1 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2127_ _0876_ _0879_ _0882_ _0884_ vssd1 vssd1 vccd1 vccd1 _0885_ sky130_fd_sc_hd__a31o_1
XFILLER_26_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2058_ _0407_ _0815_ vssd1 vssd1 vccd1 vccd1 _0816_ sky130_fd_sc_hd__nand2_4
XTAP_TAPCELL_ROW_55_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1360_ CB_0.config_dataA\[1\] vssd1 vssd1 vccd1 vccd1 _1154_ sky130_fd_sc_hd__inv_2
Xoutput70 net70 vssd1 vssd1 vccd1 vccd1 CBeast_out[3] sky130_fd_sc_hd__buf_2
Xoutput81 net81 vssd1 vssd1 vccd1 vccd1 CBnorth_out[13] sky130_fd_sc_hd__buf_2
X_3030_ clknet_leaf_10_clk _0238_ net219 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[102\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__2098__A2 net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput92 net92 vssd1 vssd1 vccd1 vccd1 SBsouth_out[10] sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_9_clk_A clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2745_ CB_0.config_dataB\[13\] net162 net265 vssd1 vssd1 vccd1 vccd1 _0281_ sky130_fd_sc_hd__mux2_1
X_2814_ clknet_leaf_1_clk _0022_ net191 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_2676_ SB0.route_sel\[76\] SB0.route_sel\[75\] net235 vssd1 vssd1 vccd1 vccd1 _0212_
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1558_ CB_1.config_dataA\[19\] CB_1.config_dataA\[18\] net128 _1308_ vssd1 vssd1
+ vccd1 vccd1 _1352_ sky130_fd_sc_hd__and4_1
X_1627_ SB0.route_sel\[26\] SB0.route_sel\[27\] vssd1 vssd1 vccd1 vccd1 _0389_ sky130_fd_sc_hd__nor2_1
X_1489_ net145 net144 vssd1 vssd1 vccd1 vccd1 _1283_ sky130_fd_sc_hd__and2b_1
XANTENNA__2089__A2 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1827__A2 net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2252__A2 net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_25_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__1460__A0 net26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2530_ LE_0A.edge_mode LE_0A.config_data\[16\] net234 vssd1 vssd1 vccd1 vccd1 _0068_
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2712__A0 CB_0.config_dataA\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1412_ SB0.route_sel\[98\] vssd1 vssd1 vccd1 vccd1 _1206_ sky130_fd_sc_hd__inv_2
X_2461_ LE_0A.dff1_out _0645_ net60 vssd1 vssd1 vccd1 vccd1 _0000_ sky130_fd_sc_hd__mux2_1
X_2392_ SB0.route_sel\[58\] _1188_ vssd1 vssd1 vccd1 vccd1 _1105_ sky130_fd_sc_hd__nor2_1
XFILLER_3_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3013_ clknet_leaf_2_clk _0221_ net197 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[85\]
+ sky130_fd_sc_hd__dfstp_1
Xclkbuf_leaf_16_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2728_ CB_0.config_dataA\[16\] CB_0.config_dataA\[15\] net265 vssd1 vssd1 vccd1 vccd1
+ _0264_ sky130_fd_sc_hd__mux2_1
X_2659_ SB0.route_sel\[59\] SB0.route_sel\[58\] net256 vssd1 vssd1 vccd1 vccd1 _0195_
+ sky130_fd_sc_hd__mux2_1
Xfanout156 CB_0.config_dataB\[18\] vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__clkbuf_2
Xfanout123 net124 vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__clkbuf_2
Xfanout167 CB_0.config_dataB\[0\] vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__buf_2
Xfanout134 CB_1.le_outB vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__buf_2
Xfanout178 CB_1.config_dataB\[16\] vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__buf_2
Xfanout189 net193 vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__clkbuf_2
Xfanout145 CB_1.config_dataA\[16\] vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__clkbuf_2
XANTENNA__1510__X _1304_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_25_Left_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1961_ net27 net28 net164 vssd1 vssd1 vccd1 vccd1 _0721_ sky130_fd_sc_hd__mux2_1
X_1892_ _1228_ _0474_ vssd1 vssd1 vccd1 vccd1 _0652_ sky130_fd_sc_hd__nand2_1
XFILLER_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2513_ net352 net57 net246 vssd1 vssd1 vccd1 vccd1 _0051_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_5_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2444_ _1206_ SB0.route_sel\[99\] SB0.route_sel\[100\] _1207_ vssd1 vssd1 vccd1 vccd1
+ _1140_ sky130_fd_sc_hd__o22a_1
X_2375_ _1330_ _0377_ _0819_ vssd1 vssd1 vccd1 vccd1 _1094_ sky130_fd_sc_hd__o21ai_1
XANTENNA__2161__A1 net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1975__A1 _1321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2748__S net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2055__Y _0813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2160_ CB_1.config_dataA\[15\] _0917_ vssd1 vssd1 vccd1 vccd1 _0918_ sky130_fd_sc_hd__or2_1
X_2091_ net141 net127 net128 net133 LEI0.config_data\[6\] LEI0.config_data\[7\] vssd1
+ vssd1 vccd1 vccd1 _0849_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_16_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1875_ _0636_ _0604_ _0602_ vssd1 vssd1 vccd1 vccd1 _0637_ sky130_fd_sc_hd__mux2_1
X_1944_ LE_0B.config_data\[4\] LE_0B.config_data\[5\] _0703_ vssd1 vssd1 vccd1 vccd1
+ _0704_ sky130_fd_sc_hd__mux2_1
X_2993_ clknet_leaf_25_clk _0201_ net197 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[65\]
+ sky130_fd_sc_hd__dfstp_1
X_2427_ _0407_ _1128_ vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__and2_1
X_2289_ _1201_ net181 CB_1.config_dataB\[15\] _1044_ net179 vssd1 vssd1 vccd1 vccd1
+ _1045_ sky130_fd_sc_hd__o2111a_1
X_2358_ _0482_ _1085_ _0484_ vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__a21o_1
XANTENNA_fanout254_X net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input27_A CBnorth_in[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1636__B1 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1591_ SB0.route_sel\[100\] SB0.route_sel\[101\] net32 vssd1 vssd1 vccd1 vccd1 _0353_
+ sky130_fd_sc_hd__a21bo_1
X_1660_ SB0.route_sel\[3\] SB0.route_sel\[2\] _0419_ _0420_ _0421_ vssd1 vssd1 vccd1
+ vccd1 _0422_ sky130_fd_sc_hd__a221o_1
XANTENNA_output95_A net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2212_ net183 _0967_ vssd1 vssd1 vccd1 vccd1 _0968_ sky130_fd_sc_hd__and2b_1
X_2143_ CB_1.config_dataA\[10\] _0900_ _0887_ _0885_ vssd1 vssd1 vccd1 vccd1 _0901_
+ sky130_fd_sc_hd__o211a_1
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2074_ _0827_ _0831_ _1237_ vssd1 vssd1 vccd1 vccd1 _0832_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_28_Left_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1858_ _0613_ _0619_ CB_0.config_dataA\[15\] _0607_ vssd1 vssd1 vccd1 vccd1 _0620_
+ sky130_fd_sc_hd__a2bb2o_1
X_1927_ _1226_ _0685_ CB_0.config_dataB\[2\] vssd1 vssd1 vccd1 vccd1 _0687_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout214_A net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2976_ clknet_leaf_22_clk _0184_ net214 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[48\]
+ sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_12_Left_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1789_ net15 net20 net173 vssd1 vssd1 vccd1 vccd1 _0551_ sky130_fd_sc_hd__mux2_1
XANTENNA__1866__A0 net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2291__A0 _0831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold92 LEI0.config_data\[13\] vssd1 vssd1 vccd1 vccd1 net364 sky130_fd_sc_hd__dlygate4sd3_1
Xhold70 _0062_ vssd1 vssd1 vccd1 vccd1 net342 sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 LE_0B.config_data\[7\] vssd1 vssd1 vccd1 vccd1 net353 sky130_fd_sc_hd__dlygate4sd3_1
X_2830_ clknet_leaf_13_clk net388 net226 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[37\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_35_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_1 CBeast_in[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2692_ SB0.route_sel\[92\] SB0.route_sel\[91\] net257 vssd1 vssd1 vccd1 vccd1 _0228_
+ sky130_fd_sc_hd__mux2_1
X_1712_ _0470_ _0471_ _0472_ _0469_ vssd1 vssd1 vccd1 vccd1 _0474_ sky130_fd_sc_hd__o31ai_2
XFILLER_6_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1643_ SB0.route_sel\[11\] SB0.route_sel\[10\] _0404_ vssd1 vssd1 vccd1 vccd1 _0405_
+ sky130_fd_sc_hd__and3_1
X_2761_ CB_1.config_dataA\[9\] net149 net260 vssd1 vssd1 vccd1 vccd1 _0297_ sky130_fd_sc_hd__mux2_1
X_1574_ _1358_ _0334_ vssd1 vssd1 vccd1 vccd1 _0336_ sky130_fd_sc_hd__nor2_1
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1848__A0 net23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2057_ _1163_ SB0.route_sel\[14\] SB0.route_sel\[9\] _1164_ _0814_ vssd1 vssd1 vccd1
+ vccd1 _0815_ sky130_fd_sc_hd__a221o_1
X_2126_ net149 _0883_ CB_1.config_dataA\[10\] vssd1 vssd1 vccd1 vccd1 _0884_ sky130_fd_sc_hd__o21ai_1
XFILLER_19_190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2959_ clknet_leaf_26_clk _0167_ net194 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[31\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_fanout217_X net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2756__S net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput82 net82 vssd1 vssd1 vccd1 vccd1 CBnorth_out[1] sky130_fd_sc_hd__buf_2
Xoutput93 net93 vssd1 vssd1 vccd1 vccd1 SBsouth_out[11] sky130_fd_sc_hd__buf_2
Xoutput71 net71 vssd1 vssd1 vccd1 vccd1 CBeast_out[4] sky130_fd_sc_hd__buf_2
XANTENNA__2098__A3 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2813_ clknet_leaf_1_clk _0021_ net191 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_2744_ net162 CB_0.config_dataB\[11\] net263 vssd1 vssd1 vccd1 vccd1 _0280_ sky130_fd_sc_hd__mux2_1
X_1626_ _0374_ _0375_ _0384_ _0387_ vssd1 vssd1 vccd1 vccd1 _0388_ sky130_fd_sc_hd__a22o_2
X_2675_ SB0.route_sel\[75\] SB0.route_sel\[74\] net235 vssd1 vssd1 vccd1 vccd1 _0211_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__2089__A3 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1488_ _1258_ _1280_ net11 vssd1 vssd1 vccd1 vccd1 _1282_ sky130_fd_sc_hd__a21o_1
X_1557_ net132 _1306_ _1348_ vssd1 vssd1 vccd1 vccd1 _1351_ sky130_fd_sc_hd__or3_1
X_2109_ net151 _0797_ _0852_ _0866_ vssd1 vssd1 vccd1 vccd1 _0867_ sky130_fd_sc_hd__a211o_1
XFILLER_36_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3089_ clknet_leaf_20_clk _0297_ net216 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[9\]
+ sky130_fd_sc_hd__dfstp_2
XTAP_TAPCELL_ROW_52_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1524__A2 _1304_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1827__A3 net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2058__Y _0816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2252__A3 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2460_ _1149_ _1150_ _0534_ vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__o21a_1
X_1411_ SB0.route_sel\[89\] vssd1 vssd1 vccd1 vccd1 _1205_ sky130_fd_sc_hd__inv_2
X_2391_ _1270_ _1104_ vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__and2_2
XANTENNA__1818__A3 _0391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3012_ clknet_leaf_2_clk _0220_ net197 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[84\]
+ sky130_fd_sc_hd__dfstp_1
X_2727_ CB_0.config_dataA\[15\] CB_0.config_dataA\[14\] net265 vssd1 vssd1 vccd1 vccd1
+ _0263_ sky130_fd_sc_hd__mux2_1
X_1609_ CB_0.config_dataA\[19\] CB_0.config_dataA\[18\] _1250_ vssd1 vssd1 vccd1 vccd1
+ _0371_ sky130_fd_sc_hd__or3_1
X_2589_ CB_1.config_dataB\[9\] CB_1.config_dataB\[8\] net266 vssd1 vssd1 vccd1 vccd1
+ _0125_ sky130_fd_sc_hd__mux2_1
X_2658_ SB0.route_sel\[58\] SB0.route_sel\[57\] net256 vssd1 vssd1 vccd1 vccd1 _0194_
+ sky130_fd_sc_hd__mux2_1
Xfanout157 CB_0.config_dataB\[17\] vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__clkbuf_2
Xfanout168 CB_0.config_dataA\[13\] vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__buf_2
Xfanout124 net126 vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__buf_1
XANTENNA__1998__X _0758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout179 CB_1.config_dataB\[13\] vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__buf_2
XANTENNA_input1_A CBeast_in[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout135 _0960_ vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__clkbuf_2
Xfanout146 CB_1.config_dataA\[12\] vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__buf_2
XANTENNA_input57_A config_data_in vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_8_clk_A clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_0_Left_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input12_X net12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1960_ net15 net20 net21 net22 net163 CB_0.config_dataB\[9\] vssd1 vssd1 vccd1 vccd1
+ _0720_ sky130_fd_sc_hd__mux4_1
X_1891_ CB_0.config_dataB\[5\] _1229_ vssd1 vssd1 vccd1 vccd1 _0651_ sky130_fd_sc_hd__nor2_1
X_2443_ SB0.route_sel\[96\] SB0.route_sel\[97\] vssd1 vssd1 vccd1 vccd1 _1139_ sky130_fd_sc_hd__or2_1
X_2512_ LE_0B.dff1_out _1247_ _1151_ vssd1 vssd1 vccd1 vccd1 _0050_ sky130_fd_sc_hd__a21o_1
XFILLER_56_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3087__SET_B net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2374_ _0399_ _1093_ _0400_ vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_62_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1975__A2 _1297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2442__X net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input4_X net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_36_Left_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2090_ _0810_ _0846_ _0847_ _1236_ vssd1 vssd1 vccd1 vccd1 _0848_ sky130_fd_sc_hd__a22o_2
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2992_ clknet_leaf_27_clk _0200_ net194 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[64\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_16_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1874_ _0635_ _0634_ _0572_ vssd1 vssd1 vccd1 vccd1 _0636_ sky130_fd_sc_hd__mux2_1
X_1943_ _0700_ _0702_ vssd1 vssd1 vccd1 vccd1 _0703_ sky130_fd_sc_hd__nand2_2
XANTENNA__1590__B1 net46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2426_ _1161_ SB0.route_sel\[10\] _1162_ SB0.route_sel\[13\] _1127_ vssd1 vssd1 vccd1
+ vccd1 _1128_ sky130_fd_sc_hd__a221o_1
X_2288_ net3 net180 vssd1 vssd1 vccd1 vccd1 _1044_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_39_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2357_ _1305_ _0456_ _0827_ vssd1 vssd1 vccd1 vccd1 _1085_ sky130_fd_sc_hd__a21o_1
XANTENNA__2759__S net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1581__A0 net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1590_ _1208_ _1209_ net46 SB0.route_sel\[101\] SB0.route_sel\[100\] vssd1 vssd1
+ vccd1 vccd1 _0352_ sky130_fd_sc_hd__o2111a_1
XFILLER_7_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2211_ net1 net6 net7 net8 net185 CB_1.config_dataB\[5\] vssd1 vssd1 vccd1 vccd1
+ _0967_ sky130_fd_sc_hd__mux4_1
X_2073_ _0469_ _0830_ vssd1 vssd1 vccd1 vccd1 _0831_ sky130_fd_sc_hd__and2_2
X_2142_ CB_1.config_dataA\[11\] _0888_ _0890_ _0899_ vssd1 vssd1 vccd1 vccd1 _0900_
+ sky130_fd_sc_hd__o211a_1
X_2975_ clknet_leaf_22_clk _0183_ net212 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[47\]
+ sky130_fd_sc_hd__dfstp_1
X_1857_ _0615_ _0617_ _0618_ vssd1 vssd1 vccd1 vccd1 _0619_ sky130_fd_sc_hd__o21a_1
X_1788_ net171 CB_0.config_dataA\[7\] vssd1 vssd1 vccd1 vccd1 _0550_ sky130_fd_sc_hd__or2_1
X_1926_ _0391_ _0447_ _1225_ vssd1 vssd1 vccd1 vccd1 _0686_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout207_A net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1866__A1 net20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2409_ _1115_ _1116_ _1342_ vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__o21a_1
XFILLER_52_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2291__A1 _0838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold82 LEI0.config_data\[32\] vssd1 vssd1 vccd1 vccd1 net354 sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 _0014_ vssd1 vssd1 vccd1 vccd1 net365 sky130_fd_sc_hd__dlygate4sd3_1
Xhold60 LE_0A.config_data\[9\] vssd1 vssd1 vccd1 vccd1 net332 sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 LE_0A.config_data\[15\] vssd1 vssd1 vccd1 vccd1 net343 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_2 net58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1793__A0 net27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2691_ SB0.route_sel\[91\] SB0.route_sel\[90\] net257 vssd1 vssd1 vccd1 vccd1 _0227_
+ sky130_fd_sc_hd__mux2_1
X_1711_ _0470_ _0471_ _0472_ _0469_ vssd1 vssd1 vccd1 vccd1 _0473_ sky130_fd_sc_hd__o31a_2
X_2760_ net148 CB_1.config_dataA\[7\] net262 vssd1 vssd1 vccd1 vccd1 _0296_ sky130_fd_sc_hd__mux2_1
X_1642_ SB0.route_sel\[12\] SB0.route_sel\[13\] net34 vssd1 vssd1 vccd1 vccd1 _0404_
+ sky130_fd_sc_hd__a21bo_1
X_1573_ SB0.route_sel\[104\] SB0.route_sel\[105\] _0332_ _0333_ vssd1 vssd1 vccd1
+ vccd1 _0335_ sky130_fd_sc_hd__a211o_1
XANTENNA__1848__A1 net24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2056_ SB0.route_sel\[12\] SB0.route_sel\[13\] vssd1 vssd1 vccd1 vccd1 _0814_ sky130_fd_sc_hd__nor2_1
X_2125_ CB_1.config_dataA\[9\] CB_1.config_dataA\[11\] vssd1 vssd1 vccd1 vccd1 _0883_
+ sky130_fd_sc_hd__nand2_1
X_1909_ CB_0.config_dataB\[7\] _0668_ vssd1 vssd1 vccd1 vccd1 _0669_ sky130_fd_sc_hd__or2_1
XFILLER_22_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2958_ clknet_leaf_26_clk _0166_ net194 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[30\]
+ sky130_fd_sc_hd__dfstp_1
X_2889_ clknet_leaf_22_clk _0097_ net215 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_32_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput83 net83 vssd1 vssd1 vccd1 vccd1 CBnorth_out[2] sky130_fd_sc_hd__buf_2
XANTENNA_input42_X net42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput94 net94 vssd1 vssd1 vccd1 vccd1 SBsouth_out[12] sky130_fd_sc_hd__buf_2
Xoutput72 net72 vssd1 vssd1 vccd1 vccd1 CBeast_out[5] sky130_fd_sc_hd__buf_2
XFILLER_63_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2743_ CB_0.config_dataB\[11\] CB_0.config_dataB\[10\] net263 vssd1 vssd1 vccd1 vccd1
+ _0279_ sky130_fd_sc_hd__mux2_1
X_2812_ clknet_leaf_3_clk net391 net201 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_16_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1625_ _0382_ _0385_ _0386_ SB0.route_sel\[24\] SB0.route_sel\[25\] vssd1 vssd1 vccd1
+ vccd1 _0387_ sky130_fd_sc_hd__o311a_1
X_2674_ SB0.route_sel\[74\] SB0.route_sel\[73\] net239 vssd1 vssd1 vccd1 vccd1 _0210_
+ sky130_fd_sc_hd__mux2_1
X_1556_ net142 net143 _1308_ vssd1 vssd1 vccd1 vccd1 _1350_ sky130_fd_sc_hd__nand3_1
XANTENNA__2191__A0 _0813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1770__B1_N net30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1487_ net178 net177 vssd1 vssd1 vccd1 vccd1 _1281_ sky130_fd_sc_hd__nand2b_1
X_2039_ _1358_ _0334_ _0796_ vssd1 vssd1 vccd1 vccd1 _0797_ sky130_fd_sc_hd__or3_4
X_2108_ net151 _0803_ vssd1 vssd1 vccd1 vccd1 _0866_ sky130_fd_sc_hd__nor2_1
X_3088_ clknet_leaf_19_clk _0296_ net218 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[8\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_52_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1410_ SB0.route_sel\[92\] vssd1 vssd1 vccd1 vccd1 _1204_ sky130_fd_sc_hd__inv_2
XANTENNA__2090__X _0848_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3011_ clknet_leaf_1_clk _0219_ net196 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[83\]
+ sky130_fd_sc_hd__dfstp_1
X_2390_ SB0.route_sel\[58\] _1188_ _1189_ SB0.route_sel\[61\] _1103_ vssd1 vssd1 vccd1
+ vccd1 _1104_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_8_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2726_ CB_0.config_dataA\[14\] net168 net253 vssd1 vssd1 vccd1 vccd1 _0262_ sky130_fd_sc_hd__mux2_1
Xfanout125 net126 vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__buf_2
X_1608_ LEI0.config_data\[2\] _0369_ vssd1 vssd1 vccd1 vccd1 _0370_ sky130_fd_sc_hd__nand2b_1
X_2588_ net182 net183 net266 vssd1 vssd1 vccd1 vccd1 _0124_ sky130_fd_sc_hd__mux2_1
Xfanout136 net141 vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__buf_2
Xfanout147 CB_1.config_dataA\[12\] vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__dlymetal6s2s_1
X_2657_ SB0.route_sel\[57\] SB0.route_sel\[56\] net255 vssd1 vssd1 vccd1 vccd1 _0193_
+ sky130_fd_sc_hd__mux2_1
X_1539_ net144 net145 vssd1 vssd1 vccd1 vccd1 _1333_ sky130_fd_sc_hd__or2_1
Xfanout158 CB_0.config_dataB\[17\] vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__buf_1
Xfanout169 CB_0.config_dataA\[12\] vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_57_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2155__A0 _0819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_16_Right_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1890_ CB_0.config_dataB\[7\] _0649_ vssd1 vssd1 vccd1 vccd1 _0650_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_25_Right_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2442_ _1138_ _0336_ vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__and2b_1
X_2511_ _0734_ _0764_ _0768_ _0774_ net60 vssd1 vssd1 vccd1 vccd1 _1151_ sky130_fd_sc_hd__o221a_1
X_2373_ _1306_ _0377_ _0816_ vssd1 vssd1 vccd1 vccd1 _1093_ sky130_fd_sc_hd__o21ai_1
XFILLER_56_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_34_Right_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2709_ SB0.route_sel\[109\] SB0.route_sel\[108\] net268 vssd1 vssd1 vccd1 vccd1 _0245_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__1975__A3 _1273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_43_Right_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_52_Right_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_61_Right_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3093__SET_B net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1942_ LEI0.config_data\[5\] _0701_ vssd1 vssd1 vccd1 vccd1 _0702_ sky130_fd_sc_hd__nand2b_2
X_2991_ clknet_leaf_23_clk _0199_ net211 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[63\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1873_ LE_0A.config_data\[1\] LE_0A.config_data\[0\] _0543_ vssd1 vssd1 vccd1 vccd1
+ _0635_ sky130_fd_sc_hd__mux2_1
X_2356_ _0526_ _1084_ _0528_ vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__a21o_1
X_2425_ SB0.route_sel\[9\] SB0.route_sel\[8\] vssd1 vssd1 vccd1 vccd1 _1127_ sky130_fd_sc_hd__nor2_1
XANTENNA__1893__A2 _0492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2287_ _1028_ _1042_ vssd1 vssd1 vccd1 vccd1 _1043_ sky130_fd_sc_hd__nor2_1
XANTENNA__1645__A2 _0397_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout187_A net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_7_clk_A clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2210_ _0827_ _0831_ _0835_ _0838_ _1244_ net184 vssd1 vssd1 vccd1 vccd1 _0966_ sky130_fd_sc_hd__mux4_1
XFILLER_38_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2072_ _1193_ SB0.route_sel\[70\] SB0.route_sel\[65\] _1194_ _0829_ vssd1 vssd1 vccd1
+ vccd1 _0830_ sky130_fd_sc_hd__a221o_1
XFILLER_19_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2141_ _0896_ _0898_ vssd1 vssd1 vccd1 vccd1 _0899_ sky130_fd_sc_hd__nor2_1
X_1925_ net15 net20 net21 net22 net167 net166 vssd1 vssd1 vccd1 vccd1 _0685_ sky130_fd_sc_hd__mux4_1
X_2974_ clknet_leaf_23_clk _0182_ net212 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[46\]
+ sky130_fd_sc_hd__dfstp_1
X_1787_ net21 _0545_ _0546_ net22 vssd1 vssd1 vccd1 vccd1 _0549_ sky130_fd_sc_hd__o22a_1
X_1856_ _1297_ _0608_ _0609_ _1273_ vssd1 vssd1 vccd1 vccd1 _0618_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_55_Left_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2339_ net124 _1345_ _1323_ vssd1 vssd1 vccd1 vccd1 _1076_ sky130_fd_sc_hd__mux2_1
XANTENNA__1866__A2 net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2448__X net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2107__A3 _0781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_2_Right_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2408_ SB0.route_sel\[36\] _1176_ SB0.route_sel\[33\] SB0.route_sel\[32\] vssd1 vssd1
+ vccd1 vccd1 _1116_ sky130_fd_sc_hd__o22ai_1
XTAP_TAPCELL_ROW_10_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold83 _0033_ vssd1 vssd1 vccd1 vccd1 net355 sky130_fd_sc_hd__dlygate4sd3_1
Xhold50 LE_0A.config_data\[8\] vssd1 vssd1 vccd1 vccd1 net322 sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 LE_1A.config_data\[11\] vssd1 vssd1 vccd1 vccd1 net333 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_output119_A net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input32_A SBsouth_in[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold94 LE_1B.config_data\[15\] vssd1 vssd1 vccd1 vccd1 net366 sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 LE_1B.config_data\[6\] vssd1 vssd1 vccd1 vccd1 net344 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_31_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2534__A net60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1572_ SB0.route_sel\[104\] SB0.route_sel\[105\] _0332_ _0333_ vssd1 vssd1 vccd1
+ vccd1 _0334_ sky130_fd_sc_hd__a211oi_2
XANTENNA__1793__A1 net28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2690_ SB0.route_sel\[90\] SB0.route_sel\[89\] net241 vssd1 vssd1 vccd1 vccd1 _0226_
+ sky130_fd_sc_hd__mux2_1
X_1710_ _1192_ SB0.route_sel\[69\] vssd1 vssd1 vccd1 vccd1 _0472_ sky130_fd_sc_hd__nor2_1
X_1641_ SB0.route_sel\[15\] SB0.route_sel\[14\] _0402_ vssd1 vssd1 vccd1 vccd1 _0403_
+ sky130_fd_sc_hd__a21bo_1
XANTENNA_3 net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1848__A2 net25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2124_ CB_1.config_dataA\[11\] _0880_ _0881_ _0877_ vssd1 vssd1 vccd1 vccd1 _0882_
+ sky130_fd_sc_hd__o22ai_1
X_2055_ _0388_ _0812_ vssd1 vssd1 vccd1 vccd1 _0813_ sky130_fd_sc_hd__nand2_2
X_1839_ _0582_ _0585_ _0590_ _1219_ vssd1 vssd1 vccd1 vccd1 _0601_ sky130_fd_sc_hd__o31a_1
X_1908_ net23 net24 net25 net26 net165 CB_0.config_dataB\[5\] vssd1 vssd1 vccd1 vccd1
+ _0668_ sky130_fd_sc_hd__mux4_1
XFILLER_22_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2888_ clknet_leaf_21_clk _0096_ net215 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_2957_ clknet_leaf_27_clk _0165_ net194 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[29\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__2887__Q LE_1A.config_data\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput84 net84 vssd1 vssd1 vccd1 vccd1 CBnorth_out[3] sky130_fd_sc_hd__buf_2
Xoutput95 net95 vssd1 vssd1 vccd1 vccd1 SBsouth_out[13] sky130_fd_sc_hd__buf_2
XANTENNA_input35_X net35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput73 net73 vssd1 vssd1 vccd1 vccd1 CBeast_out[6] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_46_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_28_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2742_ CB_0.config_dataB\[10\] CB_0.config_dataB\[9\] net252 vssd1 vssd1 vccd1 vccd1
+ _0278_ sky130_fd_sc_hd__mux2_1
X_2811_ clknet_leaf_3_clk _0019_ net201 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2191__A1 _0816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1624_ SB0.route_sel\[28\] SB0.route_sel\[29\] net36 vssd1 vssd1 vccd1 vccd1 _0386_
+ sky130_fd_sc_hd__a21boi_1
X_2673_ SB0.route_sel\[73\] SB0.route_sel\[72\] net239 vssd1 vssd1 vccd1 vccd1 _0209_
+ sky130_fd_sc_hd__mux2_1
X_1555_ net175 net176 _1305_ net5 vssd1 vssd1 vccd1 vccd1 _1349_ sky130_fd_sc_hd__a31o_1
XFILLER_39_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2107_ _0792_ _0788_ _0784_ _0781_ CB_1.config_dataA\[1\] net151 vssd1 vssd1 vccd1
+ vccd1 _0865_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_19_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_clk
+ sky130_fd_sc_hd__clkbuf_8
X_3087_ clknet_leaf_18_clk _0295_ net218 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[7\]
+ sky130_fd_sc_hd__dfstp_2
X_1486_ CB_1.config_dataB\[16\] net177 vssd1 vssd1 vccd1 vccd1 _1280_ sky130_fd_sc_hd__and2b_1
XANTENNA_fanout267_A net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2038_ _0795_ vssd1 vssd1 vccd1 vccd1 _0796_ sky130_fd_sc_hd__inv_2
XANTENNA__1524__Y _1318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3010_ clknet_leaf_2_clk _0218_ net208 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[82\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_8_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_8_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2725_ net168 CB_0.config_dataA\[12\] net253 vssd1 vssd1 vccd1 vccd1 _0261_ sky130_fd_sc_hd__mux2_1
X_2656_ SB0.route_sel\[56\] SB0.route_sel\[55\] net258 vssd1 vssd1 vccd1 vccd1 _0192_
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout126 net127 vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout159 CB_0.config_dataB\[16\] vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__clkbuf_2
Xfanout137 net140 vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__clkbuf_2
X_1607_ net136 net122 net130 net134 LEI0.config_data\[0\] LEI0.config_data\[1\] vssd1
+ vssd1 vccd1 vccd1 _0369_ sky130_fd_sc_hd__mux4_1
X_2587_ net183 CB_1.config_dataB\[6\] net264 vssd1 vssd1 vccd1 vccd1 _0123_ sky130_fd_sc_hd__mux2_1
Xfanout148 net149 vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__buf_2
X_1469_ net132 _1257_ _1259_ _1261_ _1262_ vssd1 vssd1 vccd1 vccd1 _1263_ sky130_fd_sc_hd__o32a_1
X_1538_ net144 net145 vssd1 vssd1 vccd1 vccd1 _1332_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_57_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2155__A1 _0822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3053__SET_B net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2091__A0 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output101_A net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2510_ LE_0A.dff0_out _0645_ net60 vssd1 vssd1 vccd1 vccd1 _0049_ sky130_fd_sc_hd__mux2_1
X_2441_ net119 SB0.route_sel\[110\] _1213_ SB0.route_sel\[105\] _1137_ vssd1 vssd1
+ vccd1 vccd1 _1138_ sky130_fd_sc_hd__o221a_1
X_2372_ _0437_ _1092_ _0439_ vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__a21o_1
XANTENNA__1657__B1 net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2082__A0 net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout132_A net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2708_ SB0.route_sel\[108\] SB0.route_sel\[107\] net268 vssd1 vssd1 vccd1 vccd1 _0244_
+ sky130_fd_sc_hd__mux2_1
X_2639_ SB0.route_sel\[39\] SB0.route_sel\[38\] net241 vssd1 vssd1 vccd1 vccd1 _0175_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__2598__S net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1896__A0 net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input62_A nrst vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1872_ LE_0A.config_data\[3\] LE_0A.config_data\[2\] _0543_ vssd1 vssd1 vccd1 vccd1
+ _0634_ sky130_fd_sc_hd__mux2_1
X_1941_ net136 net127 net130 net134 LEI0.config_data\[3\] LEI0.config_data\[4\] vssd1
+ vssd1 vccd1 vccd1 _0701_ sky130_fd_sc_hd__mux4_1
X_2990_ clknet_leaf_23_clk _0198_ net211 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[62\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_14_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2286_ net13 net14 net180 vssd1 vssd1 vccd1 vccd1 _1042_ sky130_fd_sc_hd__mux2_1
X_2355_ _1280_ _0456_ _0838_ vssd1 vssd1 vccd1 vccd1 _1084_ sky130_fd_sc_hd__a21o_1
X_2424_ _1125_ _1126_ _0444_ vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__o21a_1
XFILLER_37_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire121 _0411_ vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__clkbuf_2
X_2140_ net148 _0838_ _0897_ CB_1.config_dataA\[11\] CB_1.config_dataA\[9\] vssd1
+ vssd1 vccd1 vccd1 _0898_ sky130_fd_sc_hd__o2111a_1
XFILLER_34_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1442__Y _1236_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2071_ SB0.route_sel\[68\] SB0.route_sel\[69\] vssd1 vssd1 vccd1 vccd1 _0829_ sky130_fd_sc_hd__nor2_1
X_1855_ net168 _0616_ CB_0.config_dataA\[15\] vssd1 vssd1 vccd1 vccd1 _0617_ sky130_fd_sc_hd__o21ba_1
X_1924_ net121 _0430_ _1225_ vssd1 vssd1 vccd1 vccd1 _0684_ sky130_fd_sc_hd__mux2_1
X_2973_ clknet_leaf_22_clk _0181_ net212 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[45\]
+ sky130_fd_sc_hd__dfstp_1
X_1786_ _0544_ _0547_ net171 vssd1 vssd1 vccd1 vccd1 _0548_ sky130_fd_sc_hd__mux2_1
X_2338_ net139 _1075_ _1299_ vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__mux2_1
XANTENNA__1866__A3 net22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2407_ SB0.route_sel\[35\] SB0.route_sel\[34\] vssd1 vssd1 vccd1 vccd1 _1115_ sky130_fd_sc_hd__and2b_1
X_2269_ _0987_ _1023_ _1024_ vssd1 vssd1 vccd1 vccd1 _1025_ sky130_fd_sc_hd__o21ai_1
XFILLER_37_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1527__Y _1321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold40 _0079_ vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_43_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input25_A CBnorth_in[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold95 LEI0.config_data\[21\] vssd1 vssd1 vccd1 vccd1 net367 sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 LE_1B.config_data\[0\] vssd1 vssd1 vccd1 vccd1 net356 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 LE_1A.config_data\[13\] vssd1 vssd1 vccd1 vccd1 net323 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 _0106_ vssd1 vssd1 vccd1 vccd1 net334 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_16_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold73 _0314_ vssd1 vssd1 vccd1 vccd1 net345 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2534__B _0934_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1571_ CB_0.config_dataA\[19\] CB_0.config_dataA\[18\] net138 _1298_ vssd1 vssd1
+ vccd1 vccd1 _0333_ sky130_fd_sc_hd__and4_1
X_1640_ SB0.route_sel\[12\] SB0.route_sel\[13\] net48 vssd1 vssd1 vccd1 vccd1 _0402_
+ sky130_fd_sc_hd__and3_1
XFILLER_6_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_4 net75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1848__A3 net26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_6_clk_A clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2123_ net4 net5 net148 vssd1 vssd1 vccd1 vccd1 _0881_ sky130_fd_sc_hd__mux2_1
X_2054_ _1173_ SB0.route_sel\[30\] SB0.route_sel\[25\] _1175_ _0811_ vssd1 vssd1 vccd1
+ vccd1 _0812_ sky130_fd_sc_hd__a221o_1
X_1838_ _0598_ _0599_ _0593_ vssd1 vssd1 vccd1 vccd1 _0600_ sky130_fd_sc_hd__a21o_1
X_1907_ _0356_ _0358_ CB_0.config_dataB\[4\] vssd1 vssd1 vccd1 vccd1 _0667_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_32_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2956_ clknet_leaf_27_clk _0164_ net194 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[28\]
+ sky130_fd_sc_hd__dfstp_1
X_2887_ clknet_leaf_29_clk _0095_ net186 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__2497__A0 LEI0.config_data\[35\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1769_ SB0.route_sel\[87\] SB0.route_sel\[86\] _0530_ vssd1 vssd1 vccd1 vccd1 _0531_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_25_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput85 net85 vssd1 vssd1 vccd1 vccd1 CBnorth_out[4] sky130_fd_sc_hd__buf_2
XANTENNA_input28_X net28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput63 net63 vssd1 vssd1 vccd1 vccd1 CBeast_out[0] sky130_fd_sc_hd__buf_2
Xoutput96 net96 vssd1 vssd1 vccd1 vccd1 SBsouth_out[1] sky130_fd_sc_hd__buf_2
Xoutput74 net74 vssd1 vssd1 vccd1 vccd1 CBeast_out[7] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_46_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2810_ clknet_leaf_3_clk _0018_ net202 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_2741_ CB_0.config_dataB\[9\] net163 net252 vssd1 vssd1 vccd1 vccd1 _0277_ sky130_fd_sc_hd__mux2_1
XANTENNA__2412__B1 _1342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2672_ SB0.route_sel\[72\] SB0.route_sel\[71\] net239 vssd1 vssd1 vccd1 vccd1 _0208_
+ sky130_fd_sc_hd__mux2_1
X_1485_ net139 _1277_ _1275_ vssd1 vssd1 vccd1 vccd1 _1279_ sky130_fd_sc_hd__mux2_1
XANTENNA__2191__A2 _0822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1623_ _1173_ _1174_ net50 SB0.route_sel\[29\] SB0.route_sel\[28\] vssd1 vssd1 vccd1
+ vccd1 _0385_ sky130_fd_sc_hd__o2111a_1
X_1554_ net175 net176 vssd1 vssd1 vccd1 vccd1 _1348_ sky130_fd_sc_hd__nand2_1
.ends

