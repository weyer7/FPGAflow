* NGSPICE file created from fpgacell.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s4s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s4s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_1 abstract view
.subckt sky130_fd_sc_hd__clkinv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_4 abstract view
.subckt sky130_fd_sc_hd__o21ba_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_2 abstract view
.subckt sky130_fd_sc_hd__o32ai_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_4 abstract view
.subckt sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd1_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

.subckt fpgacell CBeast_in[0] CBeast_in[10] CBeast_in[11] CBeast_in[12] CBeast_in[13]
+ CBeast_in[14] CBeast_in[15] CBeast_in[1] CBeast_in[2] CBeast_in[3] CBeast_in[4]
+ CBeast_in[5] CBeast_in[6] CBeast_in[7] CBeast_in[8] CBeast_in[9] CBeast_out[0] CBeast_out[10]
+ CBeast_out[11] CBeast_out[12] CBeast_out[13] CBeast_out[14] CBeast_out[15] CBeast_out[1]
+ CBeast_out[2] CBeast_out[3] CBeast_out[4] CBeast_out[5] CBeast_out[6] CBeast_out[7]
+ CBeast_out[8] CBeast_out[9] CBnorth_in[0] CBnorth_in[10] CBnorth_in[11] CBnorth_in[12]
+ CBnorth_in[13] CBnorth_in[14] CBnorth_in[15] CBnorth_in[1] CBnorth_in[2] CBnorth_in[3]
+ CBnorth_in[4] CBnorth_in[5] CBnorth_in[6] CBnorth_in[7] CBnorth_in[8] CBnorth_in[9]
+ CBnorth_out[0] CBnorth_out[10] CBnorth_out[11] CBnorth_out[12] CBnorth_out[13] CBnorth_out[14]
+ CBnorth_out[15] CBnorth_out[1] CBnorth_out[2] CBnorth_out[3] CBnorth_out[4] CBnorth_out[5]
+ CBnorth_out[6] CBnorth_out[7] CBnorth_out[8] CBnorth_out[9] SBsouth_in[0] SBsouth_in[10]
+ SBsouth_in[11] SBsouth_in[12] SBsouth_in[13] SBsouth_in[14] SBsouth_in[15] SBsouth_in[1]
+ SBsouth_in[2] SBsouth_in[3] SBsouth_in[4] SBsouth_in[5] SBsouth_in[6] SBsouth_in[7]
+ SBsouth_in[8] SBsouth_in[9] SBsouth_out[0] SBsouth_out[10] SBsouth_out[11] SBsouth_out[12]
+ SBsouth_out[13] SBsouth_out[14] SBsouth_out[15] SBsouth_out[1] SBsouth_out[2] SBsouth_out[3]
+ SBsouth_out[4] SBsouth_out[5] SBsouth_out[6] SBsouth_out[7] SBsouth_out[8] SBsouth_out[9]
+ SBwest_in[0] SBwest_in[10] SBwest_in[11] SBwest_in[12] SBwest_in[13] SBwest_in[14]
+ SBwest_in[15] SBwest_in[1] SBwest_in[2] SBwest_in[3] SBwest_in[4] SBwest_in[5] SBwest_in[6]
+ SBwest_in[7] SBwest_in[8] SBwest_in[9] SBwest_out[0] SBwest_out[10] SBwest_out[11]
+ SBwest_out[12] SBwest_out[13] SBwest_out[14] SBwest_out[15] SBwest_out[1] SBwest_out[2]
+ SBwest_out[3] SBwest_out[4] SBwest_out[5] SBwest_out[6] SBwest_out[7] SBwest_out[8]
+ SBwest_out[9] clk config_data_in config_data_out config_en en le_clk le_en le_nrst
+ nrst vccd1 vssd1
XFILLER_54_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2106_ CB_1.config_dataB\[12\] _0735_ vssd1 vssd1 vccd1 vccd1 _0736_ sky130_fd_sc_hd__nand2_1
X_3086_ SB0.route_sel\[126\] SB0.route_sel\[125\] net298 vssd1 vssd1 vccd1 vccd1 _0254_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_37_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2037_ net165 net161 net15 vssd1 vssd1 vccd1 vccd1 _0667_ sky130_fd_sc_hd__o21ai_1
X_3155_ net170 CB_1.config_dataA\[17\] net222 vssd1 vssd1 vccd1 vccd1 _0323_ sky130_fd_sc_hd__mux2_1
X_2939_ CB_1.config_dataB\[3\] CB_1.config_dataB\[4\] net225 vssd1 vssd1 vccd1 vccd1
+ _0107_ sky130_fd_sc_hd__mux2_1
XANTENNA__2954__A1 CB_1.config_dataB\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_15_Left_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2182__A2 net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2642__A0 _0956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2237__A3 _0865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2158__C1 _0755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1684__A1 _1521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2228__A3 net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3301__SET_B net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2655_ _1280_ _1281_ net146 vssd1 vssd1 vccd1 vccd1 _1282_ sky130_fd_sc_hd__o21ba_1
XANTENNA_clone35_B1 _0470_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1606_ SB0.route_sel\[11\] vssd1 vssd1 vccd1 vccd1 _1444_ sky130_fd_sc_hd__inv_2
XFILLER_8_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2724_ SB0.route_sel\[34\] _1432_ SB0.route_sel\[37\] _1433_ _1331_ vssd1 vssd1 vccd1
+ vccd1 _1332_ sky130_fd_sc_hd__a221o_1
XANTENNA__3113__A1 CB_0.config_dataB\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2586_ LE_0A.config_data\[7\] LE_0A.config_data\[6\] _1180_ vssd1 vssd1 vccd1 vccd1
+ _1213_ sky130_fd_sc_hd__mux2_1
X_3207_ clknet_leaf_5_clk _0027_ net256 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clone51_C1 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout149 net150 vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__buf_8
XANTENNA__2737__X net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3138_ CB_0.config_dataB\[24\] CB_1.config_dataA\[0\] net230 vssd1 vssd1 vccd1 vccd1
+ _0306_ sky130_fd_sc_hd__mux2_1
X_3069_ SB0.route_sel\[109\] SB0.route_sel\[108\] net300 vssd1 vssd1 vccd1 vccd1 _0237_
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold170 LEI0.config_data\[29\] vssd1 vssd1 vccd1 vccd1 net480 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_0_Left_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_31_clk_A clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2440_ net142 net155 LEI0.config_data\[27\] vssd1 vssd1 vccd1 vccd1 _1068_ sky130_fd_sc_hd__mux2_1
X_2371_ SB0.route_sel\[70\] SB0.route_sel\[71\] vssd1 vssd1 vccd1 vccd1 _0999_ sky130_fd_sc_hd__nand2b_1
XANTENNA__2449__A3 net26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clone46_C1 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2638_ net31 net32 net18 net19 net187 net186 vssd1 vssd1 vccd1 vccd1 _1265_ sky130_fd_sc_hd__mux4_1
X_2569_ _0991_ _0994_ net191 vssd1 vssd1 vccd1 vccd1 _1196_ sky130_fd_sc_hd__mux2_1
X_2707_ _1320_ _1549_ vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__and2_4
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_36_Left_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_45_Left_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input55_A SBwest_in[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1940_ SB0.route_sel\[104\] SB0.route_sel\[105\] _0569_ _0568_ vssd1 vssd1 vccd1
+ vccd1 _0570_ sky130_fd_sc_hd__a211o_4
X_1871_ CB_0.config_dataA\[23\] CB_0.config_dataA\[22\] vssd1 vssd1 vccd1 vccd1 _0501_
+ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_54_Left_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3472_ clknet_leaf_4_clk _0292_ net262 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[11\]
+ sky130_fd_sc_hd__dfstp_1
X_2423_ _0956_ net339 CB_0.config_dataB\[5\] vssd1 vssd1 vccd1 vccd1 _1051_ sky130_fd_sc_hd__mux2_1
XANTENNA_clone32_A1 _0393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_63_Left_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2354_ _0367_ _0358_ _0981_ net305 vssd1 vssd1 vccd1 vccd1 _0982_ sky130_fd_sc_hd__a211o_4
X_2285_ net171 net170 vssd1 vssd1 vccd1 vccd1 _0914_ sky130_fd_sc_hd__nor2_2
XFILLER_64_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2358__A2 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input2_X net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2294__A1 net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2597__A2 net25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input58_X net58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2070_ net198 _0698_ _0699_ vssd1 vssd1 vccd1 vccd1 _0700_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_3_Left_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_64_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2972_ SB0.route_sel\[12\] SB0.route_sel\[11\] net292 vssd1 vssd1 vccd1 vccd1 _0140_
+ sky130_fd_sc_hd__mux2_1
X_1854_ CB_0.config_dataA\[23\] CB_0.config_dataA\[22\] _0363_ vssd1 vssd1 vccd1 vccd1
+ _0484_ sky130_fd_sc_hd__or3_1
X_1923_ SB0.route_sel\[98\] SB0.route_sel\[99\] vssd1 vssd1 vccd1 vccd1 _0553_ sky130_fd_sc_hd__nand2_1
X_1785_ _0404_ _0410_ _0414_ SB0.route_sel\[16\] SB0.route_sel\[17\] vssd1 vssd1 vccd1
+ vccd1 _0415_ sky130_fd_sc_hd__o2111ai_2
X_3455_ clknet_leaf_10_clk _0275_ net263 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[19\]
+ sky130_fd_sc_hd__dfstp_1
X_2406_ LEI0.config_data\[15\] net147 _1033_ LEI0.config_data\[16\] vssd1 vssd1 vccd1
+ vccd1 _1034_ sky130_fd_sc_hd__o211a_1
X_3386_ clknet_leaf_4_clk _0206_ net252 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[78\]
+ sky130_fd_sc_hd__dfstp_1
X_3524_ clknet_leaf_0_clk _0344_ net241 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_2199_ _0820_ _0824_ _0827_ CB_1.config_dataA\[4\] vssd1 vssd1 vccd1 vccd1 _0828_
+ sky130_fd_sc_hd__a31o_1
XFILLER_25_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2268_ _1462_ _0886_ _0896_ _0874_ vssd1 vssd1 vccd1 vccd1 _0897_ sky130_fd_sc_hd__a31o_1
X_2337_ SB0.route_sel\[2\] SB0.route_sel\[3\] SB0.route_sel\[5\] _1449_ _0964_ vssd1
+ vssd1 vccd1 vccd1 _0965_ sky130_fd_sc_hd__o221a_1
XANTENNA__2276__A1 _0829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1808__Y _0438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold74 LE_0A.config_data\[11\] vssd1 vssd1 vccd1 vccd1 net384 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1711__B1 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input18_A CBnorth_in[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold85 _0074_ vssd1 vssd1 vccd1 vccd1 net395 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2019__A1 _0643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold96 LE_1B.config_data\[6\] vssd1 vssd1 vccd1 vccd1 net406 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2390__X _1018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3240_ clknet_leaf_7_clk _0060_ net255 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__3435__Q net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1570_ SB0.route_sel\[83\] vssd1 vssd1 vccd1 vccd1 _1408_ sky130_fd_sc_hd__inv_2
XANTENNA_5 _0338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2122_ net196 _0750_ _0751_ vssd1 vssd1 vccd1 vccd1 _0752_ sky130_fd_sc_hd__a21o_1
X_2053_ _0682_ _0494_ _1496_ vssd1 vssd1 vccd1 vccd1 _0683_ sky130_fd_sc_hd__a21bo_4
XANTENNA__2258__A1 _0449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3171_ net413 LE_1B.config_data\[8\] net202 vssd1 vssd1 vccd1 vccd1 _0339_ sky130_fd_sc_hd__mux2_1
XANTENNA__1909__X _0539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2955_ CB_1.config_dataB\[19\] CB_1.config_dataB\[20\] net223 vssd1 vssd1 vccd1 vccd1
+ _0123_ sky130_fd_sc_hd__mux2_1
X_2886_ net410 net383 net218 vssd1 vssd1 vccd1 vccd1 _0055_ sky130_fd_sc_hd__mux2_1
X_1906_ _1514_ _0501_ vssd1 vssd1 vccd1 vccd1 _0536_ sky130_fd_sc_hd__or2_1
X_1837_ _0466_ _0465_ _0460_ vssd1 vssd1 vccd1 vccd1 _0467_ sky130_fd_sc_hd__or3b_4
XANTENNA__2430__B2 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2430__A1 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1768_ net201 net200 vssd1 vssd1 vccd1 vccd1 _0398_ sky130_fd_sc_hd__nor2_1
X_3507_ clknet_leaf_23_clk _0327_ net274 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[21\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_fanout205_A net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2497__A1 net28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3438_ clknet_leaf_8_clk _0258_ net259 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[2\]
+ sky130_fd_sc_hd__dfstp_2
X_3369_ clknet_leaf_24_clk _0189_ net272 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[61\]
+ sky130_fd_sc_hd__dfstp_1
X_1699_ net46 _1535_ _1536_ vssd1 vssd1 vccd1 vccd1 _1537_ sky130_fd_sc_hd__a21oi_1
XANTENNA__1819__X _0449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput75 net75 vssd1 vssd1 vccd1 vccd1 CBeast_out[12] sky130_fd_sc_hd__buf_6
Xoutput97 net97 vssd1 vssd1 vccd1 vccd1 CBnorth_out[3] sky130_fd_sc_hd__buf_6
XANTENNA__2385__X _1013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output124_A net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput86 net86 vssd1 vssd1 vccd1 vccd1 CBeast_out[8] sky130_fd_sc_hd__buf_6
XFILLER_16_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2671_ _1296_ _0581_ vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__and2_4
X_1622_ CB_1.config_dataA\[9\] vssd1 vssd1 vccd1 vccd1 _1460_ sky130_fd_sc_hd__inv_2
X_2740_ _0425_ _1342_ vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__and2_1
XANTENNA_clone40_A1 _0562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout309 net310 vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__clkbuf_4
X_3223_ clknet_leaf_28_clk _0043_ net248 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[43\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_54_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2105_ net4 net6 net5 net7 net196 net197 vssd1 vssd1 vccd1 vccd1 _0735_ sky130_fd_sc_hd__mux4_1
X_3085_ SB0.route_sel\[125\] SB0.route_sel\[124\] net298 vssd1 vssd1 vccd1 vccd1 _0253_
+ sky130_fd_sc_hd__mux2_1
X_2036_ SB0.route_sel\[66\] SB0.route_sel\[67\] vssd1 vssd1 vccd1 vccd1 _0666_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_37_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clone49_C1 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3154_ net171 net170 net222 vssd1 vssd1 vccd1 vccd1 _0322_ sky130_fd_sc_hd__mux2_1
X_2938_ CB_1.config_dataB\[2\] CB_1.config_dataB\[3\] net225 vssd1 vssd1 vccd1 vccd1
+ _0106_ sky130_fd_sc_hd__mux2_1
XFILLER_22_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout155_A CB_0.le_outB vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2182__A3 net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2869_ net472 LEI0.config_data\[38\] net214 vssd1 vssd1 vccd1 vccd1 _0038_ sky130_fd_sc_hd__mux2_1
XANTENNA__2642__A1 _0959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrebuffer8 _0580_ vssd1 vssd1 vccd1 vccd1 net318 sky130_fd_sc_hd__dlymetal6s4s_1
XANTENNA_clkbuf_leaf_5_clk_A clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1905__B1 net22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1841__C1 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2723_ SB0.route_sel\[33\] SB0.route_sel\[32\] vssd1 vssd1 vccd1 vccd1 _1331_ sky130_fd_sc_hd__nor2_1
X_2654_ LEI0.config_data\[38\] net234 vssd1 vssd1 vccd1 vccd1 _1281_ sky130_fd_sc_hd__nand2_1
X_2585_ LEI0.config_data\[14\] net234 _1210_ _1185_ vssd1 vssd1 vccd1 vccd1 _1212_
+ sky130_fd_sc_hd__a31o_1
XANTENNA_clone35_A1 _0467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1605_ SB0.route_sel\[10\] vssd1 vssd1 vccd1 vccd1 _1443_ sky130_fd_sc_hd__inv_2
X_3137_ CB_0.config_dataB\[23\] CB_0.config_dataB\[24\] net227 vssd1 vssd1 vccd1 vccd1
+ _0305_ sky130_fd_sc_hd__mux2_1
X_3206_ clknet_leaf_5_clk _0026_ net256 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__1922__X _0552_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clone51_B1 _0370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3068_ SB0.route_sel\[108\] SB0.route_sel\[107\] net300 vssd1 vssd1 vccd1 vccd1 _0236_
+ sky130_fd_sc_hd__mux2_1
XFILLER_35_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2019_ _0643_ _0639_ _0647_ _0648_ vssd1 vssd1 vccd1 vccd1 _0649_ sky130_fd_sc_hd__a211o_1
Xhold171 LEI0.config_data\[28\] vssd1 vssd1 vccd1 vccd1 net481 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2818__B1_N _0371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold160 LE_1B.config_data\[3\] vssd1 vssd1 vccd1 vccd1 net470 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2538__S1 CB_0.config_dataA\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clone33_X net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1969__A3 net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3146__S net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2370_ _0655_ _0649_ _0997_ net307 vssd1 vssd1 vccd1 vccd1 _0998_ sky130_fd_sc_hd__a211o_4
XANTENNA__2606__A1 _1021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2606__B2 _1018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2706_ SB0.route_sel\[58\] _1420_ SB0.route_sel\[61\] _1421_ _1319_ vssd1 vssd1 vccd1
+ vccd1 _1320_ sky130_fd_sc_hd__a221o_1
X_2499_ _1125_ _1126_ _1469_ vssd1 vssd1 vccd1 vccd1 _1127_ sky130_fd_sc_hd__mux2_1
X_2637_ _1021_ _1259_ _1260_ _1018_ _1476_ vssd1 vssd1 vccd1 vccd1 _1264_ sky130_fd_sc_hd__a221o_1
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2568_ _1193_ _1194_ _1472_ vssd1 vssd1 vccd1 vccd1 _1195_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_12_Right_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_21_Right_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2376__A3 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_30_Right_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input48_A SBsouth_in[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2049__C1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2393__X _1021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1737__X _0367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1870_ _1541_ _0498_ net23 vssd1 vssd1 vccd1 vccd1 _0500_ sky130_fd_sc_hd__o21ai_1
XFILLER_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2422_ _1042_ _1045_ _1049_ CB_0.config_dataB\[8\] vssd1 vssd1 vccd1 vccd1 _1050_
+ sky130_fd_sc_hd__or4b_1
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3471_ clknet_leaf_4_clk _0291_ net261 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[10\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_clone32_A2 _0384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2353_ SB0.route_sel\[42\] SB0.route_sel\[43\] SB0.route_sel\[45\] _1429_ _0980_
+ vssd1 vssd1 vccd1 vccd1 _0981_ sky130_fd_sc_hd__o221a_1
X_2284_ net171 _0543_ net170 vssd1 vssd1 vccd1 vccd1 _0913_ sky130_fd_sc_hd__o21a_1
XFILLER_64_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1999_ _1518_ _0604_ net18 vssd1 vssd1 vccd1 vccd1 _0629_ sky130_fd_sc_hd__o21ai_1
XANTENNA_clkbuf_leaf_30_clk_A clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2597__A3 net26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2046__A2 _0665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1922_ SB0.route_sel\[96\] SB0.route_sel\[97\] _0550_ _0551_ vssd1 vssd1 vccd1 vccd1
+ _0552_ sky130_fd_sc_hd__a211o_4
XTAP_TAPCELL_ROW_29_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2283__B _0521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2971_ SB0.route_sel\[11\] SB0.route_sel\[10\] net292 vssd1 vssd1 vccd1 vccd1 _0139_
+ sky130_fd_sc_hd__mux2_1
X_1853_ _0360_ _0417_ net24 vssd1 vssd1 vccd1 vccd1 _0483_ sky130_fd_sc_hd__o21ai_1
X_1784_ SB0.route_sel\[21\] SB0.route_sel\[20\] net57 _0411_ _0413_ vssd1 vssd1 vccd1
+ vccd1 _0414_ sky130_fd_sc_hd__a41o_1
X_3523_ clknet_leaf_32_clk net428 net241 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_3454_ clknet_leaf_10_clk _0274_ net263 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[18\]
+ sky130_fd_sc_hd__dfstp_1
X_2405_ LEI0.config_data\[15\] net160 vssd1 vssd1 vccd1 vccd1 _1033_ sky130_fd_sc_hd__nand2_1
X_3385_ clknet_leaf_4_clk _0205_ net261 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[77\]
+ sky130_fd_sc_hd__dfstp_1
X_2336_ SB0.route_sel\[6\] SB0.route_sel\[7\] vssd1 vssd1 vccd1 vccd1 _0964_ sky130_fd_sc_hd__nand2b_1
XANTENNA_fanout185_A CB_0.config_dataB\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2198_ net176 _0825_ _0826_ vssd1 vssd1 vccd1 vccd1 _0827_ sky130_fd_sc_hd__a21o_1
XFILLER_25_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2267_ CB_1.config_dataA\[13\] _0889_ _0892_ _0895_ vssd1 vssd1 vccd1 vccd1 _0896_
+ sky130_fd_sc_hd__or4_1
XANTENNA_fanout238_X net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold75 _0061_ vssd1 vssd1 vccd1 vccd1 net385 sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 LE_0B.config_data\[3\] vssd1 vssd1 vccd1 vccd1 net396 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1840__X _0470_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold97 _0338_ vssd1 vssd1 vccd1 vccd1 net407 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1711__A1 _1548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2671__X net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_6 _0424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3170_ net406 LE_1B.config_data\[7\] net202 vssd1 vssd1 vccd1 vccd1 _0338_ sky130_fd_sc_hd__mux2_1
X_2121_ net359 _0729_ _0733_ net345 CB_1.config_dataB\[12\] vssd1 vssd1 vccd1 vccd1
+ _0751_ sky130_fd_sc_hd__a221o_1
XFILLER_34_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2052_ _0589_ _0681_ CB_1.config_dataB\[4\] vssd1 vssd1 vccd1 vccd1 _0682_ sky130_fd_sc_hd__a21oi_1
X_1905_ _1518_ _0498_ net22 vssd1 vssd1 vccd1 vccd1 _0535_ sky130_fd_sc_hd__o21ai_1
X_2885_ net456 net410 net218 vssd1 vssd1 vccd1 vccd1 _0054_ sky130_fd_sc_hd__mux2_1
XANTENNA_clone38_A1 _0675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2954_ CB_1.config_dataB\[18\] CB_1.config_dataB\[19\] net224 vssd1 vssd1 vccd1 vccd1
+ _0122_ sky130_fd_sc_hd__mux2_1
X_1836_ net144 _0464_ net237 vssd1 vssd1 vccd1 vccd1 _0466_ sky130_fd_sc_hd__o21ai_1
X_3506_ clknet_leaf_24_clk _0326_ net272 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[20\]
+ sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_6_Right_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1698_ SB0.route_sel\[61\] SB0.route_sel\[60\] net62 _1534_ _1527_ vssd1 vssd1 vccd1
+ vccd1 _1536_ sky130_fd_sc_hd__a41o_1
X_1767_ _0393_ _0384_ _0396_ net305 vssd1 vssd1 vccd1 vccd1 _0397_ sky130_fd_sc_hd__a211o_4
XANTENNA__2497__A2 net29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3437_ clknet_leaf_8_clk _0257_ net259 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[1\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_57_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3299_ clknet_leaf_17_clk _0119_ net283 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[16\]
+ sky130_fd_sc_hd__dfstp_1
X_2319_ LE_1A.config_data\[1\] LE_1A.config_data\[0\] _0836_ vssd1 vssd1 vccd1 vccd1
+ _0948_ sky130_fd_sc_hd__mux2_1
X_3368_ clknet_leaf_24_clk _0188_ net272 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[60\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_57_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput98 net98 vssd1 vssd1 vccd1 vccd1 CBnorth_out[4] sky130_fd_sc_hd__buf_6
Xoutput76 net76 vssd1 vssd1 vccd1 vccd1 CBeast_out[13] sky130_fd_sc_hd__buf_6
Xoutput87 net87 vssd1 vssd1 vccd1 vccd1 CBeast_out[9] sky130_fd_sc_hd__buf_6
XANTENNA_input30_A CBnorth_in[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output117_A net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_59_Right_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2561__B net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2670_ _1394_ _1395_ SB0.route_sel\[109\] _1397_ _1295_ vssd1 vssd1 vccd1 vccd1 _1296_
+ sky130_fd_sc_hd__a221o_1
X_1621_ CB_1.config_dataA\[7\] vssd1 vssd1 vccd1 vccd1 _1459_ sky130_fd_sc_hd__inv_2
XANTENNA_clone40_A2 _0552_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2104_ net349 _0729_ _0733_ net352 _1483_ vssd1 vssd1 vccd1 vccd1 _0734_ sky130_fd_sc_hd__a221o_1
X_3222_ clknet_leaf_3_clk _0042_ net253 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[42\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2479__A2 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3153_ CB_1.config_dataA\[14\] net171 net224 vssd1 vssd1 vccd1 vccd1 _0321_ sky130_fd_sc_hd__mux2_1
XFILLER_62_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2035_ SB0.route_sel\[65\] SB0.route_sel\[64\] _0664_ _0663_ vssd1 vssd1 vccd1 vccd1
+ _0665_ sky130_fd_sc_hd__a211o_4
X_3084_ SB0.route_sel\[124\] SB0.route_sel\[123\] net298 vssd1 vssd1 vccd1 vccd1 _0252_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_37_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clone49_B1 _0490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2868_ LEI0.config_data\[36\] net472 net219 vssd1 vssd1 vccd1 vccd1 _0037_ sky130_fd_sc_hd__mux2_1
X_2937_ net200 CB_1.config_dataB\[2\] net225 vssd1 vssd1 vccd1 vccd1 _0105_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout148_A net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2799_ _1376_ _0511_ _0512_ vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__a21boi_1
X_1819_ _0445_ _0439_ _0448_ net305 vssd1 vssd1 vccd1 vccd1 _0449_ sky130_fd_sc_hd__a211o_4
XANTENNA__2167__A1 _0683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2094__A0 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clone35_A2 _0461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1841__B1 _0470_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2722_ _0368_ _1330_ vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__and2_4
X_2653_ CB_0.config_dataA\[19\] _1268_ _1278_ _1279_ vssd1 vssd1 vccd1 vccd1 _1280_
+ sky130_fd_sc_hd__o31a_1
X_2584_ LEI0.config_data\[14\] net234 _1210_ _1185_ vssd1 vssd1 vccd1 vccd1 _1211_
+ sky130_fd_sc_hd__a31oi_2
XANTENNA_clone51_A1 _0367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1604_ SB0.route_sel\[9\] vssd1 vssd1 vccd1 vccd1 _1442_ sky130_fd_sc_hd__inv_2
X_3136_ CB_0.config_dataB\[22\] CB_0.config_dataB\[23\] net227 vssd1 vssd1 vccd1 vccd1
+ _0304_ sky130_fd_sc_hd__mux2_1
X_3067_ SB0.route_sel\[107\] SB0.route_sel\[106\] net299 vssd1 vssd1 vccd1 vccd1 _0235_
+ sky130_fd_sc_hd__mux2_1
X_3205_ clknet_leaf_5_clk _0025_ net256 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_2018_ SB0.route_sel\[73\] SB0.route_sel\[72\] vssd1 vssd1 vccd1 vccd1 _0648_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout220_X net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3466__SET_B net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold161 LEI0.config_data\[4\] vssd1 vssd1 vccd1 vccd1 net471 sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 LEI0.config_data\[35\] vssd1 vssd1 vccd1 vccd1 net482 sky130_fd_sc_hd__dlygate4sd3_1
Xhold150 LE_1B.config_data\[1\] vssd1 vssd1 vccd1 vccd1 net460 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_56_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2312__A1 _0899_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2636_ CB_0.config_dataA\[17\] _1262_ vssd1 vssd1 vccd1 vccd1 _1263_ sky130_fd_sc_hd__nand2_1
XANTENNA__2790__A1 _0959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clone46_A1 _1548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2705_ SB0.route_sel\[57\] SB0.route_sel\[56\] vssd1 vssd1 vccd1 vccd1 _1319_ sky130_fd_sc_hd__nor2_1
X_2498_ net17 net24 net25 net26 net179 CB_0.config_dataB\[16\] vssd1 vssd1 vccd1 vccd1
+ _1126_ sky130_fd_sc_hd__mux4_1
X_2567_ net31 net32 net18 net19 CB_0.config_dataA\[5\] CB_0.config_dataA\[6\] vssd1
+ vssd1 vccd1 vccd1 _1194_ sky130_fd_sc_hd__mux4_1
XANTENNA__2764__X net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3119_ net183 net182 net214 vssd1 vssd1 vccd1 vccd1 _0287_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_4_clk_A clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1741__C1 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2674__X net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2772__A1 _1021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2421_ _1046_ _1047_ _1048_ vssd1 vssd1 vccd1 vccd1 _1049_ sky130_fd_sc_hd__a21oi_1
X_3470_ clknet_leaf_4_clk _0290_ net261 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[9\]
+ sky130_fd_sc_hd__dfstp_1
X_2283_ net171 _0521_ vssd1 vssd1 vccd1 vccd1 _0912_ sky130_fd_sc_hd__nand2_1
X_2352_ SB0.route_sel\[46\] SB0.route_sel\[47\] vssd1 vssd1 vccd1 vccd1 _0980_ sky130_fd_sc_hd__nand2b_1
XFILLER_64_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2288__A0 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2802__B1_N _0584_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout228_A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2460__A0 net31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2619_ _1173_ _1174_ _1179_ LE_0A.config_data\[4\] vssd1 vssd1 vccd1 vccd1 _1246_
+ sky130_fd_sc_hd__a211o_1
X_1998_ _1518_ _0604_ vssd1 vssd1 vccd1 vccd1 _0628_ sky130_fd_sc_hd__or2_1
XANTENNA__2212__A0 _0637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2279__A0 net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2654__B net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2754__A1 SB0.route_sel\[120\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire146 _1256_ vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_13_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input60_A SBwest_in[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1714__C1 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout290 net302 vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_29_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1921_ net145 _0549_ net237 vssd1 vssd1 vccd1 vccd1 _0551_ sky130_fd_sc_hd__o21ai_1
X_1852_ _0359_ _0416_ vssd1 vssd1 vccd1 vccd1 _0482_ sky130_fd_sc_hd__nand2_1
X_2970_ SB0.route_sel\[10\] SB0.route_sel\[9\] net291 vssd1 vssd1 vccd1 vccd1 _0138_
+ sky130_fd_sc_hd__mux2_1
X_3453_ clknet_leaf_10_clk _0273_ net263 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[17\]
+ sky130_fd_sc_hd__dfstp_1
X_1783_ _0404_ _0412_ vssd1 vssd1 vccd1 vccd1 _0413_ sky130_fd_sc_hd__nand2_1
X_3522_ clknet_leaf_32_clk _0342_ net241 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_3384_ clknet_leaf_4_clk _0204_ net261 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[76\]
+ sky130_fd_sc_hd__dfstp_1
X_2404_ _1025_ _1026_ _1031_ vssd1 vssd1 vccd1 vccd1 _1032_ sky130_fd_sc_hd__o21ai_4
X_2266_ net172 _0893_ _0894_ vssd1 vssd1 vccd1 vccd1 _0895_ sky130_fd_sc_hd__a21oi_1
X_2335_ _0487_ _0481_ _0962_ net306 vssd1 vssd1 vccd1 vccd1 _0963_ sky130_fd_sc_hd__a211o_4
X_2197_ _0491_ _0804_ _0807_ _0471_ CB_1.config_dataA\[2\] vssd1 vssd1 vccd1 vccd1
+ _0826_ sky130_fd_sc_hd__a221o_1
XFILLER_1_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2761__Y net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold98 LE_0A.config_data\[14\] vssd1 vssd1 vccd1 vccd1 net408 sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 _0071_ vssd1 vssd1 vccd1 vccd1 net397 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1711__A2 _1539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold76 LE_1A.config_data\[0\] vssd1 vssd1 vccd1 vccd1 net386 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_43_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_7 _1539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input63_X net63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2120_ net327 net344 net197 vssd1 vssd1 vccd1 vccd1 _0750_ sky130_fd_sc_hd__mux2_1
XFILLER_3_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2051_ _0544_ _0585_ _0638_ _0680_ vssd1 vssd1 vccd1 vccd1 _0681_ sky130_fd_sc_hd__o22a_1
X_1904_ _1518_ _0498_ vssd1 vssd1 vccd1 vccd1 _0534_ sky130_fd_sc_hd__or2_1
X_2884_ net454 LE_0A.config_data\[4\] net216 vssd1 vssd1 vccd1 vccd1 _0053_ sky130_fd_sc_hd__mux2_1
XANTENNA__2415__A0 net20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1835_ net153 _0462_ _0463_ _0464_ vssd1 vssd1 vccd1 vccd1 _0465_ sky130_fd_sc_hd__o211a_1
XANTENNA_clone38_A2 _0665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2953_ CB_1.config_dataB\[17\] CB_1.config_dataB\[18\] net229 vssd1 vssd1 vccd1 vccd1
+ _0121_ sky130_fd_sc_hd__mux2_1
XANTENNA__1654__A CB_0.le_outB vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3436_ clknet_leaf_4_clk _0256_ net261 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[0\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__2469__B net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1697_ SB0.route_sel\[61\] SB0.route_sel\[60\] vssd1 vssd1 vccd1 vccd1 _1535_ sky130_fd_sc_hd__nand2_1
X_3505_ clknet_leaf_22_clk _0325_ net273 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[19\]
+ sky130_fd_sc_hd__dfstp_1
X_1766_ _1430_ SB0.route_sel\[32\] SB0.route_sel\[37\] SB0.route_sel\[36\] _0395_
+ vssd1 vssd1 vccd1 vccd1 _0396_ sky130_fd_sc_hd__o221a_1
XANTENNA__2497__A3 net30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3298_ clknet_leaf_17_clk _0118_ net279 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[15\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_fanout295_A net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2249_ net172 _0875_ _0877_ vssd1 vssd1 vccd1 vccd1 _0878_ sky130_fd_sc_hd__a21oi_1
X_2318_ LE_1A.config_data\[3\] _0836_ _0867_ _0946_ vssd1 vssd1 vccd1 vccd1 _0947_
+ sky130_fd_sc_hd__o211a_1
X_3367_ clknet_leaf_24_clk _0187_ net267 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[59\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__2185__A2 _0543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput99 net99 vssd1 vssd1 vccd1 vccd1 CBnorth_out[5] sky130_fd_sc_hd__buf_6
Xoutput88 net88 vssd1 vssd1 vccd1 vccd1 CBnorth_out[0] sky130_fd_sc_hd__buf_6
Xoutput77 net77 vssd1 vssd1 vccd1 vccd1 CBeast_out[14] sky130_fd_sc_hd__buf_6
XANTENNA_input23_A CBnorth_in[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2645__A0 net27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1620_ SB0.route_sel\[122\] vssd1 vssd1 vccd1 vccd1 _1458_ sky130_fd_sc_hd__inv_2
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3083_ SB0.route_sel\[123\] SB0.route_sel\[122\] net301 vssd1 vssd1 vccd1 vccd1 _0251_
+ sky130_fd_sc_hd__mux2_1
X_2103_ net197 net196 vssd1 vssd1 vccd1 vccd1 _0733_ sky130_fd_sc_hd__nor2_1
XFILLER_39_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3221_ clknet_leaf_3_clk _0041_ net246 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[41\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2479__A3 net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3152_ CB_1.config_dataA\[13\] CB_1.config_dataA\[14\] net224 vssd1 vssd1 vccd1 vccd1
+ _0320_ sky130_fd_sc_hd__mux2_1
X_2034_ net144 _0662_ net237 vssd1 vssd1 vccd1 vccd1 _0664_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_45_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clone49_A1 _0487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout308_A net66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2798_ _1528_ net162 _0521_ vssd1 vssd1 vccd1 vccd1 _1376_ sky130_fd_sc_hd__o21ai_1
X_2867_ net482 LEI0.config_data\[36\] net211 vssd1 vssd1 vccd1 vccd1 _0036_ sky130_fd_sc_hd__mux2_1
X_2936_ net201 net200 net225 vssd1 vssd1 vccd1 vccd1 _0104_ sky130_fd_sc_hd__mux2_1
X_1818_ _1434_ SB0.route_sel\[24\] SB0.route_sel\[29\] SB0.route_sel\[28\] _0447_
+ vssd1 vssd1 vccd1 vccd1 _0448_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout210_A net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3419_ clknet_leaf_15_clk _0239_ net281 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[111\]
+ sky130_fd_sc_hd__dfstp_1
X_1749_ SB0.route_sel\[38\] SB0.route_sel\[39\] vssd1 vssd1 vccd1 vccd1 _0379_ sky130_fd_sc_hd__nand2_1
XFILLER_53_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2007__X _0637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clone16_A net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input26_X net26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2677__X net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2094__A1 net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1841__A1 _0467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2652_ CB_0.config_dataA\[18\] CB_0.config_dataA\[17\] CB_0.config_dataA\[19\] _1260_
+ vssd1 vssd1 vccd1 vccd1 _1279_ sky130_fd_sc_hd__or4bb_1
XTAP_TAPCELL_ROW_42_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2721_ _1426_ SB0.route_sel\[40\] _1427_ SB0.route_sel\[43\] _1329_ vssd1 vssd1 vccd1
+ vccd1 _1330_ sky130_fd_sc_hd__a221o_1
X_2583_ _1199_ _1209_ _1187_ vssd1 vssd1 vccd1 vccd1 _1210_ sky130_fd_sc_hd__a21o_1
XANTENNA_clone51_A2 _0358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3204_ clknet_leaf_3_clk _0024_ net245 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_1603_ SB0.route_sel\[20\] vssd1 vssd1 vccd1 vccd1 _1441_ sky130_fd_sc_hd__inv_2
XANTENNA__2609__A0 net31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3135_ CB_0.config_dataB\[21\] CB_0.config_dataB\[22\] net226 vssd1 vssd1 vccd1 vccd1
+ _0303_ sky130_fd_sc_hd__mux2_1
X_3066_ SB0.route_sel\[106\] SB0.route_sel\[105\] net299 vssd1 vssd1 vccd1 vccd1 _0234_
+ sky130_fd_sc_hd__mux2_1
X_2017_ net48 _0645_ _0646_ vssd1 vssd1 vccd1 vccd1 _0647_ sky130_fd_sc_hd__a21oi_1
XFILLER_50_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2919_ net434 net391 net204 vssd1 vssd1 vccd1 vccd1 _0088_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_19_Left_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold162 LEI0.config_data\[37\] vssd1 vssd1 vccd1 vccd1 net472 sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 _0333_ vssd1 vssd1 vccd1 vccd1 net461 sky130_fd_sc_hd__dlygate4sd3_1
Xhold140 LEI0.config_data\[46\] vssd1 vssd1 vccd1 vccd1 net450 sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 LEI0.config_data\[22\] vssd1 vssd1 vccd1 vccd1 net483 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_56_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clone46_A2 _1539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2635_ net20 net22 net21 net23 net186 net187 vssd1 vssd1 vccd1 vccd1 _1262_ sky130_fd_sc_hd__mux4_1
X_2704_ _1318_ _0676_ vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__and2_4
X_2497_ net27 net28 net29 net30 net179 net178 vssd1 vssd1 vccd1 vccd1 _1125_ sky130_fd_sc_hd__mux4_1
XANTENNA__2542__A2 _1014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2566_ net20 net22 net21 net23 CB_0.config_dataA\[6\] CB_0.config_dataA\[5\] vssd1
+ vssd1 vccd1 vccd1 _1193_ sky130_fd_sc_hd__mux4_1
X_3118_ CB_0.config_dataB\[4\] net183 net214 vssd1 vssd1 vccd1 vccd1 _0286_ sky130_fd_sc_hd__mux2_1
X_3049_ SB0.route_sel\[89\] SB0.route_sel\[88\] net295 vssd1 vssd1 vccd1 vccd1 _0217_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_2_157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1741__B1 _0370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2049__A1 _0675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2420_ net350 _1039_ _1040_ net317 _1466_ vssd1 vssd1 vccd1 vccd1 _1048_ sky130_fd_sc_hd__a221o_1
XANTENNA__1732__B1 net28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2351_ _0975_ net347 CB_0.config_dataB\[0\] vssd1 vssd1 vccd1 vccd1 _0979_ sky130_fd_sc_hd__mux2_1
XANTENNA__2288__A1 net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1753__Y _0383_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2282_ net170 net171 vssd1 vssd1 vccd1 vccd1 _0911_ sky130_fd_sc_hd__and2b_2
XTAP_TAPCELL_ROW_50_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2212__A1 _0615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1997_ _0617_ _0621_ _0625_ _0626_ vssd1 vssd1 vccd1 vccd1 _0627_ sky130_fd_sc_hd__a211o_4
X_2618_ LEI0.config_data\[26\] net234 _1243_ _1218_ vssd1 vssd1 vccd1 vccd1 _1245_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__3083__S net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2549_ LEI0.config_data\[0\] net160 vssd1 vssd1 vccd1 vccd1 _1176_ sky130_fd_sc_hd__nand2_1
XFILLER_51_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1962__B1 net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input53_A SBwest_in[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout280 net283 vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_29_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout291 net292 vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__clkbuf_4
X_1920_ _0547_ net153 _0548_ _0549_ vssd1 vssd1 vccd1 vccd1 _0550_ sky130_fd_sc_hd__o211a_1
X_1851_ _0472_ _0476_ _0480_ SB0.route_sel\[8\] SB0.route_sel\[9\] vssd1 vssd1 vccd1
+ vccd1 _0481_ sky130_fd_sc_hd__o2111ai_4
X_3452_ clknet_leaf_10_clk _0272_ net263 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[16\]
+ sky130_fd_sc_hd__dfstp_1
X_2403_ net304 LEI0.config_data\[5\] _1028_ _1030_ vssd1 vssd1 vccd1 vccd1 _1031_
+ sky130_fd_sc_hd__or4_4
X_3383_ clknet_leaf_4_clk _0203_ net261 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[75\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_clkbuf_leaf_3_clk_A clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1782_ SB0.route_sel\[21\] SB0.route_sel\[20\] net41 vssd1 vssd1 vccd1 vccd1 _0412_
+ sky130_fd_sc_hd__a21bo_1
X_3521_ clknet_leaf_32_clk _0341_ net241 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__1705__B1 net30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2196_ _0428_ _0449_ net177 vssd1 vssd1 vccd1 vccd1 _0825_ sky130_fd_sc_hd__mux2_1
X_2265_ _0371_ _0873_ _0876_ _0397_ _1461_ vssd1 vssd1 vccd1 vccd1 _0894_ sky130_fd_sc_hd__a221o_1
X_2334_ SB0.route_sel\[10\] SB0.route_sel\[11\] SB0.route_sel\[13\] _1445_ _0961_
+ vssd1 vssd1 vccd1 vccd1 _0962_ sky130_fd_sc_hd__o221a_1
XFILLER_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold88 LE_0A.config_data\[2\] vssd1 vssd1 vccd1 vccd1 net398 sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 _0064_ vssd1 vssd1 vccd1 vccd1 net409 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold77 _0086_ vssd1 vssd1 vccd1 vccd1 net387 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_16_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2424__B2 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2424__A1 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_7_Left_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input56_X net56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_8 net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2050_ _1495_ net362 net348 _0398_ CB_1.config_dataB\[2\] vssd1 vssd1 vccd1 vccd1
+ _0680_ sky130_fd_sc_hd__a221o_1
XANTENNA__2816__B1_N _1526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2415__A1 net22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2591__A net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2952_ net194 CB_1.config_dataB\[17\] net224 vssd1 vssd1 vccd1 vccd1 _0120_ sky130_fd_sc_hd__mux2_1
XFILLER_34_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1903_ _0527_ _0523_ _0530_ _0531_ _0532_ vssd1 vssd1 vccd1 vccd1 _0533_ sky130_fd_sc_hd__a221o_1
X_2883_ net398 LE_0A.config_data\[3\] net216 vssd1 vssd1 vccd1 vccd1 _0052_ sky130_fd_sc_hd__mux2_1
X_1834_ CB_0.config_dataA\[23\] CB_0.config_dataA\[22\] _0389_ vssd1 vssd1 vccd1 vccd1
+ _0464_ sky130_fd_sc_hd__or3_1
X_1765_ SB0.route_sel\[39\] SB0.route_sel\[38\] vssd1 vssd1 vccd1 vccd1 _0395_ sky130_fd_sc_hd__nand2b_1
XANTENNA__2351__A0 _0975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3435_ clknet_leaf_12_clk _0255_ net275 vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__dfstp_2
X_3504_ clknet_leaf_24_clk _0324_ net273 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[18\]
+ sky130_fd_sc_hd__dfstp_1
X_1696_ SB0.route_sel\[63\] SB0.route_sel\[62\] vssd1 vssd1 vccd1 vccd1 _1534_ sky130_fd_sc_hd__nand2_1
X_3366_ clknet_leaf_26_clk _0186_ net267 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[58\]
+ sky130_fd_sc_hd__dfstp_1
X_3297_ clknet_leaf_16_clk _0117_ net280 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[14\]
+ sky130_fd_sc_hd__dfstp_1
X_2179_ _0659_ _0804_ _0807_ _0679_ CB_1.config_dataA\[2\] vssd1 vssd1 vccd1 vccd1
+ _0808_ sky130_fd_sc_hd__a221o_1
X_2248_ _0659_ _0873_ _0876_ _0679_ CB_1.config_dataA\[12\] vssd1 vssd1 vccd1 vccd1
+ _0877_ sky130_fd_sc_hd__a221o_1
X_2317_ _0829_ _0830_ _0835_ LE_1A.config_data\[2\] vssd1 vssd1 vccd1 vccd1 _0946_
+ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout288_A net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3449__SET_B net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput89 net89 vssd1 vssd1 vccd1 vccd1 CBnorth_out[10] sky130_fd_sc_hd__buf_6
XANTENNA__2342__A0 net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput78 net78 vssd1 vssd1 vccd1 vccd1 CBeast_out[15] sky130_fd_sc_hd__buf_6
XANTENNA__1851__Y _0481_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2645__A1 net28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input16_A CBeast_in[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_0__f_clk_X clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1908__B1 net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3220_ clknet_leaf_3_clk _0040_ net245 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[40\]
+ sky130_fd_sc_hd__dfrtp_1
X_2033_ _0660_ net151 _0661_ _0662_ vssd1 vssd1 vccd1 vccd1 _0663_ sky130_fd_sc_hd__o211a_1
X_3082_ SB0.route_sel\[122\] SB0.route_sel\[121\] net301 vssd1 vssd1 vccd1 vccd1 _0250_
+ sky130_fd_sc_hd__mux2_1
X_2102_ net197 net354 _0731_ CB_1.config_dataB\[11\] vssd1 vssd1 vccd1 vccd1 _0732_
+ sky130_fd_sc_hd__o211a_1
X_3151_ CB_1.config_dataA\[12\] CB_1.config_dataA\[13\] net225 vssd1 vssd1 vccd1 vccd1
+ _0319_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_45_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clone49_A2 _0481_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2935_ CB_1.config_dataA\[24\] CB_1.config_dataB\[0\] net222 vssd1 vssd1 vccd1 vccd1
+ _0103_ sky130_fd_sc_hd__mux2_1
X_2797_ _1375_ _0464_ _0466_ vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__a21oi_2
X_2866_ net484 net482 net211 vssd1 vssd1 vccd1 vccd1 _0035_ sky130_fd_sc_hd__mux2_1
X_1817_ SB0.route_sel\[31\] SB0.route_sel\[30\] vssd1 vssd1 vccd1 vccd1 _0447_ sky130_fd_sc_hd__nand2b_1
XANTENNA_fanout203_A net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1748_ _0374_ _0376_ _0377_ vssd1 vssd1 vccd1 vccd1 _0378_ sky130_fd_sc_hd__a21bo_1
X_1679_ CB_0.config_dataB\[23\] CB_0.config_dataB\[22\] vssd1 vssd1 vccd1 vccd1 _1517_
+ sky130_fd_sc_hd__nand2b_2
X_3418_ clknet_leaf_15_clk _0238_ net280 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[110\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__2767__Y net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input8_A CBeast_in[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3349_ clknet_leaf_28_clk _0169_ net250 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[41\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_53_251 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input19_X net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output122_A net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1841__A2 _0461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2651_ CB_0.config_dataA\[18\] _1271_ _1274_ _1277_ vssd1 vssd1 vccd1 vccd1 _1278_
+ sky130_fd_sc_hd__nor4_1
X_2582_ CB_0.config_dataA\[8\] _1202_ _1205_ _1208_ _1473_ vssd1 vssd1 vccd1 vccd1
+ _1209_ sky130_fd_sc_hd__o41a_1
X_1602_ SB0.route_sel\[19\] vssd1 vssd1 vccd1 vccd1 _1440_ sky130_fd_sc_hd__inv_2
X_2720_ SB0.route_sel\[47\] SB0.route_sel\[46\] vssd1 vssd1 vccd1 vccd1 _1329_ sky130_fd_sc_hd__nor2_1
XANTENNA__3495__SET_B net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3203_ clknet_leaf_1_clk _0023_ net245 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_4_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3134_ CB_0.config_dataB\[20\] CB_0.config_dataB\[21\] net226 vssd1 vssd1 vccd1 vccd1
+ _0302_ sky130_fd_sc_hd__mux2_1
X_3065_ SB0.route_sel\[105\] SB0.route_sel\[104\] net300 vssd1 vssd1 vccd1 vccd1 _0233_
+ sky130_fd_sc_hd__mux2_1
X_2016_ SB0.route_sel\[77\] SB0.route_sel\[76\] net64 _0644_ _0639_ vssd1 vssd1 vccd1
+ vccd1 _0646_ sky130_fd_sc_hd__a41o_1
XFILLER_27_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_30_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2918_ net440 net434 net205 vssd1 vssd1 vccd1 vccd1 _0087_ sky130_fd_sc_hd__mux2_1
Xhold141 LE_0B.config_data\[12\] vssd1 vssd1 vccd1 vccd1 net451 sky130_fd_sc_hd__dlygate4sd3_1
Xhold174 LEI0.config_data\[34\] vssd1 vssd1 vccd1 vccd1 net484 sky130_fd_sc_hd__dlygate4sd3_1
X_2849_ LEI0.config_data\[17\] LEI0.config_data\[18\] net207 vssd1 vssd1 vccd1 vccd1
+ _0018_ sky130_fd_sc_hd__mux2_1
Xhold130 LE_1A.config_data\[1\] vssd1 vssd1 vccd1 vccd1 net440 sky130_fd_sc_hd__dlygate4sd3_1
Xhold152 LEI0.config_data\[8\] vssd1 vssd1 vccd1 vccd1 net462 sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 LE_1B.config_data\[9\] vssd1 vssd1 vccd1 vccd1 net473 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_56_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_21_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__1857__X _0487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2200__Y _0829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_20_Left_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_12_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__1767__X _0397_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2527__A0 net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2634_ _1001_ _0998_ _0991_ _0994_ net187 net186 vssd1 vssd1 vccd1 vccd1 _1261_ sky130_fd_sc_hd__mux4_1
X_2565_ _1188_ _1189_ _1191_ vssd1 vssd1 vccd1 vccd1 _1192_ sky130_fd_sc_hd__a21o_1
X_2703_ _1414_ SB0.route_sel\[64\] _1416_ SB0.route_sel\[67\] _1317_ vssd1 vssd1 vccd1
+ vccd1 _1318_ sky130_fd_sc_hd__a221o_1
X_2496_ net178 _1122_ _1123_ vssd1 vssd1 vccd1 vccd1 _1124_ sky130_fd_sc_hd__a21o_1
X_3117_ CB_0.config_dataB\[3\] CB_0.config_dataB\[4\] net215 vssd1 vssd1 vccd1 vccd1
+ _0285_ sky130_fd_sc_hd__mux2_1
XFILLER_63_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3048_ SB0.route_sel\[88\] SB0.route_sel\[87\] net290 vssd1 vssd1 vccd1 vccd1 _0216_
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_2_158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1741__A1 _0367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2049__A2 _0665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2221__A2 _0543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_1_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2281_ LEI0.config_data\[43\] _0907_ _0909_ LEI0.config_data\[44\] net303 vssd1 vssd1
+ vccd1 vccd1 _0910_ sky130_fd_sc_hd__a2111oi_1
X_2350_ _1548_ _1539_ _0977_ net306 vssd1 vssd1 vccd1 vccd1 _0978_ sky130_fd_sc_hd__a211o_4
XTAP_TAPCELL_ROW_50_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1996_ SB0.route_sel\[80\] SB0.route_sel\[81\] vssd1 vssd1 vccd1 vccd1 _0626_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_15_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2617_ LEI0.config_data\[26\] net234 _1243_ _1218_ vssd1 vssd1 vccd1 vccd1 _1244_
+ sky130_fd_sc_hd__a31oi_2
X_2548_ net143 net156 LEI0.config_data\[0\] vssd1 vssd1 vccd1 vccd1 _1175_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_66_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2775__Y net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2479_ net142 net155 net150 net160 LEI0.config_data\[39\] LEI0.config_data\[40\]
+ vssd1 vssd1 vccd1 vccd1 _1107_ sky130_fd_sc_hd__mux4_1
XFILLER_18_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload0 clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload0/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout281 net283 vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__clkbuf_2
XANTENNA__2398__B net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout270 net271 vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input46_A SBsouth_in[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout292 net293 vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__clkbuf_4
XANTENNA__1714__A1 _1548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1850_ SB0.route_sel\[13\] SB0.route_sel\[12\] net56 _0477_ _0479_ vssd1 vssd1 vccd1
+ vccd1 _0480_ sky130_fd_sc_hd__a41o_1
X_1781_ SB0.route_sel\[22\] SB0.route_sel\[23\] vssd1 vssd1 vccd1 vccd1 _0411_ sky130_fd_sc_hd__nand2_1
X_3520_ clknet_leaf_32_clk net474 net241 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_3451_ clknet_leaf_10_clk _0271_ net263 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[15\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__2101__B _0521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3382_ clknet_leaf_4_clk _0202_ net261 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[74\]
+ sky130_fd_sc_hd__dfstp_1
X_2402_ LEI0.config_data\[3\] _1493_ _1029_ LEI0.config_data\[4\] vssd1 vssd1 vccd1
+ vccd1 _1030_ sky130_fd_sc_hd__o211a_1
X_2333_ SB0.route_sel\[14\] SB0.route_sel\[15\] vssd1 vssd1 vccd1 vccd1 _0961_ sky130_fd_sc_hd__nand2b_1
X_2195_ CB_1.config_dataA\[3\] _0823_ vssd1 vssd1 vccd1 vccd1 _0824_ sky130_fd_sc_hd__nor2_1
X_2264_ _1526_ _1552_ net173 vssd1 vssd1 vccd1 vccd1 _0893_ sky130_fd_sc_hd__mux2_1
XANTENNA__1780__X _0410_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout233_A net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_23_Left_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1979_ _0605_ net152 _0606_ _0608_ vssd1 vssd1 vccd1 vccd1 _0609_ sky130_fd_sc_hd__o211a_1
XANTENNA__2197__B2 _0471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2197__A1 _0491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_42_Left_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold67 LE_0A.config_data\[7\] vssd1 vssd1 vccd1 vccd1 net377 sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 _0052_ vssd1 vssd1 vccd1 vccd1 net399 sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 LE_1B.config_data\[13\] vssd1 vssd1 vccd1 vccd1 net388 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_51_Left_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_9 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_60_Left_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input49_X net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1902_ SB0.route_sel\[112\] SB0.route_sel\[113\] vssd1 vssd1 vccd1 vccd1 _0532_ sky130_fd_sc_hd__nand2_1
XANTENNA__2415__A2 net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2951_ net195 net194 net229 vssd1 vssd1 vccd1 vccd1 _0119_ sky130_fd_sc_hd__mux2_1
X_2882_ net421 net398 net216 vssd1 vssd1 vccd1 vccd1 _0051_ sky130_fd_sc_hd__mux2_1
X_1833_ _0386_ _0417_ net17 vssd1 vssd1 vccd1 vccd1 _0463_ sky130_fd_sc_hd__o21ai_1
XANTENNA__2179__A1 _0659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2179__B2 _0679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_0_clk_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3503_ clknet_leaf_24_clk _0323_ net273 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[17\]
+ sky130_fd_sc_hd__dfstp_1
X_1764_ _0393_ _0384_ net305 vssd1 vssd1 vccd1 vccd1 _0394_ sky130_fd_sc_hd__a21oi_4
X_3296_ clknet_leaf_16_clk _0116_ net280 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[13\]
+ sky130_fd_sc_hd__dfstp_1
X_3434_ clknet_leaf_12_clk _0254_ net275 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[126\]
+ sky130_fd_sc_hd__dfstp_1
X_2316_ _0942_ _0867_ _0943_ _0944_ _0898_ vssd1 vssd1 vccd1 vccd1 _0945_ sky130_fd_sc_hd__a221o_1
X_3365_ clknet_leaf_26_clk _0185_ net267 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[57\]
+ sky130_fd_sc_hd__dfstp_1
X_1695_ _1529_ _1531_ _1532_ vssd1 vssd1 vccd1 vccd1 _1533_ sky130_fd_sc_hd__a21bo_1
X_2178_ net177 net176 vssd1 vssd1 vccd1 vccd1 _0807_ sky130_fd_sc_hd__nor2_1
X_2247_ net173 net172 vssd1 vssd1 vccd1 vccd1 _0876_ sky130_fd_sc_hd__nor2_1
XANTENNA__2406__A2 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2342__A1 net24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput79 net79 vssd1 vssd1 vccd1 vccd1 CBeast_out[1] sky130_fd_sc_hd__buf_6
XFILLER_0_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2645__A2 net29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1853__B1 net24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_2_clk_A clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_19_Right_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_28_Right_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3150_ net172 CB_1.config_dataA\[12\] net225 vssd1 vssd1 vccd1 vccd1 _0318_ sky130_fd_sc_hd__mux2_1
X_2032_ _0389_ _0607_ vssd1 vssd1 vccd1 vccd1 _0662_ sky130_fd_sc_hd__or2_1
X_2101_ net197 _0521_ vssd1 vssd1 vccd1 vccd1 _0731_ sky130_fd_sc_hd__nand2_1
X_3081_ SB0.route_sel\[121\] SB0.route_sel\[120\] net298 vssd1 vssd1 vccd1 vccd1 _0249_
+ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_37_Right_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3455__SET_B net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2865_ LEI0.config_data\[33\] net484 net211 vssd1 vssd1 vccd1 vccd1 _0034_ sky130_fd_sc_hd__mux2_1
X_2934_ net69 _0802_ _1393_ vssd1 vssd1 vccd1 vccd1 _0102_ sky130_fd_sc_hd__a21oi_1
X_1678_ CB_0.config_dataB\[23\] CB_0.config_dataB\[22\] vssd1 vssd1 vccd1 vccd1 _1516_
+ sky130_fd_sc_hd__and2b_1
X_2796_ net153 _0966_ _0462_ vssd1 vssd1 vccd1 vccd1 _1375_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_46_Right_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1816_ _0439_ _0445_ net305 vssd1 vssd1 vccd1 vccd1 _0446_ sky130_fd_sc_hd__a21o_4
X_1747_ net148 _1501_ _0375_ net236 vssd1 vssd1 vccd1 vccd1 _0377_ sky130_fd_sc_hd__o31a_1
XPHY_EDGE_ROW_55_Right_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3417_ clknet_leaf_16_clk _0237_ net280 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[109\]
+ sky130_fd_sc_hd__dfstp_1
X_3279_ clknet_leaf_32_clk _0099_ net242 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_3348_ clknet_leaf_28_clk _0168_ net249 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[40\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_53_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1850__A3 net56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2800__B1_N _0543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_64_Right_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2618__A2 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clone61_X net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2079__A0 net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clone7_C1 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2251__A0 net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2650_ net186 _1275_ _1276_ vssd1 vssd1 vccd1 vccd1 _1277_ sky130_fd_sc_hd__a21oi_1
X_2581_ net190 _1206_ _1207_ vssd1 vssd1 vccd1 vccd1 _1208_ sky130_fd_sc_hd__a21oi_1
X_1601_ SB0.route_sel\[18\] vssd1 vssd1 vccd1 vccd1 _1439_ sky130_fd_sc_hd__inv_2
X_3133_ CB_0.config_dataB\[19\] CB_0.config_dataB\[20\] net226 vssd1 vssd1 vccd1 vccd1
+ _0301_ sky130_fd_sc_hd__mux2_1
X_3202_ clknet_leaf_1_clk _0022_ net244 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_3064_ SB0.route_sel\[104\] SB0.route_sel\[103\] net300 vssd1 vssd1 vccd1 vccd1 _0232_
+ sky130_fd_sc_hd__mux2_1
X_2015_ SB0.route_sel\[77\] SB0.route_sel\[76\] vssd1 vssd1 vccd1 vccd1 _0645_ sky130_fd_sc_hd__nand2_1
XANTENNA__2124__X _0754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2848_ LEI0.config_data\[16\] LEI0.config_data\[17\] net214 vssd1 vssd1 vccd1 vccd1
+ _0017_ sky130_fd_sc_hd__mux2_1
X_2917_ net386 LE_1A.config_data\[1\] net204 vssd1 vssd1 vccd1 vccd1 _0086_ sky130_fd_sc_hd__mux2_1
X_2779_ _1366_ _0652_ _0654_ vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__a21oi_4
Xhold142 _0080_ vssd1 vssd1 vccd1 vccd1 net452 sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 LE_1A.config_data\[11\] vssd1 vssd1 vccd1 vccd1 net441 sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 _0340_ vssd1 vssd1 vccd1 vccd1 net474 sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 _0008_ vssd1 vssd1 vccd1 vccd1 net463 sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 LE_1B.config_data\[11\] vssd1 vssd1 vccd1 vccd1 net485 sky130_fd_sc_hd__dlygate4sd3_1
Xhold120 _0347_ vssd1 vssd1 vccd1 vccd1 net430 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_56_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clone21_A CBeast_in[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input31_X net31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2702_ SB0.route_sel\[71\] SB0.route_sel\[70\] vssd1 vssd1 vccd1 vccd1 _1317_ sky130_fd_sc_hd__nor2_1
X_2495_ net371 _1109_ _1113_ net319 CB_0.config_dataB\[17\] vssd1 vssd1 vccd1 vccd1
+ _1123_ sky130_fd_sc_hd__a221o_1
XANTENNA__2527__A1 net24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2633_ net186 net187 vssd1 vssd1 vccd1 vccd1 _1260_ sky130_fd_sc_hd__and2b_1
X_2564_ _1018_ _1186_ _1190_ _1021_ _1472_ vssd1 vssd1 vccd1 vccd1 _1191_ sky130_fd_sc_hd__a221o_1
X_3116_ CB_0.config_dataB\[2\] CB_0.config_dataB\[3\] net215 vssd1 vssd1 vccd1 vccd1
+ _0284_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_2_159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout263_A net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3047_ SB0.route_sel\[87\] SB0.route_sel\[86\] net290 vssd1 vssd1 vccd1 vccd1 _0215_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_18_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1741__A2 _0358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2029__X _0659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2757__B2 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2205__A net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2390__C1 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2280_ LEI0.config_data\[43\] _0908_ vssd1 vssd1 vccd1 vccd1 _0909_ sky130_fd_sc_hd__nor2_1
XANTENNA__2460__A3 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2445__A0 _0956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2616_ _1475_ _1230_ _1241_ _1242_ vssd1 vssd1 vccd1 vccd1 _1243_ sky130_fd_sc_hd__a31o_1
X_1995_ net34 _0623_ _0624_ vssd1 vssd1 vccd1 vccd1 _0625_ sky130_fd_sc_hd__a21oi_1
XFILLER_20_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2547_ LEI0.config_data\[2\] net234 vssd1 vssd1 vccd1 vccd1 _1174_ sky130_fd_sc_hd__and2_2
X_2478_ LE_0B.config_data\[1\] _1032_ _1064_ _1105_ vssd1 vssd1 vccd1 vccd1 _1106_
+ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_66_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload1 clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload1/Y sky130_fd_sc_hd__clkinvlp_4
XANTENNA__1688__X _1526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout260 net264 vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__clkbuf_2
Xfanout282 net283 vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__clkbuf_4
XFILLER_46_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout271 net285 vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input39_A SBsouth_in[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout293 net296 vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__clkbuf_4
XANTENNA__1714__A2 _1539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2427__A0 net27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2978__A1 SB0.route_sel\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1780_ net320 _0408_ _0409_ _0406_ net235 vssd1 vssd1 vccd1 vccd1 _0410_ sky130_fd_sc_hd__o221a_1
XFILLER_10_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3450_ clknet_leaf_9_clk _0270_ net263 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[14\]
+ sky130_fd_sc_hd__dfstp_1
X_2332_ _0956_ net339 CB_0.config_dataB\[0\] vssd1 vssd1 vccd1 vccd1 _0960_ sky130_fd_sc_hd__mux2_1
X_2401_ LEI0.config_data\[3\] net160 vssd1 vssd1 vccd1 vccd1 _1029_ sky130_fd_sc_hd__nand2_1
X_3381_ clknet_leaf_4_clk _0201_ net262 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[73\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2363__C1 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2194_ _0821_ _0822_ CB_1.config_dataA\[2\] vssd1 vssd1 vccd1 vccd1 _0823_ sky130_fd_sc_hd__mux2_1
XFILLER_37_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2263_ _0890_ _0891_ CB_1.config_dataA\[12\] vssd1 vssd1 vccd1 vccd1 _0892_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout226_A net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1978_ _1544_ _0607_ vssd1 vssd1 vccd1 vccd1 _0608_ sky130_fd_sc_hd__or2_1
Xhold68 _0057_ vssd1 vssd1 vccd1 vccd1 net378 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 LE_0B.config_data\[10\] vssd1 vssd1 vccd1 vccd1 net389 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2354__C1 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clone1_A1 _0829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2648__A0 _0975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2881_ net464 net421 net216 vssd1 vssd1 vccd1 vccd1 _0050_ sky130_fd_sc_hd__mux2_1
X_1901_ _0528_ _0529_ _0523_ vssd1 vssd1 vccd1 vccd1 _0531_ sky130_fd_sc_hd__a21oi_1
X_1832_ _0385_ _0416_ vssd1 vssd1 vccd1 vccd1 _0462_ sky130_fd_sc_hd__nand2_1
XANTENNA__2415__A3 net23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2950_ CB_1.config_dataB\[14\] CB_1.config_dataB\[15\] net229 vssd1 vssd1 vccd1 vccd1
+ _0118_ sky130_fd_sc_hd__mux2_1
XANTENNA__2281__D1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1763_ _0392_ _0391_ _0383_ vssd1 vssd1 vccd1 vccd1 _0393_ sky130_fd_sc_hd__or3b_4
X_3433_ clknet_leaf_12_clk _0253_ net275 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[125\]
+ sky130_fd_sc_hd__dfstp_1
X_1694_ net148 _1501_ _1530_ net235 vssd1 vssd1 vccd1 vccd1 _1532_ sky130_fd_sc_hd__o31a_1
X_3502_ clknet_leaf_22_clk _0322_ net273 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[16\]
+ sky130_fd_sc_hd__dfstp_1
X_3295_ clknet_leaf_16_clk _0115_ net279 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[12\]
+ sky130_fd_sc_hd__dfstp_2
X_2246_ _0637_ _0615_ net173 vssd1 vssd1 vccd1 vccd1 _0875_ sky130_fd_sc_hd__mux2_1
X_2315_ LE_1A.config_data\[5\] _0836_ _0866_ vssd1 vssd1 vccd1 vccd1 _0944_ sky130_fd_sc_hd__o21a_1
X_3364_ clknet_leaf_26_clk _0184_ net270 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[56\]
+ sky130_fd_sc_hd__dfstp_1
X_2177_ _0637_ _0615_ net177 vssd1 vssd1 vccd1 vccd1 _0806_ sky130_fd_sc_hd__mux2_4
XFILLER_25_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout229_X net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2645__A3 net30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2342__A2 net25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input61_X net61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3080_ SB0.route_sel\[120\] SB0.route_sel\[119\] net300 vssd1 vssd1 vccd1 vccd1 _0248_
+ sky130_fd_sc_hd__mux2_1
X_2100_ CB_1.config_dataB\[13\] _1483_ CB_1.config_dataB\[14\] _0729_ vssd1 vssd1
+ vccd1 vccd1 _0730_ sky130_fd_sc_hd__and4b_1
X_2031_ _0386_ _0604_ net31 vssd1 vssd1 vccd1 vccd1 _0661_ sky130_fd_sc_hd__o21ai_1
X_2795_ _1374_ _0484_ _0486_ vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__a21oi_2
X_1815_ _0443_ _0444_ _0438_ vssd1 vssd1 vccd1 vccd1 _0445_ sky130_fd_sc_hd__or3b_4
XTAP_TAPCELL_ROW_45_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2864_ LEI0.config_data\[32\] LEI0.config_data\[33\] net211 vssd1 vssd1 vccd1 vccd1
+ _0033_ sky130_fd_sc_hd__mux2_1
X_2933_ LE_1B.dff_out net69 vssd1 vssd1 vccd1 vccd1 _1393_ sky130_fd_sc_hd__nor2_1
X_1677_ net145 _1513_ _1514_ net237 vssd1 vssd1 vccd1 vccd1 _1515_ sky130_fd_sc_hd__o31a_1
X_3416_ clknet_leaf_16_clk _0236_ net280 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[108\]
+ sky130_fd_sc_hd__dfstp_1
X_1746_ net157 net169 net165 _0375_ _1501_ vssd1 vssd1 vccd1 vccd1 _0376_ sky130_fd_sc_hd__o32a_1
X_2229_ net1 net8 net9 net10 net175 net174 vssd1 vssd1 vccd1 vccd1 _0858_ sky130_fd_sc_hd__mux4_1
X_3278_ clknet_leaf_32_clk net417 net242 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_3347_ clknet_leaf_28_clk _0167_ net249 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[39\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_fanout293_A net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input21_A CBnorth_in[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2079__A1 net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2251__A1 net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output108_A net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1762__B1 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2580_ _0963_ _1186_ _1190_ _0966_ CB_0.config_dataA\[7\] vssd1 vssd1 vccd1 vccd1
+ _1207_ sky130_fd_sc_hd__a221o_1
X_1600_ SB0.route_sel\[17\] vssd1 vssd1 vccd1 vccd1 _1438_ sky130_fd_sc_hd__inv_2
X_3132_ CB_0.config_dataB\[18\] CB_0.config_dataB\[19\] net226 vssd1 vssd1 vccd1 vccd1
+ _0300_ sky130_fd_sc_hd__mux2_1
XANTENNA__2609__A3 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3063_ SB0.route_sel\[103\] SB0.route_sel\[102\] net298 vssd1 vssd1 vccd1 vccd1 _0231_
+ sky130_fd_sc_hd__mux2_1
X_3201_ clknet_leaf_1_clk _0021_ net245 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_2014_ SB0.route_sel\[79\] SB0.route_sel\[78\] vssd1 vssd1 vccd1 vccd1 _0644_ sky130_fd_sc_hd__nand2_1
X_2778_ net329 _0998_ _0650_ vssd1 vssd1 vccd1 vccd1 _1366_ sky130_fd_sc_hd__mux2_4
XFILLER_50_278 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_2_1__f_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2847_ LEI0.config_data\[15\] LEI0.config_data\[16\] net214 vssd1 vssd1 vccd1 vccd1
+ _0016_ sky130_fd_sc_hd__mux2_1
Xhold110 LE_1A.config_data\[8\] vssd1 vssd1 vccd1 vccd1 net420 sky130_fd_sc_hd__dlygate4sd3_1
X_2916_ LE_0B.config_data\[16\] net386 net205 vssd1 vssd1 vccd1 vccd1 _0085_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout306_A net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold154 LE_0A.config_data\[0\] vssd1 vssd1 vccd1 vccd1 net464 sky130_fd_sc_hd__dlygate4sd3_1
X_1729_ CB_0.config_dataB\[21\] CB_0.config_dataB\[24\] CB_0.config_dataB\[20\] vssd1
+ vssd1 vccd1 vccd1 _0359_ sky130_fd_sc_hd__nor3b_2
Xhold165 LEI0.config_data\[1\] vssd1 vssd1 vccd1 vccd1 net475 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout296_X net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold132 LE_0B.config_data\[8\] vssd1 vssd1 vccd1 vccd1 net442 sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 LE_0B.config_data\[1\] vssd1 vssd1 vccd1 vccd1 net431 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_1_clk_A clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold176 LEI0.config_data\[10\] vssd1 vssd1 vccd1 vccd1 net486 sky130_fd_sc_hd__dlygate4sd3_1
Xhold143 LEI0.config_data\[45\] vssd1 vssd1 vccd1 vccd1 net453 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_56_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1744__B1 net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input69_A le_en vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input24_X net24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2632_ net187 net186 vssd1 vssd1 vccd1 vccd1 _1259_ sky130_fd_sc_hd__nor2_1
X_2701_ _0676_ _1316_ vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__and2_4
XANTENNA__2527__A2 net25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2494_ _0956_ net339 net179 vssd1 vssd1 vccd1 vccd1 _1122_ sky130_fd_sc_hd__mux2_1
X_2563_ net191 net190 vssd1 vssd1 vccd1 vccd1 _1190_ sky130_fd_sc_hd__nor2_1
XANTENNA__2814__B1_N _1552_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3115_ net184 CB_0.config_dataB\[2\] net215 vssd1 vssd1 vccd1 vccd1 _0283_ sky130_fd_sc_hd__mux2_1
X_3046_ SB0.route_sel\[86\] SB0.route_sel\[85\] net290 vssd1 vssd1 vccd1 vccd1 _0214_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout256_A net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2215__A1 _0659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2215__B2 _0679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout309_X net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2045__X _0675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2142__A0 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1994_ SB0.route_sel\[85\] SB0.route_sel\[84\] net50 _0622_ _0617_ vssd1 vssd1 vccd1
+ vccd1 _0624_ sky130_fd_sc_hd__a41o_1
X_2615_ CB_0.config_dataA\[13\] _1474_ CB_0.config_dataA\[14\] _1221_ vssd1 vssd1
+ vccd1 vccd1 _1242_ sky130_fd_sc_hd__and4b_1
XANTENNA__1794__X _0424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload30 clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 clkload30/Y sky130_fd_sc_hd__inv_8
XANTENNA__1956__A0 net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2546_ _1160_ _1172_ _1149_ vssd1 vssd1 vccd1 vccd1 _1173_ sky130_fd_sc_hd__o21ai_4
X_2477_ _1025_ _1026_ _1031_ LE_0B.config_data\[0\] vssd1 vssd1 vccd1 vccd1 _1105_
+ sky130_fd_sc_hd__o211a_1
XANTENNA__2133__A0 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3029_ SB0.route_sel\[69\] SB0.route_sel\[68\] net297 vssd1 vssd1 vccd1 vccd1 _0197_
+ sky130_fd_sc_hd__mux2_1
Xclkload2 clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload2/Y sky130_fd_sc_hd__inv_6
XANTENNA__3302__SET_B net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2739__A2 SB0.route_sel\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout283 net284 vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__clkbuf_2
Xfanout261 net263 vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__clkbuf_4
Xfanout294 net296 vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__clkbuf_4
Xfanout272 net273 vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__clkbuf_4
Xfanout250 net285 vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__clkbuf_2
XFILLER_61_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2427__A1 net28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2400_ LEI0.config_data\[4\] _1027_ vssd1 vssd1 vccd1 vccd1 _1028_ sky130_fd_sc_hd__nor2_1
XFILLER_24_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3380_ clknet_leaf_4_clk _0200_ net262 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[72\]
+ sky130_fd_sc_hd__dfstp_1
X_2262_ net11 net12 net13 net14 net173 CB_1.config_dataA\[11\] vssd1 vssd1 vccd1 vccd1
+ _0891_ sky130_fd_sc_hd__mux4_1
X_2331_ _0445_ _0439_ _0958_ net305 vssd1 vssd1 vccd1 vccd1 _0959_ sky130_fd_sc_hd__a211o_4
X_2193_ net11 net12 net13 net331 net177 net176 vssd1 vssd1 vccd1 vccd1 _0822_ sky130_fd_sc_hd__mux4_1
X_1977_ CB_0.config_dataA\[22\] CB_0.config_dataA\[23\] vssd1 vssd1 vccd1 vccd1 _0607_
+ sky130_fd_sc_hd__nand2b_1
XANTENNA_fanout219_A net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2529_ _1154_ _1155_ CB_0.config_dataA\[2\] vssd1 vssd1 vccd1 vccd1 _1156_ sky130_fd_sc_hd__mux2_1
XANTENNA__2354__B1 _0981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold69 LE_1B.config_data\[14\] vssd1 vssd1 vccd1 vccd1 net379 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1875__A SB0.route_sel\[120\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input51_A SBwest_in[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2648__A1 _0978_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2880_ net65 net464 net216 vssd1 vssd1 vccd1 vccd1 _0049_ sky130_fd_sc_hd__mux2_1
X_1900_ _1452_ _1453_ net38 vssd1 vssd1 vccd1 vccd1 _0530_ sky130_fd_sc_hd__o21ai_1
X_1831_ _0455_ _0451_ _0458_ _0459_ _0460_ vssd1 vssd1 vccd1 vccd1 _0461_ sky130_fd_sc_hd__a221o_1
X_1762_ net144 _0390_ net234 vssd1 vssd1 vccd1 vccd1 _0392_ sky130_fd_sc_hd__o21ai_1
X_3432_ clknet_leaf_12_clk _0252_ net275 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[124\]
+ sky130_fd_sc_hd__dfstp_1
X_1693_ net157 net169 net167 _1530_ _1501_ vssd1 vssd1 vccd1 vccd1 _1531_ sky130_fd_sc_hd__o32a_1
X_3363_ clknet_leaf_26_clk _0183_ net270 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[55\]
+ sky130_fd_sc_hd__dfstp_1
X_3501_ clknet_leaf_21_clk _0321_ net274 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[15\]
+ sky130_fd_sc_hd__dfstp_1
X_3294_ clknet_leaf_16_clk _0114_ net279 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[11\]
+ sky130_fd_sc_hd__dfstp_1
X_2176_ CB_1.config_dataA\[3\] CB_1.config_dataA\[2\] CB_1.config_dataA\[4\] _0804_
+ vssd1 vssd1 vccd1 vccd1 _0805_ sky130_fd_sc_hd__or4bb_1
X_2245_ CB_1.config_dataA\[13\] _1461_ CB_1.config_dataA\[14\] _0873_ vssd1 vssd1
+ vccd1 vccd1 _0874_ sky130_fd_sc_hd__and4b_1
X_2314_ LE_1A.config_data\[4\] net311 vssd1 vssd1 vccd1 vccd1 _0943_ sky130_fd_sc_hd__nand2b_1
XFILLER_25_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2342__A3 net26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_1_Right_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2878__A1 CB_0.config_data_inA vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2566__A0 net20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input54_X net54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2053__X _0683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2030_ net164 _0603_ vssd1 vssd1 vccd1 vccd1 _0660_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_45_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2932_ net438 LEI0.config_data_in net202 vssd1 vssd1 vccd1 vccd1 _0101_ sky130_fd_sc_hd__mux2_1
X_2794_ net153 _0963_ _0482_ vssd1 vssd1 vccd1 vccd1 _1374_ sky130_fd_sc_hd__mux2_1
X_1814_ net144 _0442_ net237 vssd1 vssd1 vccd1 vccd1 _0444_ sky130_fd_sc_hd__o21ai_1
X_2863_ net487 LEI0.config_data\[32\] net211 vssd1 vssd1 vccd1 vccd1 _0032_ sky130_fd_sc_hd__mux2_1
X_1745_ CB_1.config_dataA\[24\] CB_1.config_dataA\[21\] CB_1.config_dataA\[20\] vssd1
+ vssd1 vccd1 vccd1 _0375_ sky130_fd_sc_hd__or3_4
X_1676_ CB_0.config_dataA\[24\] CB_0.config_dataA\[20\] CB_0.config_dataA\[21\] vssd1
+ vssd1 vccd1 vccd1 _1514_ sky130_fd_sc_hd__or3b_2
X_3415_ clknet_leaf_14_clk _0235_ net280 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[107\]
+ sky130_fd_sc_hd__dfstp_1
X_3346_ clknet_leaf_28_clk _0166_ net249 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[38\]
+ sky130_fd_sc_hd__dfstp_1
X_2228_ net11 net12 net13 net14 net175 net174 vssd1 vssd1 vccd1 vccd1 _0857_ sky130_fd_sc_hd__mux4_1
XFILLER_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3277_ clknet_leaf_30_clk _0097_ net247 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_2159_ _1481_ _1482_ _0691_ vssd1 vssd1 vccd1 vccd1 _0789_ sky130_fd_sc_hd__mux2_1
XANTENNA__2548__A0 net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_39_Left_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1771__A1 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_48_Left_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input14_A CBeast_in[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2079__A2 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_57_Left_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2251__A2 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_24_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3200_ clknet_leaf_1_clk _0020_ net245 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[20\]
+ sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_66_Left_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3131_ CB_0.config_dataB\[17\] CB_0.config_dataB\[18\] net226 vssd1 vssd1 vccd1 vccd1
+ _0299_ sky130_fd_sc_hd__mux2_1
X_3062_ SB0.route_sel\[102\] SB0.route_sel\[101\] net298 vssd1 vssd1 vccd1 vccd1 _0230_
+ sky130_fd_sc_hd__mux2_1
X_2013_ _0640_ _0641_ _0642_ vssd1 vssd1 vccd1 vccd1 _0643_ sky130_fd_sc_hd__a21bo_1
Xclkbuf_leaf_15_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_35_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1797__X _0427_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2915_ LE_1A.dff_out _0950_ net69 vssd1 vssd1 vccd1 vccd1 _0084_ sky130_fd_sc_hd__mux2_1
Xhold100 LE_0A.config_data\[5\] vssd1 vssd1 vccd1 vccd1 net410 sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 LE_0A.config_data\[3\] vssd1 vssd1 vccd1 vccd1 net454 sky130_fd_sc_hd__dlygate4sd3_1
Xhold111 LE_0A.config_data\[1\] vssd1 vssd1 vccd1 vccd1 net421 sky130_fd_sc_hd__dlygate4sd3_1
X_2777_ _1365_ _0630_ _0632_ vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__a21oi_4
X_2846_ LEI0.config_data\[14\] LEI0.config_data\[15\] net214 vssd1 vssd1 vccd1 vccd1
+ _0015_ sky130_fd_sc_hd__mux2_1
XANTENNA__1986__D1 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold122 _0069_ vssd1 vssd1 vccd1 vccd1 net432 sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 LE_1A.config_data\[7\] vssd1 vssd1 vccd1 vccd1 net443 sky130_fd_sc_hd__dlygate4sd3_1
X_1728_ _1554_ _0352_ _0356_ _0357_ vssd1 vssd1 vccd1 vccd1 _0358_ sky130_fd_sc_hd__a211o_1
XANTENNA_input6_A CBeast_in[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold177 LEI0.config_data\[31\] vssd1 vssd1 vccd1 vccd1 net487 sky130_fd_sc_hd__dlygate4sd3_1
X_3329_ clknet_leaf_29_clk _0149_ net247 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[21\]
+ sky130_fd_sc_hd__dfstp_1
Xhold166 LE_1B.config_data\[10\] vssd1 vssd1 vccd1 vccd1 net476 sky130_fd_sc_hd__dlygate4sd3_1
X_1659_ SB0.route_sel\[50\] SB0.route_sel\[51\] vssd1 vssd1 vccd1 vccd1 _1497_ sky130_fd_sc_hd__nand2_1
Xhold155 LE_0B.config_data_in vssd1 vssd1 vccd1 vccd1 net465 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2331__X _0959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input17_X net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output120_A net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2631_ net187 _1014_ _1257_ net186 vssd1 vssd1 vccd1 vccd1 _1258_ sky130_fd_sc_hd__o211a_1
XANTENNA__2527__A3 net26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2562_ net191 _1014_ net190 vssd1 vssd1 vccd1 vccd1 _1189_ sky130_fd_sc_hd__o21a_1
X_2700_ _1414_ _1415_ SB0.route_sel\[69\] _1417_ _1315_ vssd1 vssd1 vccd1 vccd1 _1316_
+ sky130_fd_sc_hd__a221o_1
X_2493_ CB_0.config_dataB\[17\] _1119_ _1120_ _1112_ vssd1 vssd1 vccd1 vccd1 _1121_
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__2401__B net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_4_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_4_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3114_ net185 net184 net217 vssd1 vssd1 vccd1 vccd1 _0282_ sky130_fd_sc_hd__mux2_1
X_3045_ SB0.route_sel\[85\] SB0.route_sel\[84\] net289 vssd1 vssd1 vccd1 vccd1 _0213_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_18_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2829_ _1391_ _0453_ _0454_ vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__a21boi_2
XANTENNA_input9_X net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1662__B1 net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2236__X _0865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1956__A1 net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1993_ SB0.route_sel\[85\] SB0.route_sel\[84\] vssd1 vssd1 vccd1 vccd1 _0623_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_0_clk_A clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2614_ _1234_ _1237_ _1240_ CB_0.config_dataA\[13\] vssd1 vssd1 vccd1 vccd1 _1241_
+ sky130_fd_sc_hd__or4b_1
X_2545_ CB_0.config_dataA\[3\] _1163_ _1167_ _1171_ CB_0.config_dataA\[4\] vssd1 vssd1
+ vccd1 vccd1 _1172_ sky130_fd_sc_hd__a41o_1
Xclkload31 clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 clkload31/Y sky130_fd_sc_hd__clkinv_4
Xclkload20 clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 clkload20/Y sky130_fd_sc_hd__inv_12
XFILLER_9_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2476_ LE_0B.config_data\[3\] _1032_ _1063_ _1103_ vssd1 vssd1 vccd1 vccd1 _1104_
+ sky130_fd_sc_hd__a211o_1
XANTENNA__2133__A1 net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3028_ SB0.route_sel\[68\] SB0.route_sel\[67\] net297 vssd1 vssd1 vccd1 vccd1 _0196_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__2436__A2 net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1985__X _0615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload3 clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 clkload3/Y sky130_fd_sc_hd__clkinv_8
Xfanout240 net243 vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__clkbuf_4
Xfanout284 net285 vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__clkbuf_2
XANTENNA__2427__A2 net29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout262 net263 vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__buf_2
Xfanout295 net296 vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__buf_2
Xfanout251 net253 vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__clkbuf_4
XFILLER_27_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout273 net274 vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_2_3__f_clk_X clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2363__A1 _0633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2828__B1_N _0471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2192_ net1 net8 net9 net330 net177 net176 vssd1 vssd1 vccd1 vccd1 _0821_ sky130_fd_sc_hd__mux4_1
XFILLER_37_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2261_ net1 net8 net9 net335 net173 CB_1.config_dataA\[11\] vssd1 vssd1 vccd1 vccd1
+ _0890_ sky130_fd_sc_hd__mux4_1
X_2330_ SB0.route_sel\[26\] SB0.route_sel\[27\] SB0.route_sel\[29\] _1437_ _0957_
+ vssd1 vssd1 vccd1 vccd1 _0958_ sky130_fd_sc_hd__o221a_1
XFILLER_37_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1976_ _1541_ _0604_ net19 vssd1 vssd1 vccd1 vccd1 _0606_ sky130_fd_sc_hd__o21ai_1
X_2528_ net27 net28 net29 net30 net193 CB_0.config_dataA\[1\] vssd1 vssd1 vccd1 vccd1
+ _1155_ sky130_fd_sc_hd__mux4_1
XANTENNA__2354__A1 _0367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2459_ net20 net22 net21 net23 net180 net181 vssd1 vssd1 vccd1 vccd1 _1087_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_26_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input44_A SBsouth_in[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1761_ net152 _0387_ _0388_ _0390_ vssd1 vssd1 vccd1 vccd1 _0391_ sky130_fd_sc_hd__o211a_1
XFILLER_42_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1830_ SB0.route_sel\[1\] SB0.route_sel\[0\] vssd1 vssd1 vccd1 vccd1 _0460_ sky130_fd_sc_hd__nand2_1
X_3500_ clknet_leaf_20_clk _0320_ net274 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[14\]
+ sky130_fd_sc_hd__dfstp_1
X_3431_ clknet_leaf_12_clk _0251_ net275 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[123\]
+ sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_27_Left_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3362_ clknet_leaf_26_clk _0182_ net270 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[54\]
+ sky130_fd_sc_hd__dfstp_1
X_2313_ LE_1A.config_data\[7\] LE_1A.config_data\[6\] net311 vssd1 vssd1 vccd1 vccd1
+ _0942_ sky130_fd_sc_hd__mux2_4
X_1692_ CB_1.config_dataA\[24\] CB_1.config_dataA\[21\] CB_1.config_dataA\[20\] vssd1
+ vssd1 vccd1 vccd1 _1530_ sky130_fd_sc_hd__nand3b_4
X_2175_ net176 net177 vssd1 vssd1 vccd1 vccd1 _0804_ sky130_fd_sc_hd__and2b_1
X_3293_ clknet_leaf_18_clk _0113_ net279 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[10\]
+ sky130_fd_sc_hd__dfstp_1
X_2244_ net172 net173 vssd1 vssd1 vccd1 vccd1 _0873_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_23_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_11_Left_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2024__B1 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1959_ _1477_ _0586_ _0588_ vssd1 vssd1 vccd1 vccd1 _0589_ sky130_fd_sc_hd__a21oi_1
XFILLER_56_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1929__B1_N net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1838__B1 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2566__A1 net22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2334__X _0962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input47_X net47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clknet_0_clk sky130_fd_sc_hd__clkbuf_16
X_2931_ net445 net438 net204 vssd1 vssd1 vccd1 vccd1 _0100_ sky130_fd_sc_hd__mux2_1
X_1813_ _0440_ net151 _0441_ _0442_ vssd1 vssd1 vccd1 vccd1 _0443_ sky130_fd_sc_hd__o211a_1
X_2793_ _0422_ _1373_ vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__nor2_4
X_2862_ LEI0.config_data\[30\] net487 net211 vssd1 vssd1 vccd1 vccd1 _0031_ sky130_fd_sc_hd__mux2_1
X_1744_ net169 net165 net11 vssd1 vssd1 vccd1 vccd1 _0374_ sky130_fd_sc_hd__o21ai_1
X_3414_ clknet_leaf_14_clk _0234_ net282 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[106\]
+ sky130_fd_sc_hd__dfstp_1
X_1675_ CB_0.config_dataA\[23\] CB_0.config_dataA\[22\] vssd1 vssd1 vccd1 vccd1 _1513_
+ sky130_fd_sc_hd__nand2b_1
X_3276_ clknet_leaf_30_clk _0096_ net247 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_3345_ clknet_leaf_28_clk _0165_ net248 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[37\]
+ sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_15_Right_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout279_A net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2227_ net174 _0854_ _0855_ vssd1 vssd1 vccd1 vccd1 _0856_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_24_Right_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2089_ LEI0.config_data\[21\] net147 _0718_ LEI0.config_data\[22\] vssd1 vssd1 vccd1
+ vccd1 _0719_ sky130_fd_sc_hd__o211a_1
X_2158_ _0722_ _0785_ _0787_ _0786_ _0755_ vssd1 vssd1 vccd1 vccd1 _0788_ sky130_fd_sc_hd__o221ai_2
XANTENNA__2796__A1 _0966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout234_X net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_33_Right_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1771__A2 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2079__A3 net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clone7_A2 _0570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_42_Right_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_51_Right_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2251__A3 net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3130_ net178 CB_0.config_dataB\[17\] net226 vssd1 vssd1 vccd1 vccd1 _0298_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_60_Right_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3061_ SB0.route_sel\[101\] SB0.route_sel\[100\] net295 vssd1 vssd1 vccd1 vccd1 _0229_
+ sky130_fd_sc_hd__mux2_1
X_2012_ net149 _0349_ _0593_ net236 vssd1 vssd1 vccd1 vccd1 _0642_ sky130_fd_sc_hd__o31a_1
XANTENNA__3500__SET_B net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2778__A1 _0998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2845_ net477 LEI0.config_data\[14\] net213 vssd1 vssd1 vccd1 vccd1 _0014_ sky130_fd_sc_hd__mux2_1
X_2914_ net433 LE_0B.config_data\[16\] net208 vssd1 vssd1 vccd1 vccd1 _0083_ sky130_fd_sc_hd__mux2_1
Xhold145 _0053_ vssd1 vssd1 vccd1 vccd1 net455 sky130_fd_sc_hd__dlygate4sd3_1
X_2776_ net329 _0991_ _0628_ vssd1 vssd1 vccd1 vccd1 _1365_ sky130_fd_sc_hd__mux2_4
Xhold167 LEI0.config_data\[13\] vssd1 vssd1 vccd1 vccd1 net477 sky130_fd_sc_hd__dlygate4sd3_1
Xhold101 LE_0A.config_data\[12\] vssd1 vssd1 vccd1 vccd1 net411 sky130_fd_sc_hd__dlygate4sd3_1
X_1658_ CB_1.config_dataB\[3\] CB_1.config_dataB\[2\] CB_1.config_dataB\[4\] _1495_
+ vssd1 vssd1 vccd1 vccd1 _1496_ sky130_fd_sc_hd__or4bb_1
Xhold134 LEI0.config_data\[40\] vssd1 vssd1 vccd1 vccd1 net444 sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 LE_0B.config_data\[15\] vssd1 vssd1 vccd1 vccd1 net433 sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 LE_1A.config_data\[5\] vssd1 vssd1 vccd1 vccd1 net422 sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 LE_1B.config_data\[4\] vssd1 vssd1 vccd1 vccd1 net466 sky130_fd_sc_hd__dlygate4sd3_1
X_1727_ SB0.route_sel\[41\] SB0.route_sel\[40\] vssd1 vssd1 vccd1 vccd1 _0357_ sky130_fd_sc_hd__nand2_1
XFILLER_58_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3259_ clknet_leaf_2_clk net424 net244 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_3328_ clknet_leaf_30_clk _0148_ net247 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[20\]
+ sky130_fd_sc_hd__dfstp_1
Xhold178 LEI0.config_data\[43\] vssd1 vssd1 vccd1 vccd1 net488 sky130_fd_sc_hd__dlygate4sd3_1
X_1589_ SB0.route_sel\[42\] vssd1 vssd1 vccd1 vccd1 _1427_ sky130_fd_sc_hd__inv_2
XANTENNA__2218__A0 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_14_Left_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2506__Y _1134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2492_ net317 _1109_ _1113_ net350 _1469_ vssd1 vssd1 vccd1 vccd1 _1120_ sky130_fd_sc_hd__a221o_1
X_2630_ net187 net138 vssd1 vssd1 vccd1 vccd1 _1257_ sky130_fd_sc_hd__nand2_1
X_2561_ net191 net138 vssd1 vssd1 vccd1 vccd1 _1188_ sky130_fd_sc_hd__nand2_1
XANTENNA__2393__C1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3113_ CB_0.config_dataA\[24\] CB_0.config_dataB\[0\] net226 vssd1 vssd1 vccd1 vccd1
+ _0281_ sky130_fd_sc_hd__mux2_1
XANTENNA_clone11_C1 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3302__Q CB_1.config_dataB\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3044_ SB0.route_sel\[84\] SB0.route_sel\[83\] net289 vssd1 vssd1 vccd1 vccd1 _0212_
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout144_A CB_0.le_outA vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2828_ net165 net163 _0471_ vssd1 vssd1 vccd1 vccd1 _1391_ sky130_fd_sc_hd__o21bai_1
X_2759_ SB0.route_sel\[112\] SB0.route_sel\[113\] vssd1 vssd1 vccd1 vccd1 _1355_ sky130_fd_sc_hd__or2_1
XFILLER_48_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2611__A0 _0991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2390__A2 _0570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1956__A2 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1992_ SB0.route_sel\[87\] SB0.route_sel\[86\] vssd1 vssd1 vccd1 vccd1 _0622_ sky130_fd_sc_hd__nand2_1
Xclkload10 clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 clkload10/Y sky130_fd_sc_hd__inv_6
X_2544_ _1168_ _1169_ _1170_ vssd1 vssd1 vccd1 vccd1 _1171_ sky130_fd_sc_hd__a21o_1
X_2613_ net188 _1238_ _1239_ vssd1 vssd1 vccd1 vccd1 _1240_ sky130_fd_sc_hd__a21oi_1
XANTENNA__2366__C1 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2475_ _1025_ _1026_ _1031_ LE_0B.config_data\[2\] vssd1 vssd1 vccd1 vccd1 _1103_
+ sky130_fd_sc_hd__o211a_1
Xclkload21 clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 clkload21/Y sky130_fd_sc_hd__inv_12
XTAP_TAPCELL_ROW_66_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3027_ SB0.route_sel\[67\] SB0.route_sel\[66\] net297 vssd1 vssd1 vccd1 vccd1 _0195_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout261_A net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout147_X net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2357__C1 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload4 clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 clkload4/Y sky130_fd_sc_hd__inv_6
Xfanout263 net264 vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__clkbuf_4
Xfanout230 net231 vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__clkbuf_4
Xfanout252 net253 vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__clkbuf_4
Xfanout274 net285 vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__clkbuf_4
Xfanout241 net243 vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__clkbuf_2
Xfanout285 net71 vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__buf_2
XANTENNA__2427__A3 net30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2832__A0 LEI0.config_data\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout296 net302 vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__clkbuf_2
XANTENNA__2337__X _0965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3467__SET_B net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2363__A2 _0627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2191_ net176 _0818_ _0819_ vssd1 vssd1 vccd1 vccd1 _0820_ sky130_fd_sc_hd__a21o_1
XANTENNA__2520__C1 net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2260_ net172 _0887_ _0888_ vssd1 vssd1 vccd1 vccd1 _0889_ sky130_fd_sc_hd__a21oi_1
X_1975_ _1540_ _0603_ vssd1 vssd1 vccd1 vccd1 _0605_ sky130_fd_sc_hd__nand2_1
X_2527_ net17 net24 net25 net26 net193 net192 vssd1 vssd1 vccd1 vccd1 _1154_ sky130_fd_sc_hd__mux4_1
X_2458_ net313 _1074_ _1084_ net180 CB_0.config_dataB\[12\] vssd1 vssd1 vccd1 vccd1
+ _1086_ sky130_fd_sc_hd__a221o_1
XFILLER_29_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2354__A2 _0358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2710__X net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout264_X net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2389_ SB0.route_sel\[106\] SB0.route_sel\[107\] SB0.route_sel\[109\] _1397_ _1016_
+ vssd1 vssd1 vccd1 vccd1 _1017_ sky130_fd_sc_hd__o221a_1
XFILLER_45_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input37_A SBsouth_in[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3103__S net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2942__S net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1760_ _1513_ _0389_ vssd1 vssd1 vccd1 vccd1 _0390_ sky130_fd_sc_hd__or2_1
XANTENNA__2584__A2 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1792__B1 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1691_ net169 net167 net14 vssd1 vssd1 vccd1 vccd1 _1529_ sky130_fd_sc_hd__o21ai_1
X_3292_ clknet_leaf_18_clk _0112_ net276 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[9\]
+ sky130_fd_sc_hd__dfstp_1
X_3430_ clknet_leaf_12_clk _0250_ net275 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[122\]
+ sky130_fd_sc_hd__dfstp_1
X_3361_ clknet_leaf_26_clk _0181_ net269 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[53\]
+ sky130_fd_sc_hd__dfstp_1
X_2312_ _0899_ _0904_ _0906_ _0940_ vssd1 vssd1 vccd1 vccd1 _0941_ sky130_fd_sc_hd__o31a_1
X_2174_ _0802_ _1491_ _0803_ vssd1 vssd1 vccd1 vccd1 CB_1.le_outB sky130_fd_sc_hd__a21oi_4
X_2243_ LEI0.config_data\[31\] _0869_ _0871_ LEI0.config_data\[32\] net303 vssd1 vssd1
+ vccd1 vccd1 _0872_ sky130_fd_sc_hd__a2111oi_1
XFILLER_33_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3450__SET_B net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1889_ _0506_ _0518_ net309 vssd1 vssd1 vccd1 vccd1 _0519_ sky130_fd_sc_hd__a21oi_2
X_1958_ CB_1.config_dataB\[2\] _0587_ CB_1.config_dataB\[3\] vssd1 vssd1 vccd1 vccd1
+ _0588_ sky130_fd_sc_hd__a21bo_1
XANTENNA__1838__A1 _0467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2812__B1_N _0679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2566__A2 net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2350__X _0978_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload2_A clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3298__SET_B net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2861_ net480 LEI0.config_data\[30\] net211 vssd1 vssd1 vccd1 vccd1 _0030_ sky130_fd_sc_hd__mux2_1
X_2930_ net449 net445 net204 vssd1 vssd1 vccd1 vccd1 _0099_ sky130_fd_sc_hd__mux2_1
X_3413_ clknet_leaf_14_clk _0233_ net282 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[105\]
+ sky130_fd_sc_hd__dfstp_1
X_1812_ CB_0.config_dataA\[23\] CB_0.config_dataA\[22\] _1544_ vssd1 vssd1 vccd1 vccd1
+ _0442_ sky130_fd_sc_hd__or3_1
X_2792_ _0418_ _0956_ _0421_ _0420_ vssd1 vssd1 vccd1 vccd1 _1373_ sky130_fd_sc_hd__o211a_1
X_1674_ _1511_ vssd1 vssd1 vccd1 vccd1 _1512_ sky130_fd_sc_hd__inv_2
X_1743_ CB_1.config_dataB\[21\] CB_1.config_dataB\[20\] CB_1.config_dataB\[24\] vssd1
+ vssd1 vccd1 vccd1 _0373_ sky130_fd_sc_hd__or3_1
X_2226_ _0491_ _0842_ _0843_ _0471_ CB_1.config_dataA\[7\] vssd1 vssd1 vccd1 vccd1
+ _0855_ sky130_fd_sc_hd__a221o_1
X_3275_ clknet_leaf_30_clk net405 net247 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_3344_ clknet_leaf_28_clk _0164_ net248 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[36\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_53_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2088_ LEI0.config_data\[21\] net160 vssd1 vssd1 vccd1 vccd1 _0718_ sky130_fd_sc_hd__nand2_1
X_2157_ LE_1B.config_data\[5\] _0691_ _0723_ vssd1 vssd1 vccd1 vccd1 _0787_ sky130_fd_sc_hd__a21o_1
XFILLER_42_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2181__A0 net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2058__A net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3060_ SB0.route_sel\[100\] SB0.route_sel\[99\] net295 vssd1 vssd1 vccd1 vccd1 _0228_
+ sky130_fd_sc_hd__mux2_1
X_2011_ net158 net166 net161 _0593_ _0349_ vssd1 vssd1 vccd1 vccd1 _0641_ sky130_fd_sc_hd__o32a_1
X_2844_ LEI0.config_data\[12\] net477 net213 vssd1 vssd1 vccd1 vccd1 _0013_ sky130_fd_sc_hd__mux2_1
X_2913_ net425 net433 net208 vssd1 vssd1 vccd1 vccd1 _0082_ sky130_fd_sc_hd__mux2_1
XANTENNA__1600__A SB0.route_sel\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold146 LE_0A.config_data\[4\] vssd1 vssd1 vccd1 vccd1 net456 sky130_fd_sc_hd__dlygate4sd3_1
X_2775_ _1364_ _0608_ _0610_ vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__a21oi_4
Xhold102 _0062_ vssd1 vssd1 vccd1 vccd1 net412 sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 LEI0.config_data\[25\] vssd1 vssd1 vccd1 vccd1 net478 sky130_fd_sc_hd__dlygate4sd3_1
X_1657_ _1478_ net200 vssd1 vssd1 vccd1 vccd1 _1495_ sky130_fd_sc_hd__nor2_1
Xhold113 LE_0B.config_data\[11\] vssd1 vssd1 vccd1 vccd1 net423 sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 LE_1B.config_data\[2\] vssd1 vssd1 vccd1 vccd1 net467 sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 LE_1A.config_data\[14\] vssd1 vssd1 vccd1 vccd1 net445 sky130_fd_sc_hd__dlygate4sd3_1
Xhold179 LEI0.config_data_in vssd1 vssd1 vccd1 vccd1 net489 sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 LE_1A.config_data\[2\] vssd1 vssd1 vccd1 vccd1 net434 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1738__B1 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1726_ net44 _0354_ _0355_ vssd1 vssd1 vccd1 vccd1 _0356_ sky130_fd_sc_hd__a21oi_1
X_1588_ SB0.route_sel\[41\] vssd1 vssd1 vccd1 vccd1 _1426_ sky130_fd_sc_hd__inv_2
XANTENNA__1910__B1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3258_ clknet_leaf_2_clk net390 net244 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_3327_ clknet_leaf_30_clk _0147_ net247 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[19\]
+ sky130_fd_sc_hd__dfstp_1
X_3189_ clknet_leaf_31_clk _0009_ net242 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_2209_ net326 net155 LEI0.config_data\[18\] vssd1 vssd1 vccd1 vccd1 _0838_ sky130_fd_sc_hd__mux2_4
XANTENNA__2218__A1 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_0__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_2_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__2950__S net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output106_A net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2491_ net20 net22 net21 net23 CB_0.config_dataB\[16\] CB_0.config_dataB\[15\] vssd1
+ vssd1 vccd1 vccd1 _1119_ sky130_fd_sc_hd__mux4_1
X_2560_ _1471_ _1472_ CB_0.config_dataA\[9\] _1186_ vssd1 vssd1 vccd1 vccd1 _1187_
+ sky130_fd_sc_hd__and4_1
X_3112_ CB_0.config_dataA\[23\] CB_0.config_dataA\[24\] net227 vssd1 vssd1 vccd1 vccd1
+ _0280_ sky130_fd_sc_hd__mux2_1
XFILLER_55_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clone11_B1 _1013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3043_ SB0.route_sel\[83\] SB0.route_sel\[82\] net289 vssd1 vssd1 vccd1 vccd1 _0211_
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3021__S net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2758_ _1354_ _0519_ vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__and2b_1
XANTENNA_fanout304_A net66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2827_ net320 _0474_ _0475_ _1390_ net235 vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__o221a_1
X_1709_ net145 _1545_ net237 vssd1 vssd1 vccd1 vccd1 _1547_ sky130_fd_sc_hd__o21ai_1
X_2689_ _1308_ _0634_ vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__and2_4
XFILLER_46_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2611__A1 _0994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input67_A en vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input22_X net22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3106__S net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2945__S net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2612_ _1001_ _1220_ _1221_ _0998_ CB_0.config_dataA\[12\] vssd1 vssd1 vccd1 vccd1
+ _1239_ sky130_fd_sc_hd__a221o_1
XANTENNA__1956__A3 net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1991_ _0618_ _0619_ _0620_ vssd1 vssd1 vccd1 vccd1 _0621_ sky130_fd_sc_hd__a21bo_1
Xclkload11 clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 clkload11/Y sky130_fd_sc_hd__clkinv_8
Xclkload22 clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 clkload22/Y sky130_fd_sc_hd__inv_12
XTAP_TAPCELL_ROW_15_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2543_ _1018_ _1148_ _1151_ _1021_ _1470_ vssd1 vssd1 vccd1 vccd1 _1170_ sky130_fd_sc_hd__a221o_1
X_2474_ _1065_ _1063_ _1099_ _1101_ vssd1 vssd1 vccd1 vccd1 _1102_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_66_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3026_ SB0.route_sel\[66\] SB0.route_sel\[65\] net298 vssd1 vssd1 vccd1 vccd1 _0194_
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout254_A net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload5 clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 clkload5/Y sky130_fd_sc_hd__clkinv_8
XANTENNA_fanout307_X net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2357__B1 _0984_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout220 net221 vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__buf_2
Xfanout264 net285 vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__buf_4
Xfanout231 _1392_ vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__buf_2
Xfanout275 net284 vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__clkbuf_4
XANTENNA__2109__A0 _0615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout297 net302 vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__clkbuf_4
Xfanout253 net285 vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__buf_2
Xfanout286 net287 vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__clkbuf_4
Xfanout242 net243 vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__clkbuf_4
XFILLER_24_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2353__X _0981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2060__A2 _0683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2190_ _0371_ _0804_ _0807_ _0397_ _1450_ vssd1 vssd1 vccd1 vccd1 _0819_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_63_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1974_ CB_0.config_dataB\[22\] CB_0.config_dataB\[23\] vssd1 vssd1 vccd1 vccd1 _0604_
+ sky130_fd_sc_hd__nand2b_1
XFILLER_52_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clone17_C1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2526_ net192 _1150_ _1152_ vssd1 vssd1 vccd1 vccd1 _1153_ sky130_fd_sc_hd__a21o_1
X_2388_ SB0.route_sel\[110\] SB0.route_sel\[111\] vssd1 vssd1 vccd1 vccd1 _1016_ sky130_fd_sc_hd__nand2b_1
X_2457_ net336 _1071_ vssd1 vssd1 vccd1 vccd1 _1085_ sky130_fd_sc_hd__and2_1
XFILLER_43_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3009_ SB0.route_sel\[49\] SB0.route_sel\[48\] net292 vssd1 vssd1 vccd1 vccd1 _0177_
+ sky130_fd_sc_hd__mux2_1
XFILLER_51_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2569__A0 _0991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1690_ CB_1.config_dataB\[24\] CB_1.config_dataB\[20\] CB_1.config_dataB\[21\] vssd1
+ vssd1 vccd1 vccd1 _1528_ sky130_fd_sc_hd__nand3b_2
X_3291_ clknet_leaf_18_clk _0111_ net276 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[8\]
+ sky130_fd_sc_hd__dfstp_1
X_2311_ LEI0.config_data\[44\] net232 _0938_ _0910_ vssd1 vssd1 vccd1 vccd1 _0940_
+ sky130_fd_sc_hd__a31o_1
X_2242_ LEI0.config_data\[31\] _0870_ vssd1 vssd1 vccd1 vccd1 _0871_ sky130_fd_sc_hd__nor2_1
X_3360_ clknet_leaf_26_clk _0180_ net269 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[52\]
+ sky130_fd_sc_hd__dfstp_1
X_2173_ LE_1B.dff_out _1491_ net232 vssd1 vssd1 vccd1 vccd1 _0803_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_31_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1957_ net4 net6 net5 net7 CB_1.config_dataB\[1\] net201 vssd1 vssd1 vccd1 vccd1
+ _0587_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_23_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1888_ _0513_ _0507_ _0516_ _0517_ _0505_ vssd1 vssd1 vccd1 vccd1 _0518_ sky130_fd_sc_hd__a221o_4
X_2509_ _1098_ _1104_ _1106_ _1136_ vssd1 vssd1 vccd1 vccd1 _1137_ sky130_fd_sc_hd__a31o_1
XFILLER_56_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3489_ clknet_leaf_16_clk _0309_ net280 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[3\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__1838__A2 _0461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2566__A3 net23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1710__X _1548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2953__S net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_27_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_output136_A net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1811_ _1541_ _0417_ net26 vssd1 vssd1 vccd1 vccd1 _0441_ sky130_fd_sc_hd__o21ai_1
X_2791_ _1372_ _0442_ _0444_ vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__a21oi_4
X_2860_ net481 net480 net211 vssd1 vssd1 vccd1 vccd1 _0029_ sky130_fd_sc_hd__mux2_1
XANTENNA__2254__A2 _0543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3412_ clknet_leaf_14_clk _0232_ net282 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[104\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_7_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1742_ SB0.route_sel\[34\] SB0.route_sel\[35\] vssd1 vssd1 vccd1 vccd1 _0372_ sky130_fd_sc_hd__nand2_1
X_1673_ SB0.route_sel\[49\] SB0.route_sel\[48\] vssd1 vssd1 vccd1 vccd1 _1511_ sky130_fd_sc_hd__and2_1
XANTENNA__2190__A1 _0371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2190__B2 _0397_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2225_ _0428_ _0449_ net175 vssd1 vssd1 vccd1 vccd1 _0854_ sky130_fd_sc_hd__mux2_1
X_3274_ clknet_leaf_30_clk _0094_ net247 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_3343_ clknet_leaf_28_clk _0163_ net251 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[35\]
+ sky130_fd_sc_hd__dfstp_1
Xclkbuf_leaf_18_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_36_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2156_ _0690_ LE_1B.config_data\[4\] vssd1 vssd1 vccd1 vccd1 _0786_ sky130_fd_sc_hd__and2_4
XPHY_EDGE_ROW_5_Right_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2087_ net326 net155 LEI0.config_data\[21\] vssd1 vssd1 vccd1 vccd1 _0717_ sky130_fd_sc_hd__mux2_1
XANTENNA__2716__X net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2989_ SB0.route_sel\[29\] SB0.route_sel\[28\] net291 vssd1 vssd1 vccd1 vccd1 _0157_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__2181__A1 net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1995__A1 net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input52_X net52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2010_ net166 net161 net16 vssd1 vssd1 vccd1 vccd1 _0640_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_58_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_35_Left_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2912_ LE_0B.config_data\[13\] net425 net208 vssd1 vssd1 vccd1 vccd1 _0081_ sky130_fd_sc_hd__mux2_1
X_2774_ net329 _0994_ _0605_ vssd1 vssd1 vccd1 vccd1 _1364_ sky130_fd_sc_hd__mux2_4
XPHY_EDGE_ROW_44_Left_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2843_ LEI0.config_data\[11\] LEI0.config_data\[12\] net212 vssd1 vssd1 vccd1 vccd1
+ _0012_ sky130_fd_sc_hd__mux2_1
XANTENNA__1738__A1 _0367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1725_ SB0.route_sel\[45\] SB0.route_sel\[44\] net60 _0353_ _1554_ vssd1 vssd1 vccd1
+ vccd1 _0355_ sky130_fd_sc_hd__a41o_1
Xclkbuf_leaf_7_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_clk
+ sky130_fd_sc_hd__clkbuf_8
Xhold114 _0079_ vssd1 vssd1 vccd1 vccd1 net424 sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 LEI0.config_data\[39\] vssd1 vssd1 vccd1 vccd1 net457 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2826__B1_N _0491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold136 LE_1A.config_data\[10\] vssd1 vssd1 vccd1 vccd1 net446 sky130_fd_sc_hd__dlygate4sd3_1
Xhold125 LE_1B.config_data\[5\] vssd1 vssd1 vccd1 vccd1 net435 sky130_fd_sc_hd__dlygate4sd3_1
X_3326_ clknet_leaf_30_clk _0146_ net248 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[18\]
+ sky130_fd_sc_hd__dfstp_1
Xhold158 _0334_ vssd1 vssd1 vccd1 vccd1 net468 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3019__S net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold103 LE_1B.config_data\[7\] vssd1 vssd1 vccd1 vccd1 net413 sky130_fd_sc_hd__dlygate4sd3_1
Xhold169 LEI0.config_data\[7\] vssd1 vssd1 vccd1 vccd1 net479 sky130_fd_sc_hd__dlygate4sd3_1
X_1656_ net160 vssd1 vssd1 vccd1 vccd1 _1494_ sky130_fd_sc_hd__inv_2
X_1587_ SB0.route_sel\[52\] vssd1 vssd1 vccd1 vccd1 _1425_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout284_A net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1910__A1 _0533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_53_Left_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2139_ CB_1.config_dataB\[16\] _0767_ _0768_ vssd1 vssd1 vccd1 vccd1 _0769_ sky130_fd_sc_hd__a21oi_1
X_3257_ clknet_leaf_2_clk _0077_ net244 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_2208_ net147 net159 LEI0.config_data\[18\] vssd1 vssd1 vccd1 vccd1 _0837_ sky130_fd_sc_hd__mux2_1
X_3188_ clknet_leaf_0_clk net463 net242 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2218__A2 net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input12_A CBeast_in[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2356__X _0984_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2490_ _1114_ _1116_ _1117_ CB_0.config_dataB\[17\] vssd1 vssd1 vccd1 vccd1 _1118_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__2393__A1 _0562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3111_ CB_0.config_dataA\[22\] CB_0.config_dataA\[23\] net226 vssd1 vssd1 vccd1 vccd1
+ _0279_ sky130_fd_sc_hd__mux2_1
XANTENNA_clone11_A1 _0539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3042_ SB0.route_sel\[82\] SB0.route_sel\[81\] net289 vssd1 vssd1 vccd1 vccd1 _0210_
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1671__A3 net61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2713__Y net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1708_ _1492_ _1542_ _1543_ _1545_ vssd1 vssd1 vccd1 vccd1 _1546_ sky130_fd_sc_hd__o211a_1
X_2757_ _1455_ SB0.route_sel\[121\] SB0.route_sel\[126\] net136 _1353_ vssd1 vssd1
+ vccd1 vccd1 _1354_ sky130_fd_sc_hd__o221a_1
X_2688_ SB0.route_sel\[82\] _1408_ SB0.route_sel\[85\] _1409_ _1307_ vssd1 vssd1 vccd1
+ vccd1 _1308_ sky130_fd_sc_hd__a221o_1
X_2826_ net166 net163 _0491_ vssd1 vssd1 vccd1 vccd1 _1390_ sky130_fd_sc_hd__o21ba_1
XANTENNA_input4_A CBeast_in[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1639_ CB_1.config_dataB\[2\] vssd1 vssd1 vccd1 vccd1 _1477_ sky130_fd_sc_hd__inv_2
X_3309_ clknet_leaf_24_clk _0129_ net272 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[1\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__2439__A2 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input15_X net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3122__S net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1990_ net149 _1502_ _0593_ net236 vssd1 vssd1 vccd1 vccd1 _0620_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_15_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2542_ net193 _1014_ net192 vssd1 vssd1 vccd1 vccd1 _1169_ sky130_fd_sc_hd__o21a_1
X_2611_ _0991_ _0994_ CB_0.config_dataA\[10\] vssd1 vssd1 vccd1 vccd1 _1238_ sky130_fd_sc_hd__mux2_1
Xclkload12 clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 clkload12/Y sky130_fd_sc_hd__clkinv_1
Xclkload23 clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 clkload23/Y sky130_fd_sc_hd__bufinv_16
X_2473_ LE_0B.config_data\[5\] _1032_ _1064_ _1100_ vssd1 vssd1 vccd1 vccd1 _1101_
+ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_66_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3025_ SB0.route_sel\[65\] SB0.route_sel\[64\] net298 vssd1 vssd1 vccd1 vccd1 _0193_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__2156__B LE_1B.config_data\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload6 clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 clkload6/X sky130_fd_sc_hd__clkbuf_4
X_2809_ _1381_ _0619_ _0620_ vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__a21boi_2
XANTENNA__2357__A1 _0393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout221 net231 vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__buf_2
XANTENNA_input7_X net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout276 net284 vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__buf_2
Xfanout298 net301 vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__clkbuf_4
Xfanout254 net264 vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__clkbuf_4
XANTENNA__3496__SET_B net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout243 net285 vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__buf_2
XANTENNA__1803__X _0433_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout232 net233 vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__buf_4
Xfanout287 net288 vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__clkbuf_4
Xfanout210 net221 vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__clkbuf_4
XFILLER_42_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1973_ CB_0.config_dataB\[22\] CB_0.config_dataB\[23\] vssd1 vssd1 vccd1 vccd1 _0603_
+ sky130_fd_sc_hd__and2b_1
XANTENNA_clone17_B1 _0427_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2525_ _0982_ _1148_ _1151_ _0985_ _1470_ vssd1 vssd1 vccd1 vccd1 _1152_ sky130_fd_sc_hd__a221o_1
XANTENNA_clone33_C1 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2387_ net185 net321 net184 vssd1 vssd1 vccd1 vccd1 _1015_ sky130_fd_sc_hd__o21a_1
X_2456_ net341 net338 net181 vssd1 vssd1 vccd1 vccd1 _1084_ sky130_fd_sc_hd__mux2_1
XANTENNA__3324__Q SB0.route_sel\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2719__X net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3008_ SB0.route_sel\[48\] SB0.route_sel\[47\] net292 vssd1 vssd1 vccd1 vccd1 _0176_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__2502__A1 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2502__B2 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2569__A1 _0994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1712__A_N SB0.route_sel\[63\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3290_ clknet_leaf_18_clk _0110_ net276 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[7\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__1701__C1 _1538_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2310_ LEI0.config_data\[44\] net232 _0938_ net139 vssd1 vssd1 vccd1 vccd1 _0939_
+ sky130_fd_sc_hd__a31oi_1
X_2172_ _0788_ _0784_ _0792_ _0796_ _0801_ vssd1 vssd1 vccd1 vccd1 _0802_ sky130_fd_sc_hd__a32o_2
X_2241_ net142 net155 LEI0.config_data\[30\] vssd1 vssd1 vccd1 vccd1 _0870_ sky130_fd_sc_hd__mux2_1
XANTENNA_clone28_C1 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1887_ _0514_ _0515_ _0507_ vssd1 vssd1 vccd1 vccd1 _0517_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_31_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1956_ net15 net16 net2 net3 net201 CB_1.config_dataB\[1\] vssd1 vssd1 vccd1 vccd1
+ _0586_ sky130_fd_sc_hd__mux4_1
X_3488_ clknet_leaf_15_clk _0308_ net280 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[2\]
+ sky130_fd_sc_hd__dfstp_2
X_2508_ LEI0.config_data\[41\] _1134_ _1108_ vssd1 vssd1 vccd1 vccd1 _1136_ sky130_fd_sc_hd__a21o_1
X_2439_ LEI0.config_data\[27\] net147 _1066_ LEI0.config_data\[28\] vssd1 vssd1 vccd1
+ vccd1 _1067_ sky130_fd_sc_hd__o211a_1
XANTENNA_rebuffer15_A _0675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input42_A SBsouth_in[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output129_A net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1810_ _1540_ _0416_ vssd1 vssd1 vccd1 vccd1 _0440_ sky130_fd_sc_hd__nand2_1
X_2790_ net329 _0959_ _0440_ vssd1 vssd1 vccd1 vccd1 _1372_ sky130_fd_sc_hd__mux2_4
X_1741_ _0367_ _0358_ _0370_ net305 vssd1 vssd1 vccd1 vccd1 _0371_ sky130_fd_sc_hd__a211o_4
X_3411_ clknet_leaf_19_clk _0231_ net276 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[103\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_7_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1672_ _1508_ _1509_ _1506_ _1497_ vssd1 vssd1 vccd1 vccd1 _1510_ sky130_fd_sc_hd__a2bb2o_4
X_3342_ clknet_leaf_28_clk _0162_ net252 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[34\]
+ sky130_fd_sc_hd__dfstp_1
X_2224_ _0845_ _0848_ _0852_ CB_1.config_dataA\[8\] vssd1 vssd1 vccd1 vccd1 _0853_
+ sky130_fd_sc_hd__or4b_1
X_2155_ LE_1B.config_data\[6\] LE_1B.config_data\[7\] _0691_ vssd1 vssd1 vccd1 vccd1
+ _0785_ sky130_fd_sc_hd__mux2_1
X_3273_ clknet_leaf_30_clk _0093_ net247 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_2086_ _0703_ _0715_ _0693_ vssd1 vssd1 vccd1 vccd1 _0716_ sky130_fd_sc_hd__o21ai_4
XTAP_TAPCELL_ROW_36_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1939_ net145 _0567_ net238 vssd1 vssd1 vccd1 vccd1 _0569_ sky130_fd_sc_hd__o21ai_1
XFILLER_21_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2988_ SB0.route_sel\[28\] SB0.route_sel\[27\] net286 vssd1 vssd1 vccd1 vccd1 _0156_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__1913__C1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2181__A2 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2166__C1 _0755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_11_Right_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2090__A net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_20_Right_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3125__S net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2911_ net451 LE_0B.config_data\[13\] net206 vssd1 vssd1 vccd1 vccd1 _0080_ sky130_fd_sc_hd__mux2_1
X_2773_ _0549_ _1363_ _0551_ vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__a21oi_4
Xhold104 _0339_ vssd1 vssd1 vccd1 vccd1 net414 sky130_fd_sc_hd__dlygate4sd3_1
Xhold126 LE_1A.config_data\[4\] vssd1 vssd1 vccd1 vccd1 net436 sky130_fd_sc_hd__dlygate4sd3_1
X_1724_ SB0.route_sel\[45\] SB0.route_sel\[44\] vssd1 vssd1 vccd1 vccd1 _0354_ sky130_fd_sc_hd__nand2_1
XANTENNA__1738__A2 _0358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2842_ net486 LEI0.config_data\[11\] net204 vssd1 vssd1 vccd1 vccd1 _0011_ sky130_fd_sc_hd__mux2_1
Xhold115 LE_0B.config_data\[14\] vssd1 vssd1 vccd1 vccd1 net425 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1910__A2 _0539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold159 LEI0.config_data\[2\] vssd1 vssd1 vccd1 vccd1 net469 sky130_fd_sc_hd__dlygate4sd3_1
X_3256_ clknet_leaf_6_clk _0076_ net254 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold137 LE_0B.config_data\[2\] vssd1 vssd1 vccd1 vccd1 net447 sky130_fd_sc_hd__dlygate4sd3_1
X_1655_ net150 vssd1 vssd1 vccd1 vccd1 _1493_ sky130_fd_sc_hd__inv_2
X_3325_ clknet_leaf_28_clk _0145_ net248 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[17\]
+ sky130_fd_sc_hd__dfstp_2
Xhold148 LE_1B.config_data\[0\] vssd1 vssd1 vccd1 vccd1 net458 sky130_fd_sc_hd__dlygate4sd3_1
X_1586_ SB0.route_sel\[53\] vssd1 vssd1 vccd1 vccd1 _1424_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout277_A net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2069_ net361 _0692_ _0694_ net357 _1479_ vssd1 vssd1 vccd1 vccd1 _0699_ sky130_fd_sc_hd__a221o_1
X_2138_ net12 _0760_ _0761_ net11 CB_1.config_dataB\[18\] vssd1 vssd1 vccd1 vccd1
+ _0768_ sky130_fd_sc_hd__a221o_1
XANTENNA__2320__C1 _0899_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2207_ _0830_ _0829_ _0835_ vssd1 vssd1 vccd1 vccd1 _0836_ sky130_fd_sc_hd__a21oi_4
X_3187_ clknet_leaf_0_clk _0007_ net242 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2218__A3 net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout232_X net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2537__S0 CB_0.config_dataA\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2393__A2 _0552_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3110_ CB_0.config_dataA\[21\] CB_0.config_dataA\[22\] net226 vssd1 vssd1 vccd1 vccd1
+ _0278_ sky130_fd_sc_hd__mux2_1
XFILLER_4_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clone11_A2 _0533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3041_ SB0.route_sel\[81\] SB0.route_sel\[80\] net290 vssd1 vssd1 vccd1 vccd1 _0209_
+ sky130_fd_sc_hd__mux2_1
XFILLER_63_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2825_ net320 _0408_ _0409_ _1389_ net235 vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__o221a_4
X_1638_ CB_0.config_dataA\[17\] vssd1 vssd1 vccd1 vccd1 _1476_ sky130_fd_sc_hd__inv_2
X_1707_ _1513_ _1544_ vssd1 vssd1 vccd1 vccd1 _1545_ sky130_fd_sc_hd__or2_1
X_2756_ _1458_ SB0.route_sel\[123\] vssd1 vssd1 vccd1 vccd1 _1353_ sky130_fd_sc_hd__nand2_1
X_2687_ SB0.route_sel\[80\] SB0.route_sel\[81\] vssd1 vssd1 vccd1 vccd1 _1307_ sky130_fd_sc_hd__nor2_1
XFILLER_58_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3239_ clknet_leaf_7_clk _0059_ net258 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2136__A2 _1526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1569_ SB0.route_sel\[82\] vssd1 vssd1 vccd1 vccd1 _1407_ sky130_fd_sc_hd__inv_2
X_3308_ clknet_leaf_23_clk _0128_ net272 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[0\]
+ sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_18_Left_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2086__Y _0716_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3088__A0 CB_0.config_data_inA vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2810__B1_N _0659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output111_A net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2610_ _1235_ _1236_ _1474_ vssd1 vssd1 vccd1 vccd1 _1237_ sky130_fd_sc_hd__mux2_1
X_2541_ net193 net138 vssd1 vssd1 vccd1 vccd1 _1168_ sky130_fd_sc_hd__nand2_1
Xclkload13 clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 clkload13/Y sky130_fd_sc_hd__clkinv_2
X_2472_ _1025_ _1026_ _1031_ LE_0B.config_data\[4\] vssd1 vssd1 vccd1 vccd1 _1100_
+ sky130_fd_sc_hd__o211a_1
Xclkload24 clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 clkload24/X sky130_fd_sc_hd__clkbuf_8
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_66_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3024_ SB0.route_sel\[64\] SB0.route_sel\[63\] net289 vssd1 vssd1 vccd1 vccd1 _0192_
+ sky130_fd_sc_hd__mux2_1
Xclkload7 clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 clkload7/Y sky130_fd_sc_hd__inv_6
X_2808_ _1499_ net161 _0637_ vssd1 vssd1 vccd1 vccd1 _1381_ sky130_fd_sc_hd__o21bai_4
XANTENNA_fanout142_A net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout211 net221 vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__buf_2
Xfanout200 CB_1.config_dataB\[1\] vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__buf_2
XANTENNA__2211__D1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2739_ _1438_ SB0.route_sel\[16\] _1439_ SB0.route_sel\[19\] _1341_ vssd1 vssd1 vccd1
+ vccd1 _1342_ sky130_fd_sc_hd__a221o_1
Xfanout222 net224 vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__clkbuf_4
XANTENNA__2357__A2 _0384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout277 net284 vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__clkbuf_4
Xfanout299 net300 vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__clkbuf_4
Xfanout255 net264 vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__clkbuf_4
Xfanout233 net239 vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__clkbuf_4
Xfanout244 net246 vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_29_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout266 net268 vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__clkbuf_4
Xfanout288 net302 vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__clkbuf_2
XANTENNA__2045__A1 _0670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clone17_A1 _0424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1972_ _0590_ _0596_ _0600_ _0601_ vssd1 vssd1 vccd1 vccd1 _0602_ sky130_fd_sc_hd__a211o_4
XANTENNA__1795__B1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2524_ net193 net192 vssd1 vssd1 vccd1 vccd1 _1151_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_49_Right_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2455_ CB_0.config_dataB\[13\] _1076_ _1079_ _1082_ vssd1 vssd1 vccd1 vccd1 _1083_
+ sky130_fd_sc_hd__or4_1
XANTENNA__1617__A SB0.route_sel\[120\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clone33_B1 _0981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2386_ _0539_ _0533_ _1013_ net310 vssd1 vssd1 vccd1 vccd1 _1014_ sky130_fd_sc_hd__a211o_4
XPHY_EDGE_ROW_58_Right_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3007_ SB0.route_sel\[47\] SB0.route_sel\[46\] net292 vssd1 vssd1 vccd1 vccd1 _0175_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__2630__B net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3515__Q LE_1B.config_data\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3128__S net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2171_ _0755_ _0798_ _0800_ _0757_ _0783_ vssd1 vssd1 vccd1 vccd1 _0801_ sky130_fd_sc_hd__o32a_1
X_2240_ net147 net159 LEI0.config_data\[30\] vssd1 vssd1 vccd1 vccd1 _0869_ sky130_fd_sc_hd__mux2_1
XANTENNA_clone44_C1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1886_ SB0.route_sel\[124\] SB0.route_sel\[125\] net39 vssd1 vssd1 vccd1 vccd1 _0516_
+ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_31_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1955_ _0398_ net352 net349 _1495_ _1477_ vssd1 vssd1 vccd1 vccd1 _0585_ sky130_fd_sc_hd__a221o_1
X_3487_ clknet_leaf_15_clk _0307_ net280 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[1\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__2193__A0 net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2438_ LEI0.config_data\[27\] net160 vssd1 vssd1 vccd1 vccd1 _1066_ sky130_fd_sc_hd__nand2_1
X_2507_ _1134_ LEI0.config_data\[41\] _1108_ vssd1 vssd1 vccd1 vccd1 _1135_ sky130_fd_sc_hd__a21oi_2
X_2369_ SB0.route_sel\[74\] SB0.route_sel\[75\] SB0.route_sel\[77\] _1413_ _0996_
+ vssd1 vssd1 vccd1 vccd1 _0997_ sky130_fd_sc_hd__o221a_1
XANTENNA__2248__B2 _0679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2248__A1 _0659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1809__X _0439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2487__A1 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input35_A SBsouth_in[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_6_Left_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2551__A net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1740_ _1426_ SB0.route_sel\[40\] SB0.route_sel\[45\] SB0.route_sel\[44\] _0369_
+ vssd1 vssd1 vccd1 vccd1 _0370_ sky130_fd_sc_hd__o221a_1
X_1671_ SB0.route_sel\[53\] SB0.route_sel\[52\] net61 _1507_ _1497_ vssd1 vssd1 vccd1
+ vccd1 _1509_ sky130_fd_sc_hd__a41o_1
X_3410_ clknet_leaf_19_clk _0230_ net276 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[102\]
+ sky130_fd_sc_hd__dfstp_1
X_3272_ clknet_leaf_30_clk net382 net247 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_3341_ clknet_leaf_27_clk _0161_ net252 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[33\]
+ sky130_fd_sc_hd__dfstp_1
X_2223_ _0849_ _0850_ _0851_ vssd1 vssd1 vccd1 vccd1 _0852_ sky130_fd_sc_hd__a21oi_1
X_2085_ CB_1.config_dataB\[8\] _0707_ _0711_ _0714_ CB_1.config_dataB\[9\] vssd1 vssd1
+ vccd1 vccd1 _0715_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_36_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2154_ _0757_ _0783_ vssd1 vssd1 vccd1 vccd1 _0784_ sky130_fd_sc_hd__nor2_1
XANTENNA_clone39_C1 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2987_ SB0.route_sel\[27\] SB0.route_sel\[26\] net286 vssd1 vssd1 vccd1 vccd1 _0155_
+ sky130_fd_sc_hd__mux2_1
X_1938_ _0565_ _1492_ _0566_ _0567_ vssd1 vssd1 vccd1 vccd1 _0568_ sky130_fd_sc_hd__o211a_1
X_1869_ _1540_ _0497_ vssd1 vssd1 vccd1 vccd1 _0499_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout222_A net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2181__A3 net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_32_Left_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkload0_A clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input38_X net38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2910_ net423 LE_0B.config_data\[12\] net206 vssd1 vssd1 vccd1 vccd1 _0079_ sky130_fd_sc_hd__mux2_1
X_2841_ LEI0.config_data\[9\] net486 net205 vssd1 vssd1 vccd1 vccd1 _0010_ sky130_fd_sc_hd__mux2_1
X_2772_ net153 _1021_ _0547_ vssd1 vssd1 vccd1 vccd1 _1363_ sky130_fd_sc_hd__mux2_2
X_1654_ CB_0.le_outB vssd1 vssd1 vccd1 vccd1 _1492_ sky130_fd_sc_hd__inv_6
Xhold105 LE_0A.config_data\[15\] vssd1 vssd1 vccd1 vccd1 net415 sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 LE_0B.config_data\[7\] vssd1 vssd1 vccd1 vccd1 net448 sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 LE_0B.config_data\[0\] vssd1 vssd1 vccd1 vccd1 net437 sky130_fd_sc_hd__dlygate4sd3_1
Xhold116 _0081_ vssd1 vssd1 vccd1 vccd1 net426 sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 _0332_ vssd1 vssd1 vccd1 vccd1 net459 sky130_fd_sc_hd__dlygate4sd3_1
X_1723_ SB0.route_sel\[47\] SB0.route_sel\[46\] vssd1 vssd1 vccd1 vccd1 _0353_ sky130_fd_sc_hd__nand2_1
XFILLER_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3255_ clknet_leaf_6_clk _0075_ net254 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_1585_ SB0.route_sel\[50\] vssd1 vssd1 vccd1 vccd1 _1423_ sky130_fd_sc_hd__inv_2
X_3324_ clknet_leaf_25_clk _0144_ net266 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[16\]
+ sky130_fd_sc_hd__dfstp_2
X_2206_ LEI0.config_data\[7\] _0831_ _0834_ vssd1 vssd1 vccd1 vccd1 _0835_ sky130_fd_sc_hd__o21ba_1
X_2068_ _1526_ net356 CB_1.config_dataB\[5\] vssd1 vssd1 vccd1 vccd1 _0698_ sky130_fd_sc_hd__mux2_1
X_2137_ net13 net331 CB_1.config_dataB\[15\] vssd1 vssd1 vccd1 vccd1 _0767_ sky130_fd_sc_hd__mux2_1
X_3186_ clknet_leaf_3_clk _0006_ net245 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2743__X net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1831__C1 _0460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2653__X _1280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclone61 _0487_ _0481_ _0962_ net306 vssd1 vssd1 vccd1 vccd1 net371 sky130_fd_sc_hd__a211o_1
XANTENNA__2145__A3 _0615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3040_ SB0.route_sel\[80\] SB0.route_sel\[79\] net290 vssd1 vssd1 vccd1 vccd1 _0208_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__2302__A0 net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2824_ net168 net163 _0428_ vssd1 vssd1 vccd1 vccd1 _1389_ sky130_fd_sc_hd__o21ba_4
X_1637_ CB_0.config_dataA\[14\] vssd1 vssd1 vccd1 vccd1 _1475_ sky130_fd_sc_hd__inv_2
X_1706_ CB_0.config_dataA\[24\] CB_0.config_dataA\[21\] CB_0.config_dataA\[20\] vssd1
+ vssd1 vccd1 vccd1 _1544_ sky130_fd_sc_hd__nand3b_1
X_2755_ _1352_ _0519_ vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__and2b_1
XANTENNA_clone52_C1 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2686_ _1306_ _0612_ vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__and2_4
XFILLER_64_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3238_ clknet_leaf_7_clk net402 net258 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_1568_ SB0.route_sel\[81\] vssd1 vssd1 vccd1 vccd1 _1406_ sky130_fd_sc_hd__inv_2
X_3307_ clknet_leaf_23_clk _0127_ net273 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[24\]
+ sky130_fd_sc_hd__dfstp_1
X_3169_ net435 net406 net202 vssd1 vssd1 vccd1 vccd1 _0337_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3088__A1 CB_0.config_dataA\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output104_A net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2540_ _1166_ vssd1 vssd1 vccd1 vccd1 _1167_ sky130_fd_sc_hd__inv_2
XANTENNA__3428__Q SB0.route_sel\[120\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload14 clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 clkload14/Y sky130_fd_sc_hd__bufinv_16
X_2471_ _1096_ _1097_ _1070_ vssd1 vssd1 vccd1 vccd1 _1099_ sky130_fd_sc_hd__o21ai_1
Xclkload25 clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 clkload25/X sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_66_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3023_ SB0.route_sel\[63\] SB0.route_sel\[62\] net293 vssd1 vssd1 vccd1 vccd1 _0191_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_66_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clone47_C1 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2807_ _1380_ _0594_ _0595_ vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__a21boi_2
X_2738_ SB0.route_sel\[22\] SB0.route_sel\[23\] vssd1 vssd1 vccd1 vccd1 _1341_ sky130_fd_sc_hd__nor2_1
Xclkload8 clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 clkload8/Y sky130_fd_sc_hd__bufinv_16
XFILLER_59_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2669_ _1396_ SB0.route_sel\[107\] vssd1 vssd1 vccd1 vccd1 _1295_ sky130_fd_sc_hd__nor2_1
Xfanout256 net264 vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__clkbuf_4
Xfanout234 net239 vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__buf_2
Xfanout212 net215 vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__clkbuf_4
Xfanout245 net246 vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__clkbuf_4
Xfanout201 CB_1.config_dataB\[0\] vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__clkbuf_4
Xfanout223 net224 vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__clkbuf_2
Xfanout278 net284 vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__clkbuf_2
Xfanout289 net302 vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__clkbuf_4
Xfanout267 net268 vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__clkbuf_4
XANTENNA_clone10_A net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input65_A config_data_in vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input20_X net20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2284__A2 _0543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clone17_A2 _0415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1971_ SB0.route_sel\[88\] SB0.route_sel\[89\] vssd1 vssd1 vccd1 vccd1 _0601_ sky130_fd_sc_hd__nand2_1
XANTENNA__1795__A1 _0415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2385_ _1452_ SB0.route_sel\[117\] SB0.route_sel\[114\] SB0.route_sel\[115\] _1012_
+ vssd1 vssd1 vccd1 vccd1 _1013_ sky130_fd_sc_hd__o221a_1
X_2523_ net328 _0978_ net193 vssd1 vssd1 vccd1 vccd1 _1150_ sky130_fd_sc_hd__mux2_1
X_2454_ CB_0.config_dataB\[11\] _1080_ _1081_ vssd1 vssd1 vccd1 vccd1 _1082_ sky130_fd_sc_hd__a21oi_1
XANTENNA_clone33_A1 _0367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput1 CBeast_in[0] vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__buf_6
XFILLER_28_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3006_ SB0.route_sel\[46\] SB0.route_sel\[45\] net292 vssd1 vssd1 vccd1 vccd1 _0174_
+ sky130_fd_sc_hd__mux2_1
XFILLER_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout305_X net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2824__B1_N _0428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2549__A LEI0.config_data\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1740__X _0370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2170_ _1488_ _0690_ _0722_ _0799_ vssd1 vssd1 vccd1 vccd1 _0800_ sky130_fd_sc_hd__o211a_1
X_1954_ _0580_ _0570_ _0583_ net310 vssd1 vssd1 vccd1 vccd1 _0584_ sky130_fd_sc_hd__a211o_4
XANTENNA__3293__SET_B net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2193__A1 net12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1885_ SB0.route_sel\[124\] SB0.route_sel\[125\] net55 vssd1 vssd1 vccd1 vccd1 _0515_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_31_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3486_ clknet_leaf_15_clk _0306_ net281 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_2506_ _1133_ _1110_ net239 vssd1 vssd1 vccd1 vccd1 _1134_ sky130_fd_sc_hd__a21boi_4
X_2368_ SB0.route_sel\[78\] SB0.route_sel\[79\] vssd1 vssd1 vccd1 vccd1 _0996_ sky130_fd_sc_hd__nand2b_1
X_2437_ LE_0B.config_data\[6\] LE_0B.config_data\[7\] _1032_ vssd1 vssd1 vccd1 vccd1
+ _1065_ sky130_fd_sc_hd__mux2_1
XFILLER_56_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2746__X net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2299_ _0371_ _0911_ _0914_ _0397_ _1464_ vssd1 vssd1 vccd1 vccd1 _0928_ sky130_fd_sc_hd__a221o_1
XFILLER_24_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_22_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input28_A CBnorth_in[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2088__B net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3436__Q CB_0.config_dataA\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1670_ _1424_ _1425_ net45 vssd1 vssd1 vccd1 vccd1 _1508_ sky130_fd_sc_hd__o21a_1
X_2222_ _0584_ _0842_ _0843_ _0564_ _1459_ vssd1 vssd1 vccd1 vccd1 _0851_ sky130_fd_sc_hd__a221o_1
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3271_ clknet_leaf_31_clk _0091_ net242 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_3340_ clknet_leaf_29_clk _0160_ net249 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[32\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_53_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2084_ net198 _0712_ _0713_ vssd1 vssd1 vccd1 vccd1 _0714_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_36_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2153_ _0781_ _0782_ CB_0.config_data_inA net238 vssd1 vssd1 vccd1 vccd1 _0783_ sky130_fd_sc_hd__o211a_1
XFILLER_26_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1937_ _0363_ _0501_ vssd1 vssd1 vccd1 vccd1 _0567_ sky130_fd_sc_hd__or2_1
X_2986_ SB0.route_sel\[26\] SB0.route_sel\[25\] net286 vssd1 vssd1 vccd1 vccd1 _0154_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__1913__A1 _0539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout215_A net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1868_ CB_0.config_dataB\[23\] CB_0.config_dataB\[22\] vssd1 vssd1 vccd1 vccd1 _0498_
+ sky130_fd_sc_hd__nand2_1
Xinput70 le_nrst vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__clkbuf_2
X_1799_ SB0.route_sel\[26\] SB0.route_sel\[27\] vssd1 vssd1 vccd1 vccd1 _0429_ sky130_fd_sc_hd__nand2_1
X_3469_ clknet_leaf_5_clk _0289_ net261 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[8\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_29_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_19_clk_A clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2386__X _1014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output134_A net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2771_ _1362_ _0567_ _0569_ vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_41_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2840_ net462 LEI0.config_data\[9\] net205 vssd1 vssd1 vccd1 vccd1 _0009_ sky130_fd_sc_hd__mux2_1
X_1653_ LE_0B.config_data_in vssd1 vssd1 vccd1 vccd1 _1491_ sky130_fd_sc_hd__inv_2
Xhold106 LE_1A.config_data\[12\] vssd1 vssd1 vccd1 vccd1 net416 sky130_fd_sc_hd__dlygate4sd3_1
Xhold128 LE_1A.config_data\[15\] vssd1 vssd1 vccd1 vccd1 net438 sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 LE_1A.config_data\[13\] vssd1 vssd1 vccd1 vccd1 net449 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_9_Right_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold117 LE_1B.config_data\[12\] vssd1 vssd1 vccd1 vccd1 net427 sky130_fd_sc_hd__dlygate4sd3_1
X_1722_ _0348_ _0350_ _0351_ vssd1 vssd1 vccd1 vccd1 _0352_ sky130_fd_sc_hd__a21bo_1
X_1584_ SB0.route_sel\[49\] vssd1 vssd1 vccd1 vccd1 _1422_ sky130_fd_sc_hd__inv_2
X_3185_ clknet_leaf_5_clk _0005_ net254 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_3254_ clknet_leaf_6_clk net395 net254 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_3323_ clknet_leaf_25_clk _0143_ net266 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[15\]
+ sky130_fd_sc_hd__dfstp_1
X_2205_ net303 LEI0.config_data\[8\] _0833_ vssd1 vssd1 vccd1 vccd1 _0834_ sky130_fd_sc_hd__or3_1
X_2067_ _0695_ _0696_ vssd1 vssd1 vccd1 vccd1 _0697_ sky130_fd_sc_hd__and2b_1
X_2136_ net357 net361 _1526_ net356 net195 net194 vssd1 vssd1 vccd1 vccd1 _0766_ sky130_fd_sc_hd__mux4_1
X_2969_ SB0.route_sel\[9\] SB0.route_sel\[8\] net291 vssd1 vssd1 vccd1 vccd1 _0137_
+ sky130_fd_sc_hd__mux2_1
XFILLER_57_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_4_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclone40 _0562_ _0552_ _1020_ net309 vssd1 vssd1 vccd1 vccd1 net350 sky130_fd_sc_hd__a211o_1
Xclone51 _0367_ _0358_ _0370_ net305 vssd1 vssd1 vccd1 vccd1 net361 sky130_fd_sc_hd__a211o_1
XANTENNA__2550__A1 LEI0.config_data\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1889__B1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2557__A net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3152__S net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2302__A1 net12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2605__A2 _1014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1705_ _1517_ _1541_ net30 vssd1 vssd1 vccd1 vccd1 _1543_ sky130_fd_sc_hd__o21ai_1
X_2754_ SB0.route_sel\[120\] SB0.route_sel\[121\] _1458_ SB0.route_sel\[123\] _1351_
+ vssd1 vssd1 vccd1 vccd1 _1352_ sky130_fd_sc_hd__o221a_1
X_2823_ _1388_ _0431_ _0432_ vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__a21boi_2
X_1636_ CB_0.config_dataA\[12\] vssd1 vssd1 vccd1 vccd1 _1474_ sky130_fd_sc_hd__inv_2
X_1567_ SB0.route_sel\[92\] vssd1 vssd1 vccd1 vccd1 _1405_ sky130_fd_sc_hd__inv_2
X_2685_ SB0.route_sel\[88\] _1402_ _1403_ SB0.route_sel\[91\] _1305_ vssd1 vssd1 vccd1
+ vccd1 _1306_ sky130_fd_sc_hd__a221o_1
X_3306_ clknet_leaf_23_clk _0126_ net273 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[23\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_fanout282_A net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3237_ clknet_leaf_8_clk net378 net258 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_2119_ CB_1.config_dataB\[13\] _0748_ vssd1 vssd1 vccd1 vccd1 _0749_ sky130_fd_sc_hd__nor2_1
X_3168_ net466 net435 net202 vssd1 vssd1 vccd1 vccd1 _0336_ sky130_fd_sc_hd__mux2_1
X_3099_ net189 net188 net217 vssd1 vssd1 vccd1 vccd1 _0267_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2780__A1 _1001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input10_A CBeast_in[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload15 clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 clkload15/Y sky130_fd_sc_hd__clkinv_2
Xclkload26 clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 clkload26/Y sky130_fd_sc_hd__bufinv_16
XFILLER_13_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1727__Y _0357_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2523__A1 _0978_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3147__S net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2470_ _1096_ _1097_ _1070_ vssd1 vssd1 vccd1 vccd1 _1098_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_66_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3022_ SB0.route_sel\[62\] SB0.route_sel\[61\] net293 vssd1 vssd1 vccd1 vccd1 _0190_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_clone47_B1 _0396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1798__C1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2806_ _1528_ net161 _0615_ vssd1 vssd1 vccd1 vccd1 _1380_ sky130_fd_sc_hd__o21bai_4
X_2668_ _1293_ LE_0A.config_data\[16\] _1294_ net233 vssd1 vssd1 vccd1 vccd1 CB_0.le_outA
+ sky130_fd_sc_hd__o211a_4
Xclkload9 clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 clkload9/Y sky130_fd_sc_hd__inv_6
X_2737_ _0425_ _1340_ vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__and2_4
X_2599_ _1224_ _1225_ CB_0.config_dataA\[12\] vssd1 vssd1 vccd1 vccd1 _1226_ sky130_fd_sc_hd__mux2_1
XANTENNA_input2_A CBeast_in[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout285_X net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout279 net283 vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__clkbuf_4
Xfanout213 net215 vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__clkbuf_4
X_1619_ SB0.route_sel\[126\] vssd1 vssd1 vccd1 vccd1 _1457_ sky130_fd_sc_hd__inv_2
Xfanout246 net285 vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__buf_2
Xfanout224 net225 vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__buf_2
Xfanout202 net209 vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__clkbuf_4
Xfanout268 net285 vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__clkbuf_2
Xfanout235 net236 vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__buf_2
XANTENNA__2278__A0 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2450__A0 net27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input58_A SBwest_in[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input13_X net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1970_ net35 _0598_ _0599_ vssd1 vssd1 vccd1 vccd1 _0600_ sky130_fd_sc_hd__a21oi_1
X_2522_ CB_0.config_dataA\[3\] CB_0.config_dataA\[2\] CB_0.config_dataA\[4\] _1148_
+ vssd1 vssd1 vccd1 vccd1 _1149_ sky130_fd_sc_hd__or4bb_1
XANTENNA__1795__A2 _0424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2384_ SB0.route_sel\[118\] SB0.route_sel\[119\] vssd1 vssd1 vccd1 vccd1 _1012_ sky130_fd_sc_hd__nand2b_1
X_2453_ net343 _1071_ _1074_ net342 _1468_ vssd1 vssd1 vccd1 vccd1 _1081_ sky130_fd_sc_hd__a221o_1
XANTENNA_clone33_A2 _0358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput2 CBeast_in[10] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__buf_2
XFILLER_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3005_ SB0.route_sel\[45\] SB0.route_sel\[44\] net292 vssd1 vssd1 vccd1 vccd1 _0173_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_34_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input5_X net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1830__Y _0460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2423__A0 _0956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2549__B net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1953_ SB0.route_sel\[104\] _1395_ SB0.route_sel\[109\] SB0.route_sel\[108\] _0582_
+ vssd1 vssd1 vccd1 vccd1 _0583_ sky130_fd_sc_hd__o221a_1
X_1884_ SB0.route_sel\[126\] net136 vssd1 vssd1 vccd1 vccd1 _0514_ sky130_fd_sc_hd__nand2_1
X_2505_ CB_0.config_dataB\[18\] _1118_ _1121_ _1132_ vssd1 vssd1 vccd1 vccd1 _1133_
+ sky130_fd_sc_hd__a31o_1
X_3485_ clknet_leaf_13_clk _0305_ net278 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[24\]
+ sky130_fd_sc_hd__dfstp_2
XANTENNA__2193__A2 net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clone44_A1 _0539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2367_ net341 net338 net185 vssd1 vssd1 vccd1 vccd1 _0995_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_39_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2436_ LEI0.config_data\[17\] net233 _1062_ _1037_ vssd1 vssd1 vccd1 vccd1 _1064_
+ sky130_fd_sc_hd__a31o_1
XFILLER_29_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2298_ _1526_ _1552_ net171 vssd1 vssd1 vccd1 vccd1 _0927_ sky130_fd_sc_hd__mux2_1
XANTENNA__2350__C1 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout150_X net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1841__X _0471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output89_A net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2221_ net175 _0543_ net174 vssd1 vssd1 vccd1 vccd1 _0850_ sky130_fd_sc_hd__o21a_1
XFILLER_38_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2152_ CB_1.config_dataB\[18\] _1486_ CB_1.config_dataB\[19\] _0760_ vssd1 vssd1
+ vccd1 vccd1 _0782_ sky130_fd_sc_hd__and4b_1
X_3270_ clknet_leaf_31_clk _0090_ net242 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2635__A0 net20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2083_ net362 _0692_ _0694_ net348 CB_1.config_dataB\[7\] vssd1 vssd1 vccd1 vccd1
+ _0713_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_36_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1936_ _0360_ _0498_ net21 vssd1 vssd1 vccd1 vccd1 _0566_ sky130_fd_sc_hd__o21ai_1
X_1867_ CB_0.config_dataB\[23\] CB_0.config_dataB\[22\] vssd1 vssd1 vccd1 vccd1 _0497_
+ sky130_fd_sc_hd__and2_1
X_2985_ SB0.route_sel\[25\] SB0.route_sel\[24\] net286 vssd1 vssd1 vccd1 vccd1 _0153_
+ sky130_fd_sc_hd__mux2_1
Xinput71 nrst vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__clkbuf_1
XANTENNA__1913__A2 _0533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3468_ clknet_leaf_5_clk _0288_ net256 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[7\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_fanout208_A net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput60 SBwest_in[5] vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__buf_1
X_1798_ _0424_ _0415_ _0427_ net303 vssd1 vssd1 vccd1 vccd1 _0428_ sky130_fd_sc_hd__a211o_4
X_2419_ net183 net321 CB_0.config_dataB\[6\] vssd1 vssd1 vccd1 vccd1 _1047_ sky130_fd_sc_hd__o21a_1
XANTENNA__2626__A0 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3399_ clknet_leaf_27_clk _0219_ net269 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[91\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__2323__C1 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input40_A SBsouth_in[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output127_A net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2770_ net153 _1018_ _0565_ vssd1 vssd1 vccd1 vccd1 _1362_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_41_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1721_ net148 _1501_ _0349_ net235 vssd1 vssd1 vccd1 vccd1 _0351_ sky130_fd_sc_hd__o31a_1
Xhold129 LE_0B.config_data\[4\] vssd1 vssd1 vccd1 vccd1 net439 sky130_fd_sc_hd__dlygate4sd3_1
X_3322_ clknet_leaf_25_clk _0142_ net266 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[14\]
+ sky130_fd_sc_hd__dfstp_1
Xhold107 _0098_ vssd1 vssd1 vccd1 vccd1 net417 sky130_fd_sc_hd__dlygate4sd3_1
X_1652_ LE_1B.config_data\[11\] vssd1 vssd1 vccd1 vccd1 _1490_ sky130_fd_sc_hd__inv_2
Xhold118 _0343_ vssd1 vssd1 vccd1 vccd1 net428 sky130_fd_sc_hd__dlygate4sd3_1
X_1583_ SB0.route_sel\[60\] vssd1 vssd1 vccd1 vccd1 _1421_ sky130_fd_sc_hd__inv_2
X_3184_ clknet_leaf_6_clk _0004_ net254 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_3253_ clknet_leaf_6_clk _0073_ net254 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_2135_ CB_1.config_dataB\[16\] _0763_ _0764_ vssd1 vssd1 vccd1 vccd1 _0765_ sky130_fd_sc_hd__a21oi_1
X_2204_ LEI0.config_data\[6\] net147 _0832_ LEI0.config_data\[7\] vssd1 vssd1 vccd1
+ vccd1 _0833_ sky130_fd_sc_hd__o211a_1
XANTENNA__2608__A0 net20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2066_ net345 net359 net327 net344 net199 net198 vssd1 vssd1 vccd1 vccd1 _0696_ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout158_A net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1919_ _0389_ _0501_ vssd1 vssd1 vccd1 vccd1 _0549_ sky130_fd_sc_hd__or2_1
X_2899_ net437 net431 net206 vssd1 vssd1 vccd1 vccd1 _0068_ sky130_fd_sc_hd__mux2_1
X_2968_ SB0.route_sel\[8\] SB0.route_sel\[7\] net291 vssd1 vssd1 vccd1 vccd1 _0136_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_55_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2311__A2 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclone52 _0655_ _0649_ _0658_ net307 vssd1 vssd1 vccd1 vccd1 net362 sky130_fd_sc_hd__a211o_1
XANTENNA__2302__A2 net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1704_ _1516_ _1540_ vssd1 vssd1 vccd1 vccd1 _1542_ sky130_fd_sc_hd__nand2_1
X_2753_ _1456_ SB0.route_sel\[125\] vssd1 vssd1 vccd1 vccd1 _1351_ sky130_fd_sc_hd__nand2_1
X_2684_ SB0.route_sel\[94\] SB0.route_sel\[95\] vssd1 vssd1 vccd1 vccd1 _1305_ sky130_fd_sc_hd__nor2_1
X_2822_ net167 net163 _0449_ vssd1 vssd1 vccd1 vccd1 _1388_ sky130_fd_sc_hd__o21bai_4
X_1635_ CB_0.config_dataA\[9\] vssd1 vssd1 vccd1 vccd1 _1473_ sky130_fd_sc_hd__inv_2
XANTENNA_clone52_A1 _0655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1566_ SB0.route_sel\[91\] vssd1 vssd1 vccd1 vccd1 _1404_ sky130_fd_sc_hd__inv_2
X_3305_ clknet_leaf_23_clk _0125_ net273 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[22\]
+ sky130_fd_sc_hd__dfstp_1
X_3098_ CB_0.config_dataA\[9\] net189 net217 vssd1 vssd1 vccd1 vccd1 _0266_ sky130_fd_sc_hd__mux2_1
X_3236_ clknet_leaf_8_clk _0056_ net258 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout275_A net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2118_ _0746_ _0747_ CB_1.config_dataB\[12\] vssd1 vssd1 vccd1 vccd1 _0748_ sky130_fd_sc_hd__mux2_1
X_2049_ _0675_ _0665_ _0678_ net309 vssd1 vssd1 vccd1 vccd1 _0679_ sky130_fd_sc_hd__a211o_4
X_3167_ net470 net466 net202 vssd1 vssd1 vccd1 vccd1 _0335_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_18_clk_A clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload16 clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 clkload16/Y sky130_fd_sc_hd__inv_8
Xclkload27 clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 clkload27/Y sky130_fd_sc_hd__clkinvlp_4
XANTENNA__2332__S CB_0.config_dataB\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_41_Left_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2680__X net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_50_Left_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3021_ SB0.route_sel\[61\] SB0.route_sel\[60\] net296 vssd1 vssd1 vccd1 vccd1 _0189_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_clone47_A1 _0393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2805_ _1379_ _0555_ _0556_ vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__a21boi_2
XANTENNA__1798__B1 _0427_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1618_ SB0.route_sel\[124\] vssd1 vssd1 vccd1 vccd1 _1456_ sky130_fd_sc_hd__inv_2
XANTENNA__1934__X _0564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2667_ LE_0A.dff_out LE_0A.config_data\[16\] vssd1 vssd1 vccd1 vccd1 _1294_ sky130_fd_sc_hd__nand2b_1
X_2736_ SB0.route_sel\[18\] _1440_ SB0.route_sel\[21\] _1441_ _1339_ vssd1 vssd1 vccd1
+ vccd1 _1340_ sky130_fd_sc_hd__a221o_1
X_2598_ net27 net28 net29 net30 net189 net188 vssd1 vssd1 vccd1 vccd1 _1225_ sky130_fd_sc_hd__mux4_1
Xfanout258 net260 vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__clkbuf_4
Xfanout214 net215 vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__clkbuf_4
Xfanout225 net231 vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__buf_2
Xfanout269 net271 vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__clkbuf_4
Xfanout236 net238 vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__buf_2
X_3219_ clknet_leaf_3_clk _0039_ net245 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[39\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2749__Y net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout247 net248 vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__clkbuf_4
XANTENNA__2278__A1 net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout203 net209 vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__clkbuf_2
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3501__SET_B net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1789__B1 net25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2450__A1 net28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2521_ net192 net193 vssd1 vssd1 vccd1 vccd1 _1148_ sky130_fd_sc_hd__and2b_1
XANTENNA__1754__X _0384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2452_ net328 net347 CB_0.config_dataB\[10\] vssd1 vssd1 vccd1 vccd1 _1080_ sky130_fd_sc_hd__mux2_1
X_2383_ net185 _1010_ vssd1 vssd1 vccd1 vccd1 _1011_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_18_Right_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput3 CBeast_in[11] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_27_Right_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3004_ SB0.route_sel\[44\] SB0.route_sel\[43\] net292 vssd1 vssd1 vccd1 vccd1 _0172_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout238_A net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2196__A0 _0428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_36_Right_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2719_ _1328_ _0368_ vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__and2_4
XFILLER_59_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_45_Right_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_54_Right_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1934__B1 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input70_A le_nrst vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_63_Right_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1952_ SB0.route_sel\[111\] SB0.route_sel\[110\] vssd1 vssd1 vccd1 vccd1 _0582_ sky130_fd_sc_hd__nand2b_1
XFILLER_33_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1883_ _0509_ _0511_ _0512_ vssd1 vssd1 vccd1 vccd1 _0513_ sky130_fd_sc_hd__a21bo_1
X_3484_ clknet_leaf_13_clk _0304_ net278 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[23\]
+ sky130_fd_sc_hd__dfstp_2
X_2504_ _1131_ _1128_ _1124_ CB_0.config_dataB\[19\] vssd1 vssd1 vccd1 vccd1 _1132_
+ sky130_fd_sc_hd__a31o_1
XANTENNA_clone44_A2 _0533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2435_ LEI0.config_data\[17\] net233 _1062_ _1037_ vssd1 vssd1 vccd1 vccd1 _1063_
+ sky130_fd_sc_hd__a31oi_4
XFILLER_56_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2366_ _0611_ _0602_ _0993_ net307 vssd1 vssd1 vccd1 vccd1 _0994_ sky130_fd_sc_hd__a211o_4
X_2297_ _0916_ _0919_ _0922_ _0925_ vssd1 vssd1 vccd1 vccd1 _0926_ sky130_fd_sc_hd__a22o_1
XANTENNA__2350__B1 _0977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1861__C1 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout143_X net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout310_X net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2332__A0 _0956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2220_ net175 _0521_ vssd1 vssd1 vccd1 vccd1 _0849_ sky130_fd_sc_hd__nand2_1
X_2082_ _0615_ net312 _1480_ vssd1 vssd1 vccd1 vccd1 _0712_ sky130_fd_sc_hd__mux2_1
XFILLER_38_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2151_ CB_1.config_dataB\[17\] _0770_ _0780_ vssd1 vssd1 vccd1 vccd1 _0781_ sky130_fd_sc_hd__a21oi_1
XANTENNA__2635__A1 net22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clone39_A2 _0570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2399__A0 net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2984_ SB0.route_sel\[24\] SB0.route_sel\[23\] net286 vssd1 vssd1 vccd1 vccd1 _0152_
+ sky130_fd_sc_hd__mux2_1
X_1935_ _0359_ _0497_ vssd1 vssd1 vccd1 vccd1 _0565_ sky130_fd_sc_hd__nand2_1
X_1866_ SB0.route_sel\[124\] SB0.route_sel\[125\] _1457_ net136 _0495_ vssd1 vssd1
+ vccd1 vccd1 _0496_ sky130_fd_sc_hd__o221a_1
XANTENNA__1655__A net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput50 SBwest_in[10] vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__buf_1
X_1797_ _1438_ SB0.route_sel\[16\] SB0.route_sel\[21\] SB0.route_sel\[20\] _0426_
+ vssd1 vssd1 vccd1 vccd1 _0427_ sky130_fd_sc_hd__o221a_1
Xinput61 SBwest_in[6] vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__buf_1
X_2418_ CB_0.config_dataB\[5\] _1010_ vssd1 vssd1 vccd1 vccd1 _1046_ sky130_fd_sc_hd__nand2_1
X_3467_ clknet_leaf_5_clk _0287_ net264 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[6\]
+ sky130_fd_sc_hd__dfstp_1
X_3398_ clknet_leaf_26_clk _0218_ net270 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[90\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__2626__A1 net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2349_ SB0.route_sel\[58\] SB0.route_sel\[59\] SB0.route_sel\[61\] _1421_ _0976_
+ vssd1 vssd1 vccd1 vccd1 _0977_ sky130_fd_sc_hd__o221a_1
XPHY_EDGE_ROW_0_Right_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2013__X _0643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input33_A SBsouth_in[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2683__X net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2093__A2 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold108 LE_0A.config_data\[13\] vssd1 vssd1 vccd1 vccd1 net418 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_41_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1651_ LE_1B.config_data\[10\] vssd1 vssd1 vccd1 vccd1 _1489_ sky130_fd_sc_hd__inv_2
X_1720_ net157 net169 net166 _0349_ _1501_ vssd1 vssd1 vccd1 vccd1 _0350_ sky130_fd_sc_hd__o32a_1
X_3252_ clknet_leaf_5_clk _0072_ net254 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_3321_ clknet_leaf_25_clk _0141_ net266 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[13\]
+ sky130_fd_sc_hd__dfstp_1
X_1582_ SB0.route_sel\[59\] vssd1 vssd1 vccd1 vccd1 _1420_ sky130_fd_sc_hd__inv_2
Xhold119 LE_1B.config_data\[15\] vssd1 vssd1 vccd1 vccd1 net429 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2608__A1 net22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3183_ clknet_leaf_6_clk _0003_ net254 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_2065_ net1 net8 net9 net330 net199 net198 vssd1 vssd1 vccd1 vccd1 _0695_ sky130_fd_sc_hd__mux4_1
X_2134_ net5 _0760_ _0761_ net4 _1485_ vssd1 vssd1 vccd1 vccd1 _0764_ sky130_fd_sc_hd__a221o_1
X_2203_ LEI0.config_data\[6\] net160 vssd1 vssd1 vccd1 vccd1 _0832_ sky130_fd_sc_hd__nand2_1
XFILLER_34_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2967_ SB0.route_sel\[7\] SB0.route_sel\[6\] net291 vssd1 vssd1 vccd1 vccd1 _0135_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout220_A net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1918_ _0386_ _0498_ net20 vssd1 vssd1 vccd1 vccd1 _0548_ sky130_fd_sc_hd__o21ai_1
X_2898_ net465 net437 net206 vssd1 vssd1 vccd1 vccd1 _0067_ sky130_fd_sc_hd__mux2_1
X_1849_ _0472_ _0478_ vssd1 vssd1 vccd1 vccd1 _0479_ sky130_fd_sc_hd__nand2_1
X_3519_ clknet_leaf_32_clk net414 net240 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2311__A3 _0938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1672__X _1510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclone31 _0633_ _0627_ _0990_ net307 vssd1 vssd1 vccd1 vccd1 net341 sky130_fd_sc_hd__a211o_1
XFILLER_43_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclone20 CBeast_in[3] vssd1 vssd1 vccd1 vccd1 net330 sky130_fd_sc_hd__clkbuf_1
Xclone42 _0562_ _0552_ net308 _0546_ vssd1 vssd1 vccd1 vccd1 net352 sky130_fd_sc_hd__a211o_1
XANTENNA__3024__A1 SB0.route_sel\[63\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_20_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__3451__SET_B net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2822__B1_N _0449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input36_X net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2302__A3 net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2821_ _1387_ _0376_ _0377_ vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__a21boi_2
XFILLER_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1703_ CB_0.config_dataB\[24\] CB_0.config_dataB\[20\] CB_0.config_dataB\[21\] vssd1
+ vssd1 vccd1 vccd1 _1541_ sky130_fd_sc_hd__nand3b_2
X_1634_ CB_0.config_dataA\[7\] vssd1 vssd1 vccd1 vccd1 _1472_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_11_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_clone52_A2 _0649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2683_ _1304_ _0612_ vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__and2_4
X_2752_ _0468_ _1350_ vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__and2_4
X_3235_ clknet_leaf_8_clk _0055_ net260 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__3299__SET_B net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1565_ SB0.route_sel\[90\] vssd1 vssd1 vccd1 vccd1 _1403_ sky130_fd_sc_hd__inv_2
X_3304_ clknet_leaf_23_clk _0124_ net273 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[21\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__2483__B net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3097_ CB_0.config_dataA\[8\] CB_0.config_dataA\[9\] net217 vssd1 vssd1 vccd1 vccd1
+ _0265_ sky130_fd_sc_hd__mux2_1
X_2117_ net11 net12 net13 net331 net197 net196 vssd1 vssd1 vccd1 vccd1 _0747_ sky130_fd_sc_hd__mux4_1
X_2048_ _1414_ SB0.route_sel\[64\] SB0.route_sel\[69\] SB0.route_sel\[68\] _0677_
+ vssd1 vssd1 vccd1 vccd1 _0678_ sky130_fd_sc_hd__o221a_1
XANTENNA__2057__A2 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3166_ net467 LE_1B.config_data\[3\] net202 vssd1 vssd1 vccd1 vccd1 _0334_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout268_A net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2765__A0 CB_0.le_outB vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload28 clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 clkload28/Y sky130_fd_sc_hd__clkinv_2
Xclkload17 clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 clkload17/Y sky130_fd_sc_hd__inv_8
XTAP_TAPCELL_ROW_66_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3020_ SB0.route_sel\[60\] SB0.route_sel\[59\] net296 vssd1 vssd1 vccd1 vccd1 _0188_
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_0_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_clone47_A2 _0384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2804_ net165 net162 _0564_ vssd1 vssd1 vccd1 vccd1 _1379_ sky130_fd_sc_hd__o21bai_1
XANTENNA__1798__A1 _0424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2597_ net17 net24 net25 net26 net189 net188 vssd1 vssd1 vccd1 vccd1 _1224_ sky130_fd_sc_hd__mux4_1
X_2666_ _1283_ _1288_ _1292_ _1248_ _1284_ vssd1 vssd1 vccd1 vccd1 _1293_ sky130_fd_sc_hd__a32o_2
X_1617_ SB0.route_sel\[120\] vssd1 vssd1 vccd1 vccd1 _1455_ sky130_fd_sc_hd__inv_2
XANTENNA__1970__A1 net35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout204 net209 vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__clkbuf_4
X_2735_ SB0.route_sel\[17\] SB0.route_sel\[16\] vssd1 vssd1 vccd1 vccd1 _1339_ sky130_fd_sc_hd__nor2_1
Xfanout259 net260 vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__clkbuf_4
Xfanout226 net228 vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__clkbuf_4
Xfanout215 net221 vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__clkbuf_2
Xfanout237 net238 vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__buf_2
X_3218_ clknet_leaf_4_clk _0038_ net256 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[38\]
+ sky130_fd_sc_hd__dfrtp_1
X_3149_ net173 net172 net225 vssd1 vssd1 vccd1 vccd1 _0317_ sky130_fd_sc_hd__mux2_1
Xfanout248 net250 vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__clkbuf_4
XANTENNA__2450__A2 net29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1860__X _0490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2269__A2 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output102_A net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2977__A0 SB0.route_sel\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2451_ _1077_ _1078_ CB_0.config_dataB\[12\] vssd1 vssd1 vccd1 vccd1 _1079_ sky130_fd_sc_hd__mux2_1
X_2520_ _1146_ LE_0B.config_data\[16\] _1147_ net233 vssd1 vssd1 vccd1 vccd1 CB_0.le_outB
+ sky130_fd_sc_hd__o211a_4
Xinput4 CBeast_in[12] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__buf_2
X_2382_ _0506_ _0518_ _1009_ net309 vssd1 vssd1 vccd1 vccd1 _1010_ sky130_fd_sc_hd__a211oi_4
XANTENNA_clkbuf_leaf_17_clk_A clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3003_ SB0.route_sel\[43\] SB0.route_sel\[42\] net288 vssd1 vssd1 vccd1 vccd1 _0171_
+ sky130_fd_sc_hd__mux2_1
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_2_1__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_2_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_36_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout300_A net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2196__A1 _0449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2718_ SB0.route_sel\[42\] _1428_ SB0.route_sel\[45\] _1429_ _1327_ vssd1 vssd1 vccd1
+ vccd1 _1328_ sky130_fd_sc_hd__a221o_1
XFILLER_59_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2649_ _0985_ _1259_ _1260_ _0982_ _1476_ vssd1 vssd1 vccd1 vccd1 _1276_ sky130_fd_sc_hd__a221o_1
XFILLER_59_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1855__X _0485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1934__A1 _0562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input63_A SBwest_in[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2686__X net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1870__B1 net23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1951_ _0570_ net318 net309 vssd1 vssd1 vccd1 vccd1 _0581_ sky130_fd_sc_hd__a21oi_4
X_1882_ net149 _1530_ _0510_ net236 vssd1 vssd1 vccd1 vccd1 _0512_ sky130_fd_sc_hd__o31a_1
X_3483_ clknet_leaf_13_clk _0303_ net277 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[22\]
+ sky130_fd_sc_hd__dfstp_2
X_2503_ _1129_ net178 _1130_ vssd1 vssd1 vccd1 vccd1 _1131_ sky130_fd_sc_hd__a21o_1
X_2434_ _1467_ _1050_ _1060_ _1061_ vssd1 vssd1 vccd1 vccd1 _1062_ sky130_fd_sc_hd__a31o_1
X_2365_ SB0.route_sel\[90\] SB0.route_sel\[91\] SB0.route_sel\[93\] _1405_ _0992_
+ vssd1 vssd1 vccd1 vccd1 _0993_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_39_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2296_ CB_1.config_dataA\[16\] _0923_ _0924_ vssd1 vssd1 vccd1 vccd1 _0925_ sky130_fd_sc_hd__a21oi_1
XANTENNA__2350__A1 _1548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1861__B1 _0490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout250_A net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2169__A1 _0683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout303_X net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input66_X net66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2580__A1 _0963_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2580__B2 _0966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clone2_C1 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2081_ _0710_ vssd1 vssd1 vccd1 vccd1 _0711_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_36_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2150_ _1486_ _0779_ CB_1.config_dataB\[19\] vssd1 vssd1 vccd1 vccd1 _0780_ sky130_fd_sc_hd__a21o_1
XANTENNA__2096__A0 net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2635__A2 net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1934_ _0562_ _0552_ net308 _0546_ vssd1 vssd1 vccd1 vccd1 _0564_ sky130_fd_sc_hd__a211o_4
X_2983_ SB0.route_sel\[23\] SB0.route_sel\[22\] net286 vssd1 vssd1 vccd1 vccd1 _0151_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__1843__B1 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1865_ _1455_ SB0.route_sel\[121\] vssd1 vssd1 vccd1 vccd1 _0495_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_26_Left_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput51 SBwest_in[11] vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__buf_1
Xinput40 SBsouth_in[1] vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__clkbuf_1
X_1796_ SB0.route_sel\[23\] SB0.route_sel\[22\] vssd1 vssd1 vccd1 vccd1 _0426_ sky130_fd_sc_hd__nand2b_1
Xinput62 SBwest_in[7] vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout298_A net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2417_ _1043_ _1044_ _1466_ vssd1 vssd1 vccd1 vccd1 _1045_ sky130_fd_sc_hd__mux2_1
X_3466_ clknet_leaf_5_clk _0286_ net264 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[5\]
+ sky130_fd_sc_hd__dfstp_1
X_3397_ clknet_leaf_26_clk _0217_ net269 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[89\]
+ sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_10_Left_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2348_ SB0.route_sel\[62\] SB0.route_sel\[63\] vssd1 vssd1 vccd1 vccd1 _0976_ sky130_fd_sc_hd__nand2b_1
X_2279_ net143 net155 LEI0.config_data\[42\] vssd1 vssd1 vccd1 vccd1 _0908_ sky130_fd_sc_hd__mux2_1
XFILLER_52_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input26_A CBnorth_in[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2078__A0 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3474__SET_B net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2617__A2 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2093__A3 _0716_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output94_A net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2351__S CB_0.config_dataB\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold109 LE_0A.config_data\[9\] vssd1 vssd1 vccd1 vccd1 net419 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2002__B1 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2250__A0 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1650_ LE_1B.config_data\[9\] vssd1 vssd1 vccd1 vccd1 _1488_ sky130_fd_sc_hd__inv_2
X_1581_ SB0.route_sel\[58\] vssd1 vssd1 vccd1 vccd1 _1419_ sky130_fd_sc_hd__inv_2
X_3182_ clknet_leaf_6_clk _0002_ net255 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_3251_ clknet_leaf_3_clk net397 net246 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_3320_ clknet_leaf_25_clk _0140_ net266 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[12\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__2305__A1 _0491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2305__B2 _0471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2202_ net326 net155 LEI0.config_data\[6\] vssd1 vssd1 vccd1 vccd1 _0831_ sky130_fd_sc_hd__mux2_1
XANTENNA__2608__A2 net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2064_ net199 net198 vssd1 vssd1 vccd1 vccd1 _0694_ sky130_fd_sc_hd__nor2_1
X_2133_ net6 net7 CB_1.config_dataB\[15\] vssd1 vssd1 vccd1 vccd1 _0763_ sky130_fd_sc_hd__mux2_1
XANTENNA__1816__B1 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1917_ _0385_ _0497_ vssd1 vssd1 vccd1 vccd1 _0547_ sky130_fd_sc_hd__nand2_1
X_2897_ LE_0B.dff_out _1146_ net69 vssd1 vssd1 vccd1 vccd1 _0066_ sky130_fd_sc_hd__mux2_1
X_2966_ SB0.route_sel\[6\] SB0.route_sel\[5\] net291 vssd1 vssd1 vccd1 vccd1 _0134_
+ sky130_fd_sc_hd__mux2_1
X_3518_ clknet_leaf_32_clk net407 net240 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_1848_ SB0.route_sel\[13\] SB0.route_sel\[12\] net40 vssd1 vssd1 vccd1 vccd1 _0478_
+ sky130_fd_sc_hd__a21bo_1
X_1779_ net157 net168 net163 _0407_ _1502_ vssd1 vssd1 vccd1 vccd1 _0409_ sky130_fd_sc_hd__o32ai_2
X_3449_ clknet_leaf_9_clk _0269_ net263 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[13\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_4_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclone21 CBeast_in[7] vssd1 vssd1 vccd1 vccd1 net331 sky130_fd_sc_hd__clkbuf_1
Xclone32 _0393_ _0384_ _0984_ net305 vssd1 vssd1 vccd1 vccd1 net342 sky130_fd_sc_hd__a211o_1
Xclone10 net150 vssd1 vssd1 vccd1 vccd1 net320 sky130_fd_sc_hd__buf_6
XANTENNA__2535__B2 _1001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2535__A1 _0998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input29_X net29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output132_A net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2751_ _1446_ SB0.route_sel\[0\] _1447_ SB0.route_sel\[3\] _1349_ vssd1 vssd1 vccd1
+ vccd1 _1350_ sky130_fd_sc_hd__a221o_1
X_2820_ net169 net165 _0397_ vssd1 vssd1 vccd1 vccd1 _1387_ sky130_fd_sc_hd__o21bai_4
X_1633_ CB_0.config_dataA\[8\] vssd1 vssd1 vccd1 vccd1 _1471_ sky130_fd_sc_hd__inv_2
X_1702_ CB_0.config_dataB\[24\] CB_0.config_dataB\[20\] CB_0.config_dataB\[21\] vssd1
+ vssd1 vccd1 vccd1 _1540_ sky130_fd_sc_hd__and3b_1
XANTENNA__2774__A1 _0994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2682_ SB0.route_sel\[90\] _1404_ SB0.route_sel\[93\] _1405_ _1303_ vssd1 vssd1 vccd1
+ vccd1 _1304_ sky130_fd_sc_hd__a221o_1
X_1564_ SB0.route_sel\[89\] vssd1 vssd1 vccd1 vccd1 _1402_ sky130_fd_sc_hd__inv_2
XFILLER_66_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3234_ clknet_leaf_8_clk _0054_ net258 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_3303_ clknet_leaf_23_clk _0123_ net273 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[20\]
+ sky130_fd_sc_hd__dfstp_1
X_3165_ net460 LE_1B.config_data\[2\] net202 vssd1 vssd1 vccd1 vccd1 _0333_ sky130_fd_sc_hd__mux2_1
X_3096_ CB_0.config_dataA\[7\] CB_0.config_dataA\[8\] net217 vssd1 vssd1 vccd1 vccd1
+ _0264_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2047_ SB0.route_sel\[71\] SB0.route_sel\[70\] vssd1 vssd1 vccd1 vccd1 _0677_ sky130_fd_sc_hd__nand2b_1
X_2116_ net1 net8 net9 net330 net197 net196 vssd1 vssd1 vccd1 vccd1 _0746_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_60_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2949_ CB_1.config_dataB\[13\] CB_1.config_dataB\[14\] net230 vssd1 vssd1 vccd1 vccd1
+ _0117_ sky130_fd_sc_hd__mux2_1
XANTENNA__3087__S net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1827__C net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1683__X _1521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2019__X _0649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_13_Left_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload29 clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 clkload29/Y sky130_fd_sc_hd__bufinv_16
Xclkload18 clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 clkload18/Y sky130_fd_sc_hd__clkinv_8
XANTENNA__2689__X net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2803_ _1378_ _0573_ _0574_ vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__a21boi_2
X_2734_ _1338_ _0446_ vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__nor2_4
XANTENNA__1798__A2 _0415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout227 net228 vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__clkbuf_2
Xfanout216 net218 vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__clkbuf_4
X_1616_ SB0.route_sel\[114\] vssd1 vssd1 vccd1 vccd1 _1454_ sky130_fd_sc_hd__inv_2
X_2596_ net188 _1219_ _1222_ vssd1 vssd1 vccd1 vccd1 _1223_ sky130_fd_sc_hd__a21oi_1
X_2665_ _1212_ _1289_ _1291_ _1245_ vssd1 vssd1 vccd1 vccd1 _1292_ sky130_fd_sc_hd__a211o_1
Xfanout238 net239 vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__clkbuf_2
Xfanout205 net209 vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout280_A net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3217_ clknet_leaf_4_clk _0037_ net261 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[37\]
+ sky130_fd_sc_hd__dfrtp_1
X_3148_ CB_1.config_dataA\[9\] CB_1.config_dataA\[10\] net229 vssd1 vssd1 vccd1 vccd1
+ _0316_ sky130_fd_sc_hd__mux2_1
Xfanout249 net250 vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__clkbuf_4
X_3079_ SB0.route_sel\[119\] SB0.route_sel\[118\] net300 vssd1 vssd1 vccd1 vccd1 _0247_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__2781__Y net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2450__A3 net30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2426__A0 net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2269__A3 _0897_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2977__A1 SB0.route_sel\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2450_ net27 net28 net29 net30 net181 CB_0.config_dataB\[11\] vssd1 vssd1 vccd1 vccd1
+ _1078_ sky130_fd_sc_hd__mux4_1
X_2381_ _1456_ SB0.route_sel\[125\] SB0.route_sel\[122\] SB0.route_sel\[123\] _1008_
+ vssd1 vssd1 vccd1 vccd1 _1009_ sky130_fd_sc_hd__o221a_1
XFILLER_5_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput5 CBeast_in[13] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__buf_2
XANTENNA__1815__C_N _0438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3002_ SB0.route_sel\[42\] SB0.route_sel\[41\] net288 vssd1 vssd1 vccd1 vccd1 _0170_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_62_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1674__A _1511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2717_ SB0.route_sel\[41\] SB0.route_sel\[40\] vssd1 vssd1 vccd1 vccd1 _1327_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout283_X net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2648_ _0975_ _0978_ net187 vssd1 vssd1 vccd1 vccd1 _1275_ sky130_fd_sc_hd__mux2_1
X_2579_ _0956_ _0959_ CB_0.config_dataA\[5\] vssd1 vssd1 vccd1 vccd1 _1206_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_25_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1934__A2 _0552_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input56_A SBwest_in[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input11_X net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1950_ _0575_ _0571_ _0579_ _1395_ _1394_ vssd1 vssd1 vccd1 vccd1 _0580_ sky130_fd_sc_hd__a2111o_1
XPHY_EDGE_ROW_38_Left_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2502_ net343 _1109_ _1113_ net342 _1469_ vssd1 vssd1 vccd1 vccd1 _1130_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_47_Left_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1881_ net158 net167 net162 _0510_ _1530_ vssd1 vssd1 vccd1 vccd1 _0511_ sky130_fd_sc_hd__o32a_1
X_3482_ clknet_leaf_13_clk _0302_ net277 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[21\]
+ sky130_fd_sc_hd__dfstp_2
X_2433_ CB_0.config_dataB\[8\] _1466_ CB_0.config_dataB\[9\] _1040_ vssd1 vssd1 vccd1
+ vccd1 _1061_ sky130_fd_sc_hd__and4b_1
X_2364_ SB0.route_sel\[94\] SB0.route_sel\[95\] vssd1 vssd1 vccd1 vccd1 _0992_ sky130_fd_sc_hd__nand2b_1
XANTENNA__2335__C1 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2350__A2 _1539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2638__A0 net31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_56_Left_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2295_ net16 _0911_ _0914_ net15 CB_1.config_dataA\[17\] vssd1 vssd1 vccd1 vccd1
+ _0924_ sky130_fd_sc_hd__a221o_1
XANTENNA__1861__A1 _0487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_10 _0415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout243_A net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_65_Left_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input3_X net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_0__f_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_16_clk_A clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input59_X net59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2635__A3 net23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2080_ _0708_ _0709_ _1479_ vssd1 vssd1 vccd1 vccd1 _0710_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1933_ _0552_ _0562_ net308 vssd1 vssd1 vccd1 vccd1 _0563_ sky130_fd_sc_hd__a21oi_2
X_2982_ SB0.route_sel\[22\] SB0.route_sel\[21\] net286 vssd1 vssd1 vccd1 vccd1 _0150_
+ sky130_fd_sc_hd__mux2_1
Xinput30 CBnorth_in[7] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__buf_2
X_3465_ clknet_leaf_5_clk _0285_ net264 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[4\]
+ sky130_fd_sc_hd__dfstp_1
X_1864_ CB_1.config_dataB\[3\] _0403_ _0400_ _0493_ vssd1 vssd1 vccd1 vccd1 _0494_
+ sky130_fd_sc_hd__or4_4
Xinput52 SBwest_in[12] vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__buf_1
Xinput41 SBsouth_in[2] vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__buf_1
Xinput63 SBwest_in[8] vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__buf_1
X_1795_ _0415_ _0424_ net303 vssd1 vssd1 vccd1 vccd1 _0425_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout193_A CB_0.config_dataA\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2416_ net31 net32 net18 net19 net183 net182 vssd1 vssd1 vccd1 vccd1 _1044_ sky130_fd_sc_hd__mux4_1
X_3396_ clknet_leaf_27_clk _0216_ net253 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[88\]
+ sky130_fd_sc_hd__dfstp_1
X_2347_ _1511_ _1510_ _1522_ _0974_ vssd1 vssd1 vccd1 vccd1 _0975_ sky130_fd_sc_hd__a211o_4
X_2278_ net147 net159 LEI0.config_data\[42\] vssd1 vssd1 vccd1 vccd1 _0907_ sky130_fd_sc_hd__mux2_1
XFILLER_52_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2562__A2 _1014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3507__SET_B net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input19_A CBnorth_in[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2078__A1 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2250__A1 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1580_ SB0.route_sel\[57\] vssd1 vssd1 vccd1 vccd1 _1418_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_49_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3181_ clknet_leaf_6_clk _0001_ net255 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_2132_ net349 _0760_ _0761_ net352 _0759_ vssd1 vssd1 vccd1 vccd1 _0762_ sky130_fd_sc_hd__a221o_1
X_3250_ clknet_leaf_2_clk _0070_ net246 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_2201_ LEI0.config_data\[8\] net233 vssd1 vssd1 vccd1 vccd1 _0830_ sky130_fd_sc_hd__and2_1
XANTENNA__2608__A3 net23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2063_ CB_1.config_dataB\[8\] CB_1.config_dataB\[7\] CB_1.config_dataB\[9\] _0692_
+ vssd1 vssd1 vccd1 vccd1 _0693_ sky130_fd_sc_hd__or4bb_1
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1816__A1 _0439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2792__A2 _0956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2896_ net415 LE_0A.config_data\[16\] net212 vssd1 vssd1 vccd1 vccd1 _0065_ sky130_fd_sc_hd__mux2_1
X_1916_ SB0.route_sel\[96\] _1398_ _1401_ SB0.route_sel\[103\] _0545_ vssd1 vssd1
+ vccd1 vccd1 _0546_ sky130_fd_sc_hd__o221a_1
X_2965_ SB0.route_sel\[5\] SB0.route_sel\[4\] net293 vssd1 vssd1 vccd1 vccd1 _0133_
+ sky130_fd_sc_hd__mux2_1
X_1847_ SB0.route_sel\[15\] SB0.route_sel\[14\] vssd1 vssd1 vccd1 vccd1 _0477_ sky130_fd_sc_hd__nand2_1
X_3448_ clknet_leaf_9_clk _0268_ net260 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[12\]
+ sky130_fd_sc_hd__dfstp_1
X_3517_ clknet_leaf_32_clk _0337_ net240 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_1778_ _1502_ _0407_ vssd1 vssd1 vccd1 vccd1 _0408_ sky130_fd_sc_hd__or2_1
X_3379_ clknet_leaf_11_clk _0199_ net262 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[71\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclone11 _0539_ _0533_ _1013_ net310 vssd1 vssd1 vccd1 vccd1 net321 sky130_fd_sc_hd__a211o_1
XANTENNA__2232__B2 _0397_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclone44 _0539_ _0533_ _0542_ net309 vssd1 vssd1 vccd1 vccd1 net354 sky130_fd_sc_hd__a211o_1
Xclone33 _0367_ _0358_ _0981_ net305 vssd1 vssd1 vccd1 vccd1 net343 sky130_fd_sc_hd__a211o_1
XANTENNA__2232__A1 _0371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2299__B2 _0397_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2299__A1 _0371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2040__X _0670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output125_A net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2681_ SB0.route_sel\[88\] SB0.route_sel\[89\] vssd1 vssd1 vccd1 vccd1 _1303_ sky130_fd_sc_hd__nor2_1
X_2750_ SB0.route_sel\[7\] SB0.route_sel\[6\] vssd1 vssd1 vccd1 vccd1 _1349_ sky130_fd_sc_hd__nor2_1
X_1701_ _1527_ _1533_ _1537_ _1538_ vssd1 vssd1 vccd1 vccd1 _1539_ sky130_fd_sc_hd__a211o_1
X_1632_ CB_0.config_dataA\[2\] vssd1 vssd1 vccd1 vccd1 _1470_ sky130_fd_sc_hd__inv_2
X_1563_ SB0.route_sel\[102\] vssd1 vssd1 vccd1 vccd1 _1401_ sky130_fd_sc_hd__inv_2
X_3302_ clknet_leaf_21_clk _0122_ net274 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[19\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__1982__B1 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3233_ clknet_leaf_8_clk net455 net258 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_3095_ net190 CB_0.config_dataA\[7\] net217 vssd1 vssd1 vccd1 vccd1 _0263_ sky130_fd_sc_hd__mux2_1
X_2115_ net196 _0743_ _0744_ vssd1 vssd1 vccd1 vccd1 _0745_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_1_149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3164_ net458 LE_1B.config_data\[1\] net202 vssd1 vssd1 vccd1 vccd1 _0332_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2046_ net314 _0665_ net309 vssd1 vssd1 vccd1 vccd1 _0676_ sky130_fd_sc_hd__a21oi_4
XANTENNA_fanout156_A CB_0.le_outB vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2779__Y net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2948_ CB_1.config_dataB\[12\] CB_1.config_dataB\[13\] net230 vssd1 vssd1 vccd1 vccd1
+ _0116_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout209_X net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2125__X _0755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2879_ LE_0A.dff_out _1293_ net69 vssd1 vssd1 vccd1 vccd1 _0048_ sky130_fd_sc_hd__mux2_1
XANTENNA__2150__B1 CB_1.config_dataB\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2453__A1 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2035__X _0665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2453__B2 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload19 clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 clkload19/Y sky130_fd_sc_hd__bufinv_16
XANTENNA__2508__A2 _1134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2664_ LE_0A.config_data\[9\] _1180_ _1211_ _1290_ vssd1 vssd1 vccd1 vccd1 _1291_
+ sky130_fd_sc_hd__o211a_1
X_2802_ _1555_ net162 _0584_ vssd1 vssd1 vccd1 vccd1 _1378_ sky130_fd_sc_hd__o21bai_4
X_2733_ SB0.route_sel\[25\] _1435_ SB0.route_sel\[31\] SB0.route_sel\[30\] _1337_
+ vssd1 vssd1 vccd1 vccd1 _1338_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_14_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout217 net218 vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__clkbuf_4
Xfanout228 net231 vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__buf_2
X_1615_ SB0.route_sel\[117\] vssd1 vssd1 vccd1 vccd1 _1453_ sky130_fd_sc_hd__inv_2
X_2595_ _0966_ _1220_ _1221_ _0963_ CB_0.config_dataA\[12\] vssd1 vssd1 vccd1 vccd1
+ _1222_ sky130_fd_sc_hd__a221o_1
Xfanout239 _1504_ vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__buf_2
Xfanout206 net208 vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_65_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3078_ SB0.route_sel\[118\] SB0.route_sel\[117\] net299 vssd1 vssd1 vccd1 vccd1 _0246_
+ sky130_fd_sc_hd__mux2_1
X_3147_ CB_1.config_dataA\[8\] CB_1.config_dataA\[9\] net229 vssd1 vssd1 vccd1 vccd1
+ _0315_ sky130_fd_sc_hd__mux2_1
XFILLER_42_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3216_ clknet_leaf_3_clk _0036_ net253 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[36\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout273_A net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2029_ _0655_ _0649_ _0658_ net307 vssd1 vssd1 vccd1 vccd1 _0659_ sky130_fd_sc_hd__a211o_4
XANTENNA_fanout159_X net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2426__A1 net24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2380_ _1457_ net136 vssd1 vssd1 vccd1 vccd1 _1008_ sky130_fd_sc_hd__nand2_1
XFILLER_64_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput6 CBeast_in[14] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__buf_2
X_3001_ SB0.route_sel\[41\] SB0.route_sel\[40\] net288 vssd1 vssd1 vccd1 vccd1 _0169_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_62_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2647_ _1272_ _1273_ _1476_ vssd1 vssd1 vccd1 vccd1 _1274_ sky130_fd_sc_hd__mux2_1
X_2716_ _1523_ _1326_ vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__and2_4
X_2578_ _1203_ _1204_ _1472_ vssd1 vssd1 vccd1 vccd1 _1205_ sky130_fd_sc_hd__mux2_1
XANTENNA__2105__A0 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2656__A1 _1280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3081__A1 SB0.route_sel\[120\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_14_Right_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2592__A0 _0956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_23_Right_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input49_A SBwest_in[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_32_Right_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1880_ CB_1.config_dataA\[23\] CB_1.config_dataA\[22\] vssd1 vssd1 vccd1 vccd1 _0510_
+ sky130_fd_sc_hd__nand2_2
X_3481_ clknet_leaf_13_clk _0301_ net277 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[20\]
+ sky130_fd_sc_hd__dfstp_2
X_2501_ net328 net347 net179 vssd1 vssd1 vccd1 vccd1 _1129_ sky130_fd_sc_hd__mux2_4
X_2432_ CB_0.config_dataB\[8\] _1053_ _1056_ _1059_ vssd1 vssd1 vccd1 vccd1 _1060_
+ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_41_Right_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2363_ _0633_ _0627_ _0990_ net307 vssd1 vssd1 vccd1 vccd1 _0991_ sky130_fd_sc_hd__a211o_4
X_2294_ net2 net3 CB_1.config_dataA\[15\] vssd1 vssd1 vccd1 vccd1 _0923_ sky130_fd_sc_hd__mux2_1
XANTENNA__2820__B1_N _0397_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2335__B1 _0962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_50_Right_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1861__A2 _0481_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout236_A net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_11 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clone2_A1 _0633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2203__B net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput20 CBnorth_in[12] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__buf_2
Xinput31 CBnorth_in[8] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_44_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1932_ _0553_ _0557_ _0561_ vssd1 vssd1 vccd1 vccd1 _0562_ sky130_fd_sc_hd__a21bo_1
X_1863_ net200 _0450_ _0492_ vssd1 vssd1 vccd1 vccd1 _0493_ sky130_fd_sc_hd__a21oi_1
X_2981_ SB0.route_sel\[21\] SB0.route_sel\[20\] net286 vssd1 vssd1 vccd1 vccd1 _0149_
+ sky130_fd_sc_hd__mux2_1
X_2415_ net20 net22 net21 net23 CB_0.config_dataB\[6\] net183 vssd1 vssd1 vccd1 vccd1
+ _1043_ sky130_fd_sc_hd__mux4_1
X_1794_ _0423_ _0422_ vssd1 vssd1 vccd1 vccd1 _0424_ sky130_fd_sc_hd__or2_4
X_3464_ clknet_leaf_7_clk _0284_ net256 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[3\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__2556__A0 net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput53 SBwest_in[13] vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__clkbuf_2
Xinput64 SBwest_in[9] vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__clkbuf_1
Xinput42 SBsouth_in[3] vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__clkbuf_1
X_3395_ clknet_leaf_27_clk _0215_ net252 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[87\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__1819__C1 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2277_ LE_1A.config_data\[9\] net311 _0866_ _0905_ vssd1 vssd1 vccd1 vccd1 _0906_
+ sky130_fd_sc_hd__o211a_1
X_2346_ SB0.route_sel\[50\] SB0.route_sel\[51\] SB0.route_sel\[53\] _1425_ _0973_
+ vssd1 vssd1 vccd1 vccd1 _0974_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout239_X net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_32_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_32_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__2795__B1 _0486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2078__A2 net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2250__A2 net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_23_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__2538__A0 net20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3288__SET_B net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2200_ _0828_ _0817_ _0805_ vssd1 vssd1 vccd1 vccd1 _0829_ sky130_fd_sc_hd__o21ai_4
X_2062_ _1480_ net198 vssd1 vssd1 vccd1 vccd1 _0692_ sky130_fd_sc_hd__nor2_1
X_2131_ net194 net195 vssd1 vssd1 vccd1 vccd1 _0761_ sky130_fd_sc_hd__nor2_1
X_3180_ clknet_leaf_32_clk _0000_ net240 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_2964_ SB0.route_sel\[4\] SB0.route_sel\[3\] net293 vssd1 vssd1 vccd1 vccd1 _0132_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__1816__A2 _0445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_14_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2895_ net408 LE_0A.config_data\[15\] net213 vssd1 vssd1 vccd1 vccd1 _0064_ sky130_fd_sc_hd__mux2_1
X_1915_ SB0.route_sel\[101\] SB0.route_sel\[100\] vssd1 vssd1 vccd1 vccd1 _0545_ sky130_fd_sc_hd__or2_1
X_1777_ CB_1.config_dataA\[23\] CB_1.config_dataA\[22\] vssd1 vssd1 vccd1 vccd1 _0407_
+ sky130_fd_sc_hd__or2_2
X_1846_ net320 _0474_ _0475_ _0473_ net235 vssd1 vssd1 vccd1 vccd1 _0476_ sky130_fd_sc_hd__o221a_1
X_3447_ clknet_leaf_9_clk _0267_ net260 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[11\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_clkbuf_leaf_15_clk_A clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3378_ clknet_leaf_12_clk _0198_ net262 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[70\]
+ sky130_fd_sc_hd__dfstp_1
X_3516_ clknet_leaf_32_clk _0336_ net240 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_4_Right_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_55_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2329_ SB0.route_sel\[30\] SB0.route_sel\[31\] vssd1 vssd1 vccd1 vccd1 _0957_ sky130_fd_sc_hd__nand2b_1
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclone34 _0445_ _0439_ _0448_ net305 vssd1 vssd1 vccd1 vccd1 net344 sky130_fd_sc_hd__a211o_1
XFILLER_25_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input31_A CBnorth_in[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output118_A net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1631_ CB_0.config_dataB\[17\] vssd1 vssd1 vccd1 vccd1 _1469_ sky130_fd_sc_hd__inv_2
X_2680_ _0563_ _1302_ vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__and2_4
XFILLER_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1700_ SB0.route_sel\[57\] SB0.route_sel\[56\] vssd1 vssd1 vccd1 vccd1 _1538_ sky130_fd_sc_hd__nand2_1
X_3232_ clknet_leaf_7_clk net399 net258 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_3301_ clknet_leaf_17_clk _0121_ net279 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[18\]
+ sky130_fd_sc_hd__dfstp_1
X_1562_ SB0.route_sel\[100\] vssd1 vssd1 vccd1 vccd1 _1400_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_3_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_54_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3094_ net191 net190 net217 vssd1 vssd1 vccd1 vccd1 _0262_ sky130_fd_sc_hd__mux2_1
X_2114_ net361 _0729_ _0733_ net357 _1483_ vssd1 vssd1 vccd1 vccd1 _0744_ sky130_fd_sc_hd__a221o_1
X_2045_ _0670_ _0666_ _0674_ _1415_ _1414_ vssd1 vssd1 vccd1 vccd1 _0675_ sky130_fd_sc_hd__a2111o_1
X_3163_ LE_0A.config_data\[16\] net458 net206 vssd1 vssd1 vccd1 vccd1 _0331_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_2_2__f_clk_X clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2947_ net196 CB_1.config_dataB\[12\] net229 vssd1 vssd1 vccd1 vccd1 _0115_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout149_A net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1829_ _0456_ _0457_ _0451_ vssd1 vssd1 vccd1 vccd1 _0459_ sky130_fd_sc_hd__a21oi_1
X_2878_ net450 CB_0.config_data_inA net210 vssd1 vssd1 vccd1 vccd1 _0047_ sky130_fd_sc_hd__mux2_1
XFILLER_45_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input34_X net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2801_ _1377_ _0525_ _0526_ vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__a21boi_1
XTAP_TAPCELL_ROW_14_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1614_ SB0.route_sel\[116\] vssd1 vssd1 vccd1 vccd1 _1452_ sky130_fd_sc_hd__inv_2
X_2594_ net188 net189 vssd1 vssd1 vccd1 vccd1 _1221_ sky130_fd_sc_hd__and2b_1
X_2663_ _1173_ _1174_ _1179_ LE_0A.config_data\[8\] vssd1 vssd1 vccd1 vccd1 _1290_
+ sky130_fd_sc_hd__a211o_1
X_2732_ SB0.route_sel\[26\] SB0.route_sel\[27\] vssd1 vssd1 vccd1 vccd1 _1337_ sky130_fd_sc_hd__nand2b_1
Xfanout218 net221 vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__clkbuf_2
Xfanout229 net231 vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__clkbuf_4
XANTENNA__2548__S LEI0.config_data\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout207 net208 vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__clkbuf_4
X_3215_ clknet_leaf_3_clk _0035_ net251 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[35\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2668__C1 net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3077_ SB0.route_sel\[117\] SB0.route_sel\[116\] net299 vssd1 vssd1 vccd1 vccd1 _0245_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3146_ CB_1.config_dataA\[7\] CB_1.config_dataA\[8\] net229 vssd1 vssd1 vccd1 vccd1
+ _0314_ sky130_fd_sc_hd__mux2_1
X_2028_ _1410_ SB0.route_sel\[72\] SB0.route_sel\[77\] SB0.route_sel\[76\] _0657_
+ vssd1 vssd1 vccd1 vccd1 _0658_ sky130_fd_sc_hd__o221a_1
XANTENNA__2435__A2 net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout221_X net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2426__A2 net25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput7 CBeast_in[15] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_62_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3000_ SB0.route_sel\[40\] SB0.route_sel\[39\] net288 vssd1 vssd1 vccd1 vccd1 _0168_
+ sky130_fd_sc_hd__mux2_1
X_2646_ net17 net24 net25 net26 CB_0.config_dataA\[15\] CB_0.config_dataA\[16\] vssd1
+ vssd1 vccd1 vccd1 _1273_ sky130_fd_sc_hd__mux4_1
X_2577_ net17 net24 net25 net26 net191 net190 vssd1 vssd1 vccd1 vccd1 _1204_ sky130_fd_sc_hd__mux4_1
X_2715_ _1422_ SB0.route_sel\[48\] _1423_ SB0.route_sel\[51\] _1325_ vssd1 vssd1 vccd1
+ vccd1 _1326_ sky130_fd_sc_hd__a221o_1
XANTENNA__2105__A1 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3129_ CB_0.config_dataB\[15\] net178 net226 vssd1 vssd1 vccd1 vccd1 _0297_ sky130_fd_sc_hd__mux2_1
XFILLER_27_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2592__A1 _0959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1698__A3 net62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3480_ clknet_leaf_13_clk _0300_ net277 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[19\]
+ sky130_fd_sc_hd__dfstp_1
X_2500_ CB_0.config_dataB\[18\] _1127_ vssd1 vssd1 vccd1 vccd1 _1128_ sky130_fd_sc_hd__nor2_1
X_2431_ net182 _1057_ _1058_ vssd1 vssd1 vccd1 vccd1 _1059_ sky130_fd_sc_hd__a21oi_1
XANTENNA__2335__A1 _0487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2362_ SB0.route_sel\[82\] SB0.route_sel\[83\] SB0.route_sel\[85\] _1409_ _0989_
+ vssd1 vssd1 vccd1 vccd1 _0990_ sky130_fd_sc_hd__o221a_1
X_2293_ CB_1.config_dataA\[16\] _0920_ _0921_ vssd1 vssd1 vccd1 vccd1 _0922_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_47_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2127__A net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2574__B2 _0985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2574__A1 _0982_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout229_A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput130 net130 vssd1 vssd1 vccd1 vccd1 SBwest_out[4] sky130_fd_sc_hd__buf_8
X_2629_ LEI0.config_data\[37\] _1253_ _1255_ LEI0.config_data\[38\] net304 vssd1 vssd1
+ vccd1 vccd1 _1256_ sky130_fd_sc_hd__a2111oi_1
XANTENNA__2262__A0 net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clone2_A2 _0627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2317__A1 _0829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input61_A SBwest_in[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2980_ SB0.route_sel\[20\] SB0.route_sel\[19\] net286 vssd1 vssd1 vccd1 vccd1 _0148_
+ sky130_fd_sc_hd__mux2_1
Xinput21 CBnorth_in[13] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__clkbuf_2
Xinput32 CBnorth_in[9] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__clkbuf_2
X_1793_ _0419_ _0421_ _0420_ SB0.route_sel\[16\] SB0.route_sel\[17\] vssd1 vssd1 vccd1
+ vccd1 _0423_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_44_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput10 CBeast_in[3] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__buf_8
X_1931_ _0559_ _0560_ SB0.route_sel\[96\] SB0.route_sel\[97\] vssd1 vssd1 vccd1 vccd1
+ _0561_ sky130_fd_sc_hd__o211a_1
Xinput54 SBwest_in[14] vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__clkbuf_2
X_1862_ _0398_ net345 net359 _1495_ CB_1.config_dataB\[2\] vssd1 vssd1 vccd1 vccd1
+ _0492_ sky130_fd_sc_hd__a221o_1
Xinput43 SBsouth_in[4] vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__buf_1
Xinput65 config_data_in vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__clkbuf_1
X_3463_ clknet_leaf_7_clk _0283_ net259 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[2\]
+ sky130_fd_sc_hd__dfstp_2
X_2414_ net182 _1038_ _1041_ vssd1 vssd1 vccd1 vccd1 _1042_ sky130_fd_sc_hd__a21oi_1
X_3394_ clknet_leaf_4_clk _0214_ net252 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[86\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__1819__B1 _0448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2276_ _0829_ _0830_ _0835_ LE_1A.config_data\[8\] vssd1 vssd1 vccd1 vccd1 _0905_
+ sky130_fd_sc_hd__a211o_1
X_2345_ SB0.route_sel\[54\] SB0.route_sel\[55\] vssd1 vssd1 vccd1 vccd1 _0973_ sky130_fd_sc_hd__nand2b_1
XANTENNA__1696__A SB0.route_sel\[63\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout301_X net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2078__A3 net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2538__A1 net22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2786__A1 _0982_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2250__A3 net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2130_ net194 net195 vssd1 vssd1 vccd1 vccd1 _0760_ sky130_fd_sc_hd__and2b_1
X_2061_ _0683_ _0684_ _0689_ vssd1 vssd1 vccd1 vccd1 _0691_ sky130_fd_sc_hd__a21o_2
X_1914_ net201 net354 _0522_ net200 vssd1 vssd1 vccd1 vccd1 _0544_ sky130_fd_sc_hd__o211a_1
X_2963_ SB0.route_sel\[3\] SB0.route_sel\[2\] net293 vssd1 vssd1 vccd1 vccd1 _0131_
+ sky130_fd_sc_hd__mux2_1
X_2894_ net418 net408 net213 vssd1 vssd1 vccd1 vccd1 _0063_ sky130_fd_sc_hd__mux2_1
XANTENNA__1985__C1 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1776_ net168 net163 net9 vssd1 vssd1 vccd1 vccd1 _0406_ sky130_fd_sc_hd__o21a_1
X_3515_ clknet_leaf_32_clk _0335_ net240 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_1845_ net157 net166 net163 _0407_ _0349_ vssd1 vssd1 vccd1 vccd1 _0475_ sky130_fd_sc_hd__o32ai_2
X_3446_ clknet_leaf_9_clk _0266_ net259 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[10\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_fanout296_A net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3377_ clknet_leaf_4_clk _0197_ net262 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[69\]
+ sky130_fd_sc_hd__dfstp_1
X_2328_ _0424_ _0415_ _0955_ net303 vssd1 vssd1 vccd1 vccd1 _0956_ sky130_fd_sc_hd__a211o_4
XANTENNA__2162__C1 _0755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3294__SET_B net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2259_ _0491_ _0873_ _0876_ _0471_ CB_1.config_dataA\[12\] vssd1 vssd1 vccd1 vccd1
+ _0888_ sky130_fd_sc_hd__a221o_1
XANTENNA__2768__A1 _1014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2217__A0 net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclone35 _0467_ _0461_ _0470_ net306 vssd1 vssd1 vccd1 vccd1 net345 sky130_fd_sc_hd__a211o_1
Xclone46 _1548_ _1539_ _1551_ net306 vssd1 vssd1 vccd1 vccd1 net356 sky130_fd_sc_hd__a211o_1
XFILLER_0_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1728__C1 _0357_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input24_A CBnorth_in[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2049__X _0679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2153__C1 net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2208__A0 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1630_ CB_0.config_dataB\[12\] vssd1 vssd1 vccd1 vccd1 _1468_ sky130_fd_sc_hd__inv_2
X_3231_ clknet_leaf_8_clk _0051_ net258 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_3300_ clknet_leaf_17_clk _0120_ net279 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[17\]
+ sky130_fd_sc_hd__dfstp_1
X_1561_ SB0.route_sel\[98\] vssd1 vssd1 vccd1 vccd1 _1399_ sky130_fd_sc_hd__inv_2
X_3162_ CB_1.config_dataA\[23\] CB_1.config_dataA\[24\] net223 vssd1 vssd1 vccd1 vccd1
+ _0330_ sky130_fd_sc_hd__mux2_1
X_3093_ CB_0.config_dataA\[4\] net191 net216 vssd1 vssd1 vccd1 vccd1 _0261_ sky130_fd_sc_hd__mux2_1
X_2113_ _1526_ net356 net197 vssd1 vssd1 vccd1 vccd1 _0743_ sky130_fd_sc_hd__mux2_1
X_2044_ net47 _0672_ _0673_ vssd1 vssd1 vccd1 vccd1 _0674_ sky130_fd_sc_hd__a21oi_1
XANTENNA__1798__X _0428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2946_ net197 net196 net229 vssd1 vssd1 vccd1 vccd1 _0114_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_17_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2877_ net453 net450 net210 vssd1 vssd1 vccd1 vccd1 _0046_ sky130_fd_sc_hd__mux2_1
X_1759_ CB_0.config_dataA\[24\] CB_0.config_dataA\[21\] CB_0.config_dataA\[20\] vssd1
+ vssd1 vccd1 vccd1 _0389_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout309_A net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout211_A net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap140 _0872_ vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__clkbuf_1
X_1828_ _1448_ _1449_ net33 vssd1 vssd1 vccd1 vccd1 _0458_ sky130_fd_sc_hd__o21ai_1
XFILLER_57_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3429_ clknet_leaf_18_clk _0249_ net276 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[121\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_0_140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input27_X net27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output130_A net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_14_clk_A clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2800_ _1499_ _0508_ _0543_ vssd1 vssd1 vccd1 vccd1 _1377_ sky130_fd_sc_hd__o21bai_1
X_2731_ _1336_ _0446_ vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__nor2_8
XTAP_TAPCELL_ROW_14_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1613_ SB0.route_sel\[113\] vssd1 vssd1 vccd1 vccd1 _1451_ sky130_fd_sc_hd__inv_2
X_2593_ net189 net188 vssd1 vssd1 vccd1 vccd1 _1220_ sky130_fd_sc_hd__nor2_1
X_2662_ LE_0A.config_data\[11\] LE_0A.config_data\[10\] _1180_ vssd1 vssd1 vccd1 vccd1
+ _1289_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_29_clk_A clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout219 net221 vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__clkbuf_4
X_3145_ net174 CB_1.config_dataA\[7\] net230 vssd1 vssd1 vccd1 vccd1 _0313_ sky130_fd_sc_hd__mux2_1
Xfanout208 net209 vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__buf_2
X_3214_ clknet_leaf_3_clk _0034_ net251 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[34\]
+ sky130_fd_sc_hd__dfrtp_1
X_3076_ SB0.route_sel\[116\] SB0.route_sel\[115\] net299 vssd1 vssd1 vccd1 vccd1 _0244_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2027_ SB0.route_sel\[79\] SB0.route_sel\[78\] vssd1 vssd1 vccd1 vccd1 _0657_ sky130_fd_sc_hd__nand2b_1
X_2929_ net416 LE_1A.config_data\[13\] net204 vssd1 vssd1 vccd1 vccd1 _0098_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_17_Left_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1991__X _0621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2426__A3 net26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2347__C1 _0974_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput8 CBeast_in[1] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_62_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2714_ SB0.route_sel\[55\] SB0.route_sel\[54\] vssd1 vssd1 vccd1 vccd1 _1325_ sky130_fd_sc_hd__nor2_1
X_2645_ net27 net28 net29 net30 CB_0.config_dataA\[15\] net186 vssd1 vssd1 vccd1 vccd1
+ _1272_ sky130_fd_sc_hd__mux4_1
X_2576_ net27 net28 net29 net30 net191 net190 vssd1 vssd1 vccd1 vccd1 _1203_ sky130_fd_sc_hd__mux4_1
XANTENNA__2338__C1 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2105__A2 net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3128_ CB_0.config_dataB\[14\] net179 net219 vssd1 vssd1 vccd1 vccd1 _0296_ sky130_fd_sc_hd__mux2_1
X_3059_ SB0.route_sel\[99\] SB0.route_sel\[98\] net295 vssd1 vssd1 vccd1 vccd1 _0227_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_33_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_2_Left_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2430_ net342 _1039_ _1040_ net343 _1466_ vssd1 vssd1 vccd1 vccd1 _1058_ sky130_fd_sc_hd__a221o_1
X_2361_ SB0.route_sel\[86\] SB0.route_sel\[87\] vssd1 vssd1 vccd1 vccd1 _0989_ sky130_fd_sc_hd__nand2b_1
XANTENNA__2520__X CB_0.le_outB vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2335__A2 _0481_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2638__A3 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2292_ _0659_ _0911_ _0914_ _0679_ vssd1 vssd1 vccd1 vccd1 _0921_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_47_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2127__B CB_0.config_data_inA vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2559_ net190 net191 vssd1 vssd1 vccd1 vccd1 _1186_ sky130_fd_sc_hd__and2b_1
Xoutput131 net131 vssd1 vssd1 vccd1 vccd1 SBwest_out[5] sky130_fd_sc_hd__buf_8
X_2628_ LEI0.config_data\[37\] _1254_ vssd1 vssd1 vccd1 vccd1 _1255_ sky130_fd_sc_hd__nor2_1
Xoutput120 net120 vssd1 vssd1 vccd1 vccd1 SBwest_out[0] sky130_fd_sc_hd__buf_6
XPHY_EDGE_ROW_34_Left_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_43_Left_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2262__A1 net12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input54_A SBwest_in[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1930_ SB0.route_sel\[101\] SB0.route_sel\[100\] net52 _0558_ _0553_ vssd1 vssd1
+ vccd1 vccd1 _0560_ sky130_fd_sc_hd__a41o_1
Xinput22 CBnorth_in[14] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__buf_2
Xinput66 config_en vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__clkbuf_2
X_1792_ net144 _0420_ net234 vssd1 vssd1 vccd1 vccd1 _0422_ sky130_fd_sc_hd__o21ai_1
Xinput11 CBeast_in[4] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__buf_6
Xinput55 SBwest_in[15] vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__buf_1
Xinput44 SBsouth_in[5] vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__buf_1
Xinput33 SBsouth_in[0] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_1
X_1861_ _0487_ _0481_ _0490_ net306 vssd1 vssd1 vccd1 vccd1 _0491_ sky130_fd_sc_hd__a211o_4
XANTENNA__1764__B1 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3462_ clknet_leaf_7_clk _0282_ net259 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[1\]
+ sky130_fd_sc_hd__dfstp_1
X_2344_ _0970_ _0971_ CB_0.config_dataB\[2\] vssd1 vssd1 vccd1 vccd1 _0972_ sky130_fd_sc_hd__mux2_1
X_2413_ net313 _1039_ _1040_ net336 CB_0.config_dataB\[7\] vssd1 vssd1 vccd1 vccd1
+ _1041_ sky130_fd_sc_hd__a221o_1
X_3393_ clknet_leaf_27_clk _0213_ net252 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[85\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_52_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_35_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2275_ LE_1A.config_data\[11\] net311 _0867_ _0903_ vssd1 vssd1 vccd1 vccd1 _0904_
+ sky130_fd_sc_hd__o211a_1
XANTENNA__1819__A1 _0445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2335__X _0963_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2538__A2 net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_5_Left_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2060_ _0684_ _0683_ _0689_ vssd1 vssd1 vccd1 vccd1 _0690_ sky130_fd_sc_hd__a21oi_4
X_1913_ _0539_ _0533_ _0542_ net309 vssd1 vssd1 vccd1 vccd1 _0543_ sky130_fd_sc_hd__a211o_4
X_2893_ net411 LE_0A.config_data\[13\] net213 vssd1 vssd1 vccd1 vccd1 _0062_ sky130_fd_sc_hd__mux2_1
XANTENNA__2226__B2 _0471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2226__A1 _0491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2405__B net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2962_ SB0.route_sel\[2\] SB0.route_sel\[1\] net293 vssd1 vssd1 vccd1 vccd1 _0130_
+ sky130_fd_sc_hd__mux2_1
X_3445_ clknet_leaf_9_clk _0265_ net259 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[9\]
+ sky130_fd_sc_hd__dfstp_1
X_3514_ clknet_leaf_32_clk net468 net240 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_1775_ CB_1.config_dataB\[23\] CB_1.config_dataB\[22\] vssd1 vssd1 vccd1 vccd1 _0405_
+ sky130_fd_sc_hd__or2_1
X_1844_ _0349_ _0407_ vssd1 vssd1 vccd1 vccd1 _0474_ sky130_fd_sc_hd__or2_1
X_3376_ clknet_leaf_12_clk _0196_ net262 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[68\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_fanout289_A net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2258_ _0428_ _0449_ CB_1.config_dataA\[10\] vssd1 vssd1 vccd1 vccd1 _0887_ sky130_fd_sc_hd__mux2_1
X_2327_ SB0.route_sel\[18\] SB0.route_sel\[19\] SB0.route_sel\[21\] _1441_ _0954_
+ vssd1 vssd1 vccd1 vccd1 _0955_ sky130_fd_sc_hd__o221a_1
XANTENNA__2217__A1 net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2189_ _1526_ _1552_ net177 vssd1 vssd1 vccd1 vccd1 _0818_ sky130_fd_sc_hd__mux2_1
XFILLER_25_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1976__B1 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclone47 _0393_ _0384_ _0396_ net305 vssd1 vssd1 vccd1 vccd1 net357 sky130_fd_sc_hd__a211o_1
XANTENNA__2153__B1 CB_0.config_data_inA vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1900__B1 net38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input17_A CBnorth_in[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_31_Left_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3101__S net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2940__S net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2208__A1 net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1560_ SB0.route_sel\[97\] vssd1 vssd1 vccd1 vccd1 _1398_ sky130_fd_sc_hd__inv_2
X_3230_ clknet_leaf_8_clk _0050_ net258 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_2112_ _1483_ _0738_ _0741_ _0737_ vssd1 vssd1 vccd1 vccd1 _0742_ sky130_fd_sc_hd__a211o_1
X_3161_ CB_1.config_dataA\[22\] CB_1.config_dataA\[23\] net223 vssd1 vssd1 vccd1 vccd1
+ _0329_ sky130_fd_sc_hd__mux2_1
X_3092_ CB_0.config_dataA\[3\] CB_0.config_dataA\[4\] net218 vssd1 vssd1 vccd1 vccd1
+ _0260_ sky130_fd_sc_hd__mux2_1
XANTENNA__2447__A1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2447__B2 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2043_ SB0.route_sel\[69\] SB0.route_sel\[68\] net63 _0671_ _0666_ vssd1 vssd1 vccd1
+ vccd1 _0673_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_60_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2945_ CB_1.config_dataB\[9\] CB_1.config_dataB\[10\] net229 vssd1 vssd1 vccd1 vccd1
+ _0113_ sky130_fd_sc_hd__mux2_1
X_1827_ SB0.route_sel\[5\] SB0.route_sel\[4\] net49 vssd1 vssd1 vccd1 vccd1 _0457_
+ sky130_fd_sc_hd__and3_1
X_2876_ LEI0.config_data\[44\] net453 net210 vssd1 vssd1 vccd1 vccd1 _0045_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_17_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3428_ clknet_leaf_15_clk _0248_ net281 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[120\]
+ sky130_fd_sc_hd__dfstp_1
X_1758_ _1517_ _0386_ net27 vssd1 vssd1 vccd1 vccd1 _0388_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout204_A net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1689_ SB0.route_sel\[58\] SB0.route_sel\[59\] vssd1 vssd1 vccd1 vccd1 _1527_ sky130_fd_sc_hd__nand2_1
XANTENNA__1725__A3 net60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap141 _0840_ vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__buf_1
XFILLER_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input9_A CBeast_in[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3359_ clknet_leaf_26_clk _0179_ net269 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[51\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_51_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1884__B net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clone9_X net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output123_A net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2601__A1 _0985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2601__B2 _0982_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2661_ _1212_ _1285_ _1287_ _1244_ vssd1 vssd1 vccd1 vccd1 _1288_ sky130_fd_sc_hd__a211o_1
X_2730_ _1434_ _1435_ _1335_ vssd1 vssd1 vccd1 vccd1 _1336_ sky130_fd_sc_hd__a21oi_1
X_2592_ _0956_ _0959_ net189 vssd1 vssd1 vccd1 vccd1 _1219_ sky130_fd_sc_hd__mux2_1
XANTENNA__2117__A0 net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1612_ CB_1.config_dataA\[2\] vssd1 vssd1 vccd1 vccd1 _1450_ sky130_fd_sc_hd__inv_2
Xfanout209 net221 vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__clkbuf_2
X_3075_ SB0.route_sel\[115\] SB0.route_sel\[114\] net299 vssd1 vssd1 vccd1 vccd1 _0243_
+ sky130_fd_sc_hd__mux2_1
X_3144_ CB_1.config_dataA\[5\] CB_1.config_dataA\[6\] net230 vssd1 vssd1 vccd1 vccd1
+ _0312_ sky130_fd_sc_hd__mux2_1
XFILLER_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3213_ clknet_leaf_3_clk _0033_ net251 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[33\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_65_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2026_ _0655_ _0649_ net307 vssd1 vssd1 vccd1 vccd1 _0656_ sky130_fd_sc_hd__a21oi_2
X_2859_ LEI0.config_data\[27\] net481 net207 vssd1 vssd1 vccd1 vccd1 _0028_ sky130_fd_sc_hd__mux2_1
X_2928_ net441 net416 net210 vssd1 vssd1 vccd1 vccd1 _0097_ sky130_fd_sc_hd__mux2_1
XFILLER_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2108__A0 net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_2_3__f_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2831__A1 LEI0.config_data\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2347__B1 _1522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput9 CBeast_in[2] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__buf_6
XFILLER_32_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2644_ net186 _1269_ _1270_ vssd1 vssd1 vccd1 vccd1 _1271_ sky130_fd_sc_hd__a21oi_1
X_2713_ _1323_ _1324_ _1523_ vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__a21boi_4
X_2575_ net190 _1200_ _1201_ vssd1 vssd1 vccd1 vccd1 _1202_ sky130_fd_sc_hd__a21oi_1
XANTENNA__2338__B1 _0965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2105__A3 net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3127_ CB_0.config_dataB\[13\] CB_0.config_dataB\[14\] net220 vssd1 vssd1 vccd1 vccd1
+ _0295_ sky130_fd_sc_hd__mux2_1
XFILLER_42_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3058_ SB0.route_sel\[98\] SB0.route_sel\[97\] net298 vssd1 vssd1 vccd1 vccd1 _0226_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout271_A net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2577__A0 net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2009_ SB0.route_sel\[74\] SB0.route_sel\[75\] vssd1 vssd1 vccd1 vccd1 _0639_ sky130_fd_sc_hd__nand2_1
XFILLER_23_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1785__D1 SB0.route_sel\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_13_clk_A clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2338__X _0966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clone32_X net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_28_clk_A clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2360_ CB_0.config_dataB\[3\] _0972_ _0987_ _0969_ vssd1 vssd1 vccd1 vccd1 _0988_
+ sky130_fd_sc_hd__and4bb_1
X_2291_ _0637_ _0615_ CB_1.config_dataA\[15\] vssd1 vssd1 vccd1 vccd1 _0920_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_10_Right_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput121 net121 vssd1 vssd1 vccd1 vccd1 SBwest_out[10] sky130_fd_sc_hd__buf_8
Xoutput132 net132 vssd1 vssd1 vccd1 vccd1 SBwest_out[6] sky130_fd_sc_hd__buf_6
X_2627_ net142 net156 LEI0.config_data\[36\] vssd1 vssd1 vccd1 vccd1 _1254_ sky130_fd_sc_hd__mux2_1
Xoutput110 net110 vssd1 vssd1 vccd1 vccd1 SBsouth_out[15] sky130_fd_sc_hd__buf_6
X_2489_ net31 _1113_ _1115_ net178 vssd1 vssd1 vccd1 vccd1 _1117_ sky130_fd_sc_hd__a22oi_1
X_2558_ LEI0.config_data\[13\] _1183_ _1184_ vssd1 vssd1 vccd1 vccd1 _1185_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_38_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1997__X _0627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout274_X net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2798__B1 _0521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2262__A2 net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input47_A SBsouth_in[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3104__S net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2943__S net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1860_ _1442_ SB0.route_sel\[8\] SB0.route_sel\[13\] SB0.route_sel\[12\] _0489_ vssd1
+ vssd1 vccd1 vccd1 _0490_ sky130_fd_sc_hd__o221a_1
Xclkbuf_leaf_26_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_clk
+ sky130_fd_sc_hd__clkbuf_8
Xinput23 CBnorth_in[15] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__buf_2
Xinput67 en vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__clkbuf_1
X_3461_ clknet_leaf_13_clk _0281_ net278 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_1791_ _0417_ _1518_ net151 vssd1 vssd1 vccd1 vccd1 _0421_ sky130_fd_sc_hd__or3_4
Xinput12 CBeast_in[5] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__buf_6
XANTENNA__1764__A1 _0393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput34 SBsouth_in[10] vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__buf_1
Xinput45 SBsouth_in[6] vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__buf_1
Xinput56 SBwest_in[1] vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__buf_1
X_2343_ net27 net28 net29 net30 net185 net184 vssd1 vssd1 vccd1 vccd1 _0971_ sky130_fd_sc_hd__mux4_1
X_2412_ net182 net183 vssd1 vssd1 vccd1 vccd1 _1040_ sky130_fd_sc_hd__and2b_1
X_3392_ clknet_leaf_27_clk _0212_ net252 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[84\]
+ sky130_fd_sc_hd__dfstp_1
X_2274_ _0829_ _0830_ _0835_ LE_1A.config_data\[10\] vssd1 vssd1 vccd1 vccd1 _0903_
+ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_17_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_25_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1819__A2 _0439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout234_A net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1989_ net157 net168 _0591_ _0593_ _1502_ vssd1 vssd1 vccd1 vccd1 _0619_ sky130_fd_sc_hd__o32a_1
XFILLER_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1691__B1 net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2538__A3 net23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2171__B2 _0783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2171__A1 _0755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_62_Left_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1912_ SB0.route_sel\[112\] _1451_ SB0.route_sel\[116\] SB0.route_sel\[117\] _0541_
+ vssd1 vssd1 vccd1 vccd1 _0542_ sky130_fd_sc_hd__o221a_1
X_2892_ net384 LE_0A.config_data\[12\] net213 vssd1 vssd1 vccd1 vccd1 _0061_ sky130_fd_sc_hd__mux2_1
X_2961_ SB0.route_sel\[1\] SB0.route_sel\[0\] net293 vssd1 vssd1 vccd1 vccd1 _0129_
+ sky130_fd_sc_hd__mux2_1
X_1843_ net166 _0405_ net8 vssd1 vssd1 vccd1 vccd1 _0473_ sky130_fd_sc_hd__o21a_1
X_3444_ clknet_leaf_7_clk _0264_ net259 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[8\]
+ sky130_fd_sc_hd__dfstp_1
Xclkbuf_leaf_6_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_clk
+ sky130_fd_sc_hd__clkbuf_8
X_3513_ clknet_leaf_32_clk net461 net240 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_1774_ SB0.route_sel\[18\] SB0.route_sel\[19\] vssd1 vssd1 vccd1 vccd1 _0404_ sky130_fd_sc_hd__and2_1
X_3375_ clknet_leaf_11_clk _0195_ net261 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[67\]
+ sky130_fd_sc_hd__dfstp_1
X_2257_ _0878_ _0881_ _0885_ CB_1.config_dataA\[13\] vssd1 vssd1 vccd1 vccd1 _0886_
+ sky130_fd_sc_hd__or4b_1
X_2326_ SB0.route_sel\[22\] SB0.route_sel\[23\] vssd1 vssd1 vccd1 vccd1 _0954_ sky130_fd_sc_hd__nand2b_1
XANTENNA__2217__A2 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2188_ _0812_ _0809_ _0816_ CB_1.config_dataA\[3\] vssd1 vssd1 vccd1 vccd1 _0817_
+ sky130_fd_sc_hd__and4bb_1
Xclone26 _0655_ _0649_ _0997_ net307 vssd1 vssd1 vccd1 vccd1 net336 sky130_fd_sc_hd__a211o_1
Xclone37 _1548_ _1539_ _0977_ net306 vssd1 vssd1 vccd1 vccd1 net347 sky130_fd_sc_hd__a211o_1
XFILLER_16_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2346__X _0974_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3091_ CB_0.config_dataA\[2\] CB_0.config_dataA\[3\] net217 vssd1 vssd1 vccd1 vccd1
+ _0259_ sky130_fd_sc_hd__mux2_1
X_2111_ net196 _0739_ _0740_ vssd1 vssd1 vccd1 vccd1 _0741_ sky130_fd_sc_hd__a21oi_1
X_2042_ SB0.route_sel\[69\] SB0.route_sel\[68\] vssd1 vssd1 vccd1 vccd1 _0672_ sky130_fd_sc_hd__nand2_1
X_3160_ CB_1.config_dataA\[21\] CB_1.config_dataA\[22\] net223 vssd1 vssd1 vccd1 vccd1
+ _0328_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_8_Right_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2944_ CB_1.config_dataB\[8\] CB_1.config_dataB\[9\] net228 vssd1 vssd1 vccd1 vccd1
+ _0112_ sky130_fd_sc_hd__mux2_1
X_1826_ SB0.route_sel\[7\] SB0.route_sel\[6\] vssd1 vssd1 vccd1 vccd1 _0456_ sky130_fd_sc_hd__nand2_1
X_2875_ net488 LEI0.config_data\[44\] net210 vssd1 vssd1 vccd1 vccd1 _0044_ sky130_fd_sc_hd__mux2_1
X_3427_ clknet_leaf_15_clk _0247_ net281 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[119\]
+ sky130_fd_sc_hd__dfstp_1
Xmax_cap164 _0385_ vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__clkbuf_1
X_1757_ _1516_ net164 vssd1 vssd1 vccd1 vccd1 _0387_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_39_Right_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3358_ clknet_leaf_26_clk _0178_ net269 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[50\]
+ sky130_fd_sc_hd__dfstp_1
X_1688_ _1510_ _1511_ _1522_ _1525_ vssd1 vssd1 vccd1 vccd1 _1526_ sky130_fd_sc_hd__a211o_2
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3289_ clknet_leaf_19_clk _0109_ net276 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[6\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__1894__B1 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2309_ _1463_ _1464_ CB_1.config_dataA\[19\] _0911_ _0937_ vssd1 vssd1 vccd1 vccd1
+ _0938_ sky130_fd_sc_hd__a41o_1
XANTENNA__1949__A1 net37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_48_Right_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2071__A0 net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_57_Right_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1737__C_N _0357_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_66_Right_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2951__S net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output116_A net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2660_ LE_0A.config_data\[13\] _1180_ _1211_ _1286_ vssd1 vssd1 vccd1 vccd1 _1287_
+ sky130_fd_sc_hd__o211a_1
X_1611_ SB0.route_sel\[4\] vssd1 vssd1 vccd1 vccd1 _1449_ sky130_fd_sc_hd__inv_2
XANTENNA__2117__A1 net12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2591_ net310 LEI0.config_data\[26\] _1217_ _1215_ vssd1 vssd1 vccd1 vccd1 _1218_
+ sky130_fd_sc_hd__nor4_4
X_3212_ clknet_leaf_28_clk _0032_ net251 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[32\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_65_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3074_ SB0.route_sel\[114\] SB0.route_sel\[113\] net299 vssd1 vssd1 vccd1 vccd1 _0242_
+ sky130_fd_sc_hd__mux2_1
X_3143_ CB_1.config_dataA\[4\] net175 net230 vssd1 vssd1 vccd1 vccd1 _0311_ sky130_fd_sc_hd__mux2_1
X_2025_ _0653_ _0654_ _0648_ vssd1 vssd1 vccd1 vccd1 _0655_ sky130_fd_sc_hd__or3b_4
XFILLER_35_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2927_ net446 net441 net210 vssd1 vssd1 vccd1 vccd1 _0096_ sky130_fd_sc_hd__mux2_1
X_2789_ _1371_ _0390_ _0392_ vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__a21oi_4
X_2858_ LEI0.config_data\[26\] LEI0.config_data\[27\] net214 vssd1 vssd1 vccd1 vccd1
+ _0027_ sky130_fd_sc_hd__mux2_1
X_1809_ _0429_ _0433_ _0437_ _0438_ vssd1 vssd1 vccd1 vccd1 _0439_ sky130_fd_sc_hd__a211o_1
XANTENNA__2108__A1 net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2056__B net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2595__B2 _0963_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2595__A1 _0966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3107__S net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2347__A1 _1511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2946__S net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1858__B1 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3452__SET_B net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2643_ _0966_ _1259_ _1260_ _0963_ CB_0.config_dataA\[17\] vssd1 vssd1 vccd1 vccd1
+ _1270_ sky130_fd_sc_hd__a221o_1
X_2574_ _0982_ _1186_ _1190_ _0985_ _1472_ vssd1 vssd1 vccd1 vccd1 _1201_ sky130_fd_sc_hd__a221o_1
XANTENNA__2338__A1 _0467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2712_ _1423_ SB0.route_sel\[51\] _1424_ SB0.route_sel\[52\] vssd1 vssd1 vccd1 vccd1
+ _1324_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout264_A net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3126_ CB_0.config_dataB\[12\] CB_0.config_dataB\[13\] net220 vssd1 vssd1 vccd1 vccd1
+ _0294_ sky130_fd_sc_hd__mux2_1
X_3057_ SB0.route_sel\[97\] SB0.route_sel\[96\] net298 vssd1 vssd1 vccd1 vccd1 _0225_
+ sky130_fd_sc_hd__mux2_1
X_2008_ net201 net312 _0616_ net200 vssd1 vssd1 vccd1 vccd1 _0638_ sky130_fd_sc_hd__o211a_1
XANTENNA__2604__B net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2577__A1 net24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2026__B1 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1785__C1 SB0.route_sel\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2354__X _0982_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2290_ net170 _0917_ _0918_ vssd1 vssd1 vccd1 vccd1 _0919_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_47_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clone18_C1 _0974_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1767__C1 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput100 net100 vssd1 vssd1 vccd1 vccd1 CBnorth_out[6] sky130_fd_sc_hd__buf_6
Xoutput122 net122 vssd1 vssd1 vccd1 vccd1 SBwest_out[11] sky130_fd_sc_hd__buf_8
Xoutput133 net133 vssd1 vssd1 vccd1 vccd1 SBwest_out[7] sky130_fd_sc_hd__buf_8
X_2557_ net310 LEI0.config_data\[14\] _1182_ vssd1 vssd1 vccd1 vccd1 _1184_ sky130_fd_sc_hd__or3_1
X_2626_ net147 net159 LEI0.config_data\[36\] vssd1 vssd1 vccd1 vccd1 _1253_ sky130_fd_sc_hd__mux2_1
Xoutput111 net111 vssd1 vssd1 vccd1 vccd1 SBsouth_out[1] sky130_fd_sc_hd__buf_6
X_2488_ net32 _1109_ vssd1 vssd1 vccd1 vccd1 _1116_ sky130_fd_sc_hd__nand2_1
XFILLER_28_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3109_ CB_0.config_dataA\[20\] CB_0.config_dataA\[21\] net227 vssd1 vssd1 vccd1 vccd1
+ _0277_ sky130_fd_sc_hd__mux2_1
XFILLER_55_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_38_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2262__A3 net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2349__X _0977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1790_ CB_0.config_dataA\[23\] CB_0.config_dataA\[22\] _1514_ vssd1 vssd1 vccd1 vccd1
+ _0420_ sky130_fd_sc_hd__or3_2
Xinput13 CBeast_in[6] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_44_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1700__Y _1538_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput24 CBnorth_in[1] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__buf_2
X_3460_ clknet_leaf_13_clk _0280_ net278 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[24\]
+ sky130_fd_sc_hd__dfstp_1
X_2411_ net183 net182 vssd1 vssd1 vccd1 vccd1 _1039_ sky130_fd_sc_hd__nor2_1
X_3391_ clknet_leaf_28_clk _0211_ net252 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[83\]
+ sky130_fd_sc_hd__dfstp_1
Xinput35 SBsouth_in[11] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__buf_1
Xinput46 SBsouth_in[7] vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__clkbuf_1
Xinput68 le_clk vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__buf_1
Xinput57 SBwest_in[2] vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__buf_1
XANTENNA__1764__A2 _0384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2342_ net17 net24 net25 net26 net185 net184 vssd1 vssd1 vccd1 vccd1 _0970_ sky130_fd_sc_hd__mux4_1
X_2273_ _0867_ _0868_ _0900_ _0901_ _0898_ vssd1 vssd1 vccd1 vccd1 _0902_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout227_A net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_12_clk_A clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1988_ net168 net161 net2 vssd1 vssd1 vccd1 vccd1 _0618_ sky130_fd_sc_hd__o21ai_1
XANTENNA__2154__B _0783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2609_ net31 net32 net18 net19 CB_0.config_dataA\[10\] CB_0.config_dataA\[11\] vssd1
+ vssd1 vccd1 vccd1 _1236_ sky130_fd_sc_hd__mux4_1
XFILLER_57_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_27_clk_A clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_2_2__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_2_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
Xfanout190 CB_0.config_dataA\[6\] vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__clkbuf_2
XANTENNA__2459__A0 net20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2954__S net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2960_ SB0.route_sel\[0\] CB_1.config_dataB\[24\] net293 vssd1 vssd1 vccd1 vccd1
+ _0128_ sky130_fd_sc_hd__mux2_1
XFILLER_63_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1911_ SB0.route_sel\[119\] SB0.route_sel\[118\] vssd1 vssd1 vccd1 vccd1 _0541_ sky130_fd_sc_hd__nand2b_1
X_2891_ net393 net384 net213 vssd1 vssd1 vccd1 vccd1 _0060_ sky130_fd_sc_hd__mux2_1
X_1773_ _0401_ _0402_ CB_1.config_dataB\[2\] vssd1 vssd1 vccd1 vccd1 _0403_ sky130_fd_sc_hd__mux2_4
X_1842_ SB0.route_sel\[10\] SB0.route_sel\[11\] vssd1 vssd1 vccd1 vccd1 _0472_ sky130_fd_sc_hd__and2_1
X_3443_ clknet_leaf_7_clk _0263_ net259 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[7\]
+ sky130_fd_sc_hd__dfstp_1
X_3374_ clknet_leaf_12_clk _0194_ net275 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[66\]
+ sky130_fd_sc_hd__dfstp_1
X_3512_ clknet_leaf_32_clk net459 net241 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_57_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2187_ _0813_ _0814_ _0815_ vssd1 vssd1 vccd1 vccd1 _0816_ sky130_fd_sc_hd__a21o_1
X_2325_ CB_0.config_dataB\[3\] CB_0.config_dataB\[2\] CB_0.config_dataB\[4\] _0952_
+ vssd1 vssd1 vccd1 vccd1 _0953_ sky130_fd_sc_hd__or4bb_1
XANTENNA_clone31_C1 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2256_ _0883_ _0884_ vssd1 vssd1 vccd1 vccd1 _0885_ sky130_fd_sc_hd__nor2_1
XANTENNA__2217__A3 net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclone16 net143 vssd1 vssd1 vccd1 vccd1 net326 sky130_fd_sc_hd__buf_6
XANTENNA__2386__C1 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclone38 _0675_ _0665_ _0678_ net309 vssd1 vssd1 vccd1 vccd1 net348 sky130_fd_sc_hd__a211o_1
Xclone49 _0487_ _0481_ _0490_ net306 vssd1 vssd1 vccd1 vccd1 net359 sky130_fd_sc_hd__a211o_1
XFILLER_56_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_54_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input62_X net62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3090_ net192 CB_0.config_dataA\[2\] net218 vssd1 vssd1 vccd1 vccd1 _0258_ sky130_fd_sc_hd__mux2_1
XFILLER_47_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2110_ net362 _0729_ _0733_ net348 CB_1.config_dataB\[12\] vssd1 vssd1 vccd1 vccd1
+ _0740_ sky130_fd_sc_hd__a221o_1
X_2041_ SB0.route_sel\[71\] SB0.route_sel\[70\] vssd1 vssd1 vccd1 vccd1 _0671_ sky130_fd_sc_hd__nand2_1
X_2943_ CB_1.config_dataB\[7\] CB_1.config_dataB\[8\] net228 vssd1 vssd1 vccd1 vccd1
+ _0111_ sky130_fd_sc_hd__mux2_1
XFILLER_22_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1756_ CB_0.config_dataB\[21\] CB_0.config_dataB\[20\] CB_0.config_dataB\[24\] vssd1
+ vssd1 vccd1 vccd1 _0386_ sky130_fd_sc_hd__or3_2
XANTENNA_clone26_C1 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1825_ _0452_ _0453_ _0454_ vssd1 vssd1 vccd1 vccd1 _0455_ sky130_fd_sc_hd__a21bo_1
X_2874_ LEI0.config_data\[42\] net488 net210 vssd1 vssd1 vccd1 vccd1 _0043_ sky130_fd_sc_hd__mux2_1
X_3426_ clknet_leaf_15_clk _0246_ net281 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[118\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_fanout294_A net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3357_ clknet_leaf_25_clk _0177_ net268 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[49\]
+ sky130_fd_sc_hd__dfstp_1
X_2308_ CB_1.config_dataA\[18\] _0926_ _0936_ CB_1.config_dataA\[19\] vssd1 vssd1
+ vccd1 vccd1 _0937_ sky130_fd_sc_hd__a211oi_1
X_1687_ _1422_ SB0.route_sel\[48\] SB0.route_sel\[53\] SB0.route_sel\[52\] _1524_
+ vssd1 vssd1 vccd1 vccd1 _1525_ sky130_fd_sc_hd__o221a_1
X_3288_ clknet_leaf_18_clk _0108_ net279 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[5\]
+ sky130_fd_sc_hd__dfstp_1
X_2239_ LE_1A.config_data\[15\] LE_1A.config_data\[14\] _0836_ vssd1 vssd1 vccd1 vccd1
+ _0868_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2071__A1 net12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3227__Q CB_0.config_data_inA vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input22_A CBnorth_in[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3087__A0 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2357__X _0985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2126__A2 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output109_A net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output90_A net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2590_ LEI0.config_data\[25\] _1216_ vssd1 vssd1 vccd1 vccd1 _1217_ sky130_fd_sc_hd__nor2_1
X_1610_ SB0.route_sel\[5\] vssd1 vssd1 vccd1 vccd1 _1448_ sky130_fd_sc_hd__inv_2
X_3142_ CB_1.config_dataA\[3\] CB_1.config_dataA\[4\] net230 vssd1 vssd1 vccd1 vccd1
+ _0310_ sky130_fd_sc_hd__mux2_1
XANTENNA__2117__A2 net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3211_ clknet_leaf_28_clk _0031_ net251 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_65_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3073_ SB0.route_sel\[113\] SB0.route_sel\[112\] net299 vssd1 vssd1 vccd1 vccd1 _0241_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__3475__SET_B net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2024_ net144 _0652_ net234 vssd1 vssd1 vccd1 vccd1 _0654_ sky130_fd_sc_hd__o21ai_1
XANTENNA__2708__A SB0.route_sel\[63\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2857_ net478 LEI0.config_data\[26\] net214 vssd1 vssd1 vccd1 vccd1 _0026_ sky130_fd_sc_hd__mux2_1
X_2926_ net404 LE_1A.config_data\[10\] net210 vssd1 vssd1 vccd1 vccd1 _0095_ sky130_fd_sc_hd__mux2_1
X_2788_ net152 _0985_ _0387_ vssd1 vssd1 vccd1 vccd1 _1371_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout307_A net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1808_ SB0.route_sel\[25\] SB0.route_sel\[24\] vssd1 vssd1 vccd1 vccd1 _0438_ sky130_fd_sc_hd__nand2_1
X_1739_ SB0.route_sel\[47\] SB0.route_sel\[46\] vssd1 vssd1 vccd1 vccd1 _0369_ sky130_fd_sc_hd__nand2b_1
XFILLER_58_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2108__A2 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3409_ clknet_leaf_19_clk _0229_ net271 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[101\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__2292__B2 _0679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2292__A1 _0659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2044__A1 net47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2347__A2 _1510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input25_X net25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3123__S net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1858__A1 _0481_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2711_ SB0.route_sel\[49\] SB0.route_sel\[48\] vssd1 vssd1 vccd1 vccd1 _1323_ sky130_fd_sc_hd__or2_1
X_2642_ _0956_ _0959_ net187 vssd1 vssd1 vccd1 vccd1 _1269_ sky130_fd_sc_hd__mux2_1
X_2573_ _0975_ _0978_ net191 vssd1 vssd1 vccd1 vccd1 _1200_ sky130_fd_sc_hd__mux2_1
XANTENNA__2338__A2 _0461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3125_ net180 CB_0.config_dataB\[12\] net219 vssd1 vssd1 vccd1 vccd1 _0293_ sky130_fd_sc_hd__mux2_1
X_3056_ SB0.route_sel\[96\] SB0.route_sel\[95\] net295 vssd1 vssd1 vccd1 vccd1 _0224_
+ sky130_fd_sc_hd__mux2_1
X_2007_ _0633_ _0627_ _0636_ net307 vssd1 vssd1 vccd1 vccd1 _0637_ sky130_fd_sc_hd__a211o_4
XTAP_TAPCELL_ROW_25_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2725__X net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2274__A1 _0829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2577__A2 net25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2026__A1 _0655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2909_ net389 LE_0B.config_data\[11\] net206 vssd1 vssd1 vccd1 vccd1 _0078_ sky130_fd_sc_hd__mux2_1
XANTENNA__2017__A1 net48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2265__B2 _0397_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2265__A1 _0371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2370__X _0998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1776__B1 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1714__X _1552_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clone18_B1 _1522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1767__B1 _0396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput101 net101 vssd1 vssd1 vccd1 vccd1 CBnorth_out[7] sky130_fd_sc_hd__buf_6
Xoutput123 net123 vssd1 vssd1 vccd1 vccd1 SBwest_out[12] sky130_fd_sc_hd__buf_6
X_2487_ net18 net19 net179 vssd1 vssd1 vccd1 vccd1 _1115_ sky130_fd_sc_hd__mux2_1
X_2625_ LE_0A.config_data\[1\] _1180_ _1211_ _1251_ vssd1 vssd1 vccd1 vccd1 _1252_
+ sky130_fd_sc_hd__o211a_1
Xoutput134 net134 vssd1 vssd1 vccd1 vccd1 SBwest_out[8] sky130_fd_sc_hd__buf_8
X_2556_ net143 net156 LEI0.config_data\[12\] vssd1 vssd1 vccd1 vccd1 _1183_ sky130_fd_sc_hd__mux2_1
XANTENNA_clone34_C1 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput112 net112 vssd1 vssd1 vccd1 vccd1 SBsouth_out[2] sky130_fd_sc_hd__buf_4
XANTENNA__3325__Q SB0.route_sel\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3108_ CB_0.config_dataA\[19\] CB_0.config_dataA\[20\] net227 vssd1 vssd1 vccd1 vccd1
+ _0276_ sky130_fd_sc_hd__mux2_1
XANTENNA__2495__B2 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2495__A1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3039_ SB0.route_sel\[79\] SB0.route_sel\[78\] net290 vssd1 vssd1 vccd1 vccd1 _0207_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__1758__B1 net27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput25 CBnorth_in[2] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__buf_2
Xinput14 CBeast_in[7] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__buf_8
Xinput36 SBsouth_in[12] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__buf_1
X_2341_ net184 _0960_ _0968_ vssd1 vssd1 vccd1 vccd1 _0969_ sky130_fd_sc_hd__a21o_1
X_2410_ net341 net338 net183 vssd1 vssd1 vccd1 vccd1 _1038_ sky130_fd_sc_hd__mux2_1
X_3390_ clknet_leaf_3_clk _0210_ net251 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[82\]
+ sky130_fd_sc_hd__dfstp_1
Xinput58 SBwest_in[3] vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__buf_1
Xinput69 le_en vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__clkbuf_2
Xinput47 SBsouth_in[8] vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__dlymetal6s2s_1
X_2272_ LE_1A.config_data\[13\] net311 _0866_ vssd1 vssd1 vccd1 vccd1 _0901_ sky130_fd_sc_hd__o21a_1
XFILLER_60_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2229__A1 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clone29_C1 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1988__B1 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1987_ SB0.route_sel\[82\] SB0.route_sel\[83\] vssd1 vssd1 vccd1 vccd1 _0617_ sky130_fd_sc_hd__nand2_1
X_2608_ net20 net22 net21 net23 CB_0.config_dataA\[11\] CB_0.config_dataA\[10\] vssd1
+ vssd1 vccd1 vccd1 _1235_ sky130_fd_sc_hd__mux4_1
X_2539_ _1164_ _1165_ CB_0.config_dataA\[2\] vssd1 vssd1 vccd1 vccd1 _1166_ sky130_fd_sc_hd__mux2_1
XFILLER_51_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input52_A SBwest_in[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout191 CB_0.config_dataA\[5\] vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__buf_2
XANTENNA__2459__A1 net22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout180 CB_0.config_dataB\[11\] vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1910_ _0533_ _0539_ net309 vssd1 vssd1 vccd1 vccd1 _0540_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_57_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2890_ net419 net393 net216 vssd1 vssd1 vccd1 vccd1 _0059_ sky130_fd_sc_hd__mux2_1
XFILLER_34_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1772_ net11 net12 net13 net14 net201 net200 vssd1 vssd1 vccd1 vccd1 _0402_ sky130_fd_sc_hd__mux4_2
X_3511_ clknet_leaf_1_clk _0331_ net244 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_1841_ _0467_ _0461_ _0470_ net306 vssd1 vssd1 vccd1 vccd1 _0471_ sky130_fd_sc_hd__a211o_4
X_3442_ clknet_leaf_7_clk _0262_ net259 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[6\]
+ sky130_fd_sc_hd__dfstp_1
X_2324_ net184 net185 vssd1 vssd1 vccd1 vccd1 _0952_ sky130_fd_sc_hd__and2b_1
X_3373_ clknet_leaf_11_clk _0193_ net275 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[65\]
+ sky130_fd_sc_hd__dfstp_1
X_2186_ _0584_ _0804_ _0807_ _0564_ _1450_ vssd1 vssd1 vccd1 vccd1 _0815_ sky130_fd_sc_hd__a221o_1
X_2255_ _0584_ _0873_ _0876_ _0564_ _1461_ vssd1 vssd1 vccd1 vccd1 _0884_ sky130_fd_sc_hd__a221o_1
Xclone28 _0611_ _0602_ _0993_ net307 vssd1 vssd1 vccd1 vccd1 net338 sky130_fd_sc_hd__a211o_1
Xclone39 _0580_ _0570_ _0583_ net310 vssd1 vssd1 vccd1 vccd1 net349 sky130_fd_sc_hd__a211o_1
Xclone17 _0424_ _0415_ _0427_ net303 vssd1 vssd1 vccd1 vccd1 net327 sky130_fd_sc_hd__a211o_1
XANTENNA__2386__B1 _1013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Left_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2377__A0 net20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3126__S net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input55_X net55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_11_clk_A clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2040_ _0667_ _0668_ _0669_ vssd1 vssd1 vccd1 vccd1 _0670_ sky130_fd_sc_hd__a21bo_1
XFILLER_62_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2942_ net198 CB_1.config_dataB\[7\] net228 vssd1 vssd1 vccd1 vccd1 _0110_ sky130_fd_sc_hd__mux2_1
X_2873_ LEI0.config_data\[41\] LEI0.config_data\[42\] net211 vssd1 vssd1 vccd1 vccd1
+ _0042_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_26_clk_A clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1755_ CB_0.config_dataB\[21\] CB_0.config_dataB\[20\] CB_0.config_dataB\[24\] vssd1
+ vssd1 vccd1 vccd1 _0385_ sky130_fd_sc_hd__nor3_1
X_1824_ net148 _0375_ _0407_ net235 vssd1 vssd1 vccd1 vccd1 _0454_ sky130_fd_sc_hd__o31a_1
X_1686_ SB0.route_sel\[55\] SB0.route_sel\[54\] vssd1 vssd1 vccd1 vccd1 _1524_ sky130_fd_sc_hd__nand2b_1
X_3425_ clknet_leaf_15_clk _0245_ net281 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[117\]
+ sky130_fd_sc_hd__dfstp_1
X_3287_ clknet_leaf_19_clk _0107_ net276 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[4\]
+ sky130_fd_sc_hd__dfstp_1
X_3356_ clknet_leaf_25_clk _0176_ net268 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[48\]
+ sky130_fd_sc_hd__dfstp_1
X_2307_ _0932_ _0935_ _1463_ _0929_ vssd1 vssd1 vccd1 vccd1 _0936_ sky130_fd_sc_hd__and4bb_1
X_2238_ LEI0.config_data\[20\] net233 _0865_ _0840_ vssd1 vssd1 vccd1 vccd1 _0867_
+ sky130_fd_sc_hd__a31o_1
XFILLER_53_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2169_ _0683_ _0684_ _0689_ _1487_ vssd1 vssd1 vccd1 vccd1 _0799_ sky130_fd_sc_hd__a211o_1
XANTENNA__2071__A2 net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2126__A3 net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input15_A CBeast_in[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1886__B1_N net39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2598__A0 net27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2373__X _1001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3508__SET_B net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3141_ CB_1.config_dataA\[2\] CB_1.config_dataA\[3\] net230 vssd1 vssd1 vccd1 vccd1
+ _0309_ sky130_fd_sc_hd__mux2_1
XANTENNA_max_cap138_X net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3210_ clknet_leaf_3_clk _0030_ net251 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3072_ SB0.route_sel\[112\] SB0.route_sel\[111\] net299 vssd1 vssd1 vccd1 vccd1 _0240_
+ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_59_Left_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2023_ net151 _0650_ _0651_ _0652_ vssd1 vssd1 vccd1 vccd1 _0653_ sky130_fd_sc_hd__o211a_1
XFILLER_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clone37_C1 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2856_ LEI0.config_data\[24\] net478 net214 vssd1 vssd1 vccd1 vccd1 _0025_ sky130_fd_sc_hd__mux2_1
XANTENNA__2589__A0 net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1807_ net42 _0435_ _0436_ vssd1 vssd1 vccd1 vccd1 _0437_ sky130_fd_sc_hd__a21oi_1
X_2925_ net420 net404 net210 vssd1 vssd1 vccd1 vccd1 _0094_ sky130_fd_sc_hd__mux2_1
X_2787_ _1370_ _0364_ _0366_ vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__a21oi_2
XANTENNA__2108__A3 net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3408_ clknet_leaf_19_clk _0228_ net271 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[100\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_2_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout202_A net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1738_ _0367_ _0358_ net305 vssd1 vssd1 vccd1 vccd1 _0368_ sky130_fd_sc_hd__a21oi_2
X_1669_ SB0.route_sel\[55\] SB0.route_sel\[54\] vssd1 vssd1 vccd1 vccd1 _1507_ sky130_fd_sc_hd__nand2_1
XANTENNA_input7_A CBeast_in[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3339_ clknet_leaf_29_clk _0159_ net249 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[31\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__2029__C1 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1858__A2 _0487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output121_A net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2710_ _1549_ _1322_ vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__and2_4
X_2641_ _1258_ _1264_ _1267_ _1263_ CB_0.config_dataA\[18\] vssd1 vssd1 vccd1 vccd1
+ _1268_ sky130_fd_sc_hd__o2111a_1
X_2572_ _1471_ _1195_ _1198_ _1192_ vssd1 vssd1 vccd1 vccd1 _1199_ sky130_fd_sc_hd__or4b_1
X_3124_ net181 net180 net219 vssd1 vssd1 vccd1 vccd1 _0292_ sky130_fd_sc_hd__mux2_1
XANTENNA__2438__B net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3055_ SB0.route_sel\[95\] SB0.route_sel\[94\] net295 vssd1 vssd1 vccd1 vccd1 _0223_
+ sky130_fd_sc_hd__mux2_1
XFILLER_35_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2026__A2 _0649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2006_ SB0.route_sel\[80\] _1406_ SB0.route_sel\[85\] SB0.route_sel\[84\] _0635_
+ vssd1 vssd1 vccd1 vccd1 _0636_ sky130_fd_sc_hd__o221a_1
XFILLER_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2577__A3 net26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2908_ net400 net389 net206 vssd1 vssd1 vccd1 vccd1 _0077_ sky130_fd_sc_hd__mux2_1
X_2839_ LEI0.config_data\[7\] net462 net205 vssd1 vssd1 vccd1 vccd1 _0008_ sky130_fd_sc_hd__mux2_1
XANTENNA__2348__B SB0.route_sel\[63\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_22_Left_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_29_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2624_ _1173_ _1174_ _1179_ LE_0A.config_data\[0\] vssd1 vssd1 vccd1 vccd1 _1251_
+ sky130_fd_sc_hd__a211o_1
XANTENNA_clone18_A1 _1510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1767__A1 _0393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput102 net102 vssd1 vssd1 vccd1 vccd1 CBnorth_out[8] sky130_fd_sc_hd__buf_6
Xoutput124 net124 vssd1 vssd1 vccd1 vccd1 SBwest_out[13] sky130_fd_sc_hd__buf_8
X_2486_ net313 net336 net341 net338 net179 net178 vssd1 vssd1 vccd1 vccd1 _1114_ sky130_fd_sc_hd__mux4_1
Xoutput135 net135 vssd1 vssd1 vccd1 vccd1 SBwest_out[9] sky130_fd_sc_hd__buf_8
XANTENNA__2192__A1 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2555_ LEI0.config_data\[12\] _1493_ _1181_ LEI0.config_data\[13\] vssd1 vssd1 vccd1
+ vccd1 _1182_ sky130_fd_sc_hd__o211a_1
XANTENNA_clone34_B1 _0448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput113 net113 vssd1 vssd1 vccd1 vccd1 SBsouth_out[3] sky130_fd_sc_hd__buf_6
X_3107_ CB_0.config_dataA\[18\] CB_0.config_dataA\[19\] net220 vssd1 vssd1 vccd1 vccd1
+ _0275_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_38_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3038_ SB0.route_sel\[78\] SB0.route_sel\[77\] net289 vssd1 vssd1 vccd1 vccd1 _0206_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_21_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2955__A0 CB_1.config_dataB\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1815__X _0445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2238__A2 net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput26 CBnorth_in[3] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__buf_2
XANTENNA__2541__B net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput15 CBeast_in[8] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__buf_2
Xinput59 SBwest_in[4] vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__buf_1
Xinput48 SBsouth_in[9] vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput37 SBsouth_in[13] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__buf_1
X_2340_ _0952_ net371 net319 _0967_ CB_0.config_dataB\[2\] vssd1 vssd1 vccd1 vccd1
+ _0968_ sky130_fd_sc_hd__a221o_1
X_2271_ LE_1A.config_data\[12\] _0836_ vssd1 vssd1 vccd1 vccd1 _0900_ sky130_fd_sc_hd__nand2b_1
XANTENNA__2229__A2 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1685__B1 _1522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clone29_B1 _0958_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1986_ _0602_ _0611_ _0614_ _1478_ net307 vssd1 vssd1 vccd1 vccd1 _0616_ sky130_fd_sc_hd__a2111o_1
Xclkbuf_leaf_9_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2607_ _1232_ _1233_ vssd1 vssd1 vccd1 vccd1 _1234_ sky130_fd_sc_hd__nor2_1
X_2538_ net20 net22 net21 net23 net192 CB_0.config_dataA\[0\] vssd1 vssd1 vccd1 vccd1
+ _1165_ sky130_fd_sc_hd__mux4_1
X_2469_ LEI0.config_data\[29\] net233 vssd1 vssd1 vccd1 vccd1 _1097_ sky130_fd_sc_hd__nand2_1
XFILLER_28_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1903__A1 _0527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input45_A SBsouth_in[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout192 CB_0.config_dataA\[1\] vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_57_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2459__A2 net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout181 CB_0.config_dataB\[10\] vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__buf_2
Xfanout170 CB_1.config_dataA\[16\] vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__buf_2
XANTENNA__2631__A2 _1014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1840_ _1446_ SB0.route_sel\[0\] SB0.route_sel\[5\] SB0.route_sel\[4\] _0469_ vssd1
+ vssd1 vccd1 vccd1 _0470_ sky130_fd_sc_hd__o221a_1
X_3441_ clknet_leaf_8_clk _0261_ net260 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[5\]
+ sky130_fd_sc_hd__dfstp_1
X_1771_ net1 net8 net9 net10 net201 net200 vssd1 vssd1 vccd1 vccd1 _0401_ sky130_fd_sc_hd__mux4_2
X_3510_ clknet_leaf_23_clk _0330_ net274 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[24\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_8_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2147__A1 net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clone31_A1 _0633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3372_ clknet_leaf_27_clk _0192_ net252 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[64\]
+ sky130_fd_sc_hd__dfstp_1
X_2254_ net173 _0543_ _0882_ net172 vssd1 vssd1 vccd1 vccd1 _0883_ sky130_fd_sc_hd__o211a_1
XANTENNA__2147__B2 net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2323_ _0950_ LEI0.config_data_in _0951_ net232 vssd1 vssd1 vccd1 vccd1 CB_1.le_outA
+ sky130_fd_sc_hd__o211a_1
X_2185_ net177 _0543_ net176 vssd1 vssd1 vccd1 vccd1 _0814_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_40_Left_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_25_Left_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2386__A1 _0539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclone18 _1510_ _1511_ _1522_ _0974_ vssd1 vssd1 vccd1 vccd1 net328 sky130_fd_sc_hd__a211o_4
Xclone29 _0445_ _0439_ _0958_ net305 vssd1 vssd1 vccd1 vccd1 net339 sky130_fd_sc_hd__a211o_1
XFILLER_33_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1969_ SB0.route_sel\[93\] SB0.route_sel\[92\] net51 _0597_ _0590_ vssd1 vssd1 vccd1
+ vccd1 _0599_ sky130_fd_sc_hd__a41o_1
XANTENNA_fanout232_A net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2138__B2 net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2138__A1 net12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2377__A1 net22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input48_X net48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2301__A1 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clone26_A1 _0655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2941_ net199 net198 net228 vssd1 vssd1 vccd1 vccd1 _0109_ sky130_fd_sc_hd__mux2_1
XFILLER_30_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2872_ net444 LEI0.config_data\[41\] net208 vssd1 vssd1 vccd1 vccd1 _0041_ sky130_fd_sc_hd__mux2_1
X_1823_ net157 net165 net163 _0407_ _0375_ vssd1 vssd1 vccd1 vccd1 _0453_ sky130_fd_sc_hd__o32a_1
X_3424_ clknet_leaf_15_clk _0244_ net281 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[116\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_clone42_B1 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1685_ _1510_ _1511_ _1522_ vssd1 vssd1 vccd1 vccd1 _1523_ sky130_fd_sc_hd__a21oi_1
X_1754_ _0372_ _0378_ _0382_ _0383_ vssd1 vssd1 vccd1 vccd1 _0384_ sky130_fd_sc_hd__a211o_1
XANTENNA__1913__X _0543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3286_ clknet_leaf_19_clk _0106_ net270 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[3\]
+ sky130_fd_sc_hd__dfstp_1
X_3355_ clknet_leaf_25_clk _0175_ net267 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[47\]
+ sky130_fd_sc_hd__dfstp_1
X_2306_ net170 _0933_ _0934_ vssd1 vssd1 vccd1 vccd1 _0935_ sky130_fd_sc_hd__a21oi_1
XANTENNA__1879__B1 net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2237_ LEI0.config_data\[20\] net232 _0865_ net141 vssd1 vssd1 vccd1 vccd1 _0866_
+ sky130_fd_sc_hd__a31oi_4
XFILLER_53_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2099_ _1484_ net196 vssd1 vssd1 vccd1 vccd1 _0729_ sky130_fd_sc_hd__nor2_1
XFILLER_38_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2168_ _1490_ _0690_ _0723_ _0797_ vssd1 vssd1 vccd1 vccd1 _0798_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_17_Right_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2531__B2 _0966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2531__A1 _0963_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_26_Right_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2784__B1_N _0975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2598__A1 net28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_35_Right_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2770__A1 _1018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2830__A net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3071_ SB0.route_sel\[111\] SB0.route_sel\[110\] net299 vssd1 vssd1 vccd1 vccd1 _0239_
+ sky130_fd_sc_hd__mux2_1
X_3140_ net176 CB_1.config_dataA\[2\] net230 vssd1 vssd1 vccd1 vccd1 _0308_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_44_Right_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_53_Right_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2022_ _0363_ _0607_ vssd1 vssd1 vccd1 vccd1 _0652_ sky130_fd_sc_hd__or2_1
XFILLER_50_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2786_ net152 _0982_ _0361_ vssd1 vssd1 vccd1 vccd1 _1370_ sky130_fd_sc_hd__mux2_1
XANTENNA_clone37_B1 _0977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2855_ LEI0.config_data\[23\] LEI0.config_data\[24\] net207 vssd1 vssd1 vccd1 vccd1
+ _0024_ sky130_fd_sc_hd__mux2_1
X_2924_ net443 net420 net210 vssd1 vssd1 vccd1 vccd1 _0093_ sky130_fd_sc_hd__mux2_1
X_1806_ SB0.route_sel\[29\] SB0.route_sel\[28\] net58 _0434_ _0429_ vssd1 vssd1 vccd1
+ vccd1 _0436_ sky130_fd_sc_hd__a41o_1
XPHY_EDGE_ROW_62_Right_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1737_ _0366_ _0365_ _0357_ vssd1 vssd1 vccd1 vccd1 _0367_ sky130_fd_sc_hd__or3b_4
X_3407_ clknet_leaf_19_clk _0227_ net271 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[99\]
+ sky130_fd_sc_hd__dfstp_1
X_3338_ clknet_leaf_29_clk _0158_ net249 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[30\]
+ sky130_fd_sc_hd__dfstp_1
X_1599_ SB0.route_sel\[28\] vssd1 vssd1 vccd1 vccd1 _1437_ sky130_fd_sc_hd__inv_2
X_1668_ _1500_ _1503_ _1505_ vssd1 vssd1 vccd1 vccd1 _1506_ sky130_fd_sc_hd__a21bo_1
X_3269_ clknet_leaf_32_clk net392 net242 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_11_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_10_clk_A clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1818__X _0448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_25_clk_A clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2640_ _1261_ _1266_ CB_0.config_dataA\[17\] vssd1 vssd1 vccd1 vccd1 _1267_ sky130_fd_sc_hd__a21o_1
XANTENNA__1728__X _0358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2571_ net190 _1196_ _1197_ vssd1 vssd1 vccd1 vccd1 _1198_ sky130_fd_sc_hd__a21oi_1
XFILLER_4_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3123_ CB_0.config_dataB\[9\] net181 net219 vssd1 vssd1 vccd1 vccd1 _0291_ sky130_fd_sc_hd__mux2_1
X_3054_ SB0.route_sel\[94\] SB0.route_sel\[93\] net295 vssd1 vssd1 vccd1 vccd1 _0222_
+ sky130_fd_sc_hd__mux2_1
X_2005_ SB0.route_sel\[87\] SB0.route_sel\[86\] vssd1 vssd1 vccd1 vccd1 _0635_ sky130_fd_sc_hd__nand2b_1
XANTENNA__2735__A SB0.route_sel\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout145_A CB_0.le_outA vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2907_ net442 net400 net212 vssd1 vssd1 vccd1 vccd1 _0076_ sky130_fd_sc_hd__mux2_1
X_2769_ _1361_ _0536_ _0538_ vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__a21oi_4
XFILLER_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1785__A2 _0410_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2838_ LEI0.config_data\[6\] net479 net205 vssd1 vssd1 vccd1 vccd1 _0007_ sky130_fd_sc_hd__mux2_1
XANTENNA__2498__A0 net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clone20_A CBeast_in[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input30_X net30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clone18_A2 _1511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput103 net103 vssd1 vssd1 vccd1 vccd1 CBnorth_out[9] sky130_fd_sc_hd__buf_6
Xoutput125 net125 vssd1 vssd1 vccd1 vccd1 SBwest_out[14] sky130_fd_sc_hd__buf_6
X_2623_ LE_0A.config_data\[3\] _1180_ _1212_ _1249_ vssd1 vssd1 vccd1 vccd1 _1250_
+ sky130_fd_sc_hd__o211a_1
X_2554_ LEI0.config_data\[12\] CB_1.le_outB vssd1 vssd1 vccd1 vccd1 _1181_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_30_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clone34_A1 _0445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput114 net114 vssd1 vssd1 vccd1 vccd1 SBsouth_out[4] sky130_fd_sc_hd__buf_8
XANTENNA__1767__A2 _0384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2485_ net179 net178 vssd1 vssd1 vccd1 vccd1 _1113_ sky130_fd_sc_hd__nor2_1
XANTENNA__2192__A2 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput136 net136 vssd1 vssd1 vccd1 vccd1 config_data_out sky130_fd_sc_hd__buf_2
X_3106_ CB_0.config_dataA\[17\] CB_0.config_dataA\[18\] net220 vssd1 vssd1 vccd1 vccd1
+ _0274_ sky130_fd_sc_hd__mux2_1
XANTENNA__2184__B _0521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout262_A net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3037_ SB0.route_sel\[77\] SB0.route_sel\[76\] net289 vssd1 vssd1 vccd1 vccd1 _0205_
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2752__X net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2506__B1_N net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1831__X _0461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1997__A2 _0621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2238__A3 _0865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput27 CBnorth_in[4] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__buf_2
Xinput16 CBeast_in[9] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__buf_2
Xinput38 SBsouth_in[14] vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput49 SBwest_in[0] vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__buf_1
XFILLER_6_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2270_ LEI0.config_data\[32\] net232 _0897_ _0872_ vssd1 vssd1 vccd1 vccd1 _0899_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__2634__A0 _1001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_35_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1685__A1 _1510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2331__C1 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1741__X _0371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clone29_A1 _0445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1985_ _0611_ _0602_ _0614_ net307 vssd1 vssd1 vccd1 vccd1 _0615_ sky130_fd_sc_hd__a211o_4
X_2537_ net31 net32 net18 net19 CB_0.config_dataA\[0\] CB_0.config_dataA\[1\] vssd1
+ vssd1 vccd1 vccd1 _1164_ sky130_fd_sc_hd__mux4_1
X_2606_ _1021_ _1220_ _1221_ _1018_ _1474_ vssd1 vssd1 vccd1 vccd1 _1233_ sky130_fd_sc_hd__a221o_1
XANTENNA_clone61_C1 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2468_ _1083_ _1095_ _1072_ vssd1 vssd1 vccd1 vccd1 _1096_ sky130_fd_sc_hd__a21oi_1
X_2399_ net143 net156 LEI0.config_data\[3\] vssd1 vssd1 vccd1 vccd1 _1027_ sky130_fd_sc_hd__mux2_1
XFILLER_28_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input38_A SBsouth_in[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout193 CB_0.config_dataA\[0\] vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__buf_2
XANTENNA__2459__A3 net23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout182 CB_0.config_dataB\[6\] vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__buf_2
Xfanout160 CB_1.le_outB vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__clkbuf_4
Xfanout171 CB_1.config_dataA\[15\] vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__buf_2
XFILLER_42_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1770_ net200 _1553_ _0399_ vssd1 vssd1 vccd1 vccd1 _0400_ sky130_fd_sc_hd__a21oi_1
X_3440_ clknet_leaf_8_clk _0260_ net260 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[4\]
+ sky130_fd_sc_hd__dfstp_1
X_3371_ clknet_leaf_24_clk _0191_ net268 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[63\]
+ sky130_fd_sc_hd__dfstp_1
X_2184_ net177 _0521_ vssd1 vssd1 vccd1 vccd1 _0813_ sky130_fd_sc_hd__nand2_1
XANTENNA_clone31_A2 _0627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2253_ net173 _0521_ vssd1 vssd1 vccd1 vccd1 _0882_ sky130_fd_sc_hd__nand2_1
X_2322_ LE_1A.dff_out LEI0.config_data_in vssd1 vssd1 vccd1 vccd1 _0951_ sky130_fd_sc_hd__nand2b_1
XANTENNA__2386__A2 _0533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1899_ SB0.route_sel\[116\] SB0.route_sel\[117\] net54 vssd1 vssd1 vccd1 vccd1 _0529_
+ sky130_fd_sc_hd__and3_1
Xclone19 net152 vssd1 vssd1 vccd1 vccd1 net329 sky130_fd_sc_hd__clkbuf_1
XANTENNA_fanout225_A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1968_ SB0.route_sel\[93\] SB0.route_sel\[92\] vssd1 vssd1 vccd1 vccd1 _0598_ sky130_fd_sc_hd__nand2_1
XFILLER_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_3_165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclone1 _0829_ _0830_ _0835_ vssd1 vssd1 vccd1 vccd1 net311 sky130_fd_sc_hd__a21oi_4
XANTENNA__2310__A2 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3023__A0 SB0.route_sel\[63\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2377__A2 net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2547__B net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2065__A1 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2940_ CB_1.config_dataB\[4\] net199 net229 vssd1 vssd1 vccd1 vccd1 _0108_ sky130_fd_sc_hd__mux2_1
XFILLER_22_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2301__A2 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clone26_A2 _0649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2871_ net457 net444 net208 vssd1 vssd1 vccd1 vccd1 _0040_ sky130_fd_sc_hd__mux2_1
X_1822_ _0373_ _0405_ net1 vssd1 vssd1 vccd1 vccd1 _0452_ sky130_fd_sc_hd__o21ai_1
X_1753_ SB0.route_sel\[33\] SB0.route_sel\[32\] vssd1 vssd1 vccd1 vccd1 _0383_ sky130_fd_sc_hd__nand2_1
X_3423_ clknet_leaf_15_clk _0243_ net282 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[115\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_clone42_A1 _0562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1684_ _1521_ _1512_ net308 vssd1 vssd1 vccd1 vccd1 _1522_ sky130_fd_sc_hd__a21o_4
X_3354_ clknet_leaf_25_clk _0174_ net266 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[46\]
+ sky130_fd_sc_hd__dfstp_1
X_2236_ _0853_ _0863_ _0864_ vssd1 vssd1 vccd1 vccd1 _0865_ sky130_fd_sc_hd__a21o_2
X_3285_ clknet_leaf_19_clk _0105_ net270 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[2\]
+ sky130_fd_sc_hd__dfstp_2
XTAP_TAPCELL_ROW_0_135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2167_ _0683_ _0684_ _0689_ _1489_ vssd1 vssd1 vccd1 vccd1 _0797_ sky130_fd_sc_hd__a211o_1
X_2305_ _0491_ _0911_ _0914_ _0471_ CB_1.config_dataA\[17\] vssd1 vssd1 vccd1 vccd1
+ _0934_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_51_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2098_ LEI0.config_data\[34\] _0726_ _0727_ vssd1 vssd1 vccd1 vccd1 _0728_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_0_146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout228_X net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2295__B2 net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2295__A1 net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2598__A2 net29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2830__B net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1666__A_N net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input60_X net60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3070_ SB0.route_sel\[110\] SB0.route_sel\[109\] net300 vssd1 vssd1 vccd1 vccd1 _0238_
+ sky130_fd_sc_hd__mux2_1
X_2021_ _0360_ _0604_ net32 vssd1 vssd1 vccd1 vccd1 _0651_ sky130_fd_sc_hd__o21ai_1
XANTENNA__2286__B2 _0564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2286__A1 _0584_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3153__S net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clone37_A1 _1548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2923_ net381 LE_1A.config_data\[7\] net204 vssd1 vssd1 vccd1 vccd1 _0092_ sky130_fd_sc_hd__mux2_1
X_2785_ _1369_ _1520_ _1515_ vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__a21boi_2
X_1736_ net144 _0364_ net237 vssd1 vssd1 vccd1 vccd1 _0366_ sky130_fd_sc_hd__o21ai_1
X_2854_ net483 LEI0.config_data\[23\] net207 vssd1 vssd1 vccd1 vccd1 _0023_ sky130_fd_sc_hd__mux2_1
X_1805_ SB0.route_sel\[29\] SB0.route_sel\[28\] vssd1 vssd1 vccd1 vccd1 _0435_ sky130_fd_sc_hd__nand2_1
X_3406_ clknet_leaf_19_clk _0226_ net275 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[98\]
+ sky130_fd_sc_hd__dfstp_1
X_3337_ clknet_leaf_25_clk _0157_ net266 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[29\]
+ sky130_fd_sc_hd__dfstp_1
X_1598_ SB0.route_sel\[27\] vssd1 vssd1 vccd1 vccd1 _1436_ sky130_fd_sc_hd__inv_2
X_1667_ _1502_ _1501_ net320 net235 vssd1 vssd1 vccd1 vccd1 _1505_ sky130_fd_sc_hd__o31a_1
X_2219_ _0846_ _0847_ CB_1.config_dataA\[7\] vssd1 vssd1 vccd1 vccd1 _0848_ sky130_fd_sc_hd__mux2_1
XANTENNA__2755__X net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2029__A1 _0655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3199_ clknet_leaf_3_clk _0019_ net245 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_3268_ clknet_leaf_31_clk _0088_ net242 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_11_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input20_A CBnorth_in[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3295__SET_B net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output107_A net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2570_ _0998_ _1186_ _1190_ _1001_ CB_0.config_dataA\[7\] vssd1 vssd1 vccd1 vccd1
+ _1197_ sky130_fd_sc_hd__a221o_1
XANTENNA__3148__S net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1951__B1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3122_ CB_0.config_dataB\[8\] CB_0.config_dataB\[9\] net219 vssd1 vssd1 vccd1 vccd1
+ _0290_ sky130_fd_sc_hd__mux2_1
XFILLER_4_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2004_ _0633_ _0627_ net307 vssd1 vssd1 vccd1 vccd1 _0634_ sky130_fd_sc_hd__a21oi_2
X_3053_ SB0.route_sel\[93\] SB0.route_sel\[92\] net294 vssd1 vssd1 vccd1 vccd1 _0221_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__2259__B2 _0471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2259__A1 _0491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3180__Q LEI0.config_data\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2735__B SB0.route_sel\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2906_ net448 net442 net212 vssd1 vssd1 vccd1 vccd1 _0075_ sky130_fd_sc_hd__mux2_1
X_2768_ net153 _1014_ _0534_ vssd1 vssd1 vccd1 vccd1 _1361_ sky130_fd_sc_hd__mux2_2
X_2699_ _1416_ SB0.route_sel\[67\] vssd1 vssd1 vccd1 vccd1 _1315_ sky130_fd_sc_hd__nor2_1
X_2837_ LEI0.config_data\[5\] LEI0.config_data\[6\] net207 vssd1 vssd1 vccd1 vccd1
+ _0006_ sky130_fd_sc_hd__mux2_1
XANTENNA__1942__B1 net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout305_A net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1719_ CB_1.config_dataA\[24\] CB_1.config_dataA\[21\] CB_1.config_dataA\[20\] vssd1
+ vssd1 vccd1 vccd1 _0349_ sky130_fd_sc_hd__or3b_4
XANTENNA__2498__A1 net24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2380__B net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2489__A1 net31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1933__B1 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input68_A le_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input23_X net23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput126 net126 vssd1 vssd1 vccd1 vccd1 SBwest_out[15] sky130_fd_sc_hd__buf_6
X_2622_ _1173_ _1174_ _1179_ LE_0A.config_data\[2\] vssd1 vssd1 vccd1 vccd1 _1249_
+ sky130_fd_sc_hd__a211o_1
X_2553_ _1173_ _1174_ _1179_ vssd1 vssd1 vccd1 vccd1 _1180_ sky130_fd_sc_hd__a21oi_4
XANTENNA__2177__A0 _0637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clone34_A2 _0439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1924__B1 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput104 net104 vssd1 vssd1 vccd1 vccd1 SBsouth_out[0] sky130_fd_sc_hd__buf_6
Xoutput115 net115 vssd1 vssd1 vccd1 vccd1 SBsouth_out[5] sky130_fd_sc_hd__buf_8
X_3105_ net186 CB_0.config_dataA\[17\] net220 vssd1 vssd1 vccd1 vccd1 _0273_ sky130_fd_sc_hd__mux2_1
X_2484_ net179 net321 _1111_ net178 vssd1 vssd1 vccd1 vccd1 _1112_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout255_A net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3036_ SB0.route_sel\[76\] SB0.route_sel\[75\] net297 vssd1 vssd1 vccd1 vccd1 _0204_
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout308_X net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_24_clk_A clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1930__A3 net52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2340__B1 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2643__A1 _0966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2643__B2 _0963_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput28 CBnorth_in[5] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__buf_2
Xinput17 CBnorth_in[0] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__buf_2
XFILLER_52_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput39 SBsouth_in[15] vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2331__B1 _0958_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2634__A1 _0998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clone29_A2 _0439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1685__A2 _1511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1763__C_N _0383_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1984_ SB0.route_sel\[88\] _1402_ SB0.route_sel\[93\] SB0.route_sel\[92\] _0613_
+ vssd1 vssd1 vccd1 vccd1 _0614_ sky130_fd_sc_hd__o221a_1
X_2605_ net189 _1014_ _1231_ net188 vssd1 vssd1 vccd1 vccd1 _1232_ sky130_fd_sc_hd__o211a_1
X_2536_ net192 _1161_ _1162_ vssd1 vssd1 vccd1 vccd1 _1163_ sky130_fd_sc_hd__a21o_1
X_2467_ CB_0.config_dataB\[13\] _1090_ _1094_ CB_0.config_dataB\[14\] vssd1 vssd1
+ vccd1 vccd1 _1095_ sky130_fd_sc_hd__a31oi_1
XANTENNA_clone61_B1 _0962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2398_ LEI0.config_data\[5\] net233 vssd1 vssd1 vccd1 vccd1 _1026_ sky130_fd_sc_hd__nand2_2
XANTENNA__1932__X _0562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout160_X net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3019_ SB0.route_sel\[59\] SB0.route_sel\[58\] net296 vssd1 vssd1 vccd1 vccd1 _0187_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__2003__X _0633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout183 CB_0.config_dataB\[5\] vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__buf_2
Xfanout172 CB_1.config_dataA\[11\] vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__buf_2
Xfanout161 _0591_ vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__buf_2
Xfanout150 CB_1.le_outA vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__buf_8
XFILLER_59_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_57_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout194 CB_1.config_dataB\[16\] vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__buf_2
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2092__A2 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2321_ _0939_ _0949_ _0945_ _0941_ _0902_ vssd1 vssd1 vccd1 vccd1 _0950_ sky130_fd_sc_hd__a32o_1
XFILLER_6_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3370_ clknet_leaf_24_clk _0190_ net268 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[62\]
+ sky130_fd_sc_hd__dfstp_1
X_2183_ _0810_ _0811_ CB_1.config_dataA\[2\] vssd1 vssd1 vccd1 vccd1 _0812_ sky130_fd_sc_hd__mux2_1
X_2252_ _0879_ _0880_ _1461_ vssd1 vssd1 vccd1 vccd1 _0881_ sky130_fd_sc_hd__mux2_1
XFILLER_2_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2304__A0 _0428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1898_ SB0.route_sel\[118\] SB0.route_sel\[119\] vssd1 vssd1 vccd1 vccd1 _0528_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout218_A net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1967_ SB0.route_sel\[94\] SB0.route_sel\[95\] vssd1 vssd1 vccd1 vccd1 _0597_ sky130_fd_sc_hd__nand2_1
XANTENNA__2758__X net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2519_ LE_0B.dff_out LE_0B.config_data\[16\] vssd1 vssd1 vccd1 vccd1 _1147_ sky130_fd_sc_hd__nand2b_1
X_3499_ clknet_leaf_26_clk _0319_ net270 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[13\]
+ sky130_fd_sc_hd__dfstp_1
Xclone2 _0633_ _0627_ _0636_ net307 vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_3_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2310__A3 _0938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1837__X _0467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2534__A0 _0991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2377__A3 net23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input50_A SBwest_in[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2668__X CB_0.le_outA vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2065__A2 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2870_ LEI0.config_data\[38\] net457 net207 vssd1 vssd1 vccd1 vccd1 _0039_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_10_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1683_ _1520_ _1519_ _1515_ vssd1 vssd1 vccd1 vccd1 _1521_ sky130_fd_sc_hd__a21bo_1
X_1821_ SB0.route_sel\[2\] SB0.route_sel\[3\] vssd1 vssd1 vccd1 vccd1 _0451_ sky130_fd_sc_hd__nand2_1
X_1752_ net43 _0380_ _0381_ vssd1 vssd1 vccd1 vccd1 _0382_ sky130_fd_sc_hd__a21oi_1
X_3422_ clknet_leaf_14_clk _0242_ net282 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[114\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_clone42_A2 _0552_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3284_ clknet_leaf_19_clk _0104_ net270 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[1\]
+ sky130_fd_sc_hd__dfstp_1
X_3353_ clknet_leaf_25_clk _0173_ net266 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[45\]
+ sky130_fd_sc_hd__dfstp_1
X_2304_ _0428_ _0449_ net171 vssd1 vssd1 vccd1 vccd1 _0933_ sky130_fd_sc_hd__mux2_1
X_2235_ CB_1.config_dataA\[8\] _1459_ CB_1.config_dataA\[9\] _0842_ vssd1 vssd1 vccd1
+ vccd1 _0864_ sky130_fd_sc_hd__and4b_1
X_2097_ net304 LEI0.config_data\[35\] vssd1 vssd1 vccd1 vccd1 _0727_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_0_147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2166_ _0722_ _0793_ _0794_ _0795_ _0755_ vssd1 vssd1 vccd1 vccd1 _0796_ sky130_fd_sc_hd__o221ai_1
XTAP_TAPCELL_ROW_51_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_3_Right_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2999_ SB0.route_sel\[39\] SB0.route_sel\[38\] net287 vssd1 vssd1 vccd1 vccd1 _0167_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2598__A3 net30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input53_X net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2020_ _0359_ _0603_ vssd1 vssd1 vccd1 vccd1 _0650_ sky130_fd_sc_hd__nand2_1
XANTENNA_clone37_A2 _1539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2922_ net422 net381 net204 vssd1 vssd1 vccd1 vccd1 _0091_ sky130_fd_sc_hd__mux2_1
X_2853_ LEI0.config_data\[21\] net483 net206 vssd1 vssd1 vccd1 vccd1 _0022_ sky130_fd_sc_hd__mux2_1
X_1735_ net152 _0361_ _0362_ _0364_ vssd1 vssd1 vccd1 vccd1 _0365_ sky130_fd_sc_hd__o211a_1
X_2784_ _1517_ _1518_ _0975_ vssd1 vssd1 vccd1 vccd1 _1369_ sky130_fd_sc_hd__o21bai_1
X_1666_ net310 net255 vssd1 vssd1 vccd1 vccd1 _1504_ sky130_fd_sc_hd__and2b_1
X_1804_ SB0.route_sel\[31\] SB0.route_sel\[30\] vssd1 vssd1 vccd1 vccd1 _0434_ sky130_fd_sc_hd__nand2_1
XANTENNA__1940__X _0570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_37_Left_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3405_ clknet_leaf_12_clk _0225_ net275 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[97\]
+ sky130_fd_sc_hd__dfstp_1
X_3336_ clknet_leaf_29_clk _0156_ net266 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[28\]
+ sky130_fd_sc_hd__dfstp_1
X_1597_ SB0.route_sel\[24\] vssd1 vssd1 vccd1 vccd1 _1435_ sky130_fd_sc_hd__inv_2
X_3267_ clknet_leaf_31_clk _0087_ net243 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_2218_ net4 net6 net5 net7 net174 CB_1.config_dataA\[5\] vssd1 vssd1 vccd1 vccd1
+ _0847_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_46_Left_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2149_ _0771_ _0774_ _0775_ _0778_ vssd1 vssd1 vccd1 vccd1 _0779_ sky130_fd_sc_hd__a22o_1
XANTENNA__2029__A2 _0649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3198_ clknet_leaf_3_clk _0018_ net245 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_55_Left_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input13_A CBeast_in[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_64_Left_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2976__A0 SB0.route_sel\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1951__A1 _0570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3461__Q CB_0.config_dataB\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3121_ CB_0.config_dataB\[7\] CB_0.config_dataB\[8\] net219 vssd1 vssd1 vccd1 vccd1
+ _0289_ sky130_fd_sc_hd__mux2_1
X_2003_ _0631_ _0632_ _0626_ vssd1 vssd1 vccd1 vccd1 _0633_ sky130_fd_sc_hd__or3b_4
X_3052_ SB0.route_sel\[92\] SB0.route_sel\[91\] net294 vssd1 vssd1 vccd1 vccd1 _0220_
+ sky130_fd_sc_hd__mux2_1
X_2905_ net394 LE_0B.config_data\[7\] net212 vssd1 vssd1 vccd1 vccd1 _0074_ sky130_fd_sc_hd__mux2_1
X_2836_ net471 LEI0.config_data\[5\] net212 vssd1 vssd1 vccd1 vccd1 _0005_ sky130_fd_sc_hd__mux2_1
X_2767_ _0502_ _1360_ _0504_ vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__a21oi_2
X_2698_ _0656_ _1314_ vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__and2_4
X_1649_ LE_1B.config_data\[8\] vssd1 vssd1 vccd1 vccd1 _1487_ sky130_fd_sc_hd__inv_2
X_1718_ net169 net166 net12 vssd1 vssd1 vccd1 vccd1 _0348_ sky130_fd_sc_hd__o21ai_1
XANTENNA__2498__A2 net25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input5_A CBeast_in[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3319_ clknet_leaf_25_clk _0139_ net267 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[11\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__3371__Q SB0.route_sel\[63\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2186__B2 _0564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2186__A1 _0584_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1933__A1 _0552_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input16_X net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2483_ net179 net138 vssd1 vssd1 vccd1 vccd1 _1111_ sky130_fd_sc_hd__nand2_1
X_2621_ _1212_ _1213_ _1247_ _1244_ vssd1 vssd1 vccd1 vccd1 _1248_ sky130_fd_sc_hd__a211o_1
X_2552_ LEI0.config_data\[1\] _1175_ _1178_ vssd1 vssd1 vccd1 vccd1 _1179_ sky130_fd_sc_hd__o21ba_2
XANTENNA__2177__A1 _0615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput127 net127 vssd1 vssd1 vccd1 vccd1 SBwest_out[1] sky130_fd_sc_hd__buf_6
Xoutput105 net105 vssd1 vssd1 vccd1 vccd1 SBsouth_out[10] sky130_fd_sc_hd__buf_8
Xoutput116 net116 vssd1 vssd1 vccd1 vccd1 SBsouth_out[6] sky130_fd_sc_hd__clkbuf_4
X_3104_ CB_0.config_dataA\[15\] CB_0.config_dataA\[16\] net219 vssd1 vssd1 vccd1 vccd1
+ _0272_ sky130_fd_sc_hd__mux2_1
X_3035_ SB0.route_sel\[75\] SB0.route_sel\[74\] net297 vssd1 vssd1 vccd1 vccd1 _0203_
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1688__B1 _1522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2819_ _1386_ _0350_ _0351_ vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__a21boi_2
Xfanout310 net66 vssd1 vssd1 vccd1 vccd1 net310 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input8_X net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput18 CBnorth_in[10] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_2
XFILLER_54_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput29 CBnorth_in[6] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__buf_2
XFILLER_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2331__A1 _0445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2634__A2 _0991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2604_ net189 net138 vssd1 vssd1 vccd1 vccd1 _1231_ sky130_fd_sc_hd__nand2_1
X_1983_ SB0.route_sel\[95\] SB0.route_sel\[94\] vssd1 vssd1 vccd1 vccd1 _0613_ sky130_fd_sc_hd__nand2b_1
X_2535_ _0998_ _1148_ _1151_ _1001_ CB_0.config_dataA\[2\] vssd1 vssd1 vccd1 vccd1
+ _1162_ sky130_fd_sc_hd__a221o_1
XANTENNA__2570__A1 _0998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2570__B2 _1001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2466_ _1085_ _1086_ _1092_ _1093_ vssd1 vssd1 vccd1 vccd1 _1094_ sky130_fd_sc_hd__o22a_1
XANTENNA_clone61_A1 _0487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2397_ _1024_ _0988_ _0953_ vssd1 vssd1 vccd1 vccd1 _1025_ sky130_fd_sc_hd__o21a_4
X_3018_ SB0.route_sel\[58\] SB0.route_sel\[57\] net293 vssd1 vssd1 vccd1 vccd1 _0186_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__1833__B1 net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2010__B1 net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout184 CB_0.config_dataB\[1\] vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_49_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout151 net152 vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__buf_8
Xfanout195 CB_1.config_dataB\[15\] vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__buf_2
Xfanout162 _0508_ vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__buf_2
Xfanout173 CB_1.config_dataA\[10\] vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2092__A3 _0716_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2251_ net15 net16 net2 net3 CB_1.config_dataA\[10\] net172 vssd1 vssd1 vccd1 vccd1
+ _0880_ sky130_fd_sc_hd__mux4_1
X_2320_ _0866_ _0948_ _0947_ _0899_ vssd1 vssd1 vccd1 vccd1 _0949_ sky130_fd_sc_hd__a211o_1
X_2182_ net4 net6 net5 net7 CB_1.config_dataA\[1\] CB_1.config_dataA\[0\] vssd1 vssd1
+ vccd1 vccd1 _0811_ sky130_fd_sc_hd__mux4_1
XANTENNA__2068__A0 _1526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_23_clk_A clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2304__A1 _0449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1966_ _0592_ _0594_ _0595_ vssd1 vssd1 vccd1 vccd1 _0596_ sky130_fd_sc_hd__a21bo_1
X_1897_ _0524_ _0525_ _0526_ vssd1 vssd1 vccd1 vccd1 _0527_ sky130_fd_sc_hd__a21bo_1
XANTENNA__1656__A net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2240__A0 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2543__B2 _1021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2543__A1 _1018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2449_ net17 net24 net25 net26 net181 net180 vssd1 vssd1 vccd1 vccd1 _1077_ sky130_fd_sc_hd__mux4_1
XANTENNA__3082__S net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2518_ _1135_ _1141_ _1145_ _1102_ _1137_ vssd1 vssd1 vccd1 vccd1 _1146_ sky130_fd_sc_hd__o32a_4
X_3498_ clknet_leaf_26_clk _0318_ net270 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[12\]
+ sky130_fd_sc_hd__dfstp_1
Xclone3 _0675_ _0665_ _1000_ net309 vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_3_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2782__A1 _0978_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2231__A0 _1526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2534__A1 _0994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input43_A SBsouth_in[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2298__A0 _1526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1820_ net327 net344 CB_1.config_dataB\[0\] vssd1 vssd1 vccd1 vccd1 _0450_ sky130_fd_sc_hd__mux2_1
XFILLER_15_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3421_ clknet_leaf_14_clk _0241_ net282 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[113\]
+ sky130_fd_sc_hd__dfstp_1
X_1682_ _1492_ _1517_ _1518_ _1513_ _1514_ vssd1 vssd1 vccd1 vccd1 _1520_ sky130_fd_sc_hd__o32a_1
XPHY_EDGE_ROW_29_Left_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1751_ SB0.route_sel\[37\] SB0.route_sel\[36\] net59 _0379_ _0372_ vssd1 vssd1 vccd1
+ vccd1 _0381_ sky130_fd_sc_hd__a41o_1
XANTENNA__2525__A1 _0982_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2525__B2 _0985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1763__X _0393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2234_ CB_1.config_dataA\[8\] _0856_ _0859_ _0862_ _1460_ vssd1 vssd1 vccd1 vccd1
+ _0863_ sky130_fd_sc_hd__o41a_1
X_3352_ clknet_leaf_25_clk _0172_ net266 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[44\]
+ sky130_fd_sc_hd__dfstp_1
X_3283_ clknet_leaf_24_clk _0103_ net272 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_2303_ _0930_ _0931_ CB_1.config_dataA\[17\] vssd1 vssd1 vccd1 vccd1 _0932_ sky130_fd_sc_hd__mux2_1
X_2096_ net143 net155 LEI0.config_data\[33\] vssd1 vssd1 vccd1 vccd1 _0726_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2165_ LE_1B.config_data\[13\] _0691_ _0723_ vssd1 vssd1 vccd1 vccd1 _0795_ sky130_fd_sc_hd__a21o_1
X_1949_ net37 _0577_ _0578_ vssd1 vssd1 vccd1 vccd1 _0579_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout230_A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2998_ SB0.route_sel\[38\] SB0.route_sel\[37\] net287 vssd1 vssd1 vccd1 vccd1 _0166_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1673__X _1511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2507__A1 _1134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_13_Right_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2783_ _1545_ _1368_ _1547_ vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__a21oi_2
XPHY_EDGE_ROW_22_Right_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2852_ LEI0.config_data\[20\] LEI0.config_data\[21\] net207 vssd1 vssd1 vccd1 vccd1
+ _0021_ sky130_fd_sc_hd__mux2_1
X_2921_ net436 net422 net204 vssd1 vssd1 vccd1 vccd1 _0090_ sky130_fd_sc_hd__mux2_1
XANTENNA__1797__A2 SB0.route_sel\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1803_ _0430_ _0431_ _0432_ vssd1 vssd1 vccd1 vccd1 _0433_ sky130_fd_sc_hd__a21bo_1
XANTENNA__1954__C1 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1734_ _1513_ _0363_ vssd1 vssd1 vccd1 vccd1 _0364_ sky130_fd_sc_hd__or2_1
X_3404_ clknet_leaf_27_clk _0224_ net271 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[96\]
+ sky130_fd_sc_hd__dfstp_1
X_1596_ SB0.route_sel\[25\] vssd1 vssd1 vccd1 vccd1 _1434_ sky130_fd_sc_hd__inv_2
X_1665_ net157 net169 net168 _1501_ _1502_ vssd1 vssd1 vccd1 vccd1 _1503_ sky130_fd_sc_hd__o32a_1
XANTENNA_fanout278_A net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2217_ net15 net16 net2 net3 net175 CB_1.config_dataA\[6\] vssd1 vssd1 vccd1 vccd1
+ _0846_ sky130_fd_sc_hd__mux4_1
XFILLER_38_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3197_ clknet_leaf_5_clk _0017_ net256 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_31_Right_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3335_ clknet_leaf_29_clk _0155_ net249 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[27\]
+ sky130_fd_sc_hd__dfstp_1
X_3266_ clknet_leaf_32_clk net387 net242 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_2148_ net194 _0776_ _0777_ vssd1 vssd1 vccd1 vccd1 _0778_ sky130_fd_sc_hd__a21oi_1
X_2079_ net15 net16 net2 net3 net199 CB_1.config_dataB\[6\] vssd1 vssd1 vccd1 vccd1
+ _0709_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_40_Right_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout233_X net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2370__C1 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3120_ net182 CB_0.config_dataB\[7\] net214 vssd1 vssd1 vccd1 vccd1 _0288_ sky130_fd_sc_hd__mux2_1
X_3051_ SB0.route_sel\[91\] SB0.route_sel\[90\] net294 vssd1 vssd1 vccd1 vccd1 _0219_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__2416__A0 net31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2002_ net144 _0630_ net234 vssd1 vssd1 vccd1 vccd1 _0632_ sky130_fd_sc_hd__o21ai_1
X_2766_ _1359_ vssd1 vssd1 vccd1 vccd1 _1360_ sky130_fd_sc_hd__inv_2
X_2835_ LEI0.config_data\[3\] net471 net212 vssd1 vssd1 vccd1 vccd1 _0004_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_0_clk_X clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2904_ net403 net394 net212 vssd1 vssd1 vccd1 vccd1 _0073_ sky130_fd_sc_hd__mux2_1
XANTENNA__2498__A3 net26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1579_ SB0.route_sel\[68\] vssd1 vssd1 vccd1 vccd1 _1417_ sky130_fd_sc_hd__inv_2
X_1648_ CB_1.config_dataB\[17\] vssd1 vssd1 vccd1 vccd1 _1486_ sky130_fd_sc_hd__inv_2
X_2697_ _1410_ SB0.route_sel\[72\] _1411_ SB0.route_sel\[75\] _1313_ vssd1 vssd1 vccd1
+ vccd1 _1314_ sky130_fd_sc_hd__a221o_1
X_3318_ clknet_leaf_24_clk _0138_ net267 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[10\]
+ sky130_fd_sc_hd__dfstp_1
X_1717_ CB_1.config_dataB\[21\] CB_1.config_dataB\[24\] CB_1.config_dataB\[20\] vssd1
+ vssd1 vccd1 vccd1 _1555_ sky130_fd_sc_hd__or3b_2
X_3249_ clknet_leaf_2_clk net432 net246 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_16_Left_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3080__A0 SB0.route_sel\[120\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1933__A2 _0562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1861__X _0491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2646__A0 net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2620_ LE_0A.config_data\[5\] _1180_ _1211_ _1246_ vssd1 vssd1 vccd1 vccd1 _1247_
+ sky130_fd_sc_hd__o211a_1
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2482_ CB_0.config_dataB\[18\] CB_0.config_dataB\[17\] CB_0.config_dataB\[19\] _1109_
+ vssd1 vssd1 vccd1 vccd1 _1110_ sky130_fd_sc_hd__or4bb_1
Xoutput128 net128 vssd1 vssd1 vccd1 vccd1 SBwest_out[2] sky130_fd_sc_hd__buf_4
X_2551_ net310 LEI0.config_data\[2\] _1177_ vssd1 vssd1 vccd1 vccd1 _1178_ sky130_fd_sc_hd__or3_1
Xoutput117 net117 vssd1 vssd1 vccd1 vccd1 SBsouth_out[7] sky130_fd_sc_hd__buf_8
Xoutput106 net106 vssd1 vssd1 vccd1 vccd1 SBsouth_out[11] sky130_fd_sc_hd__buf_8
X_3103_ CB_0.config_dataA\[14\] net187 net219 vssd1 vssd1 vccd1 vccd1 _0271_ sky130_fd_sc_hd__mux2_1
XANTENNA__1837__C_N _0460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3034_ SB0.route_sel\[74\] SB0.route_sel\[73\] net297 vssd1 vssd1 vccd1 vccd1 _0202_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__1688__A1 _1510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout143_A CB_0.le_outA vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout310_A net66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2749_ _1347_ _1348_ _0468_ vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__a21boi_4
X_2818_ net169 net166 _0371_ vssd1 vssd1 vccd1 vccd1 _1386_ sky130_fd_sc_hd__o21bai_4
Xfanout300 net301 vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__buf_2
XANTENNA__2340__A2 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_1_Left_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput19 CBnorth_in[11] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__buf_2
XFILLER_10_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2331__A2 _0439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2634__A3 _0994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1982_ _0611_ _0602_ net307 vssd1 vssd1 vccd1 vccd1 _0612_ sky130_fd_sc_hd__a21oi_4
X_2603_ CB_0.config_dataA\[13\] _1223_ _1226_ _1229_ vssd1 vssd1 vccd1 vccd1 _1230_
+ sky130_fd_sc_hd__or4_1
X_2534_ _0991_ _0994_ net193 vssd1 vssd1 vccd1 vccd1 _1161_ sky130_fd_sc_hd__mux2_1
XANTENNA__1766__X _0396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2465_ net317 _1071_ _1074_ net350 _1468_ vssd1 vssd1 vccd1 vccd1 _1093_ sky130_fd_sc_hd__a221o_1
X_2396_ CB_0.config_dataB\[3\] _1003_ _1007_ _1023_ CB_0.config_dataB\[4\] vssd1 vssd1
+ vccd1 vccd1 _1024_ sky130_fd_sc_hd__a41o_1
XANTENNA_clone61_A2 _0481_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout260_A net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3017_ SB0.route_sel\[57\] SB0.route_sel\[56\] net292 vssd1 vssd1 vccd1 vccd1 _0185_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__3453__SET_B net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2243__D1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout185 CB_0.config_dataB\[0\] vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__buf_2
Xfanout152 _1492_ vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__buf_8
Xfanout174 CB_1.config_dataA\[6\] vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__buf_2
Xfanout196 CB_1.config_dataB\[11\] vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout163 _0405_ vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__buf_2
XANTENNA_clone3_C1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2250_ net4 net6 net5 net7 net172 net173 vssd1 vssd1 vccd1 vccd1 _0879_ sky130_fd_sc_hd__mux4_1
X_2181_ net15 net16 net2 net3 net177 CB_1.config_dataA\[1\] vssd1 vssd1 vccd1 vccd1
+ _0810_ sky130_fd_sc_hd__mux4_1
X_1965_ net149 _1530_ _0593_ net236 vssd1 vssd1 vccd1 vccd1 _0595_ sky130_fd_sc_hd__o31a_1
XANTENNA__2240__A1 net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2517_ _1063_ _1142_ _1144_ _1098_ vssd1 vssd1 vccd1 vccd1 _1145_ sky130_fd_sc_hd__o211a_1
X_1896_ net149 _1502_ _0510_ net236 vssd1 vssd1 vccd1 vccd1 _0526_ sky130_fd_sc_hd__o31a_1
X_3497_ clknet_leaf_19_clk _0317_ net270 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[11\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_56_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2379_ _1006_ vssd1 vssd1 vccd1 vccd1 _1007_ sky130_fd_sc_hd__inv_2
X_2448_ net180 _1073_ _1075_ vssd1 vssd1 vccd1 vccd1 _1076_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_3_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout263_X net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2231__A1 _1552_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input36_A SBsouth_in[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2298__A1 _1552_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2222__A1 _0584_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_4_Left_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1750_ SB0.route_sel\[37\] SB0.route_sel\[36\] vssd1 vssd1 vccd1 vccd1 _0380_ sky130_fd_sc_hd__nand2_1
X_3420_ clknet_leaf_14_clk _0240_ net282 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[112\]
+ sky130_fd_sc_hd__dfstp_1
X_1681_ _1517_ _1518_ net29 vssd1 vssd1 vccd1 vccd1 _1519_ sky130_fd_sc_hd__o21ai_1
Xmax_cap138 _1010_ vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__clkbuf_2
XANTENNA__2222__B2 _0564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3351_ clknet_leaf_29_clk _0171_ net250 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[43\]
+ sky130_fd_sc_hd__dfstp_1
X_2233_ net174 _0860_ _0861_ vssd1 vssd1 vccd1 vccd1 _0862_ sky130_fd_sc_hd__a21oi_1
XANTENNA__2289__A1 net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2289__B2 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2164_ LE_1B.config_data\[12\] _0690_ vssd1 vssd1 vccd1 vccd1 _0794_ sky130_fd_sc_hd__and2_1
X_2302_ net11 net12 net13 net14 net171 net170 vssd1 vssd1 vccd1 vccd1 _0931_ sky130_fd_sc_hd__mux4_1
X_3282_ net68 _0102_ net70 vssd1 vssd1 vccd1 vccd1 LE_1B.dff_out sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_51_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2095_ LEI0.config_data\[34\] _0724_ vssd1 vssd1 vccd1 vccd1 _0725_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_0_138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1954__X _0584_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1948_ SB0.route_sel\[109\] SB0.route_sel\[108\] net53 _0576_ _0571_ vssd1 vssd1
+ vccd1 vccd1 _0578_ sky130_fd_sc_hd__a41o_1
X_1879_ net167 net162 net7 vssd1 vssd1 vccd1 vccd1 _0509_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout223_A net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2997_ SB0.route_sel\[37\] SB0.route_sel\[36\] net287 vssd1 vssd1 vccd1 vccd1 _0165_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2025__X _0655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_22_clk_A clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_30_Left_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2695__X net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1715__A0 _1526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input39_X net39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_2_3__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_2_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_50_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2920_ net391 LE_1A.config_data\[4\] net204 vssd1 vssd1 vccd1 vccd1 _0089_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkload1_A clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1733_ CB_0.config_dataA\[24\] CB_0.config_dataA\[21\] CB_0.config_dataA\[20\] vssd1
+ vssd1 vccd1 vccd1 _0363_ sky130_fd_sc_hd__or3b_1
X_2782_ _1492_ _0978_ _1542_ vssd1 vssd1 vccd1 vccd1 _1368_ sky130_fd_sc_hd__mux2_1
X_1802_ net148 _1530_ _0407_ net235 vssd1 vssd1 vccd1 vccd1 _0432_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_13_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2851_ LEI0.config_data\[19\] LEI0.config_data\[20\] net207 vssd1 vssd1 vccd1 vccd1
+ _0020_ sky130_fd_sc_hd__mux2_1
X_3403_ clknet_leaf_27_clk _0223_ net269 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[95\]
+ sky130_fd_sc_hd__dfstp_1
X_3334_ clknet_leaf_29_clk _0154_ net249 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[26\]
+ sky130_fd_sc_hd__dfstp_1
X_1664_ CB_1.config_dataA\[24\] CB_1.config_dataA\[20\] CB_1.config_dataA\[21\] vssd1
+ vssd1 vccd1 vccd1 _1502_ sky130_fd_sc_hd__or3b_4
X_1595_ SB0.route_sel\[36\] vssd1 vssd1 vccd1 vccd1 _1433_ sky130_fd_sc_hd__inv_2
XFILLER_53_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2216_ net174 _0841_ _0844_ vssd1 vssd1 vccd1 vccd1 _0845_ sky130_fd_sc_hd__a21oi_1
X_3196_ clknet_leaf_5_clk _0016_ net256 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_2147_ net16 _0760_ _0761_ net15 _1485_ vssd1 vssd1 vccd1 vccd1 _0777_ sky130_fd_sc_hd__a221o_1
X_3265_ clknet_leaf_0_clk _0085_ net243 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_41_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2078_ net4 net6 net5 net7 CB_1.config_dataB\[6\] net199 vssd1 vssd1 vccd1 vccd1
+ _0708_ sky130_fd_sc_hd__mux4_1
XANTENNA__3088__S net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1684__X _1522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2189__A0 _1526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1936__B1 net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2001_ _0628_ net151 _0629_ _0630_ vssd1 vssd1 vccd1 vccd1 _0631_ sky130_fd_sc_hd__o211a_1
XANTENNA__2113__A0 _1526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3050_ SB0.route_sel\[90\] SB0.route_sel\[89\] net295 vssd1 vssd1 vccd1 vccd1 _0218_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_61_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2903_ net439 net403 net212 vssd1 vssd1 vccd1 vccd1 _0072_ sky130_fd_sc_hd__mux2_1
X_2765_ CB_0.le_outB _1010_ _0499_ vssd1 vssd1 vccd1 vccd1 _1359_ sky130_fd_sc_hd__mux2_2
X_2834_ net469 LEI0.config_data\[3\] net212 vssd1 vssd1 vccd1 vccd1 _0003_ sky130_fd_sc_hd__mux2_1
X_2696_ SB0.route_sel\[79\] SB0.route_sel\[78\] vssd1 vssd1 vccd1 vccd1 _1313_ sky130_fd_sc_hd__nor2_1
X_1716_ SB0.route_sel\[42\] SB0.route_sel\[43\] vssd1 vssd1 vccd1 vccd1 _1554_ sky130_fd_sc_hd__nand2_1
X_1578_ SB0.route_sel\[66\] vssd1 vssd1 vccd1 vccd1 _1416_ sky130_fd_sc_hd__inv_2
X_1647_ CB_1.config_dataB\[18\] vssd1 vssd1 vccd1 vccd1 _1485_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout290_A net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3317_ clknet_leaf_24_clk _0137_ net267 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[9\]
+ sky130_fd_sc_hd__dfstp_2
XANTENNA__2655__A1 _1280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3248_ clknet_leaf_2_clk _0068_ net244 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_3179_ net429 LE_0B.config_data_in net206 vssd1 vssd1 vccd1 vccd1 _0347_ sky130_fd_sc_hd__mux2_1
XFILLER_41_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1918__B1 net20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2646__A1 net24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2343__A0 net27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2550_ LEI0.config_data\[0\] _1493_ _1176_ LEI0.config_data\[1\] vssd1 vssd1 vccd1
+ vccd1 _1177_ sky130_fd_sc_hd__o211a_1
Xoutput107 net107 vssd1 vssd1 vccd1 vccd1 SBsouth_out[12] sky130_fd_sc_hd__buf_6
XFILLER_9_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2481_ net178 CB_0.config_dataB\[15\] vssd1 vssd1 vccd1 vccd1 _1109_ sky130_fd_sc_hd__and2b_1
Xoutput129 net129 vssd1 vssd1 vccd1 vccd1 SBwest_out[3] sky130_fd_sc_hd__buf_8
Xoutput118 net118 vssd1 vssd1 vccd1 vccd1 SBsouth_out[8] sky130_fd_sc_hd__buf_8
XANTENNA__1688__A2 _1511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3102_ CB_0.config_dataA\[13\] CB_0.config_dataA\[14\] net220 vssd1 vssd1 vccd1 vccd1
+ _0270_ sky130_fd_sc_hd__mux2_1
XANTENNA__2637__B2 _1018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2637__A1 _1021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3033_ SB0.route_sel\[73\] SB0.route_sel\[72\] net297 vssd1 vssd1 vccd1 vccd1 _0201_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_46_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2573__A0 _0975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2679_ SB0.route_sel\[96\] _1398_ _1399_ SB0.route_sel\[99\] _1301_ vssd1 vssd1 vccd1
+ vccd1 _1302_ sky130_fd_sc_hd__a221o_1
X_2748_ _1447_ SB0.route_sel\[3\] _1448_ SB0.route_sel\[4\] vssd1 vssd1 vccd1 vccd1
+ _1348_ sky130_fd_sc_hd__o22a_1
X_2817_ _1503_ _1385_ _1505_ vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__a21boi_1
XANTENNA_fanout303_A net66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3476__SET_B net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2777__Y net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout301 net302 vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__clkbuf_2
XFILLER_27_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1856__Y _0486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input66_A config_en vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input21_X net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1981_ _0609_ _0610_ _0601_ vssd1 vssd1 vccd1 vccd1 _0611_ sky130_fd_sc_hd__or3b_4
X_2602_ net188 _1227_ _1228_ vssd1 vssd1 vccd1 vccd1 _1229_ sky130_fd_sc_hd__a21oi_1
X_2533_ CB_0.config_dataA\[3\] _1156_ _1159_ _1153_ vssd1 vssd1 vccd1 vccd1 _1160_
+ sky130_fd_sc_hd__and4bb_1
X_2464_ net181 net321 _1091_ net180 vssd1 vssd1 vccd1 vccd1 _1092_ sky130_fd_sc_hd__o211a_1
X_2395_ _1011_ _1015_ _1022_ vssd1 vssd1 vccd1 vccd1 _1023_ sky130_fd_sc_hd__a21o_1
XFILLER_28_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout253_A net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3016_ SB0.route_sel\[56\] SB0.route_sel\[55\] net294 vssd1 vssd1 vccd1 vccd1 _0184_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout306_X net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_31_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_2_1__f_clk_X clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout186 CB_0.config_dataA\[16\] vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__buf_2
Xfanout175 CB_1.config_dataA\[5\] vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__clkbuf_4
Xfanout153 _1492_ vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__buf_2
Xfanout197 CB_1.config_dataB\[10\] vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1809__C1 _0438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout142 net143 vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__buf_8
XFILLER_42_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_22_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_15_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2537__A0 net31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2698__X net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2180_ _0806_ net176 _0808_ vssd1 vssd1 vccd1 vccd1 _0809_ sky130_fd_sc_hd__a21oi_2
Xclkbuf_leaf_13_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1895_ net158 net168 _0508_ _0510_ _1502_ vssd1 vssd1 vccd1 vccd1 _0525_ sky130_fd_sc_hd__o32a_1
X_1964_ net158 net167 _0591_ _0593_ _1530_ vssd1 vssd1 vccd1 vccd1 _0594_ sky130_fd_sc_hd__o32a_1
XANTENNA__2528__A0 net27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2447_ net371 _1071_ _1074_ net319 CB_0.config_dataB\[12\] vssd1 vssd1 vccd1 vccd1
+ _1075_ sky130_fd_sc_hd__a221o_1
X_2516_ LE_0B.config_data\[9\] _1032_ _1064_ _1143_ vssd1 vssd1 vccd1 vccd1 _1144_
+ sky130_fd_sc_hd__a211o_1
X_3496_ clknet_leaf_20_clk _0316_ net279 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[10\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_56_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2378_ _1004_ _1005_ CB_0.config_dataB\[2\] vssd1 vssd1 vccd1 vccd1 _1006_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_3_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_19_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input29_A CBnorth_in[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1680_ CB_0.config_dataB\[20\] CB_0.config_dataB\[24\] CB_0.config_dataB\[21\] vssd1
+ vssd1 vccd1 vccd1 _1518_ sky130_fd_sc_hd__or3b_4
X_2301_ net1 net8 net9 net335 net171 net170 vssd1 vssd1 vccd1 vccd1 _0930_ sky130_fd_sc_hd__mux4_1
X_3350_ clknet_leaf_29_clk _0170_ net250 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[42\]
+ sky130_fd_sc_hd__dfstp_1
Xmax_cap139 _0910_ vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__clkbuf_1
X_2232_ _0371_ _0842_ _0843_ _0397_ _1459_ vssd1 vssd1 vccd1 vccd1 _0861_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_2_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_clk
+ sky130_fd_sc_hd__clkbuf_8
X_3281_ clknet_leaf_32_clk _0101_ net240 vssd1 vssd1 vccd1 vccd1 LEI0.config_data_in
+ sky130_fd_sc_hd__dfrtp_1
X_2163_ LE_1B.config_data\[14\] LE_1B.config_data\[15\] _0691_ vssd1 vssd1 vccd1 vccd1
+ _0793_ sky130_fd_sc_hd__mux2_1
XFILLER_61_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2094_ net147 net159 LEI0.config_data\[33\] vssd1 vssd1 vccd1 vccd1 _0724_ sky130_fd_sc_hd__mux2_1
XFILLER_21_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1947_ SB0.route_sel\[109\] SB0.route_sel\[108\] vssd1 vssd1 vccd1 vccd1 _0577_ sky130_fd_sc_hd__nand2_1
X_1878_ CB_1.config_dataB\[23\] CB_1.config_dataB\[22\] vssd1 vssd1 vccd1 vccd1 _0508_
+ sky130_fd_sc_hd__nand2_1
X_2996_ SB0.route_sel\[36\] SB0.route_sel\[35\] net287 vssd1 vssd1 vccd1 vccd1 _0164_
+ sky130_fd_sc_hd__mux2_1
X_3479_ clknet_leaf_13_clk _0299_ net277 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[18\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_8_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2204__A2 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output135_A net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2201__B net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clone9_C1 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2850_ LEI0.config_data\[18\] LEI0.config_data\[19\] net207 vssd1 vssd1 vccd1 vccd1
+ _0019_ sky130_fd_sc_hd__mux2_1
X_1732_ _1517_ _0360_ net28 vssd1 vssd1 vccd1 vccd1 _0362_ sky130_fd_sc_hd__o21ai_1
X_2781_ _1367_ _0662_ _0664_ vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__a21oi_4
X_1801_ net157 net167 net163 _0407_ _1530_ vssd1 vssd1 vccd1 vccd1 _0431_ sky130_fd_sc_hd__o32a_1
X_1663_ CB_1.config_dataA\[23\] CB_1.config_dataA\[22\] vssd1 vssd1 vccd1 vccd1 _1501_
+ sky130_fd_sc_hd__nand2b_2
XTAP_TAPCELL_ROW_13_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3402_ clknet_leaf_27_clk _0222_ net269 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[94\]
+ sky130_fd_sc_hd__dfstp_1
X_3333_ clknet_leaf_29_clk _0153_ net249 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[25\]
+ sky130_fd_sc_hd__dfstp_1
X_3264_ net68 _0084_ net70 vssd1 vssd1 vccd1 vccd1 LE_1A.dff_out sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_7_Right_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1594_ SB0.route_sel\[35\] vssd1 vssd1 vccd1 vccd1 _1432_ sky130_fd_sc_hd__inv_2
X_2215_ _0659_ _0842_ _0843_ _0679_ CB_1.config_dataA\[7\] vssd1 vssd1 vccd1 vccd1
+ _0844_ sky130_fd_sc_hd__a221o_1
X_2077_ _0705_ _0706_ vssd1 vssd1 vccd1 vccd1 _0707_ sky130_fd_sc_hd__or2_1
XFILLER_38_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3195_ clknet_leaf_5_clk _0015_ net256 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_2146_ net2 net3 net195 vssd1 vssd1 vccd1 vccd1 _0776_ sky130_fd_sc_hd__mux2_1
X_2979_ SB0.route_sel\[19\] SB0.route_sel\[18\] net286 vssd1 vssd1 vccd1 vccd1 _0147_
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout219_X net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2370__A1 _0655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2189__A1 _1552_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_33_Left_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3300__SET_B net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input51_X net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2000_ _1514_ _0607_ vssd1 vssd1 vccd1 vccd1 _0630_ sky130_fd_sc_hd__or2_1
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_61_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2833_ net475 net469 net213 vssd1 vssd1 vccd1 vccd1 _0002_ sky130_fd_sc_hd__mux2_1
XFILLER_43_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2902_ net396 LE_0B.config_data\[4\] net208 vssd1 vssd1 vccd1 vccd1 _0071_ sky130_fd_sc_hd__mux2_1
X_2764_ _1358_ _0540_ vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__and2_4
X_1646_ net197 vssd1 vssd1 vccd1 vccd1 _1484_ sky130_fd_sc_hd__inv_2
X_2695_ _1312_ _0656_ vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__and2_4
X_1715_ _1526_ net356 net201 vssd1 vssd1 vccd1 vccd1 _1553_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout283_A net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1577_ SB0.route_sel\[64\] vssd1 vssd1 vccd1 vccd1 _1415_ sky130_fd_sc_hd__inv_2
X_3247_ clknet_leaf_1_clk _0067_ net244 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_21_clk_A clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3316_ clknet_leaf_24_clk _0136_ net267 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[8\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_66_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2129_ net195 net354 _0758_ net194 vssd1 vssd1 vccd1 vccd1 _0759_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_24_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3178_ net379 LE_1B.config_data\[15\] net206 vssd1 vssd1 vccd1 vccd1 _0346_ sky130_fd_sc_hd__mux2_1
XANTENNA__1710__C_N _1538_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2343__A1 net28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2646__A2 net25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input11_A CBeast_in[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2031__B1 net31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2480_ net304 LEI0.config_data\[41\] _1107_ vssd1 vssd1 vccd1 vccd1 _1108_ sky130_fd_sc_hd__nor3b_1
Xoutput119 net119 vssd1 vssd1 vccd1 vccd1 SBsouth_out[9] sky130_fd_sc_hd__buf_8
Xoutput108 net108 vssd1 vssd1 vccd1 vccd1 SBsouth_out[13] sky130_fd_sc_hd__buf_8
Xoutput90 net90 vssd1 vssd1 vccd1 vccd1 CBnorth_out[11] sky130_fd_sc_hd__buf_6
X_3101_ CB_0.config_dataA\[12\] CB_0.config_dataA\[13\] net220 vssd1 vssd1 vccd1 vccd1
+ _0269_ sky130_fd_sc_hd__mux2_1
X_3032_ SB0.route_sel\[72\] SB0.route_sel\[71\] net297 vssd1 vssd1 vccd1 vccd1 _0200_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_38_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2816_ _1498_ net168 _1526_ vssd1 vssd1 vccd1 vccd1 _1385_ sky130_fd_sc_hd__o21bai_1
Xfanout302 net67 vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__clkbuf_4
XANTENNA__2573__A1 _0978_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1629_ CB_0.config_dataB\[9\] vssd1 vssd1 vccd1 vccd1 _1467_ sky130_fd_sc_hd__inv_2
X_2678_ SB0.route_sel\[102\] SB0.route_sel\[103\] vssd1 vssd1 vccd1 vccd1 _1301_ sky130_fd_sc_hd__nor2_1
XANTENNA__3509__SET_B net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2747_ SB0.route_sel\[1\] SB0.route_sel\[0\] vssd1 vssd1 vccd1 vccd1 _1347_ sky130_fd_sc_hd__or2_1
XANTENNA_input3_A CBeast_in[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2564__A1 _1018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2564__B2 _1021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input59_A SBwest_in[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input14_X net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1980_ net144 _0608_ net237 vssd1 vssd1 vccd1 vccd1 _0610_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_43_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2601_ _0985_ _1220_ _1221_ _0982_ _1474_ vssd1 vssd1 vccd1 vccd1 _1228_ sky130_fd_sc_hd__a221o_1
X_2532_ net192 _1157_ _1158_ vssd1 vssd1 vccd1 vccd1 _1159_ sky130_fd_sc_hd__a21o_1
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2463_ net181 _1010_ vssd1 vssd1 vccd1 vccd1 _1091_ sky130_fd_sc_hd__nand2_1
XANTENNA__2004__B1 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2394_ _0952_ net317 net350 _0967_ _1465_ vssd1 vssd1 vccd1 vccd1 _1022_ sky130_fd_sc_hd__a221o_1
X_3015_ SB0.route_sel\[55\] SB0.route_sel\[54\] net294 vssd1 vssd1 vccd1 vccd1 _0183_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__2491__A0 net20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout246_A net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2794__A1 _0963_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input6_X net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout165 _0373_ vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__buf_2
XANTENNA__1754__C1 _0383_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout143 CB_0.le_outA vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__buf_8
Xfanout187 CB_0.config_dataA\[15\] vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__buf_2
Xfanout176 CB_1.config_dataA\[1\] vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__buf_2
Xfanout198 CB_1.config_dataB\[6\] vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__buf_2
XANTENNA__2309__X _0938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clone3_A1 _0675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2225__A0 _0428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2528__A1 net28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2776__A1 _0991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1894_ net168 net162 net6 vssd1 vssd1 vccd1 vccd1 _0524_ sky130_fd_sc_hd__o21ai_1
X_1963_ CB_1.config_dataA\[22\] CB_1.config_dataA\[23\] vssd1 vssd1 vccd1 vccd1 _0593_
+ sky130_fd_sc_hd__nand2b_2
X_3495_ clknet_leaf_18_clk _0315_ net279 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[9\]
+ sky130_fd_sc_hd__dfstp_1
X_2446_ net181 net180 vssd1 vssd1 vccd1 vccd1 _1074_ sky130_fd_sc_hd__nor2_1
X_2515_ _1025_ _1026_ _1031_ LE_0B.config_data\[8\] vssd1 vssd1 vccd1 vccd1 _1143_
+ sky130_fd_sc_hd__o211a_1
X_2377_ net20 net22 net21 net23 CB_0.config_dataB\[1\] net185 vssd1 vssd1 vccd1 vccd1
+ _1005_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_54_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1806__A3 net58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2231_ _1526_ _1552_ net175 vssd1 vssd1 vccd1 vccd1 _0860_ sky130_fd_sc_hd__mux2_1
X_3280_ clknet_leaf_32_clk _0100_ net240 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_2300_ net170 _0927_ _0928_ vssd1 vssd1 vccd1 vccd1 _0929_ sky130_fd_sc_hd__a21o_1
X_2162_ _0723_ _0789_ _0790_ _0791_ _0755_ vssd1 vssd1 vccd1 vccd1 _0792_ sky130_fd_sc_hd__a221o_1
X_2093_ LEI0.config_data\[23\] net232 _0716_ _0721_ vssd1 vssd1 vccd1 vccd1 _0723_
+ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_51_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2995_ SB0.route_sel\[35\] SB0.route_sel\[34\] net289 vssd1 vssd1 vccd1 vccd1 _0163_
+ sky130_fd_sc_hd__mux2_1
X_1946_ SB0.route_sel\[110\] SB0.route_sel\[111\] vssd1 vssd1 vccd1 vccd1 _0576_ sky130_fd_sc_hd__nand2_1
X_1877_ SB0.route_sel\[122\] SB0.route_sel\[123\] vssd1 vssd1 vccd1 vccd1 _0507_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout209_A net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3478_ clknet_leaf_13_clk _0298_ net277 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[17\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__2382__C1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2429_ net328 net347 CB_0.config_dataB\[5\] vssd1 vssd1 vccd1 vccd1 _1057_ sky130_fd_sc_hd__mux2_1
XFILLER_44_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold156_A LE_1B.config_data\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2373__C1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input41_A SBsouth_in[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output128_A net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clone9_B1 _0965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1800_ net167 net163 net335 vssd1 vssd1 vccd1 vccd1 _0430_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_13_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2600__A0 _0975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1731_ _1516_ _0359_ vssd1 vssd1 vccd1 vccd1 _0361_ sky130_fd_sc_hd__nand2_1
XANTENNA__1954__A2 _0570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2780_ net329 _1001_ _0660_ vssd1 vssd1 vccd1 vccd1 _1367_ sky130_fd_sc_hd__mux2_4
X_1662_ _1498_ net168 net13 vssd1 vssd1 vccd1 vccd1 _1500_ sky130_fd_sc_hd__o21ai_1
X_3401_ clknet_leaf_27_clk _0221_ net269 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[93\]
+ sky130_fd_sc_hd__dfstp_1
X_3194_ clknet_leaf_7_clk _0014_ net256 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_2214_ net175 net174 vssd1 vssd1 vccd1 vccd1 _0843_ sky130_fd_sc_hd__nor2_1
X_3263_ clknet_leaf_1_clk _0083_ net246 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_3332_ clknet_leaf_29_clk _0152_ net249 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[24\]
+ sky130_fd_sc_hd__dfstp_1
X_1593_ SB0.route_sel\[34\] vssd1 vssd1 vccd1 vccd1 _1431_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2076_ net349 _0692_ _0694_ net352 _1479_ vssd1 vssd1 vccd1 vccd1 _0706_ sky130_fd_sc_hd__a221o_1
X_2145_ net348 net362 net312 _0615_ net195 net194 vssd1 vssd1 vccd1 vccd1 _0775_ sky130_fd_sc_hd__mux4_1
X_1929_ SB0.route_sel\[101\] SB0.route_sel\[100\] net36 vssd1 vssd1 vccd1 vccd1 _0559_
+ sky130_fd_sc_hd__a21boi_1
X_2978_ SB0.route_sel\[18\] SB0.route_sel\[17\] net287 vssd1 vssd1 vccd1 vccd1 _0146_
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2370__A2 _0649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold90 LE_0B.config_data\[9\] vssd1 vssd1 vccd1 vccd1 net400 sky130_fd_sc_hd__dlygate4sd3_1
X_2763_ SB0.route_sel\[112\] _1451_ _1454_ SB0.route_sel\[115\] _1357_ vssd1 vssd1
+ vccd1 vccd1 _1358_ sky130_fd_sc_hd__a221o_1
XANTENNA__2416__A3 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2832_ LEI0.config_data\[0\] net475 net213 vssd1 vssd1 vccd1 vccd1 _0001_ sky130_fd_sc_hd__mux2_1
XFILLER_31_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2901_ net447 net396 net207 vssd1 vssd1 vccd1 vccd1 _0070_ sky130_fd_sc_hd__mux2_1
XANTENNA__1785__Y _0415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1645_ CB_1.config_dataB\[12\] vssd1 vssd1 vccd1 vccd1 _1483_ sky130_fd_sc_hd__inv_2
X_1576_ SB0.route_sel\[65\] vssd1 vssd1 vccd1 vccd1 _1414_ sky130_fd_sc_hd__inv_2
X_2694_ SB0.route_sel\[74\] _1412_ SB0.route_sel\[77\] _1413_ _1311_ vssd1 vssd1 vccd1
+ vccd1 _1312_ sky130_fd_sc_hd__a221o_1
XANTENNA__2808__B1_N _0637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1714_ _1548_ _1539_ _1551_ net306 vssd1 vssd1 vccd1 vccd1 _1552_ sky130_fd_sc_hd__a211o_4
XANTENNA_fanout276_A net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3246_ net68 _0066_ net70 vssd1 vssd1 vccd1 vccd1 LE_0B.dff_out sky130_fd_sc_hd__dfrtp_1
X_3315_ clknet_leaf_25_clk _0135_ net267 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[7\]
+ sky130_fd_sc_hd__dfstp_1
X_3177_ net388 net379 net203 vssd1 vssd1 vccd1 vccd1 _0345_ sky130_fd_sc_hd__mux2_1
X_2128_ net195 _0521_ vssd1 vssd1 vccd1 vccd1 _0758_ sky130_fd_sc_hd__nand2_1
XFILLER_34_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2059_ LEI0.config_data\[10\] _0685_ _0688_ vssd1 vssd1 vccd1 vccd1 _0689_ sky130_fd_sc_hd__o21ba_1
XANTENNA_fanout231_X net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2343__A2 net29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2328__C1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2646__A3 net26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput109 net109 vssd1 vssd1 vccd1 vccd1 SBsouth_out[14] sky130_fd_sc_hd__buf_6
Xoutput91 net91 vssd1 vssd1 vccd1 vccd1 CBnorth_out[12] sky130_fd_sc_hd__buf_6
X_3100_ net188 CB_0.config_dataA\[12\] net217 vssd1 vssd1 vccd1 vccd1 _0268_ sky130_fd_sc_hd__mux2_1
X_3031_ SB0.route_sel\[71\] SB0.route_sel\[70\] net297 vssd1 vssd1 vccd1 vccd1 _0199_
+ sky130_fd_sc_hd__mux2_1
Xoutput80 net80 vssd1 vssd1 vccd1 vccd1 CBeast_out[2] sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_38_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2746_ _0488_ _1346_ vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__and2_4
XFILLER_8_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2815_ _1384_ _1531_ _1532_ vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__a21boi_2
X_1559_ SB0.route_sel\[108\] vssd1 vssd1 vccd1 vccd1 _1397_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_52_Left_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1628_ CB_0.config_dataB\[7\] vssd1 vssd1 vccd1 vccd1 _1466_ sky130_fd_sc_hd__inv_2
X_2677_ _1300_ _0563_ vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__and2b_1
Xfanout303 net66 vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__buf_2
X_3229_ clknet_leaf_8_clk _0049_ net258 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_61_Left_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout279_X net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2261__A1 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1772__A0 net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2330__X _0958_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output110_A net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2600_ _0975_ _0978_ net189 vssd1 vssd1 vccd1 vccd1 _1227_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_43_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2004__A1 _0633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_20_clk_A clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2531_ _0963_ _1148_ _1151_ _0966_ CB_0.config_dataA\[2\] vssd1 vssd1 vccd1 vccd1
+ _1158_ sky130_fd_sc_hd__a221o_1
X_2462_ _1089_ vssd1 vssd1 vccd1 vccd1 _1090_ sky130_fd_sc_hd__inv_2
X_2393_ _0562_ _0552_ _1020_ net309 vssd1 vssd1 vccd1 vccd1 _1021_ sky130_fd_sc_hd__a211o_4
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3014_ SB0.route_sel\[54\] SB0.route_sel\[53\] net294 vssd1 vssd1 vccd1 vccd1 _0182_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__2491__A1 net22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2729_ SB0.route_sel\[26\] _1436_ SB0.route_sel\[29\] _1437_ vssd1 vssd1 vccd1 vccd1
+ _1335_ sky130_fd_sc_hd__a22o_1
Xfanout188 CB_0.config_dataA\[11\] vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__buf_2
Xfanout177 CB_1.config_dataA\[0\] vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__clkbuf_4
Xfanout144 CB_0.le_outA vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__clkbuf_4
Xfanout199 CB_1.config_dataB\[5\] vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__clkbuf_4
Xfanout166 _1555_ vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__buf_2
Xfanout155 CB_0.le_outB vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_29_Right_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_38_Right_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input71_A nrst vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clone3_A2 _0665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2220__B _0521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_47_Right_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_56_Right_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2225__A1 _0449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_90 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1962_ net167 net161 net3 vssd1 vssd1 vccd1 vccd1 _0592_ sky130_fd_sc_hd__o21ai_1
X_1893_ SB0.route_sel\[114\] SB0.route_sel\[115\] vssd1 vssd1 vccd1 vccd1 _0523_ sky130_fd_sc_hd__nand2_1
XANTENNA__2528__A2 net29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_65_Right_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2376_ net31 net32 net18 net19 net185 net184 vssd1 vssd1 vccd1 vccd1 _1004_ sky130_fd_sc_hd__mux4_1
X_3494_ clknet_leaf_18_clk _0314_ net279 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[8\]
+ sky130_fd_sc_hd__dfstp_1
X_2445_ _0956_ net339 CB_0.config_dataB\[10\] vssd1 vssd1 vccd1 vccd1 _1073_ sky130_fd_sc_hd__mux2_1
X_2514_ LE_0B.config_data\[10\] LE_0B.config_data\[11\] _1032_ vssd1 vssd1 vccd1 vccd1
+ _1142_ sky130_fd_sc_hd__mux2_1
XANTENNA__1751__A3 net59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclone7 net318 _0570_ _1017_ net310 vssd1 vssd1 vccd1 vccd1 net317 sky130_fd_sc_hd__a211o_1
XFILLER_47_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1718__B1 net12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2230_ _0857_ _0858_ _1459_ vssd1 vssd1 vccd1 vccd1 _0859_ sky130_fd_sc_hd__mux2_1
X_2161_ LE_1B.config_data\[1\] _0691_ _0723_ vssd1 vssd1 vccd1 vccd1 _0791_ sky130_fd_sc_hd__a21oi_1
XANTENNA_clkbuf_2_2__f_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2092_ LEI0.config_data\[23\] net232 _0716_ _0721_ vssd1 vssd1 vccd1 vccd1 _0722_
+ sky130_fd_sc_hd__a31oi_2
X_1945_ _0572_ _0573_ _0574_ vssd1 vssd1 vccd1 vccd1 _0575_ sky130_fd_sc_hd__a21bo_1
XANTENNA__1957__A0 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2994_ SB0.route_sel\[34\] SB0.route_sel\[33\] net289 vssd1 vssd1 vccd1 vccd1 _0162_
+ sky130_fd_sc_hd__mux2_1
X_1876_ _0503_ _0504_ _0505_ vssd1 vssd1 vccd1 vccd1 _0506_ sky130_fd_sc_hd__or3b_4
XTAP_TAPCELL_ROW_8_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3477_ clknet_leaf_13_clk _0297_ net277 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[16\]
+ sky130_fd_sc_hd__dfstp_1
X_2359_ net184 _0979_ _0986_ vssd1 vssd1 vccd1 vccd1 _0987_ sky130_fd_sc_hd__a21o_1
X_2428_ _1054_ _1055_ CB_0.config_dataB\[7\] vssd1 vssd1 vccd1 vccd1 _1056_ sky130_fd_sc_hd__mux2_1
XANTENNA__1890__A net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_8_Left_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clone9_A1 _0467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input34_A SBsouth_in[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1939__B1 net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1730_ CB_0.config_dataB\[21\] CB_0.config_dataB\[24\] CB_0.config_dataB\[20\] vssd1
+ vssd1 vccd1 vccd1 _0360_ sky130_fd_sc_hd__or3b_2
XANTENNA__2600__A1 _0978_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3400_ clknet_leaf_26_clk _0220_ net269 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[92\]
+ sky130_fd_sc_hd__dfstp_1
X_1661_ CB_1.config_dataB\[20\] CB_1.config_dataB\[24\] CB_1.config_dataB\[21\] vssd1
+ vssd1 vccd1 vccd1 _1499_ sky130_fd_sc_hd__or3b_2
X_3331_ clknet_leaf_29_clk _0151_ net248 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[23\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_7_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1592_ SB0.route_sel\[33\] vssd1 vssd1 vccd1 vccd1 _1430_ sky130_fd_sc_hd__inv_2
XFILLER_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2213_ net174 CB_1.config_dataA\[5\] vssd1 vssd1 vccd1 vccd1 _0842_ sky130_fd_sc_hd__and2b_1
X_3193_ clknet_leaf_6_clk _0013_ net255 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_2144_ net194 _0772_ _0773_ vssd1 vssd1 vccd1 vccd1 _0774_ sky130_fd_sc_hd__a21oi_1
X_3262_ clknet_leaf_1_clk _0082_ net246 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_64_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2075_ net199 net354 _0704_ net198 vssd1 vssd1 vccd1 vccd1 _0705_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout221_A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1928_ SB0.route_sel\[102\] SB0.route_sel\[103\] vssd1 vssd1 vccd1 vccd1 _0558_ sky130_fd_sc_hd__nand2_1
XFILLER_30_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1859_ SB0.route_sel\[15\] SB0.route_sel\[14\] vssd1 vssd1 vccd1 vccd1 _0489_ sky130_fd_sc_hd__nand2b_1
X_2977_ SB0.route_sel\[17\] SB0.route_sel\[16\] net287 vssd1 vssd1 vccd1 vccd1 _0145_
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1891__Y _0521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2649__B2 _0982_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2649__A1 _0985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input37_X net37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold91 LE_0A.config_data\[8\] vssd1 vssd1 vccd1 vccd1 net401 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_35_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2900_ net431 LE_0B.config_data\[2\] net208 vssd1 vssd1 vccd1 vccd1 _0069_ sky130_fd_sc_hd__mux2_1
Xhold80 _0078_ vssd1 vssd1 vccd1 vccd1 net390 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1857__C1 _0486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2762_ SB0.route_sel\[118\] SB0.route_sel\[119\] vssd1 vssd1 vccd1 vccd1 _1357_ sky130_fd_sc_hd__nor2_1
XFILLER_31_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2831_ net489 LEI0.config_data\[0\] net202 vssd1 vssd1 vccd1 vccd1 _0000_ sky130_fd_sc_hd__mux2_1
X_1713_ _1418_ SB0.route_sel\[56\] SB0.route_sel\[61\] SB0.route_sel\[60\] _1550_
+ vssd1 vssd1 vccd1 vccd1 _1551_ sky130_fd_sc_hd__o221a_1
XANTENNA__3465__SET_B net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2693_ SB0.route_sel\[73\] SB0.route_sel\[72\] vssd1 vssd1 vccd1 vccd1 _1311_ sky130_fd_sc_hd__nor2_1
X_1575_ SB0.route_sel\[76\] vssd1 vssd1 vccd1 vccd1 _1413_ sky130_fd_sc_hd__inv_2
X_1644_ LE_1B.config_data\[3\] vssd1 vssd1 vccd1 vccd1 _1482_ sky130_fd_sc_hd__inv_2
X_3314_ clknet_leaf_24_clk _0134_ net267 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[6\]
+ sky130_fd_sc_hd__dfstp_1
Xrebuffer12 net323 vssd1 vssd1 vccd1 vccd1 net322 sky130_fd_sc_hd__clkbuf_2
X_3245_ clknet_leaf_6_clk _0065_ net254 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_3176_ net427 net388 net203 vssd1 vssd1 vccd1 vccd1 _0344_ sky130_fd_sc_hd__mux2_1
X_2127_ net303 CB_0.config_data_inA _0756_ vssd1 vssd1 vccd1 vccd1 _0757_ sky130_fd_sc_hd__nor3b_1
XTAP_TAPCELL_ROW_24_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2058_ net303 LEI0.config_data\[11\] _0687_ vssd1 vssd1 vccd1 vccd1 _0688_ sky130_fd_sc_hd__or3_1
XANTENNA__2576__A0 net27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2153__X _0783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout224_X net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2343__A3 net30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2328__X _0956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2567__A0 net31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput92 net92 vssd1 vssd1 vccd1 vccd1 CBnorth_out[13] sky130_fd_sc_hd__buf_6
X_3030_ SB0.route_sel\[70\] SB0.route_sel\[69\] net297 vssd1 vssd1 vccd1 vccd1 _0198_
+ sky130_fd_sc_hd__mux2_1
Xoutput81 net81 vssd1 vssd1 vccd1 vccd1 CBeast_out[3] sky130_fd_sc_hd__buf_6
XANTENNA_clkbuf_leaf_9_clk_A clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2270__A2 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2701__X net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2676_ SB0.route_sel\[96\] SB0.route_sel\[97\] _1399_ SB0.route_sel\[99\] _1299_
+ vssd1 vssd1 vccd1 vccd1 _1300_ sky130_fd_sc_hd__o221a_1
XANTENNA__2007__C1 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2745_ _1442_ SB0.route_sel\[8\] _1443_ SB0.route_sel\[11\] _1345_ vssd1 vssd1 vccd1
+ vccd1 _1346_ sky130_fd_sc_hd__a221o_1
X_2814_ net169 net167 _1552_ vssd1 vssd1 vccd1 vccd1 _1384_ sky130_fd_sc_hd__o21bai_4
X_1558_ SB0.route_sel\[106\] vssd1 vssd1 vccd1 vccd1 _1396_ sky130_fd_sc_hd__inv_2
X_1627_ CB_0.config_dataB\[2\] vssd1 vssd1 vccd1 vccd1 _1465_ sky130_fd_sc_hd__inv_2
Xfanout304 net66 vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__clkbuf_2
XANTENNA__2089__A2 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3228_ net68 _0048_ net70 vssd1 vssd1 vccd1 vccd1 LE_0A.dff_out sky130_fd_sc_hd__dfrtp_1
X_3159_ CB_1.config_dataA\[20\] CB_1.config_dataA\[21\] net223 vssd1 vssd1 vccd1 vccd1
+ _0327_ sky130_fd_sc_hd__mux2_1
XFILLER_52_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2261__A2 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1772__A1 net12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output103_A net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_25_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__1897__X _0527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2530_ _0956_ _0959_ net193 vssd1 vssd1 vccd1 vccd1 _1157_ sky130_fd_sc_hd__mux2_1
XANTENNA__2004__A2 _0627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_21_Left_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2461_ _1087_ _1088_ _1468_ vssd1 vssd1 vccd1 vccd1 _1089_ sky130_fd_sc_hd__mux2_1
X_2392_ SB0.route_sel\[98\] SB0.route_sel\[99\] SB0.route_sel\[101\] _1400_ _1019_
+ vssd1 vssd1 vccd1 vccd1 _1020_ sky130_fd_sc_hd__o221a_1
XANTENNA__2491__A2 net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2128__B _0521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3013_ SB0.route_sel\[53\] SB0.route_sel\[52\] net294 vssd1 vssd1 vccd1 vccd1 _0181_
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_16_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_51_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2659_ _1173_ _1174_ _1179_ LE_0A.config_data\[12\] vssd1 vssd1 vccd1 vccd1 _1286_
+ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout301_A net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2728_ _0394_ _1334_ vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__and2_4
Xfanout178 CB_0.config_dataB\[16\] vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__buf_2
Xfanout189 CB_0.config_dataA\[10\] vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__buf_2
Xfanout145 CB_0.le_outA vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__clkbuf_2
Xfanout156 CB_0.le_outB vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout167 _1528_ vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_57_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1809__A2 _0433_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2537__A3 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input64_A SBwest_in[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1681__B1 net29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1892_ _0506_ _0518_ _0520_ _1478_ vssd1 vssd1 vccd1 vccd1 _0522_ sky130_fd_sc_hd__a211o_1
X_1961_ CB_1.config_dataB\[22\] CB_1.config_dataB\[23\] vssd1 vssd1 vccd1 vccd1 _0591_
+ sky130_fd_sc_hd__nand2b_1
XANTENNA__2528__A3 net30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3493_ clknet_leaf_14_clk _0313_ net282 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[7\]
+ sky130_fd_sc_hd__dfstp_1
X_2513_ _1063_ _1138_ _1140_ _1099_ vssd1 vssd1 vccd1 vccd1 _1141_ sky130_fd_sc_hd__o211a_1
X_2444_ CB_0.config_dataB\[13\] _1468_ CB_0.config_dataB\[14\] _1071_ vssd1 vssd1
+ vccd1 vccd1 _1072_ sky130_fd_sc_hd__and4b_1
X_2375_ net184 _0995_ _1002_ vssd1 vssd1 vccd1 vccd1 _1003_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_5_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_2_161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2207__A2 _0829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2143__A1 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2160_ LE_1B.config_data\[0\] _0690_ vssd1 vssd1 vccd1 vccd1 _0790_ sky130_fd_sc_hd__nand2_1
X_2091_ LEI0.config_data\[22\] _0717_ _0720_ vssd1 vssd1 vccd1 vccd1 _0721_ sky130_fd_sc_hd__o21ba_1
X_1875_ SB0.route_sel\[120\] SB0.route_sel\[121\] vssd1 vssd1 vccd1 vccd1 _0505_ sky130_fd_sc_hd__nand2_1
X_1944_ net149 _0349_ _0510_ net236 vssd1 vssd1 vccd1 vccd1 _0574_ sky130_fd_sc_hd__o31a_1
XANTENNA__1957__A1 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2993_ SB0.route_sel\[33\] SB0.route_sel\[32\] net289 vssd1 vssd1 vccd1 vccd1 _0161_
+ sky130_fd_sc_hd__mux2_1
X_3476_ clknet_leaf_10_clk _0296_ net264 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[15\]
+ sky130_fd_sc_hd__dfstp_1
X_2427_ net27 net28 net29 net30 net183 net182 vssd1 vssd1 vccd1 vccd1 _1055_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_24_Left_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2358_ _0952_ net343 net342 _0967_ _1465_ vssd1 vssd1 vccd1 vccd1 _0986_ sky130_fd_sc_hd__a221o_1
X_2289_ net5 _0911_ _0914_ net4 _1464_ vssd1 vssd1 vccd1 vccd1 _0918_ sky130_fd_sc_hd__a221o_1
XANTENNA__2134__B2 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2134__A1 net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2373__A1 _0675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input27_A CBnorth_in[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3102__S net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clone9_A2 _0461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2941__S net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3330_ clknet_leaf_30_clk _0150_ net247 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[22\]
+ sky130_fd_sc_hd__dfstp_1
X_1591_ SB0.route_sel\[44\] vssd1 vssd1 vccd1 vccd1 _1429_ sky130_fd_sc_hd__inv_2
X_1660_ CB_1.config_dataB\[23\] CB_1.config_dataB\[22\] vssd1 vssd1 vccd1 vccd1 _1498_
+ sky130_fd_sc_hd__nand2b_1
XANTENNA__2116__A1 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2212_ _0637_ _0615_ net175 vssd1 vssd1 vccd1 vccd1 _0841_ sky130_fd_sc_hd__mux2_1
X_3192_ clknet_leaf_5_clk _0012_ net254 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_2143_ net8 _0760_ _0761_ net1 CB_1.config_dataB\[18\] vssd1 vssd1 vccd1 vccd1 _0773_
+ sky130_fd_sc_hd__a221o_1
X_3261_ clknet_leaf_2_clk net426 net246 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_64_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2704__X net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2074_ _0506_ _0518_ _0520_ _1480_ vssd1 vssd1 vccd1 vccd1 _0704_ sky130_fd_sc_hd__a211o_1
X_1927_ _0554_ _0555_ _0556_ vssd1 vssd1 vccd1 vccd1 _0557_ sky130_fd_sc_hd__a21bo_1
X_2976_ SB0.route_sel\[16\] SB0.route_sel\[15\] net291 vssd1 vssd1 vccd1 vccd1 _0144_
+ sky130_fd_sc_hd__mux2_1
X_1858_ _0481_ _0487_ net306 vssd1 vssd1 vccd1 vccd1 _0488_ sky130_fd_sc_hd__a21oi_2
X_3459_ clknet_leaf_14_clk _0279_ net278 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[23\]
+ sky130_fd_sc_hd__dfstp_1
X_1789_ _1518_ _0417_ net25 vssd1 vssd1 vccd1 vccd1 _0419_ sky130_fd_sc_hd__o21ai_1
XFILLER_29_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2291__A0 _0637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold92 _0058_ vssd1 vssd1 vccd1 vccd1 net402 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_output133_A net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold81 LE_1A.config_data\[3\] vssd1 vssd1 vccd1 vccd1 net391 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1857__B1 _0485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold70 _0346_ vssd1 vssd1 vccd1 vccd1 net380 sky130_fd_sc_hd__dlygate4sd3_1
X_2830_ net302 net310 vssd1 vssd1 vccd1 vccd1 _1392_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_61_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_1 CBnorth_in[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2761_ _1355_ _1356_ _0540_ vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__a21boi_4
X_2692_ _0634_ _1310_ vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__and2_4
X_1643_ LE_1B.config_data\[2\] vssd1 vssd1 vccd1 vccd1 _1481_ sky130_fd_sc_hd__inv_2
X_1712_ SB0.route_sel\[63\] SB0.route_sel\[62\] vssd1 vssd1 vccd1 vccd1 _1550_ sky130_fd_sc_hd__nand2b_1
X_3244_ clknet_leaf_6_clk net409 net255 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_1574_ SB0.route_sel\[75\] vssd1 vssd1 vccd1 vccd1 _1412_ sky130_fd_sc_hd__inv_2
X_3313_ clknet_leaf_24_clk _0133_ net272 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[5\]
+ sky130_fd_sc_hd__dfstp_1
Xrebuffer13 net324 vssd1 vssd1 vccd1 vccd1 net323 sky130_fd_sc_hd__clkbuf_2
X_3175_ LE_1B.config_data\[11\] net427 net203 vssd1 vssd1 vccd1 vccd1 _0343_ sky130_fd_sc_hd__mux2_1
X_2057_ LEI0.config_data\[9\] net147 _0686_ LEI0.config_data\[10\] vssd1 vssd1 vccd1
+ vccd1 _0687_ sky130_fd_sc_hd__o211a_1
X_2126_ net326 net155 net150 net160 LEI0.config_data\[45\] LEI0.config_data\[46\]
+ vssd1 vssd1 vccd1 vccd1 _0756_ sky130_fd_sc_hd__mux4_1
XFILLER_41_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2959_ CB_1.config_dataB\[23\] CB_1.config_dataB\[24\] net222 vssd1 vssd1 vccd1 vccd1
+ _0127_ sky130_fd_sc_hd__mux2_1
XANTENNA__2576__A1 net28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2328__A1 _0424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2264__A0 _1526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput93 net93 vssd1 vssd1 vccd1 vccd1 CBnorth_out[14] sky130_fd_sc_hd__buf_6
Xoutput82 net82 vssd1 vssd1 vccd1 vccd1 CBeast_out[4] sky130_fd_sc_hd__buf_6
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2813_ _1383_ _0668_ _0669_ vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__a21boi_2
XANTENNA__2270__A3 _0897_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2675_ SB0.route_sel\[101\] _1400_ vssd1 vssd1 vccd1 vccd1 _1299_ sky130_fd_sc_hd__nand2_1
X_2744_ SB0.route_sel\[15\] SB0.route_sel\[14\] vssd1 vssd1 vccd1 vccd1 _1345_ sky130_fd_sc_hd__nor2_1
X_1626_ CB_1.config_dataA\[17\] vssd1 vssd1 vccd1 vccd1 _1464_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout281_A net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1557_ SB0.route_sel\[105\] vssd1 vssd1 vccd1 vccd1 _1395_ sky130_fd_sc_hd__inv_2
Xfanout305 net308 vssd1 vssd1 vccd1 vccd1 net305 sky130_fd_sc_hd__clkbuf_4
X_3227_ clknet_leaf_28_clk _0047_ net251 vssd1 vssd1 vccd1 vccd1 CB_0.config_data_inA
+ sky130_fd_sc_hd__dfrtp_2
X_3089_ net193 net192 net217 vssd1 vssd1 vccd1 vccd1 _0257_ sky130_fd_sc_hd__mux2_1
XANTENNA__2494__A0 _0956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2109_ _0615_ net312 _1484_ vssd1 vssd1 vccd1 vccd1 _0739_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_37_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2246__A0 _0637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3158_ CB_1.config_dataA\[19\] CB_1.config_dataA\[20\] net222 vssd1 vssd1 vccd1 vccd1
+ _0326_ sky130_fd_sc_hd__mux2_1
XANTENNA__1772__A2 net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2788__A1 _0985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2460_ net31 net32 net18 net19 net181 net180 vssd1 vssd1 vccd1 vccd1 _1088_ sky130_fd_sc_hd__mux4_1
Xrebuffer4 net315 vssd1 vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__clkbuf_2
X_2391_ _1401_ SB0.route_sel\[103\] vssd1 vssd1 vccd1 vccd1 _1019_ sky130_fd_sc_hd__nand2_1
XFILLER_3_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2491__A3 net23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2228__A0 net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3012_ SB0.route_sel\[52\] SB0.route_sel\[51\] net294 vssd1 vssd1 vccd1 vccd1 _0180_
+ sky130_fd_sc_hd__mux2_1
XFILLER_51_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3020__S net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2658_ LE_0A.config_data\[15\] LE_0A.config_data\[14\] _1180_ vssd1 vssd1 vccd1 vccd1
+ _1285_ sky130_fd_sc_hd__mux2_1
X_2589_ net143 net156 LEI0.config_data\[24\] vssd1 vssd1 vccd1 vccd1 _1216_ sky130_fd_sc_hd__mux2_1
X_1609_ SB0.route_sel\[2\] vssd1 vssd1 vccd1 vccd1 _1447_ sky130_fd_sc_hd__inv_2
X_2727_ _1430_ SB0.route_sel\[32\] _1431_ SB0.route_sel\[35\] _1333_ vssd1 vssd1 vccd1
+ vccd1 _1334_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout284_X net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout179 CB_0.config_dataB\[15\] vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__buf_2
XANTENNA_input1_A CBeast_in[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout157 net159 vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__buf_2
Xfanout168 _1499_ vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__buf_2
XFILLER_63_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2054__B net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_8_clk_A clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input57_A SBwest_in[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3105__S net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input12_X net12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2944__S net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1701__X _1539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1891_ _0518_ _0506_ _0520_ vssd1 vssd1 vccd1 vccd1 _0521_ sky130_fd_sc_hd__a21oi_4
X_1960_ SB0.route_sel\[90\] SB0.route_sel\[91\] vssd1 vssd1 vccd1 vccd1 _0590_ sky130_fd_sc_hd__nand2_1
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3492_ clknet_leaf_16_clk _0312_ net282 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[6\]
+ sky130_fd_sc_hd__dfstp_1
X_2443_ net180 CB_0.config_dataB\[10\] vssd1 vssd1 vccd1 vccd1 _1071_ sky130_fd_sc_hd__and2b_1
X_2512_ LE_0B.config_data\[13\] _1032_ _1064_ _1139_ vssd1 vssd1 vccd1 vccd1 _1140_
+ sky130_fd_sc_hd__a211o_1
XFILLER_5_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2449__A0 net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2374_ _0952_ net336 net313 _0967_ CB_0.config_dataB\[2\] vssd1 vssd1 vccd1 vccd1
+ _1002_ sky130_fd_sc_hd__a221o_1
Xclone9 _0467_ _0461_ _0965_ net306 vssd1 vssd1 vccd1 vccd1 net319 sky130_fd_sc_hd__a211o_1
XANTENNA__2707__X net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_49_Left_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input4_X net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_58_Left_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2806__B1_N _0615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2090_ net303 LEI0.config_data\[23\] _0719_ vssd1 vssd1 vccd1 vccd1 _0720_ sky130_fd_sc_hd__or3_1
XFILLER_21_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2992_ SB0.route_sel\[32\] SB0.route_sel\[31\] net287 vssd1 vssd1 vccd1 vccd1 _0160_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_16_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1874_ net145 _0502_ net237 vssd1 vssd1 vccd1 vccd1 _0504_ sky130_fd_sc_hd__o21ai_1
X_1943_ net158 net166 net162 _0510_ _0349_ vssd1 vssd1 vccd1 vccd1 _0573_ sky130_fd_sc_hd__o32a_1
XANTENNA__1957__A2 net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3475_ clknet_leaf_10_clk _0295_ net264 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[14\]
+ sky130_fd_sc_hd__dfstp_1
X_2426_ net17 net24 net25 net26 net183 net182 vssd1 vssd1 vccd1 vccd1 _1054_ sky130_fd_sc_hd__mux4_1
X_2288_ net6 net7 CB_1.config_dataA\[15\] vssd1 vssd1 vccd1 vccd1 _0917_ sky130_fd_sc_hd__mux2_1
X_2357_ _0393_ _0384_ _0984_ net305 vssd1 vssd1 vccd1 vccd1 _0985_ sky130_fd_sc_hd__a211o_4
XTAP_TAPCELL_ROW_50_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2373__A2 _0665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2125__A2 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2347__X _0975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2061__A1 _0683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2116__A2 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3260_ clknet_leaf_2_clk net452 net244 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_1590_ SB0.route_sel\[43\] vssd1 vssd1 vccd1 vccd1 _1428_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2073_ CB_1.config_dataB\[7\] _0697_ _0700_ _0702_ vssd1 vssd1 vccd1 vccd1 _0703_
+ sky130_fd_sc_hd__o211a_1
X_2142_ net9 net330 net195 vssd1 vssd1 vccd1 vccd1 _0772_ sky130_fd_sc_hd__mux2_1
X_3191_ clknet_leaf_0_clk _0011_ net243 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_2211_ LEI0.config_data\[19\] _0837_ LEI0.config_data\[20\] _0839_ net303 vssd1 vssd1
+ vccd1 vccd1 _0840_ sky130_fd_sc_hd__a2111oi_4
X_2975_ SB0.route_sel\[15\] SB0.route_sel\[14\] net291 vssd1 vssd1 vccd1 vccd1 _0143_
+ sky130_fd_sc_hd__mux2_1
X_1788_ _1518_ _0417_ vssd1 vssd1 vccd1 vccd1 _0418_ sky130_fd_sc_hd__nor2_1
X_1926_ net149 _0375_ _0510_ net236 vssd1 vssd1 vccd1 vccd1 _0556_ sky130_fd_sc_hd__o31a_1
X_1857_ SB0.route_sel\[9\] SB0.route_sel\[8\] _0485_ _0486_ vssd1 vssd1 vccd1 vccd1
+ _0487_ sky130_fd_sc_hd__a211o_4
X_3527_ clknet_leaf_1_clk net430 net244 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data_in
+ sky130_fd_sc_hd__dfrtp_1
X_3458_ clknet_leaf_13_clk _0278_ net277 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[22\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_39_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2409_ _1035_ LEI0.config_data\[16\] _1036_ vssd1 vssd1 vccd1 vccd1 _1037_ sky130_fd_sc_hd__o21ba_4
X_3389_ clknet_leaf_3_clk _0209_ net253 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[81\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__1866__B2 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2291__A1 _0615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1885__C net55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output126_A net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3494__SET_B net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold93 LE_0B.config_data\[5\] vssd1 vssd1 vccd1 vccd1 net403 sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 _0089_ vssd1 vssd1 vccd1 vccd1 net392 sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 LE_1A.config_data\[6\] vssd1 vssd1 vccd1 vccd1 net381 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_61_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2952__S net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2760_ SB0.route_sel\[116\] _1453_ _1454_ SB0.route_sel\[115\] vssd1 vssd1 vccd1
+ vccd1 _1356_ sky130_fd_sc_hd__o22a_1
XANTENNA__1793__B1 SB0.route_sel\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2585__A2 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1642_ net199 vssd1 vssd1 vccd1 vccd1 _1480_ sky130_fd_sc_hd__inv_2
X_2691_ SB0.route_sel\[80\] _1406_ _1407_ SB0.route_sel\[83\] _1309_ vssd1 vssd1 vccd1
+ vccd1 _1310_ sky130_fd_sc_hd__a221o_1
XANTENNA_2 SBwest_in[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1711_ _1548_ _1539_ net305 vssd1 vssd1 vccd1 vccd1 _1549_ sky130_fd_sc_hd__a21oi_2
X_3243_ clknet_leaf_6_clk _0063_ net255 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_1573_ SB0.route_sel\[74\] vssd1 vssd1 vccd1 vccd1 _1411_ sky130_fd_sc_hd__inv_2
X_3312_ clknet_leaf_23_clk _0132_ net272 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[4\]
+ sky130_fd_sc_hd__dfstp_1
Xrebuffer14 net325 vssd1 vssd1 vccd1 vccd1 net324 sky130_fd_sc_hd__clkbuf_1
Xrebuffer25 net10 vssd1 vssd1 vccd1 vccd1 net335 sky130_fd_sc_hd__dlygate4sd1_1
X_2125_ LEI0.config_data\[35\] net239 _0754_ _0728_ _0725_ vssd1 vssd1 vccd1 vccd1
+ _0755_ sky130_fd_sc_hd__a32o_2
X_3174_ net476 net485 net203 vssd1 vssd1 vccd1 vccd1 _0342_ sky130_fd_sc_hd__mux2_1
X_2056_ LEI0.config_data\[9\] net160 vssd1 vssd1 vccd1 vccd1 _0686_ sky130_fd_sc_hd__nand2_1
XFILLER_19_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1909_ _0538_ _0537_ _0532_ vssd1 vssd1 vccd1 vccd1 _0539_ sky130_fd_sc_hd__or3b_4
XANTENNA__2576__A2 net29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout157_A net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2958_ CB_1.config_dataB\[22\] CB_1.config_dataB\[23\] net222 vssd1 vssd1 vccd1 vccd1
+ _0126_ sky130_fd_sc_hd__mux2_1
X_2889_ net401 LE_0A.config_data\[9\] net216 vssd1 vssd1 vccd1 vccd1 _0058_ sky130_fd_sc_hd__mux2_1
XANTENNA__2328__A2 _0415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2264__A1 _1552_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput94 net94 vssd1 vssd1 vccd1 vccd1 CBnorth_out[15] sky130_fd_sc_hd__buf_6
XANTENNA__2947__S net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput72 net72 vssd1 vssd1 vccd1 vccd1 CBeast_out[0] sky130_fd_sc_hd__buf_6
Xoutput83 net83 vssd1 vssd1 vccd1 vccd1 CBeast_out[5] sky130_fd_sc_hd__buf_6
XANTENNA__2255__A1 _0584_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2007__A1 _0633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2255__B2 _0564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2812_ _0373_ net161 _0679_ vssd1 vssd1 vccd1 vccd1 _1383_ sky130_fd_sc_hd__o21bai_4
X_2743_ _1344_ _0488_ vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__and2_4
X_2674_ _1298_ _0581_ vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__and2_4
X_1556_ SB0.route_sel\[104\] vssd1 vssd1 vccd1 vccd1 _1394_ sky130_fd_sc_hd__inv_2
X_1625_ CB_1.config_dataA\[18\] vssd1 vssd1 vccd1 vccd1 _1463_ sky130_fd_sc_hd__inv_2
XANTENNA__2270__X _0899_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout274_A net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout306 net308 vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__buf_2
X_3157_ CB_1.config_dataA\[18\] CB_1.config_dataA\[19\] net222 vssd1 vssd1 vccd1 vccd1
+ _0325_ sky130_fd_sc_hd__mux2_1
X_3226_ clknet_leaf_28_clk _0046_ net248 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[46\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_54_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2108_ net15 net16 net2 net3 CB_1.config_dataB\[10\] CB_1.config_dataB\[11\] vssd1
+ vssd1 vccd1 vccd1 _0738_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_37_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3088_ CB_0.config_data_inA CB_0.config_dataA\[0\] net219 vssd1 vssd1 vccd1 vccd1
+ _0256_ sky130_fd_sc_hd__mux2_1
XANTENNA__2246__A1 _0615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2039_ _0375_ net149 _0593_ net235 vssd1 vssd1 vccd1 vccd1 _0669_ sky130_fd_sc_hd__o31a_1
XANTENNA__2182__A0 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1772__A3 net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrebuffer5 net316 vssd1 vssd1 vccd1 vccd1 net315 sky130_fd_sc_hd__clkbuf_1
X_2390_ _0580_ _0570_ _1017_ net310 vssd1 vssd1 vccd1 vccd1 _1018_ sky130_fd_sc_hd__a211o_4
XANTENNA__2173__B1 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3011_ SB0.route_sel\[51\] SB0.route_sel\[50\] net294 vssd1 vssd1 vccd1 vccd1 _0179_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_59_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2228__A1 net12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2726_ SB0.route_sel\[38\] SB0.route_sel\[39\] vssd1 vssd1 vccd1 vccd1 _1333_ sky130_fd_sc_hd__nor2_1
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2657_ _1245_ _1250_ _1252_ _1282_ vssd1 vssd1 vccd1 vccd1 _1284_ sky130_fd_sc_hd__o31a_1
X_2588_ LEI0.config_data\[24\] _1493_ _1214_ LEI0.config_data\[25\] vssd1 vssd1 vccd1
+ vccd1 _1215_ sky130_fd_sc_hd__o211a_1
Xfanout147 _1493_ vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__buf_2
X_1608_ SB0.route_sel\[1\] vssd1 vssd1 vccd1 vccd1 _1446_ sky130_fd_sc_hd__inv_2
X_3209_ clknet_leaf_3_clk _0029_ net251 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_27_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout158 net159 vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__clkbuf_2
Xfanout169 _1498_ vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__buf_2
XFILLER_27_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3121__S net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_16_Right_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1890_ net309 _0496_ vssd1 vssd1 vccd1 vccd1 _0520_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_25_Right_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3491_ clknet_leaf_16_clk _0311_ net282 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[5\]
+ sky130_fd_sc_hd__dfstp_1
X_2373_ _0675_ _0665_ _1000_ net309 vssd1 vssd1 vccd1 vccd1 _1001_ sky130_fd_sc_hd__a211o_4
XANTENNA__2146__A0 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2442_ net304 LEI0.config_data\[29\] _1067_ _1069_ vssd1 vssd1 vccd1 vccd1 _1070_
+ sky130_fd_sc_hd__or4_1
X_2511_ _1025_ _1026_ _1031_ LE_0B.config_data\[12\] vssd1 vssd1 vccd1 vccd1 _1139_
+ sky130_fd_sc_hd__o211a_1
XFILLER_56_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2449__A1 net24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_34_Right_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout237_A net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_43_Right_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2709_ _1418_ SB0.route_sel\[56\] _1419_ SB0.route_sel\[59\] _1321_ vssd1 vssd1 vccd1
+ vccd1 _1322_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_52_Right_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2137__A0 net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_61_Right_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2612__A1 _1001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2612__B2 _0998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2376__A0 net31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1942_ net166 net162 net5 vssd1 vssd1 vccd1 vccd1 _0572_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2991_ SB0.route_sel\[31\] SB0.route_sel\[30\] net287 vssd1 vssd1 vccd1 vccd1 _0159_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_16_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1873_ net153 _0499_ _0500_ _0502_ vssd1 vssd1 vccd1 vccd1 _0503_ sky130_fd_sc_hd__o211a_1
XANTENNA__1957__A3 net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3474_ clknet_leaf_11_clk _0294_ net263 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[13\]
+ sky130_fd_sc_hd__dfstp_1
X_2425_ net182 _1051_ _1052_ vssd1 vssd1 vccd1 vccd1 _1053_ sky130_fd_sc_hd__a21oi_1
XANTENNA_clone32_C1 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2356_ SB0.route_sel\[34\] SB0.route_sel\[35\] SB0.route_sel\[37\] _1433_ _0983_
+ vssd1 vssd1 vccd1 vccd1 _0984_ sky130_fd_sc_hd__o221a_1
X_2287_ _0912_ _0913_ _0915_ vssd1 vssd1 vccd1 vccd1 _0916_ sky130_fd_sc_hd__a21o_1
XANTENNA__1948__A3 net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_7_clk_A clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2358__B1 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2530__A0 _0956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2125__A3 _0754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2363__X _0991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3454__SET_B net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2597__A0 net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2210_ _0838_ LEI0.config_data\[19\] vssd1 vssd1 vccd1 vccd1 _0839_ sky130_fd_sc_hd__nor2_4
X_3190_ clknet_leaf_0_clk _0010_ net243 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_64_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2072_ CB_1.config_dataB\[7\] _0701_ CB_1.config_dataB\[8\] vssd1 vssd1 vccd1 vccd1
+ _0702_ sky130_fd_sc_hd__a21oi_1
X_2141_ net345 net359 net327 net344 net195 net194 vssd1 vssd1 vccd1 vccd1 _0771_ sky130_fd_sc_hd__mux4_1
XFILLER_34_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1925_ net158 net165 net162 _0510_ _0375_ vssd1 vssd1 vccd1 vccd1 _0555_ sky130_fd_sc_hd__o32a_1
X_2974_ SB0.route_sel\[14\] SB0.route_sel\[13\] net291 vssd1 vssd1 vccd1 vccd1 _0142_
+ sky130_fd_sc_hd__mux2_1
X_1787_ CB_0.config_dataB\[23\] CB_0.config_dataB\[22\] vssd1 vssd1 vccd1 vccd1 _0417_
+ sky130_fd_sc_hd__or2_2
X_1856_ net144 _0484_ net237 vssd1 vssd1 vccd1 vccd1 _0486_ sky130_fd_sc_hd__o21ai_2
XANTENNA__2152__C CB_1.config_dataB\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3526_ clknet_leaf_1_clk net380 net244 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_3457_ clknet_leaf_13_clk _0277_ net277 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[21\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_57_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2339_ net185 CB_0.config_dataB\[1\] vssd1 vssd1 vccd1 vccd1 _0967_ sky130_fd_sc_hd__nor2_1
XFILLER_39_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2408_ net304 LEI0.config_data\[17\] _1034_ vssd1 vssd1 vccd1 vccd1 _1036_ sky130_fd_sc_hd__or3_1
X_3388_ clknet_leaf_3_clk _0208_ net253 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[80\]
+ sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_2_Right_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2579__A0 _0956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input32_A CBnorth_in[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold83 LE_0A.config_data\[10\] vssd1 vssd1 vccd1 vccd1 net393 sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 _0092_ vssd1 vssd1 vccd1 vccd1 net382 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_output119_A net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold94 LE_1A.config_data\[9\] vssd1 vssd1 vccd1 vccd1 net404 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2253__B _0521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1710_ _1547_ _1546_ _1538_ vssd1 vssd1 vccd1 vccd1 _1548_ sky130_fd_sc_hd__or3b_4
XANTENNA__1793__B2 SB0.route_sel\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1641_ CB_1.config_dataB\[7\] vssd1 vssd1 vccd1 vccd1 _1479_ sky130_fd_sc_hd__inv_2
X_1572_ SB0.route_sel\[73\] vssd1 vssd1 vccd1 vccd1 _1410_ sky130_fd_sc_hd__inv_2
X_2690_ SB0.route_sel\[87\] SB0.route_sel\[86\] vssd1 vssd1 vccd1 vccd1 _1309_ sky130_fd_sc_hd__nor2_1
X_3311_ clknet_leaf_23_clk _0131_ net272 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[3\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_3 _0333_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3242_ clknet_leaf_7_clk net412 net255 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_2124_ _0742_ _0753_ _0730_ vssd1 vssd1 vccd1 vccd1 _0754_ sky130_fd_sc_hd__a21o_1
XANTENNA__2268__X _0897_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3173_ net473 net476 net203 vssd1 vssd1 vccd1 vccd1 _0341_ sky130_fd_sc_hd__mux2_1
Xrebuffer15 _0675_ vssd1 vssd1 vccd1 vccd1 net325 sky130_fd_sc_hd__clkbuf_1
X_2055_ net326 net155 LEI0.config_data\[9\] vssd1 vssd1 vccd1 vccd1 _0685_ sky130_fd_sc_hd__mux2_1
XFILLER_19_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1908_ net145 _0536_ net238 vssd1 vssd1 vccd1 vccd1 _0538_ sky130_fd_sc_hd__o21ai_1
XANTENNA__2576__A3 net30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2888_ net377 LE_0A.config_data\[8\] net216 vssd1 vssd1 vccd1 vccd1 _0057_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_32_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1839_ SB0.route_sel\[7\] SB0.route_sel\[6\] vssd1 vssd1 vccd1 vccd1 _0469_ sky130_fd_sc_hd__nand2b_1
X_2957_ CB_1.config_dataB\[21\] CB_1.config_dataB\[22\] net222 vssd1 vssd1 vccd1 vccd1
+ _0125_ sky130_fd_sc_hd__mux2_1
X_3509_ clknet_leaf_23_clk _0329_ net274 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[23\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_17_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2567__A3 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput95 net95 vssd1 vssd1 vccd1 vccd1 CBnorth_out[1] sky130_fd_sc_hd__buf_6
XFILLER_48_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3124__S net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput73 net73 vssd1 vssd1 vccd1 vccd1 CBeast_out[10] sky130_fd_sc_hd__buf_6
XANTENNA_input35_X net35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput84 net84 vssd1 vssd1 vccd1 vccd1 CBeast_out[6] sky130_fd_sc_hd__buf_2
XFILLER_56_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_28_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__2007__A2 _0627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2811_ _1382_ _0641_ _0642_ vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__a21boi_2
XANTENNA_clkbuf_leaf_32_clk_A clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2742_ SB0.route_sel\[10\] _1444_ SB0.route_sel\[13\] _1445_ _1343_ vssd1 vssd1 vccd1
+ vccd1 _1344_ sky130_fd_sc_hd__a221o_1
XANTENNA__3510__SET_B net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2673_ SB0.route_sel\[104\] _1395_ _1396_ SB0.route_sel\[107\] _1297_ vssd1 vssd1
+ vccd1 vccd1 _1298_ sky130_fd_sc_hd__a221o_1
Xfanout307 net308 vssd1 vssd1 vccd1 vccd1 net307 sky130_fd_sc_hd__buf_2
X_1624_ CB_1.config_dataA\[14\] vssd1 vssd1 vccd1 vccd1 _1462_ sky130_fd_sc_hd__inv_2
XFILLER_54_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clone40_C1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2107_ _0732_ _0734_ _0736_ CB_1.config_dataB\[13\] vssd1 vssd1 vccd1 vccd1 _0737_
+ sky130_fd_sc_hd__o211ai_1
X_3087_ net136 SB0.route_sel\[126\] net301 vssd1 vssd1 vccd1 vccd1 _0255_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_37_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_19_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_clk
+ sky130_fd_sc_hd__clkbuf_8
X_3156_ CB_1.config_dataA\[17\] CB_1.config_dataA\[18\] net222 vssd1 vssd1 vccd1 vccd1
+ _0324_ sky130_fd_sc_hd__mux2_1
X_3225_ clknet_leaf_31_clk _0045_ net248 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[45\]
+ sky130_fd_sc_hd__dfrtp_1
X_2038_ net157 net165 net161 _0593_ _0375_ vssd1 vssd1 vccd1 vccd1 _0668_ sky130_fd_sc_hd__o32a_1
XANTENNA__2182__A1 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2237__A2 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrebuffer6 net322 vssd1 vssd1 vccd1 vccd1 net316 sky130_fd_sc_hd__clkbuf_1
XANTENNA__1684__B1 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3010_ SB0.route_sel\[50\] SB0.route_sel\[49\] net294 vssd1 vssd1 vccd1 vccd1 _0178_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__2228__A2 net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_8_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2656_ _1280_ _1281_ net146 vssd1 vssd1 vccd1 vccd1 _1283_ sky130_fd_sc_hd__o21bai_1
XANTENNA_clone35_C1 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2725_ _1332_ _0394_ vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__and2_4
X_2587_ CB_1.le_outB LEI0.config_data\[24\] vssd1 vssd1 vccd1 vccd1 _1214_ sky130_fd_sc_hd__nand2_2
XANTENNA__2868__S net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout159 _1494_ vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__buf_2
X_1607_ SB0.route_sel\[12\] vssd1 vssd1 vccd1 vccd1 _1445_ sky130_fd_sc_hd__inv_2
Xfanout148 net150 vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__buf_8
X_3139_ CB_1.config_dataA\[0\] net176 net230 vssd1 vssd1 vccd1 vccd1 _0307_ sky130_fd_sc_hd__mux2_1
X_3208_ clknet_leaf_3_clk _0028_ net245 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_50_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2366__X _0994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3490_ clknet_leaf_16_clk _0310_ net280 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[4\]
+ sky130_fd_sc_hd__dfstp_1
X_2510_ LE_0B.config_data\[14\] LE_0B.config_data\[15\] _1032_ vssd1 vssd1 vccd1 vccd1
+ _1138_ sky130_fd_sc_hd__mux2_1
X_2372_ SB0.route_sel\[66\] SB0.route_sel\[67\] SB0.route_sel\[69\] _1417_ _0999_
+ vssd1 vssd1 vccd1 vccd1 _1000_ sky130_fd_sc_hd__o221a_1
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2441_ LEI0.config_data\[28\] _1068_ vssd1 vssd1 vccd1 vccd1 _1069_ sky130_fd_sc_hd__nor2_1
XANTENNA__2146__A1 net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2449__A2 net25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2082__A0 _0615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2639_ _1265_ vssd1 vssd1 vccd1 vccd1 _1266_ sky130_fd_sc_hd__inv_2
X_2708_ SB0.route_sel\[63\] SB0.route_sel\[62\] vssd1 vssd1 vccd1 vccd1 _1321_ sky130_fd_sc_hd__nor2_1
XFILLER_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input62_A SBwest_in[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1941_ SB0.route_sel\[106\] SB0.route_sel\[107\] vssd1 vssd1 vccd1 vccd1 _0571_ sky130_fd_sc_hd__nand2_1
XANTENNA__1811__B1 net26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1872_ _1544_ _0501_ vssd1 vssd1 vccd1 vccd1 _0502_ sky130_fd_sc_hd__or2_1
X_2990_ SB0.route_sel\[30\] SB0.route_sel\[29\] net287 vssd1 vssd1 vccd1 vccd1 _0158_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_16_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3473_ clknet_leaf_11_clk _0293_ net262 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[12\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__1903__X _0533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2424_ net319 _1039_ _1040_ net371 CB_0.config_dataB\[7\] vssd1 vssd1 vccd1 vccd1
+ _1052_ sky130_fd_sc_hd__a221o_1
XANTENNA_clone32_B1 _0984_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2286_ _0584_ _0911_ _0914_ _0564_ vssd1 vssd1 vccd1 vccd1 _0915_ sky130_fd_sc_hd__a22o_1
X_2355_ SB0.route_sel\[38\] SB0.route_sel\[39\] vssd1 vssd1 vccd1 vccd1 _0983_ sky130_fd_sc_hd__nand2b_1
XFILLER_52_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout302_X net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1899__C net54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2530__A1 _0959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2294__A0 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2597__A1 net24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2046__B1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3127__S net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2140_ _0762_ _0765_ _0766_ _0769_ vssd1 vssd1 vccd1 vccd1 _0770_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_64_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2071_ net11 net12 net13 net331 net199 net198 vssd1 vssd1 vccd1 vccd1 _0701_ sky130_fd_sc_hd__mux4_1
XFILLER_38_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_28_Left_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1855_ net153 _0482_ _0483_ _0484_ vssd1 vssd1 vccd1 vccd1 _0485_ sky130_fd_sc_hd__o211a_4
X_1924_ net165 net162 net4 vssd1 vssd1 vccd1 vccd1 _0554_ sky130_fd_sc_hd__o21ai_1
X_2973_ SB0.route_sel\[13\] SB0.route_sel\[12\] net291 vssd1 vssd1 vccd1 vccd1 _0141_
+ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_12_Left_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2037__B1 net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3456_ clknet_leaf_13_clk _0276_ net277 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[20\]
+ sky130_fd_sc_hd__dfstp_1
X_1786_ CB_0.config_dataB\[23\] CB_0.config_dataB\[22\] vssd1 vssd1 vccd1 vccd1 _0416_
+ sky130_fd_sc_hd__nor2_1
X_3525_ clknet_leaf_1_clk _0345_ net241 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout297_A net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2407_ net142 net156 LEI0.config_data\[15\] vssd1 vssd1 vccd1 vccd1 _1035_ sky130_fd_sc_hd__mux2_4
X_3387_ clknet_leaf_4_clk _0207_ net252 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[79\]
+ sky130_fd_sc_hd__dfstp_1
X_2338_ _0467_ _0461_ _0965_ net306 vssd1 vssd1 vccd1 vccd1 _0966_ sky130_fd_sc_hd__a211o_4
X_2269_ LEI0.config_data\[32\] net232 _0897_ net140 vssd1 vssd1 vccd1 vccd1 _0898_
+ sky130_fd_sc_hd__a31oi_2
XANTENNA__2579__A1 _0959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2043__A3 net63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold73 LE_0A.config_data\[6\] vssd1 vssd1 vccd1 vccd1 net383 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input25_A CBnorth_in[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold84 LE_0B.config_data\[6\] vssd1 vssd1 vccd1 vccd1 net394 sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 _0095_ vssd1 vssd1 vccd1 vccd1 net405 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_31_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1640_ net201 vssd1 vssd1 vccd1 vccd1 _1478_ sky130_fd_sc_hd__inv_2
X_1571_ SB0.route_sel\[84\] vssd1 vssd1 vccd1 vccd1 _1409_ sky130_fd_sc_hd__inv_2
X_3310_ clknet_leaf_24_clk _0130_ net272 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[2\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_4 _0334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3241_ clknet_leaf_6_clk net385 net255 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_2123_ _0745_ _0749_ _0752_ CB_1.config_dataB\[14\] vssd1 vssd1 vccd1 vccd1 _0753_
+ sky130_fd_sc_hd__a31oi_1
XANTENNA_clkbuf_leaf_6_clk_A clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2258__A0 _0428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3172_ LE_1B.config_data\[8\] net473 net203 vssd1 vssd1 vccd1 vccd1 _0340_ sky130_fd_sc_hd__mux2_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clone38_C1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2054_ LEI0.config_data\[11\] net232 vssd1 vssd1 vccd1 vccd1 _0684_ sky130_fd_sc_hd__and2_4
X_1907_ net153 _0534_ _0535_ _0536_ vssd1 vssd1 vccd1 vccd1 _0537_ sky130_fd_sc_hd__o211a_1
X_2887_ net383 net377 net216 vssd1 vssd1 vccd1 vccd1 _0056_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_32_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2956_ CB_1.config_dataB\[20\] CB_1.config_dataB\[21\] net222 vssd1 vssd1 vccd1 vccd1
+ _0124_ sky130_fd_sc_hd__mux2_1
X_1838_ _0467_ _0461_ net306 vssd1 vssd1 vccd1 vccd1 _0468_ sky130_fd_sc_hd__a21oi_4
XANTENNA__2731__Y net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2497__A0 net27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3439_ clknet_leaf_8_clk _0259_ net259 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[3\]
+ sky130_fd_sc_hd__dfstp_1
X_1769_ _1495_ net361 net357 _0398_ _1477_ vssd1 vssd1 vccd1 vccd1 _0399_ sky130_fd_sc_hd__a221o_1
X_3508_ clknet_leaf_23_clk _0328_ net274 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[22\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_57_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput96 net96 vssd1 vssd1 vccd1 vccd1 CBnorth_out[2] sky130_fd_sc_hd__buf_6
XANTENNA_input28_X net28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output131_A net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput74 net74 vssd1 vssd1 vccd1 vccd1 CBeast_out[11] sky130_fd_sc_hd__buf_6
XANTENNA__2804__B1_N _0564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput85 net85 vssd1 vssd1 vccd1 vccd1 CBeast_out[7] sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_46_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2672_ SB0.route_sel\[110\] SB0.route_sel\[111\] vssd1 vssd1 vccd1 vccd1 _1297_ sky130_fd_sc_hd__nor2_1
XFILLER_31_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2810_ _1555_ net161 _0659_ vssd1 vssd1 vccd1 vccd1 _1382_ sky130_fd_sc_hd__o21bai_4
X_2741_ SB0.route_sel\[9\] SB0.route_sel\[8\] vssd1 vssd1 vccd1 vccd1 _1343_ sky130_fd_sc_hd__nor2_1
Xfanout308 net66 vssd1 vssd1 vccd1 vccd1 net308 sky130_fd_sc_hd__clkbuf_2
X_1623_ CB_1.config_dataA\[12\] vssd1 vssd1 vccd1 vccd1 _1461_ sky130_fd_sc_hd__inv_2
X_3224_ clknet_leaf_30_clk _0044_ net248 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[44\]
+ sky130_fd_sc_hd__dfrtp_1
.ends

