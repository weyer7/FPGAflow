VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fpga
  CLASS BLOCK ;
  FOREIGN fpga ;
  ORIGIN -8.000 -8.000 ;
  SIZE 453.000 BY 455.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 239.930 459.000 240.210 463.000 ;
    END
  END clk
  PIN config_data_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 8.000 232.440 12.000 233.040 ;
    END
  END config_data_in
  PIN config_data_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 457.000 239.240 461.000 239.840 ;
    END
  END config_data_out
  PIN config_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 249.590 459.000 249.870 463.000 ;
    END
  END config_en
  PIN io_east_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 457.000 144.040 461.000 144.640 ;
    END
  END io_east_in[0]
  PIN io_east_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 457.000 198.440 461.000 199.040 ;
    END
  END io_east_in[10]
  PIN io_east_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 457.000 205.240 461.000 205.840 ;
    END
  END io_east_in[11]
  PIN io_east_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 457.000 208.640 461.000 209.240 ;
    END
  END io_east_in[12]
  PIN io_east_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 457.000 215.440 461.000 216.040 ;
    END
  END io_east_in[13]
  PIN io_east_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.090 8.000 8.370 12.000 ;
    END
  END io_east_in[14]
  PIN io_east_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.310 8.000 11.590 12.000 ;
    END
  END io_east_in[15]
  PIN io_east_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 457.000 331.040 461.000 331.640 ;
    END
  END io_east_in[16]
  PIN io_east_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 457.000 337.840 461.000 338.440 ;
    END
  END io_east_in[17]
  PIN io_east_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 457.000 341.240 461.000 341.840 ;
    END
  END io_east_in[18]
  PIN io_east_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 457.000 348.040 461.000 348.640 ;
    END
  END io_east_in[19]
  PIN io_east_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 457.000 150.840 461.000 151.440 ;
    END
  END io_east_in[1]
  PIN io_east_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 457.000 351.440 461.000 352.040 ;
    END
  END io_east_in[20]
  PIN io_east_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 457.000 358.240 461.000 358.840 ;
    END
  END io_east_in[21]
  PIN io_east_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 457.000 365.040 461.000 365.640 ;
    END
  END io_east_in[22]
  PIN io_east_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 457.000 368.440 461.000 369.040 ;
    END
  END io_east_in[23]
  PIN io_east_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 457.000 375.240 461.000 375.840 ;
    END
  END io_east_in[24]
  PIN io_east_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 457.000 378.640 461.000 379.240 ;
    END
  END io_east_in[25]
  PIN io_east_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 457.000 385.440 461.000 386.040 ;
    END
  END io_east_in[26]
  PIN io_east_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 457.000 392.240 461.000 392.840 ;
    END
  END io_east_in[27]
  PIN io_east_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 457.000 395.640 461.000 396.240 ;
    END
  END io_east_in[28]
  PIN io_east_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 457.000 402.440 461.000 403.040 ;
    END
  END io_east_in[29]
  PIN io_east_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 457.000 154.240 461.000 154.840 ;
    END
  END io_east_in[2]
  PIN io_east_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.530 8.000 14.810 12.000 ;
    END
  END io_east_in[30]
  PIN io_east_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.750 8.000 18.030 12.000 ;
    END
  END io_east_in[31]
  PIN io_east_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 457.000 161.040 461.000 161.640 ;
    END
  END io_east_in[3]
  PIN io_east_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 457.000 164.440 461.000 165.040 ;
    END
  END io_east_in[4]
  PIN io_east_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 457.000 171.240 461.000 171.840 ;
    END
  END io_east_in[5]
  PIN io_east_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 457.000 178.040 461.000 178.640 ;
    END
  END io_east_in[6]
  PIN io_east_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 457.000 181.440 461.000 182.040 ;
    END
  END io_east_in[7]
  PIN io_east_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 457.000 188.240 461.000 188.840 ;
    END
  END io_east_in[8]
  PIN io_east_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 457.000 191.640 461.000 192.240 ;
    END
  END io_east_in[9]
  PIN io_east_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 457.000 69.240 461.000 69.840 ;
    END
  END io_east_out[0]
  PIN io_east_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 457.000 123.640 461.000 124.240 ;
    END
  END io_east_out[10]
  PIN io_east_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 457.000 127.040 461.000 127.640 ;
    END
  END io_east_out[11]
  PIN io_east_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 457.000 133.840 461.000 134.440 ;
    END
  END io_east_out[12]
  PIN io_east_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 457.000 137.240 461.000 137.840 ;
    END
  END io_east_out[13]
  PIN io_east_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 8.000 222.240 12.000 222.840 ;
    END
  END io_east_out[14]
  PIN io_east_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 8.000 246.040 12.000 246.640 ;
    END
  END io_east_out[15]
  PIN io_east_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 457.000 256.240 461.000 256.840 ;
    END
  END io_east_out[16]
  PIN io_east_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 457.000 259.640 461.000 260.240 ;
    END
  END io_east_out[17]
  PIN io_east_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 457.000 266.440 461.000 267.040 ;
    END
  END io_east_out[18]
  PIN io_east_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 457.000 269.840 461.000 270.440 ;
    END
  END io_east_out[19]
  PIN io_east_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 457.000 72.640 461.000 73.240 ;
    END
  END io_east_out[1]
  PIN io_east_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 457.000 276.640 461.000 277.240 ;
    END
  END io_east_out[20]
  PIN io_east_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 457.000 283.440 461.000 284.040 ;
    END
  END io_east_out[21]
  PIN io_east_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 457.000 286.840 461.000 287.440 ;
    END
  END io_east_out[22]
  PIN io_east_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 457.000 293.640 461.000 294.240 ;
    END
  END io_east_out[23]
  PIN io_east_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 457.000 297.040 461.000 297.640 ;
    END
  END io_east_out[24]
  PIN io_east_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 457.000 303.840 461.000 304.440 ;
    END
  END io_east_out[25]
  PIN io_east_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 457.000 310.640 461.000 311.240 ;
    END
  END io_east_out[26]
  PIN io_east_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 457.000 314.040 461.000 314.640 ;
    END
  END io_east_out[27]
  PIN io_east_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 457.000 320.840 461.000 321.440 ;
    END
  END io_east_out[28]
  PIN io_east_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 457.000 324.240 461.000 324.840 ;
    END
  END io_east_out[29]
  PIN io_east_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 457.000 79.440 461.000 80.040 ;
    END
  END io_east_out[2]
  PIN io_east_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 8.000 167.840 12.000 168.440 ;
    END
  END io_east_out[30]
  PIN io_east_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 8.000 229.040 12.000 229.640 ;
    END
  END io_east_out[31]
  PIN io_east_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 457.000 82.840 461.000 83.440 ;
    END
  END io_east_out[3]
  PIN io_east_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 457.000 89.640 461.000 90.240 ;
    END
  END io_east_out[4]
  PIN io_east_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 457.000 96.440 461.000 97.040 ;
    END
  END io_east_out[5]
  PIN io_east_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 457.000 99.840 461.000 100.440 ;
    END
  END io_east_out[6]
  PIN io_east_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 457.000 106.640 461.000 107.240 ;
    END
  END io_east_out[7]
  PIN io_east_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 457.000 110.040 461.000 110.640 ;
    END
  END io_east_out[8]
  PIN io_east_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 457.000 116.840 461.000 117.440 ;
    END
  END io_east_out[9]
  PIN io_north_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 78.930 459.000 79.210 463.000 ;
    END
  END io_north_in[0]
  PIN io_north_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 133.670 459.000 133.950 463.000 ;
    END
  END io_north_in[10]
  PIN io_north_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 136.890 459.000 137.170 463.000 ;
    END
  END io_north_in[11]
  PIN io_north_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 143.330 459.000 143.610 463.000 ;
    END
  END io_north_in[12]
  PIN io_north_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 149.770 459.000 150.050 463.000 ;
    END
  END io_north_in[13]
  PIN io_north_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.970 8.000 21.250 12.000 ;
    END
  END io_north_in[14]
  PIN io_north_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.190 8.000 24.470 12.000 ;
    END
  END io_north_in[15]
  PIN io_north_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 262.470 459.000 262.750 463.000 ;
    END
  END io_north_in[16]
  PIN io_north_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 268.910 459.000 269.190 463.000 ;
    END
  END io_north_in[17]
  PIN io_north_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 272.130 459.000 272.410 463.000 ;
    END
  END io_north_in[18]
  PIN io_north_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 278.570 459.000 278.850 463.000 ;
    END
  END io_north_in[19]
  PIN io_north_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 82.150 459.000 82.430 463.000 ;
    END
  END io_north_in[1]
  PIN io_north_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 285.010 459.000 285.290 463.000 ;
    END
  END io_north_in[20]
  PIN io_north_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 291.450 459.000 291.730 463.000 ;
    END
  END io_north_in[21]
  PIN io_north_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 294.670 459.000 294.950 463.000 ;
    END
  END io_north_in[22]
  PIN io_north_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 301.110 459.000 301.390 463.000 ;
    END
  END io_north_in[23]
  PIN io_north_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 307.550 459.000 307.830 463.000 ;
    END
  END io_north_in[24]
  PIN io_north_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 310.770 459.000 311.050 463.000 ;
    END
  END io_north_in[25]
  PIN io_north_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 317.210 459.000 317.490 463.000 ;
    END
  END io_north_in[26]
  PIN io_north_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 323.650 459.000 323.930 463.000 ;
    END
  END io_north_in[27]
  PIN io_north_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 330.090 459.000 330.370 463.000 ;
    END
  END io_north_in[28]
  PIN io_north_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 333.310 459.000 333.590 463.000 ;
    END
  END io_north_in[29]
  PIN io_north_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 88.590 459.000 88.870 463.000 ;
    END
  END io_north_in[2]
  PIN io_north_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.410 8.000 27.690 12.000 ;
    END
  END io_north_in[30]
  PIN io_north_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.630 8.000 30.910 12.000 ;
    END
  END io_north_in[31]
  PIN io_north_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 95.030 459.000 95.310 463.000 ;
    END
  END io_north_in[3]
  PIN io_north_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 98.250 459.000 98.530 463.000 ;
    END
  END io_north_in[4]
  PIN io_north_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 104.690 459.000 104.970 463.000 ;
    END
  END io_north_in[5]
  PIN io_north_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 111.130 459.000 111.410 463.000 ;
    END
  END io_north_in[6]
  PIN io_north_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 117.570 459.000 117.850 463.000 ;
    END
  END io_north_in[7]
  PIN io_north_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 120.790 459.000 121.070 463.000 ;
    END
  END io_north_in[8]
  PIN io_north_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 127.230 459.000 127.510 463.000 ;
    END
  END io_north_in[9]
  PIN io_north_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 156.210 459.000 156.490 463.000 ;
    END
  END io_north_out[0]
  PIN io_north_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 210.950 459.000 211.230 463.000 ;
    END
  END io_north_out[10]
  PIN io_north_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 214.170 459.000 214.450 463.000 ;
    END
  END io_north_out[11]
  PIN io_north_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 220.610 459.000 220.890 463.000 ;
    END
  END io_north_out[12]
  PIN io_north_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 227.050 459.000 227.330 463.000 ;
    END
  END io_north_out[13]
  PIN io_north_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.790 459.000 282.070 463.000 ;
    END
  END io_north_out[14]
  PIN io_north_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 457.000 344.640 461.000 345.240 ;
    END
  END io_north_out[15]
  PIN io_north_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 339.750 459.000 340.030 463.000 ;
    END
  END io_north_out[16]
  PIN io_north_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 346.190 459.000 346.470 463.000 ;
    END
  END io_north_out[17]
  PIN io_north_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 349.410 459.000 349.690 463.000 ;
    END
  END io_north_out[18]
  PIN io_north_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 355.850 459.000 356.130 463.000 ;
    END
  END io_north_out[19]
  PIN io_north_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 159.430 459.000 159.710 463.000 ;
    END
  END io_north_out[1]
  PIN io_north_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 362.290 459.000 362.570 463.000 ;
    END
  END io_north_out[20]
  PIN io_north_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 368.730 459.000 369.010 463.000 ;
    END
  END io_north_out[21]
  PIN io_north_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 371.950 459.000 372.230 463.000 ;
    END
  END io_north_out[22]
  PIN io_north_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 378.390 459.000 378.670 463.000 ;
    END
  END io_north_out[23]
  PIN io_north_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 384.830 459.000 385.110 463.000 ;
    END
  END io_north_out[24]
  PIN io_north_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 388.050 459.000 388.330 463.000 ;
    END
  END io_north_out[25]
  PIN io_north_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 394.490 459.000 394.770 463.000 ;
    END
  END io_north_out[26]
  PIN io_north_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 400.930 459.000 401.210 463.000 ;
    END
  END io_north_out[27]
  PIN io_north_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 407.370 459.000 407.650 463.000 ;
    END
  END io_north_out[28]
  PIN io_north_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 410.590 459.000 410.870 463.000 ;
    END
  END io_north_out[29]
  PIN io_north_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 165.870 459.000 166.150 463.000 ;
    END
  END io_north_out[2]
  PIN io_north_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 457.000 232.440 461.000 233.040 ;
    END
  END io_north_out[30]
  PIN io_north_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.230 459.000 288.510 463.000 ;
    END
  END io_north_out[31]
  PIN io_north_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 172.310 459.000 172.590 463.000 ;
    END
  END io_north_out[3]
  PIN io_north_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 175.530 459.000 175.810 463.000 ;
    END
  END io_north_out[4]
  PIN io_north_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 181.970 459.000 182.250 463.000 ;
    END
  END io_north_out[5]
  PIN io_north_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 188.410 459.000 188.690 463.000 ;
    END
  END io_north_out[6]
  PIN io_north_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 194.850 459.000 195.130 463.000 ;
    END
  END io_north_out[7]
  PIN io_north_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 198.070 459.000 198.350 463.000 ;
    END
  END io_north_out[8]
  PIN io_north_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 204.510 459.000 204.790 463.000 ;
    END
  END io_north_out[9]
  PIN io_south_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 156.210 8.000 156.490 12.000 ;
    END
  END io_south_in[0]
  PIN io_south_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 210.950 8.000 211.230 12.000 ;
    END
  END io_south_in[10]
  PIN io_south_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 214.170 8.000 214.450 12.000 ;
    END
  END io_south_in[11]
  PIN io_south_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 220.610 8.000 220.890 12.000 ;
    END
  END io_south_in[12]
  PIN io_south_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 227.050 8.000 227.330 12.000 ;
    END
  END io_south_in[13]
  PIN io_south_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.850 8.000 34.130 12.000 ;
    END
  END io_south_in[14]
  PIN io_south_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.070 8.000 37.350 12.000 ;
    END
  END io_south_in[15]
  PIN io_south_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 339.750 8.000 340.030 12.000 ;
    END
  END io_south_in[16]
  PIN io_south_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 346.190 8.000 346.470 12.000 ;
    END
  END io_south_in[17]
  PIN io_south_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 349.410 8.000 349.690 12.000 ;
    END
  END io_south_in[18]
  PIN io_south_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 355.850 8.000 356.130 12.000 ;
    END
  END io_south_in[19]
  PIN io_south_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 159.430 8.000 159.710 12.000 ;
    END
  END io_south_in[1]
  PIN io_south_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 362.290 8.000 362.570 12.000 ;
    END
  END io_south_in[20]
  PIN io_south_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 368.730 8.000 369.010 12.000 ;
    END
  END io_south_in[21]
  PIN io_south_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 371.950 8.000 372.230 12.000 ;
    END
  END io_south_in[22]
  PIN io_south_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 378.390 8.000 378.670 12.000 ;
    END
  END io_south_in[23]
  PIN io_south_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 384.830 8.000 385.110 12.000 ;
    END
  END io_south_in[24]
  PIN io_south_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 388.050 8.000 388.330 12.000 ;
    END
  END io_south_in[25]
  PIN io_south_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 394.490 8.000 394.770 12.000 ;
    END
  END io_south_in[26]
  PIN io_south_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 400.930 8.000 401.210 12.000 ;
    END
  END io_south_in[27]
  PIN io_south_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 407.370 8.000 407.650 12.000 ;
    END
  END io_south_in[28]
  PIN io_south_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 410.590 8.000 410.870 12.000 ;
    END
  END io_south_in[29]
  PIN io_south_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 165.870 8.000 166.150 12.000 ;
    END
  END io_south_in[2]
  PIN io_south_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.290 8.000 40.570 12.000 ;
    END
  END io_south_in[30]
  PIN io_south_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.510 8.000 43.790 12.000 ;
    END
  END io_south_in[31]
  PIN io_south_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 172.310 8.000 172.590 12.000 ;
    END
  END io_south_in[3]
  PIN io_south_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 175.530 8.000 175.810 12.000 ;
    END
  END io_south_in[4]
  PIN io_south_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 181.970 8.000 182.250 12.000 ;
    END
  END io_south_in[5]
  PIN io_south_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 188.410 8.000 188.690 12.000 ;
    END
  END io_south_in[6]
  PIN io_south_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 194.850 8.000 195.130 12.000 ;
    END
  END io_south_in[7]
  PIN io_south_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 198.070 8.000 198.350 12.000 ;
    END
  END io_south_in[8]
  PIN io_south_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 204.510 8.000 204.790 12.000 ;
    END
  END io_south_in[9]
  PIN io_south_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 78.930 8.000 79.210 12.000 ;
    END
  END io_south_out[0]
  PIN io_south_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 133.670 8.000 133.950 12.000 ;
    END
  END io_south_out[10]
  PIN io_south_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 136.890 8.000 137.170 12.000 ;
    END
  END io_south_out[11]
  PIN io_south_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 143.330 8.000 143.610 12.000 ;
    END
  END io_south_out[12]
  PIN io_south_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 149.770 8.000 150.050 12.000 ;
    END
  END io_south_out[13]
  PIN io_south_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 457.000 242.640 461.000 243.240 ;
    END
  END io_south_out[14]
  PIN io_south_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 8.000 212.040 12.000 212.640 ;
    END
  END io_south_out[15]
  PIN io_south_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 262.470 8.000 262.750 12.000 ;
    END
  END io_south_out[16]
  PIN io_south_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 268.910 8.000 269.190 12.000 ;
    END
  END io_south_out[17]
  PIN io_south_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 272.130 8.000 272.410 12.000 ;
    END
  END io_south_out[18]
  PIN io_south_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 278.570 8.000 278.850 12.000 ;
    END
  END io_south_out[19]
  PIN io_south_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 82.150 8.000 82.430 12.000 ;
    END
  END io_south_out[1]
  PIN io_south_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 285.010 8.000 285.290 12.000 ;
    END
  END io_south_out[20]
  PIN io_south_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 291.450 8.000 291.730 12.000 ;
    END
  END io_south_out[21]
  PIN io_south_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 294.670 8.000 294.950 12.000 ;
    END
  END io_south_out[22]
  PIN io_south_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 301.110 8.000 301.390 12.000 ;
    END
  END io_south_out[23]
  PIN io_south_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 307.550 8.000 307.830 12.000 ;
    END
  END io_south_out[24]
  PIN io_south_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 310.770 8.000 311.050 12.000 ;
    END
  END io_south_out[25]
  PIN io_south_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 317.210 8.000 317.490 12.000 ;
    END
  END io_south_out[26]
  PIN io_south_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 323.650 8.000 323.930 12.000 ;
    END
  END io_south_out[27]
  PIN io_south_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 330.090 8.000 330.370 12.000 ;
    END
  END io_south_out[28]
  PIN io_south_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 333.310 8.000 333.590 12.000 ;
    END
  END io_south_out[29]
  PIN io_south_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 88.590 8.000 88.870 12.000 ;
    END
  END io_south_out[2]
  PIN io_south_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 457.000 246.040 461.000 246.640 ;
    END
  END io_south_out[30]
  PIN io_south_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 457.000 263.040 461.000 263.640 ;
    END
  END io_south_out[31]
  PIN io_south_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 95.030 8.000 95.310 12.000 ;
    END
  END io_south_out[3]
  PIN io_south_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 98.250 8.000 98.530 12.000 ;
    END
  END io_south_out[4]
  PIN io_south_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 104.690 8.000 104.970 12.000 ;
    END
  END io_south_out[5]
  PIN io_south_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 111.130 8.000 111.410 12.000 ;
    END
  END io_south_out[6]
  PIN io_south_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 117.570 8.000 117.850 12.000 ;
    END
  END io_south_out[7]
  PIN io_south_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 120.790 8.000 121.070 12.000 ;
    END
  END io_south_out[8]
  PIN io_south_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 127.230 8.000 127.510 12.000 ;
    END
  END io_south_out[9]
  PIN io_west_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 69.240 12.000 69.840 ;
    END
  END io_west_in[0]
  PIN io_west_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 123.640 12.000 124.240 ;
    END
  END io_west_in[10]
  PIN io_west_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 127.040 12.000 127.640 ;
    END
  END io_west_in[11]
  PIN io_west_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 133.840 12.000 134.440 ;
    END
  END io_west_in[12]
  PIN io_west_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 137.240 12.000 137.840 ;
    END
  END io_west_in[13]
  PIN io_west_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.730 8.000 47.010 12.000 ;
    END
  END io_west_in[14]
  PIN io_west_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.950 8.000 50.230 12.000 ;
    END
  END io_west_in[15]
  PIN io_west_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 256.240 12.000 256.840 ;
    END
  END io_west_in[16]
  PIN io_west_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 259.640 12.000 260.240 ;
    END
  END io_west_in[17]
  PIN io_west_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 263.040 12.000 263.640 ;
    END
  END io_west_in[18]
  PIN io_west_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 266.440 12.000 267.040 ;
    END
  END io_west_in[19]
  PIN io_west_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 72.640 12.000 73.240 ;
    END
  END io_west_in[1]
  PIN io_west_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 276.640 12.000 277.240 ;
    END
  END io_west_in[20]
  PIN io_west_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 283.440 12.000 284.040 ;
    END
  END io_west_in[21]
  PIN io_west_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 286.840 12.000 287.440 ;
    END
  END io_west_in[22]
  PIN io_west_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 293.640 12.000 294.240 ;
    END
  END io_west_in[23]
  PIN io_west_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 297.040 12.000 297.640 ;
    END
  END io_west_in[24]
  PIN io_west_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 303.840 12.000 304.440 ;
    END
  END io_west_in[25]
  PIN io_west_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 310.640 12.000 311.240 ;
    END
  END io_west_in[26]
  PIN io_west_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 314.040 12.000 314.640 ;
    END
  END io_west_in[27]
  PIN io_west_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 320.840 12.000 321.440 ;
    END
  END io_west_in[28]
  PIN io_west_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 324.240 12.000 324.840 ;
    END
  END io_west_in[29]
  PIN io_west_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 79.440 12.000 80.040 ;
    END
  END io_west_in[2]
  PIN io_west_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.170 8.000 53.450 12.000 ;
    END
  END io_west_in[30]
  PIN io_west_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.390 8.000 56.670 12.000 ;
    END
  END io_west_in[31]
  PIN io_west_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 82.840 12.000 83.440 ;
    END
  END io_west_in[3]
  PIN io_west_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 89.640 12.000 90.240 ;
    END
  END io_west_in[4]
  PIN io_west_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 96.440 12.000 97.040 ;
    END
  END io_west_in[5]
  PIN io_west_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 99.840 12.000 100.440 ;
    END
  END io_west_in[6]
  PIN io_west_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 106.640 12.000 107.240 ;
    END
  END io_west_in[7]
  PIN io_west_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 110.040 12.000 110.640 ;
    END
  END io_west_in[8]
  PIN io_west_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 116.840 12.000 117.440 ;
    END
  END io_west_in[9]
  PIN io_west_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 144.040 12.000 144.640 ;
    END
  END io_west_out[0]
  PIN io_west_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 198.440 12.000 199.040 ;
    END
  END io_west_out[10]
  PIN io_west_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 205.240 12.000 205.840 ;
    END
  END io_west_out[11]
  PIN io_west_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 208.640 12.000 209.240 ;
    END
  END io_west_out[12]
  PIN io_west_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 215.440 12.000 216.040 ;
    END
  END io_west_out[13]
  PIN io_west_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.490 459.000 233.770 463.000 ;
    END
  END io_west_out[14]
  PIN io_west_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 8.000 269.840 12.000 270.440 ;
    END
  END io_west_out[15]
  PIN io_west_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 331.040 12.000 331.640 ;
    END
  END io_west_out[16]
  PIN io_west_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 337.840 12.000 338.440 ;
    END
  END io_west_out[17]
  PIN io_west_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 341.240 12.000 341.840 ;
    END
  END io_west_out[18]
  PIN io_west_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 348.040 12.000 348.640 ;
    END
  END io_west_out[19]
  PIN io_west_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 150.840 12.000 151.440 ;
    END
  END io_west_out[1]
  PIN io_west_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 351.440 12.000 352.040 ;
    END
  END io_west_out[20]
  PIN io_west_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 358.240 12.000 358.840 ;
    END
  END io_west_out[21]
  PIN io_west_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 365.040 12.000 365.640 ;
    END
  END io_west_out[22]
  PIN io_west_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 368.440 12.000 369.040 ;
    END
  END io_west_out[23]
  PIN io_west_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 375.240 12.000 375.840 ;
    END
  END io_west_out[24]
  PIN io_west_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 378.640 12.000 379.240 ;
    END
  END io_west_out[25]
  PIN io_west_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 385.440 12.000 386.040 ;
    END
  END io_west_out[26]
  PIN io_west_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 392.240 12.000 392.840 ;
    END
  END io_west_out[27]
  PIN io_west_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 395.640 12.000 396.240 ;
    END
  END io_west_out[28]
  PIN io_west_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 402.440 12.000 403.040 ;
    END
  END io_west_out[29]
  PIN io_west_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 154.240 12.000 154.840 ;
    END
  END io_west_out[2]
  PIN io_west_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 8.000 273.240 12.000 273.840 ;
    END
  END io_west_out[30]
  PIN io_west_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 8.000 218.840 12.000 219.440 ;
    END
  END io_west_out[31]
  PIN io_west_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 161.040 12.000 161.640 ;
    END
  END io_west_out[3]
  PIN io_west_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 164.440 12.000 165.040 ;
    END
  END io_west_out[4]
  PIN io_west_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 171.240 12.000 171.840 ;
    END
  END io_west_out[5]
  PIN io_west_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 178.040 12.000 178.640 ;
    END
  END io_west_out[6]
  PIN io_west_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 181.440 12.000 182.040 ;
    END
  END io_west_out[7]
  PIN io_west_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 188.240 12.000 188.840 ;
    END
  END io_west_out[8]
  PIN io_west_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 191.640 12.000 192.240 ;
    END
  END io_west_out[9]
  PIN le_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 62.830 8.000 63.110 12.000 ;
    END
  END le_clk
  PIN le_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 69.270 8.000 69.550 12.000 ;
    END
  END le_en
  PIN le_nrst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 72.490 8.000 72.770 12.000 ;
    END
  END le_nrst
  PIN nrst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 243.150 459.000 243.430 463.000 ;
    END
  END nrst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 16.780 16.880 18.380 453.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 16.780 16.880 452.420 18.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 16.780 452.080 452.420 453.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 450.820 16.880 452.420 453.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 93.580 13.580 95.180 44.635 ;
    END
    PORT
      LAYER met4 ;
        RECT 93.580 428.005 95.180 456.980 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.580 13.580 190.180 44.635 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.580 428.005 190.180 456.980 ;
    END
    PORT
      LAYER met4 ;
        RECT 283.580 13.580 285.180 44.635 ;
    END
    PORT
      LAYER met4 ;
        RECT 283.580 428.005 285.180 456.980 ;
    END
    PORT
      LAYER met4 ;
        RECT 378.580 13.580 380.180 44.635 ;
    END
    PORT
      LAYER met4 ;
        RECT 378.580 428.005 380.180 456.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 13.480 93.680 455.720 95.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 13.480 188.680 455.720 190.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 13.480 283.680 455.720 285.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 13.480 378.680 455.720 380.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 29.740 35.120 31.340 435.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 435.460 35.120 437.060 435.440 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 13.480 13.580 15.080 456.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 13.480 13.580 455.720 15.180 ;
    END
    PORT
      LAYER met5 ;
        RECT 13.480 455.380 455.720 456.980 ;
    END
    PORT
      LAYER met4 ;
        RECT 454.120 13.580 455.720 456.980 ;
    END
    PORT
      LAYER met4 ;
        RECT 96.880 13.580 98.480 44.635 ;
    END
    PORT
      LAYER met4 ;
        RECT 96.880 428.005 98.480 456.980 ;
    END
    PORT
      LAYER met4 ;
        RECT 191.880 13.580 193.480 44.635 ;
    END
    PORT
      LAYER met4 ;
        RECT 191.880 428.005 193.480 456.980 ;
    END
    PORT
      LAYER met4 ;
        RECT 286.880 13.580 288.480 44.635 ;
    END
    PORT
      LAYER met4 ;
        RECT 286.880 428.005 288.480 456.980 ;
    END
    PORT
      LAYER met4 ;
        RECT 381.880 13.580 383.480 44.635 ;
    END
    PORT
      LAYER met4 ;
        RECT 381.880 428.005 383.480 456.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 13.480 96.980 455.720 98.580 ;
    END
    PORT
      LAYER met5 ;
        RECT 13.480 191.980 455.720 193.580 ;
    END
    PORT
      LAYER met5 ;
        RECT 13.480 286.980 455.720 288.580 ;
    END
    PORT
      LAYER met5 ;
        RECT 13.480 381.980 455.720 383.580 ;
    END
    PORT
      LAYER met4 ;
        RECT 33.420 35.120 35.020 435.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 439.140 35.120 440.740 435.440 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 24.190 24.395 445.010 446.270 ;
      LAYER li1 ;
        RECT 24.380 24.395 444.820 446.165 ;
      LAYER met1 ;
        RECT 12.670 24.240 450.910 446.320 ;
      LAYER met2 ;
        RECT 12.690 458.720 78.650 459.000 ;
        RECT 79.490 458.720 81.870 459.000 ;
        RECT 82.710 458.720 88.310 459.000 ;
        RECT 89.150 458.720 94.750 459.000 ;
        RECT 95.590 458.720 97.970 459.000 ;
        RECT 98.810 458.720 104.410 459.000 ;
        RECT 105.250 458.720 110.850 459.000 ;
        RECT 111.690 458.720 117.290 459.000 ;
        RECT 118.130 458.720 120.510 459.000 ;
        RECT 121.350 458.720 126.950 459.000 ;
        RECT 127.790 458.720 133.390 459.000 ;
        RECT 134.230 458.720 136.610 459.000 ;
        RECT 137.450 458.720 143.050 459.000 ;
        RECT 143.890 458.720 149.490 459.000 ;
        RECT 150.330 458.720 155.930 459.000 ;
        RECT 156.770 458.720 159.150 459.000 ;
        RECT 159.990 458.720 165.590 459.000 ;
        RECT 166.430 458.720 172.030 459.000 ;
        RECT 172.870 458.720 175.250 459.000 ;
        RECT 176.090 458.720 181.690 459.000 ;
        RECT 182.530 458.720 188.130 459.000 ;
        RECT 188.970 458.720 194.570 459.000 ;
        RECT 195.410 458.720 197.790 459.000 ;
        RECT 198.630 458.720 204.230 459.000 ;
        RECT 205.070 458.720 210.670 459.000 ;
        RECT 211.510 458.720 213.890 459.000 ;
        RECT 214.730 458.720 220.330 459.000 ;
        RECT 221.170 458.720 226.770 459.000 ;
        RECT 227.610 458.720 233.210 459.000 ;
        RECT 234.050 458.720 239.650 459.000 ;
        RECT 240.490 458.720 242.870 459.000 ;
        RECT 243.710 458.720 249.310 459.000 ;
        RECT 250.150 458.720 262.190 459.000 ;
        RECT 263.030 458.720 268.630 459.000 ;
        RECT 269.470 458.720 271.850 459.000 ;
        RECT 272.690 458.720 278.290 459.000 ;
        RECT 279.130 458.720 281.510 459.000 ;
        RECT 282.350 458.720 284.730 459.000 ;
        RECT 285.570 458.720 287.950 459.000 ;
        RECT 288.790 458.720 291.170 459.000 ;
        RECT 292.010 458.720 294.390 459.000 ;
        RECT 295.230 458.720 300.830 459.000 ;
        RECT 301.670 458.720 307.270 459.000 ;
        RECT 308.110 458.720 310.490 459.000 ;
        RECT 311.330 458.720 316.930 459.000 ;
        RECT 317.770 458.720 323.370 459.000 ;
        RECT 324.210 458.720 329.810 459.000 ;
        RECT 330.650 458.720 333.030 459.000 ;
        RECT 333.870 458.720 339.470 459.000 ;
        RECT 340.310 458.720 345.910 459.000 ;
        RECT 346.750 458.720 349.130 459.000 ;
        RECT 349.970 458.720 355.570 459.000 ;
        RECT 356.410 458.720 362.010 459.000 ;
        RECT 362.850 458.720 368.450 459.000 ;
        RECT 369.290 458.720 371.670 459.000 ;
        RECT 372.510 458.720 378.110 459.000 ;
        RECT 378.950 458.720 384.550 459.000 ;
        RECT 385.390 458.720 387.770 459.000 ;
        RECT 388.610 458.720 394.210 459.000 ;
        RECT 395.050 458.720 400.650 459.000 ;
        RECT 401.490 458.720 407.090 459.000 ;
        RECT 407.930 458.720 410.310 459.000 ;
        RECT 411.150 458.720 450.890 459.000 ;
        RECT 12.690 12.280 450.890 458.720 ;
        RECT 12.690 12.000 14.250 12.280 ;
        RECT 15.090 12.000 17.470 12.280 ;
        RECT 18.310 12.000 20.690 12.280 ;
        RECT 21.530 12.000 23.910 12.280 ;
        RECT 24.750 12.000 27.130 12.280 ;
        RECT 27.970 12.000 30.350 12.280 ;
        RECT 31.190 12.000 33.570 12.280 ;
        RECT 34.410 12.000 36.790 12.280 ;
        RECT 37.630 12.000 40.010 12.280 ;
        RECT 40.850 12.000 43.230 12.280 ;
        RECT 44.070 12.000 46.450 12.280 ;
        RECT 47.290 12.000 49.670 12.280 ;
        RECT 50.510 12.000 52.890 12.280 ;
        RECT 53.730 12.000 56.110 12.280 ;
        RECT 56.950 12.000 62.550 12.280 ;
        RECT 63.390 12.000 68.990 12.280 ;
        RECT 69.830 12.000 72.210 12.280 ;
        RECT 73.050 12.000 78.650 12.280 ;
        RECT 79.490 12.000 81.870 12.280 ;
        RECT 82.710 12.000 88.310 12.280 ;
        RECT 89.150 12.000 94.750 12.280 ;
        RECT 95.590 12.000 97.970 12.280 ;
        RECT 98.810 12.000 104.410 12.280 ;
        RECT 105.250 12.000 110.850 12.280 ;
        RECT 111.690 12.000 117.290 12.280 ;
        RECT 118.130 12.000 120.510 12.280 ;
        RECT 121.350 12.000 126.950 12.280 ;
        RECT 127.790 12.000 133.390 12.280 ;
        RECT 134.230 12.000 136.610 12.280 ;
        RECT 137.450 12.000 143.050 12.280 ;
        RECT 143.890 12.000 149.490 12.280 ;
        RECT 150.330 12.000 155.930 12.280 ;
        RECT 156.770 12.000 159.150 12.280 ;
        RECT 159.990 12.000 165.590 12.280 ;
        RECT 166.430 12.000 172.030 12.280 ;
        RECT 172.870 12.000 175.250 12.280 ;
        RECT 176.090 12.000 181.690 12.280 ;
        RECT 182.530 12.000 188.130 12.280 ;
        RECT 188.970 12.000 194.570 12.280 ;
        RECT 195.410 12.000 197.790 12.280 ;
        RECT 198.630 12.000 204.230 12.280 ;
        RECT 205.070 12.000 210.670 12.280 ;
        RECT 211.510 12.000 213.890 12.280 ;
        RECT 214.730 12.000 220.330 12.280 ;
        RECT 221.170 12.000 226.770 12.280 ;
        RECT 227.610 12.000 262.190 12.280 ;
        RECT 263.030 12.000 268.630 12.280 ;
        RECT 269.470 12.000 271.850 12.280 ;
        RECT 272.690 12.000 278.290 12.280 ;
        RECT 279.130 12.000 284.730 12.280 ;
        RECT 285.570 12.000 291.170 12.280 ;
        RECT 292.010 12.000 294.390 12.280 ;
        RECT 295.230 12.000 300.830 12.280 ;
        RECT 301.670 12.000 307.270 12.280 ;
        RECT 308.110 12.000 310.490 12.280 ;
        RECT 311.330 12.000 316.930 12.280 ;
        RECT 317.770 12.000 323.370 12.280 ;
        RECT 324.210 12.000 329.810 12.280 ;
        RECT 330.650 12.000 333.030 12.280 ;
        RECT 333.870 12.000 339.470 12.280 ;
        RECT 340.310 12.000 345.910 12.280 ;
        RECT 346.750 12.000 349.130 12.280 ;
        RECT 349.970 12.000 355.570 12.280 ;
        RECT 356.410 12.000 362.010 12.280 ;
        RECT 362.850 12.000 368.450 12.280 ;
        RECT 369.290 12.000 371.670 12.280 ;
        RECT 372.510 12.000 378.110 12.280 ;
        RECT 378.950 12.000 384.550 12.280 ;
        RECT 385.390 12.000 387.770 12.280 ;
        RECT 388.610 12.000 394.210 12.280 ;
        RECT 395.050 12.000 400.650 12.280 ;
        RECT 401.490 12.000 407.090 12.280 ;
        RECT 407.930 12.000 410.310 12.280 ;
        RECT 411.150 12.000 450.890 12.280 ;
      LAYER met3 ;
        RECT 12.000 403.440 457.000 446.245 ;
        RECT 12.400 402.040 456.600 403.440 ;
        RECT 12.000 396.640 457.000 402.040 ;
        RECT 12.400 395.240 456.600 396.640 ;
        RECT 12.000 393.240 457.000 395.240 ;
        RECT 12.400 391.840 456.600 393.240 ;
        RECT 12.000 386.440 457.000 391.840 ;
        RECT 12.400 385.040 456.600 386.440 ;
        RECT 12.000 379.640 457.000 385.040 ;
        RECT 12.400 378.240 456.600 379.640 ;
        RECT 12.000 376.240 457.000 378.240 ;
        RECT 12.400 374.840 456.600 376.240 ;
        RECT 12.000 369.440 457.000 374.840 ;
        RECT 12.400 368.040 456.600 369.440 ;
        RECT 12.000 366.040 457.000 368.040 ;
        RECT 12.400 364.640 456.600 366.040 ;
        RECT 12.000 359.240 457.000 364.640 ;
        RECT 12.400 357.840 456.600 359.240 ;
        RECT 12.000 352.440 457.000 357.840 ;
        RECT 12.400 351.040 456.600 352.440 ;
        RECT 12.000 349.040 457.000 351.040 ;
        RECT 12.400 347.640 456.600 349.040 ;
        RECT 12.000 345.640 457.000 347.640 ;
        RECT 12.000 344.240 456.600 345.640 ;
        RECT 12.000 342.240 457.000 344.240 ;
        RECT 12.400 340.840 456.600 342.240 ;
        RECT 12.000 338.840 457.000 340.840 ;
        RECT 12.400 337.440 456.600 338.840 ;
        RECT 12.000 332.040 457.000 337.440 ;
        RECT 12.400 330.640 456.600 332.040 ;
        RECT 12.000 325.240 457.000 330.640 ;
        RECT 12.400 323.840 456.600 325.240 ;
        RECT 12.000 321.840 457.000 323.840 ;
        RECT 12.400 320.440 456.600 321.840 ;
        RECT 12.000 315.040 457.000 320.440 ;
        RECT 12.400 313.640 456.600 315.040 ;
        RECT 12.000 311.640 457.000 313.640 ;
        RECT 12.400 310.240 456.600 311.640 ;
        RECT 12.000 304.840 457.000 310.240 ;
        RECT 12.400 303.440 456.600 304.840 ;
        RECT 12.000 298.040 457.000 303.440 ;
        RECT 12.400 296.640 456.600 298.040 ;
        RECT 12.000 294.640 457.000 296.640 ;
        RECT 12.400 293.240 456.600 294.640 ;
        RECT 12.000 287.840 457.000 293.240 ;
        RECT 12.400 286.440 456.600 287.840 ;
        RECT 12.000 284.440 457.000 286.440 ;
        RECT 12.400 283.040 456.600 284.440 ;
        RECT 12.000 277.640 457.000 283.040 ;
        RECT 12.400 276.240 456.600 277.640 ;
        RECT 12.000 274.240 457.000 276.240 ;
        RECT 12.400 272.840 457.000 274.240 ;
        RECT 12.000 270.840 457.000 272.840 ;
        RECT 12.400 269.440 456.600 270.840 ;
        RECT 12.000 267.440 457.000 269.440 ;
        RECT 12.400 266.040 456.600 267.440 ;
        RECT 12.000 264.040 457.000 266.040 ;
        RECT 12.400 262.640 456.600 264.040 ;
        RECT 12.000 260.640 457.000 262.640 ;
        RECT 12.400 259.240 456.600 260.640 ;
        RECT 12.000 257.240 457.000 259.240 ;
        RECT 12.400 255.840 456.600 257.240 ;
        RECT 12.000 247.040 457.000 255.840 ;
        RECT 12.400 245.640 456.600 247.040 ;
        RECT 12.000 243.640 457.000 245.640 ;
        RECT 12.000 242.240 456.600 243.640 ;
        RECT 12.000 240.240 457.000 242.240 ;
        RECT 12.000 238.840 456.600 240.240 ;
        RECT 12.000 233.440 457.000 238.840 ;
        RECT 12.400 232.040 456.600 233.440 ;
        RECT 12.000 230.040 457.000 232.040 ;
        RECT 12.400 228.640 457.000 230.040 ;
        RECT 12.000 223.240 457.000 228.640 ;
        RECT 12.400 221.840 457.000 223.240 ;
        RECT 12.000 219.840 457.000 221.840 ;
        RECT 12.400 218.440 457.000 219.840 ;
        RECT 12.000 216.440 457.000 218.440 ;
        RECT 12.400 215.040 456.600 216.440 ;
        RECT 12.000 213.040 457.000 215.040 ;
        RECT 12.400 211.640 457.000 213.040 ;
        RECT 12.000 209.640 457.000 211.640 ;
        RECT 12.400 208.240 456.600 209.640 ;
        RECT 12.000 206.240 457.000 208.240 ;
        RECT 12.400 204.840 456.600 206.240 ;
        RECT 12.000 199.440 457.000 204.840 ;
        RECT 12.400 198.040 456.600 199.440 ;
        RECT 12.000 192.640 457.000 198.040 ;
        RECT 12.400 191.240 456.600 192.640 ;
        RECT 12.000 189.240 457.000 191.240 ;
        RECT 12.400 187.840 456.600 189.240 ;
        RECT 12.000 182.440 457.000 187.840 ;
        RECT 12.400 181.040 456.600 182.440 ;
        RECT 12.000 179.040 457.000 181.040 ;
        RECT 12.400 177.640 456.600 179.040 ;
        RECT 12.000 172.240 457.000 177.640 ;
        RECT 12.400 170.840 456.600 172.240 ;
        RECT 12.000 168.840 457.000 170.840 ;
        RECT 12.400 167.440 457.000 168.840 ;
        RECT 12.000 165.440 457.000 167.440 ;
        RECT 12.400 164.040 456.600 165.440 ;
        RECT 12.000 162.040 457.000 164.040 ;
        RECT 12.400 160.640 456.600 162.040 ;
        RECT 12.000 155.240 457.000 160.640 ;
        RECT 12.400 153.840 456.600 155.240 ;
        RECT 12.000 151.840 457.000 153.840 ;
        RECT 12.400 150.440 456.600 151.840 ;
        RECT 12.000 145.040 457.000 150.440 ;
        RECT 12.400 143.640 456.600 145.040 ;
        RECT 12.000 138.240 457.000 143.640 ;
        RECT 12.400 136.840 456.600 138.240 ;
        RECT 12.000 134.840 457.000 136.840 ;
        RECT 12.400 133.440 456.600 134.840 ;
        RECT 12.000 128.040 457.000 133.440 ;
        RECT 12.400 126.640 456.600 128.040 ;
        RECT 12.000 124.640 457.000 126.640 ;
        RECT 12.400 123.240 456.600 124.640 ;
        RECT 12.000 117.840 457.000 123.240 ;
        RECT 12.400 116.440 456.600 117.840 ;
        RECT 12.000 111.040 457.000 116.440 ;
        RECT 12.400 109.640 456.600 111.040 ;
        RECT 12.000 107.640 457.000 109.640 ;
        RECT 12.400 106.240 456.600 107.640 ;
        RECT 12.000 100.840 457.000 106.240 ;
        RECT 12.400 99.440 456.600 100.840 ;
        RECT 12.000 97.440 457.000 99.440 ;
        RECT 12.400 96.040 456.600 97.440 ;
        RECT 12.000 90.640 457.000 96.040 ;
        RECT 12.400 89.240 456.600 90.640 ;
        RECT 12.000 83.840 457.000 89.240 ;
        RECT 12.400 82.440 456.600 83.840 ;
        RECT 12.000 80.440 457.000 82.440 ;
        RECT 12.400 79.040 456.600 80.440 ;
        RECT 12.000 73.640 457.000 79.040 ;
        RECT 12.400 72.240 456.600 73.640 ;
        RECT 12.000 70.240 457.000 72.240 ;
        RECT 12.400 68.840 456.600 70.240 ;
        RECT 12.000 24.315 457.000 68.840 ;
      LAYER met4 ;
        RECT 51.215 54.640 412.320 417.705 ;
      LAYER met5 ;
        RECT 52.420 385.180 416.940 416.540 ;
        RECT 52.420 290.180 416.940 377.080 ;
        RECT 52.420 195.180 416.940 282.080 ;
        RECT 52.420 100.180 416.940 187.080 ;
        RECT 52.420 54.640 416.940 92.080 ;
  END
END fpga
END LIBRARY

