VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO outel8227
  CLASS BLOCK ;
  FOREIGN outel8227 ;
  ORIGIN 0.000 0.000 ;
  SIZE 188.475 BY 199.195 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 187.920 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 187.920 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END clk
  PIN cs
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END cs
  PIN dataBusIn[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 184.475 119.040 188.475 119.640 ;
    END
  END dataBusIn[0]
  PIN dataBusIn[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 184.475 125.840 188.475 126.440 ;
    END
  END dataBusIn[1]
  PIN dataBusIn[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 184.475 132.640 188.475 133.240 ;
    END
  END dataBusIn[2]
  PIN dataBusIn[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 184.475 136.040 188.475 136.640 ;
    END
  END dataBusIn[3]
  PIN dataBusIn[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 184.475 112.240 188.475 112.840 ;
    END
  END dataBusIn[4]
  PIN dataBusIn[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 184.475 115.640 188.475 116.240 ;
    END
  END dataBusIn[5]
  PIN dataBusIn[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 184.475 129.240 188.475 129.840 ;
    END
  END dataBusIn[6]
  PIN dataBusIn[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 184.475 122.440 188.475 123.040 ;
    END
  END dataBusIn[7]
  PIN dataBusOut[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END dataBusOut[0]
  PIN dataBusOut[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END dataBusOut[1]
  PIN dataBusOut[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END dataBusOut[2]
  PIN dataBusOut[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END dataBusOut[3]
  PIN dataBusOut[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END dataBusOut[4]
  PIN dataBusOut[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END dataBusOut[5]
  PIN dataBusOut[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END dataBusOut[6]
  PIN dataBusOut[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END dataBusOut[7]
  PIN dataBusSelect
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END dataBusSelect
  PIN gpio[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 64.490 195.195 64.770 199.195 ;
    END
  END gpio[0]
  PIN gpio[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 61.270 195.195 61.550 199.195 ;
    END
  END gpio[10]
  PIN gpio[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 41.950 195.195 42.230 199.195 ;
    END
  END gpio[11]
  PIN gpio[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 54.830 195.195 55.110 199.195 ;
    END
  END gpio[12]
  PIN gpio[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 48.390 195.195 48.670 199.195 ;
    END
  END gpio[13]
  PIN gpio[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 29.070 195.195 29.350 199.195 ;
    END
  END gpio[14]
  PIN gpio[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 32.290 195.195 32.570 199.195 ;
    END
  END gpio[15]
  PIN gpio[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END gpio[16]
  PIN gpio[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END gpio[17]
  PIN gpio[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END gpio[18]
  PIN gpio[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER met3 ;
        RECT 184.475 105.440 188.475 106.040 ;
    END
  END gpio[19]
  PIN gpio[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 45.170 195.195 45.450 199.195 ;
    END
  END gpio[1]
  PIN gpio[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.621000 ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END gpio[20]
  PIN gpio[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.120500 ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 184.475 102.040 188.475 102.640 ;
    END
  END gpio[21]
  PIN gpio[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.237500 ;
    ANTENNADIFFAREA 1.075200 ;
    PORT
      LAYER met3 ;
        RECT 184.475 108.840 188.475 109.440 ;
    END
  END gpio[22]
  PIN gpio[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END gpio[23]
  PIN gpio[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 4.000 ;
    END
  END gpio[24]
  PIN gpio[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END gpio[25]
  PIN gpio[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 106.350 195.195 106.630 199.195 ;
    END
  END gpio[2]
  PIN gpio[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 51.610 195.195 51.890 199.195 ;
    END
  END gpio[3]
  PIN gpio[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END gpio[4]
  PIN gpio[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END gpio[5]
  PIN gpio[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 38.730 195.195 39.010 199.195 ;
    END
  END gpio[6]
  PIN gpio[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END gpio[7]
  PIN gpio[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 58.050 195.195 58.330 199.195 ;
    END
  END gpio[8]
  PIN gpio[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 35.510 195.195 35.790 199.195 ;
    END
  END gpio[9]
  PIN nrst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 184.475 17.040 188.475 17.640 ;
    END
  END nrst
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 182.810 187.870 ;
      LAYER li1 ;
        RECT 5.520 10.795 182.620 187.765 ;
      LAYER met1 ;
        RECT 4.670 10.640 183.930 187.920 ;
      LAYER met2 ;
        RECT 4.690 194.915 28.790 195.570 ;
        RECT 29.630 194.915 32.010 195.570 ;
        RECT 32.850 194.915 35.230 195.570 ;
        RECT 36.070 194.915 38.450 195.570 ;
        RECT 39.290 194.915 41.670 195.570 ;
        RECT 42.510 194.915 44.890 195.570 ;
        RECT 45.730 194.915 48.110 195.570 ;
        RECT 48.950 194.915 51.330 195.570 ;
        RECT 52.170 194.915 54.550 195.570 ;
        RECT 55.390 194.915 57.770 195.570 ;
        RECT 58.610 194.915 60.990 195.570 ;
        RECT 61.830 194.915 64.210 195.570 ;
        RECT 65.050 194.915 106.070 195.570 ;
        RECT 106.910 194.915 183.910 195.570 ;
        RECT 4.690 4.280 183.910 194.915 ;
        RECT 4.690 4.000 57.770 4.280 ;
        RECT 58.610 4.000 60.990 4.280 ;
        RECT 61.830 4.000 64.210 4.280 ;
        RECT 65.050 4.000 67.430 4.280 ;
        RECT 68.270 4.000 70.650 4.280 ;
        RECT 71.490 4.000 73.870 4.280 ;
        RECT 74.710 4.000 77.090 4.280 ;
        RECT 77.930 4.000 80.310 4.280 ;
        RECT 81.150 4.000 83.530 4.280 ;
        RECT 84.370 4.000 86.750 4.280 ;
        RECT 87.590 4.000 93.190 4.280 ;
        RECT 94.030 4.000 118.950 4.280 ;
        RECT 119.790 4.000 122.170 4.280 ;
        RECT 123.010 4.000 125.390 4.280 ;
        RECT 126.230 4.000 183.910 4.280 ;
      LAYER met3 ;
        RECT 3.070 181.240 185.570 187.845 ;
        RECT 4.400 179.840 185.570 181.240 ;
        RECT 3.070 157.440 185.570 179.840 ;
        RECT 4.400 156.040 185.570 157.440 ;
        RECT 3.070 154.040 185.570 156.040 ;
        RECT 4.400 152.640 185.570 154.040 ;
        RECT 3.070 147.240 185.570 152.640 ;
        RECT 4.400 145.840 185.570 147.240 ;
        RECT 3.070 137.040 185.570 145.840 ;
        RECT 3.070 135.640 184.075 137.040 ;
        RECT 3.070 133.640 185.570 135.640 ;
        RECT 3.070 132.240 184.075 133.640 ;
        RECT 3.070 130.240 185.570 132.240 ;
        RECT 3.070 128.840 184.075 130.240 ;
        RECT 3.070 126.840 185.570 128.840 ;
        RECT 3.070 125.440 184.075 126.840 ;
        RECT 3.070 123.440 185.570 125.440 ;
        RECT 3.070 122.040 184.075 123.440 ;
        RECT 3.070 120.040 185.570 122.040 ;
        RECT 3.070 118.640 184.075 120.040 ;
        RECT 3.070 116.640 185.570 118.640 ;
        RECT 3.070 115.240 184.075 116.640 ;
        RECT 3.070 113.240 185.570 115.240 ;
        RECT 3.070 111.840 184.075 113.240 ;
        RECT 3.070 109.840 185.570 111.840 ;
        RECT 3.070 108.440 184.075 109.840 ;
        RECT 3.070 106.440 185.570 108.440 ;
        RECT 3.070 105.040 184.075 106.440 ;
        RECT 3.070 103.040 185.570 105.040 ;
        RECT 3.070 101.640 184.075 103.040 ;
        RECT 3.070 21.440 185.570 101.640 ;
        RECT 4.400 20.040 185.570 21.440 ;
        RECT 3.070 18.040 185.570 20.040 ;
        RECT 3.070 16.640 184.075 18.040 ;
        RECT 3.070 9.015 185.570 16.640 ;
      LAYER met4 ;
        RECT 23.295 26.695 23.940 177.985 ;
        RECT 26.340 26.695 174.240 177.985 ;
        RECT 176.640 26.695 177.540 177.985 ;
        RECT 179.940 26.695 185.545 177.985 ;
  END
END outel8227
END LIBRARY

