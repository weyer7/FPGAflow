VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fpga
  CLASS BLOCK ;
  FOREIGN fpga ;
  ORIGIN 0.000 0.000 ;
  SIZE 1200.000 BY 1200.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.540 10.640 333.140 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 485.140 10.640 486.740 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.740 10.640 640.340 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 792.340 10.640 793.940 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 945.940 10.640 947.540 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1099.540 10.640 1101.140 1188.880 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1188.880 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1156.040 4.000 1156.640 ;
    END
  END clk
  PIN config_data
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1149.240 4.000 1149.840 ;
    END
  END config_data
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1152.640 4.000 1153.240 ;
    END
  END en
  PIN io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1084.640 4.000 1085.240 ;
    END
  END io[0]
  PIN io[100]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 550.840 4.000 551.440 ;
    END
  END io[100]
  PIN io[101]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 853.440 4.000 854.040 ;
    END
  END io[101]
  PIN io[102]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 802.440 4.000 803.040 ;
    END
  END io[102]
  PIN io[103]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 873.840 4.000 874.440 ;
    END
  END io[103]
  PIN io[104]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 856.840 4.000 857.440 ;
    END
  END io[104]
  PIN io[105]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 561.040 4.000 561.640 ;
    END
  END io[105]
  PIN io[106]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 799.040 4.000 799.640 ;
    END
  END io[106]
  PIN io[107]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 618.840 4.000 619.440 ;
    END
  END io[107]
  PIN io[108]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 870.440 4.000 871.040 ;
    END
  END io[108]
  PIN io[109]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.953500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 826.240 4.000 826.840 ;
    END
  END io[109]
  PIN io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 975.840 4.000 976.440 ;
    END
  END io[10]
  PIN io[110]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 877.240 4.000 877.840 ;
    END
  END io[110]
  PIN io[111]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met2 ;
        RECT 370.390 1196.000 370.670 1200.000 ;
    END
  END io[111]
  PIN io[112]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met2 ;
        RECT 363.950 1196.000 364.230 1200.000 ;
    END
  END io[112]
  PIN io[113]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met2 ;
        RECT 412.250 1196.000 412.530 1200.000 ;
    END
  END io[113]
  PIN io[114]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met2 ;
        RECT 347.850 1196.000 348.130 1200.000 ;
    END
  END io[114]
  PIN io[115]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met2 ;
        RECT 415.470 1196.000 415.750 1200.000 ;
    END
  END io[115]
  PIN io[116]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met2 ;
        RECT 351.070 1196.000 351.350 1200.000 ;
    END
  END io[116]
  PIN io[117]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met2 ;
        RECT 389.710 1196.000 389.990 1200.000 ;
    END
  END io[117]
  PIN io[118]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met2 ;
        RECT 354.290 1196.000 354.570 1200.000 ;
    END
  END io[118]
  PIN io[119]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met2 ;
        RECT 325.310 1196.000 325.590 1200.000 ;
    END
  END io[119]
  PIN io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1074.440 4.000 1075.040 ;
    END
  END io[11]
  PIN io[120]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met2 ;
        RECT 305.990 1196.000 306.270 1200.000 ;
    END
  END io[120]
  PIN io[121]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met2 ;
        RECT 280.230 1196.000 280.510 1200.000 ;
    END
  END io[121]
  PIN io[122]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met2 ;
        RECT 251.250 1196.000 251.530 1200.000 ;
    END
  END io[122]
  PIN io[123]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met2 ;
        RECT 215.830 1196.000 216.110 1200.000 ;
    END
  END io[123]
  PIN io[124]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.953500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met2 ;
        RECT 212.610 1196.000 212.890 1200.000 ;
    END
  END io[124]
  PIN io[125]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.953500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met2 ;
        RECT 209.390 1196.000 209.670 1200.000 ;
    END
  END io[125]
  PIN io[126]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.953500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met2 ;
        RECT 180.410 1196.000 180.690 1200.000 ;
    END
  END io[126]
  PIN io[127]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met2 ;
        RECT 167.530 1196.000 167.810 1200.000 ;
    END
  END io[127]
  PIN io[128]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1050.640 4.000 1051.240 ;
    END
  END io[128]
  PIN io[129]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met2 ;
        RECT 170.750 1196.000 171.030 1200.000 ;
    END
  END io[129]
  PIN io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.000100 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 979.240 4.000 979.840 ;
    END
  END io[12]
  PIN io[130]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met2 ;
        RECT 183.630 1196.000 183.910 1200.000 ;
    END
  END io[130]
  PIN io[131]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1016.640 4.000 1017.240 ;
    END
  END io[131]
  PIN io[132]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.813000 ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1020.040 4.000 1020.640 ;
    END
  END io[132]
  PIN io[133]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1023.440 4.000 1024.040 ;
    END
  END io[133]
  PIN io[134]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1006.440 4.000 1007.040 ;
    END
  END io[134]
  PIN io[135]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 992.840 4.000 993.440 ;
    END
  END io[135]
  PIN io[136]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1026.840 4.000 1027.440 ;
    END
  END io[136]
  PIN io[137]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1077.840 4.000 1078.440 ;
    END
  END io[137]
  PIN io[138]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 938.440 4.000 939.040 ;
    END
  END io[138]
  PIN io[139]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 904.440 4.000 905.040 ;
    END
  END io[139]
  PIN io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.130600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1081.240 4.000 1081.840 ;
    END
  END io[13]
  PIN io[140]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1115.240 4.000 1115.840 ;
    END
  END io[140]
  PIN io[141]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.481500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 901.040 4.000 901.640 ;
    END
  END io[141]
  PIN io[142]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met2 ;
        RECT 302.770 1196.000 303.050 1200.000 ;
    END
  END io[142]
  PIN io[143]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met2 ;
        RECT 225.490 1196.000 225.770 1200.000 ;
    END
  END io[143]
  PIN io[144]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 822.840 4.000 823.440 ;
    END
  END io[144]
  PIN io[145]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 867.040 4.000 867.640 ;
    END
  END io[145]
  PIN io[146]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met2 ;
        RECT 264.130 1196.000 264.410 1200.000 ;
    END
  END io[146]
  PIN io[147]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1043.840 4.000 1044.440 ;
    END
  END io[147]
  PIN io[148]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1111.840 4.000 1112.440 ;
    END
  END io[148]
  PIN io[149]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1139.040 4.000 1139.640 ;
    END
  END io[149]
  PIN io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met2 ;
        RECT 190.070 1196.000 190.350 1200.000 ;
    END
  END io[14]
  PIN io[150]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 805.840 4.000 806.440 ;
    END
  END io[150]
  PIN io[151]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 768.440 4.000 769.040 ;
    END
  END io[151]
  PIN io[152]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 608.640 4.000 609.240 ;
    END
  END io[152]
  PIN io[153]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 554.240 4.000 554.840 ;
    END
  END io[153]
  PIN io[154]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 669.840 4.000 670.440 ;
    END
  END io[154]
  PIN io[155]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 693.640 4.000 694.240 ;
    END
  END io[155]
  PIN io[156]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 697.040 4.000 697.640 ;
    END
  END io[156]
  PIN io[157]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 567.840 4.000 568.440 ;
    END
  END io[157]
  PIN io[158]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 700.440 4.000 701.040 ;
    END
  END io[158]
  PIN io[159]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 666.440 4.000 667.040 ;
    END
  END io[159]
  PIN io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 955.440 4.000 956.040 ;
    END
  END io[15]
  PIN io[160]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 625.640 4.000 626.240 ;
    END
  END io[160]
  PIN io[161]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 792.240 4.000 792.840 ;
    END
  END io[161]
  PIN io[162]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 629.040 4.000 629.640 ;
    END
  END io[162]
  PIN io[163]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 839.840 4.000 840.440 ;
    END
  END io[163]
  PIN io[164]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 809.240 4.000 809.840 ;
    END
  END io[164]
  PIN io[165]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 850.040 4.000 850.640 ;
    END
  END io[165]
  PIN io[166]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 819.440 4.000 820.040 ;
    END
  END io[166]
  PIN io[167]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1145.840 4.000 1146.440 ;
    END
  END io[167]
  PIN io[168]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 829.640 4.000 830.240 ;
    END
  END io[168]
  PIN io[169]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 731.040 4.000 731.640 ;
    END
  END io[169]
  PIN io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1088.040 4.000 1088.640 ;
    END
  END io[16]
  PIN io[170]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 557.640 4.000 558.240 ;
    END
  END io[170]
  PIN io[171]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 741.240 4.000 741.840 ;
    END
  END io[171]
  PIN io[172]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 836.440 4.000 837.040 ;
    END
  END io[172]
  PIN io[173]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 785.440 4.000 786.040 ;
    END
  END io[173]
  PIN io[174]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 860.240 4.000 860.840 ;
    END
  END io[174]
  PIN io[175]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1135.640 4.000 1136.240 ;
    END
  END io[175]
  PIN io[176]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met2 ;
        RECT 367.170 1196.000 367.450 1200.000 ;
    END
  END io[176]
  PIN io[177]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met2 ;
        RECT 409.030 1196.000 409.310 1200.000 ;
    END
  END io[177]
  PIN io[178]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met2 ;
        RECT 373.610 1196.000 373.890 1200.000 ;
    END
  END io[178]
  PIN io[179]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met2 ;
        RECT 418.690 1196.000 418.970 1200.000 ;
    END
  END io[179]
  PIN io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1067.640 4.000 1068.240 ;
    END
  END io[17]
  PIN io[180]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met2 ;
        RECT 341.410 1196.000 341.690 1200.000 ;
    END
  END io[180]
  PIN io[181]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met2 ;
        RECT 386.490 1196.000 386.770 1200.000 ;
    END
  END io[181]
  PIN io[182]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met2 ;
        RECT 331.750 1196.000 332.030 1200.000 ;
    END
  END io[182]
  PIN io[183]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met2 ;
        RECT 322.090 1196.000 322.370 1200.000 ;
    END
  END io[183]
  PIN io[184]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met2 ;
        RECT 299.550 1196.000 299.830 1200.000 ;
    END
  END io[184]
  PIN io[185]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met2 ;
        RECT 277.010 1196.000 277.290 1200.000 ;
    END
  END io[185]
  PIN io[186]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met2 ;
        RECT 254.470 1196.000 254.750 1200.000 ;
    END
  END io[186]
  PIN io[187]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met2 ;
        RECT 244.810 1196.000 245.090 1200.000 ;
    END
  END io[187]
  PIN io[188]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met2 ;
        RECT 231.930 1196.000 232.210 1200.000 ;
    END
  END io[188]
  PIN io[189]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met2 ;
        RECT 222.270 1196.000 222.550 1200.000 ;
    END
  END io[189]
  PIN io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 948.640 4.000 949.240 ;
    END
  END io[18]
  PIN io[190]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met2 ;
        RECT 177.190 1196.000 177.470 1200.000 ;
    END
  END io[190]
  PIN io[191]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.986500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met2 ;
        RECT 206.170 1196.000 206.450 1200.000 ;
    END
  END io[191]
  PIN io[192]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.392800 ;
    ANTENNADIFFAREA 5.302800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 965.640 4.000 966.240 ;
    END
  END io[192]
  PIN io[193]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 962.240 4.000 962.840 ;
    END
  END io[193]
  PIN io[194]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.392800 ;
    ANTENNADIFFAREA 5.302800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1037.040 4.000 1037.640 ;
    END
  END io[194]
  PIN io[195]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 996.240 4.000 996.840 ;
    END
  END io[195]
  PIN io[196]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.392800 ;
    ANTENNADIFFAREA 5.302800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 989.440 4.000 990.040 ;
    END
  END io[196]
  PIN io[197]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 952.040 4.000 952.640 ;
    END
  END io[197]
  PIN io[198]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.392800 ;
    ANTENNADIFFAREA 5.302800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1101.640 4.000 1102.240 ;
    END
  END io[198]
  PIN io[199]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 935.040 4.000 935.640 ;
    END
  END io[199]
  PIN io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.121600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1060.840 4.000 1061.440 ;
    END
  END io[19]
  PIN io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met2 ;
        RECT 296.330 1196.000 296.610 1200.000 ;
    END
  END io[1]
  PIN io[200]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.392800 ;
    ANTENNADIFFAREA 5.302800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 982.640 4.000 983.240 ;
    END
  END io[200]
  PIN io[201]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1091.440 4.000 1092.040 ;
    END
  END io[201]
  PIN io[202]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.392800 ;
    ANTENNADIFFAREA 5.302800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1108.440 4.000 1109.040 ;
    END
  END io[202]
  PIN io[203]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1094.840 4.000 1095.440 ;
    END
  END io[203]
  PIN io[204]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.392800 ;
    ANTENNADIFFAREA 5.302800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 918.040 4.000 918.640 ;
    END
  END io[204]
  PIN io[205]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.070300 ;
    ANTENNADIFFAREA 7.476300 ;
    PORT
      LAYER met2 ;
        RECT 260.910 1196.000 261.190 1200.000 ;
    END
  END io[205]
  PIN io[206]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.392800 ;
    ANTENNADIFFAREA 5.302800 ;
    PORT
      LAYER met2 ;
        RECT 257.690 1196.000 257.970 1200.000 ;
    END
  END io[206]
  PIN io[207]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met2 ;
        RECT 289.890 1196.000 290.170 1200.000 ;
    END
  END io[207]
  PIN io[208]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.392800 ;
    ANTENNADIFFAREA 5.302800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 884.040 4.000 884.640 ;
    END
  END io[208]
  PIN io[209]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 673.240 4.000 673.840 ;
    END
  END io[209]
  PIN io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 945.240 4.000 945.840 ;
    END
  END io[20]
  PIN io[210]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.392800 ;
    ANTENNADIFFAREA 5.302800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 887.440 4.000 888.040 ;
    END
  END io[210]
  PIN io[211]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.121600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 748.040 4.000 748.640 ;
    END
  END io[211]
  PIN io[212]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.392800 ;
    ANTENNADIFFAREA 5.302800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 894.240 4.000 894.840 ;
    END
  END io[212]
  PIN io[213]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 724.240 4.000 724.840 ;
    END
  END io[213]
  PIN io[214]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.392800 ;
    ANTENNADIFFAREA 5.302800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1142.440 4.000 1143.040 ;
    END
  END io[214]
  PIN io[215]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.121600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 690.240 4.000 690.840 ;
    END
  END io[215]
  PIN io[216]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.392800 ;
    ANTENNADIFFAREA 5.302800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.040 4.000 578.640 ;
    END
  END io[216]
  PIN io[217]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 646.040 4.000 646.640 ;
    END
  END io[217]
  PIN io[218]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.392800 ;
    ANTENNADIFFAREA 5.302800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 591.640 4.000 592.240 ;
    END
  END io[218]
  PIN io[219]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.840 4.000 653.440 ;
    END
  END io[219]
  PIN io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1064.240 4.000 1064.840 ;
    END
  END io[21]
  PIN io[220]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.392800 ;
    ANTENNADIFFAREA 5.302800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 601.840 4.000 602.440 ;
    END
  END io[220]
  PIN io[221]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 598.440 4.000 599.040 ;
    END
  END io[221]
  PIN io[222]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.392800 ;
    ANTENNADIFFAREA 5.302800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 744.640 4.000 745.240 ;
    END
  END io[222]
  PIN io[223]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 656.240 4.000 656.840 ;
    END
  END io[223]
  PIN io[224]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.392800 ;
    ANTENNADIFFAREA 5.302800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 758.240 4.000 758.840 ;
    END
  END io[224]
  PIN io[225]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 778.640 4.000 779.240 ;
    END
  END io[225]
  PIN io[226]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.392800 ;
    ANTENNADIFFAREA 5.302800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 612.040 4.000 612.640 ;
    END
  END io[226]
  PIN io[227]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 782.040 4.000 782.640 ;
    END
  END io[227]
  PIN io[228]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.392800 ;
    ANTENNADIFFAREA 5.302800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 775.240 4.000 775.840 ;
    END
  END io[228]
  PIN io[229]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 751.440 4.000 752.040 ;
    END
  END io[229]
  PIN io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1098.240 4.000 1098.840 ;
    END
  END io[22]
  PIN io[230]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.392800 ;
    ANTENNADIFFAREA 5.302800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 588.240 4.000 588.840 ;
    END
  END io[230]
  PIN io[231]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 788.840 4.000 789.440 ;
    END
  END io[231]
  PIN io[232]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.392800 ;
    ANTENNADIFFAREA 5.302800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 761.640 4.000 762.240 ;
    END
  END io[232]
  PIN io[233]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 754.840 4.000 755.440 ;
    END
  END io[233]
  PIN io[234]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.392800 ;
    ANTENNADIFFAREA 5.302800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 663.040 4.000 663.640 ;
    END
  END io[234]
  PIN io[235]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 714.040 4.000 714.640 ;
    END
  END io[235]
  PIN io[236]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.392800 ;
    ANTENNADIFFAREA 5.302800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 833.040 4.000 833.640 ;
    END
  END io[236]
  PIN io[237]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 571.240 4.000 571.840 ;
    END
  END io[237]
  PIN io[238]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.392800 ;
    ANTENNADIFFAREA 5.302800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 846.640 4.000 847.240 ;
    END
  END io[238]
  PIN io[239]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 659.640 4.000 660.240 ;
    END
  END io[239]
  PIN io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.121600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1071.040 4.000 1071.640 ;
    END
  END io[23]
  PIN io[240]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.392800 ;
    ANTENNADIFFAREA 5.302800 ;
    PORT
      LAYER met2 ;
        RECT 344.630 1196.000 344.910 1200.000 ;
    END
  END io[240]
  PIN io[241]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met2 ;
        RECT 434.790 1196.000 435.070 1200.000 ;
    END
  END io[241]
  PIN io[242]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.392800 ;
    ANTENNADIFFAREA 5.302800 ;
    PORT
      LAYER met2 ;
        RECT 334.970 1196.000 335.250 1200.000 ;
    END
  END io[242]
  PIN io[243]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met2 ;
        RECT 431.570 1196.000 431.850 1200.000 ;
    END
  END io[243]
  PIN io[244]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.392800 ;
    ANTENNADIFFAREA 5.302800 ;
    PORT
      LAYER met2 ;
        RECT 338.190 1196.000 338.470 1200.000 ;
    END
  END io[244]
  PIN io[245]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met2 ;
        RECT 428.350 1196.000 428.630 1200.000 ;
    END
  END io[245]
  PIN io[246]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.392800 ;
    ANTENNADIFFAREA 5.302800 ;
    PORT
      LAYER met2 ;
        RECT 328.530 1196.000 328.810 1200.000 ;
    END
  END io[246]
  PIN io[247]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met2 ;
        RECT 425.130 1196.000 425.410 1200.000 ;
    END
  END io[247]
  PIN io[248]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.392800 ;
    ANTENNADIFFAREA 5.302800 ;
    PORT
      LAYER met2 ;
        RECT 283.450 1196.000 283.730 1200.000 ;
    END
  END io[248]
  PIN io[249]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met2 ;
        RECT 293.110 1196.000 293.390 1200.000 ;
    END
  END io[249]
  PIN io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1105.040 4.000 1105.640 ;
    END
  END io[24]
  PIN io[250]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.392800 ;
    ANTENNADIFFAREA 5.302800 ;
    PORT
      LAYER met2 ;
        RECT 273.790 1196.000 274.070 1200.000 ;
    END
  END io[250]
  PIN io[251]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met2 ;
        RECT 267.350 1196.000 267.630 1200.000 ;
    END
  END io[251]
  PIN io[252]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.392800 ;
    ANTENNADIFFAREA 5.302800 ;
    PORT
      LAYER met2 ;
        RECT 248.030 1196.000 248.310 1200.000 ;
    END
  END io[252]
  PIN io[253]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met2 ;
        RECT 270.570 1196.000 270.850 1200.000 ;
    END
  END io[253]
  PIN io[254]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.392800 ;
    ANTENNADIFFAREA 5.302800 ;
    PORT
      LAYER met2 ;
        RECT 186.850 1196.000 187.130 1200.000 ;
    END
  END io[254]
  PIN io[255]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met2 ;
        RECT 241.590 1196.000 241.870 1200.000 ;
    END
  END io[255]
  PIN io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 649.440 4.000 650.040 ;
    END
  END io[25]
  PIN io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 574.640 4.000 575.240 ;
    END
  END io[26]
  PIN io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 615.440 4.000 616.040 ;
    END
  END io[27]
  PIN io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 717.440 4.000 718.040 ;
    END
  END io[28]
  PIN io[29]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 686.840 4.000 687.440 ;
    END
  END io[29]
  PIN io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1047.240 4.000 1047.840 ;
    END
  END io[2]
  PIN io[30]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 720.840 4.000 721.440 ;
    END
  END io[30]
  PIN io[31]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 639.240 4.000 639.840 ;
    END
  END io[31]
  PIN io[32]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 581.440 4.000 582.040 ;
    END
  END io[32]
  PIN io[33]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1125.440 4.000 1126.040 ;
    END
  END io[33]
  PIN io[34]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 642.640 4.000 643.240 ;
    END
  END io[34]
  PIN io[35]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 914.640 4.000 915.240 ;
    END
  END io[35]
  PIN io[36]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.000100 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 595.040 4.000 595.640 ;
    END
  END io[36]
  PIN io[37]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 911.240 4.000 911.840 ;
    END
  END io[37]
  PIN io[38]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 676.640 4.000 677.240 ;
    END
  END io[38]
  PIN io[39]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 907.840 4.000 908.440 ;
    END
  END io[39]
  PIN io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met2 ;
        RECT 196.510 1196.000 196.790 1200.000 ;
    END
  END io[3]
  PIN io[40]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1118.640 4.000 1119.240 ;
    END
  END io[40]
  PIN io[41]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 584.840 4.000 585.440 ;
    END
  END io[41]
  PIN io[42]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1132.240 4.000 1132.840 ;
    END
  END io[42]
  PIN io[43]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 710.640 4.000 711.240 ;
    END
  END io[43]
  PIN io[44]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.000100 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 890.840 4.000 891.440 ;
    END
  END io[44]
  PIN io[45]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 635.840 4.000 636.440 ;
    END
  END io[45]
  PIN io[46]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 897.640 4.000 898.240 ;
    END
  END io[46]
  PIN io[47]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 707.240 4.000 707.840 ;
    END
  END io[47]
  PIN io[48]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met2 ;
        RECT 360.730 1196.000 361.010 1200.000 ;
    END
  END io[48]
  PIN io[49]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met2 ;
        RECT 421.910 1196.000 422.190 1200.000 ;
    END
  END io[49]
  PIN io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.000100 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1040.440 4.000 1041.040 ;
    END
  END io[4]
  PIN io[50]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met2 ;
        RECT 357.510 1196.000 357.790 1200.000 ;
    END
  END io[50]
  PIN io[51]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met2 ;
        RECT 405.810 1196.000 406.090 1200.000 ;
    END
  END io[51]
  PIN io[52]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.000100 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met2 ;
        RECT 318.870 1196.000 319.150 1200.000 ;
    END
  END io[52]
  PIN io[53]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met2 ;
        RECT 402.590 1196.000 402.870 1200.000 ;
    END
  END io[53]
  PIN io[54]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met2 ;
        RECT 315.650 1196.000 315.930 1200.000 ;
    END
  END io[54]
  PIN io[55]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met2 ;
        RECT 399.370 1196.000 399.650 1200.000 ;
    END
  END io[55]
  PIN io[56]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met2 ;
        RECT 199.730 1196.000 200.010 1200.000 ;
    END
  END io[56]
  PIN io[57]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met2 ;
        RECT 286.670 1196.000 286.950 1200.000 ;
    END
  END io[57]
  PIN io[58]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met2 ;
        RECT 228.710 1196.000 228.990 1200.000 ;
    END
  END io[58]
  PIN io[59]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met2 ;
        RECT 238.370 1196.000 238.650 1200.000 ;
    END
  END io[59]
  PIN io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1054.040 4.000 1054.640 ;
    END
  END io[5]
  PIN io[60]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.000100 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met2 ;
        RECT 193.290 1196.000 193.570 1200.000 ;
    END
  END io[60]
  PIN io[61]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met2 ;
        RECT 235.150 1196.000 235.430 1200.000 ;
    END
  END io[61]
  PIN io[62]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met2 ;
        RECT 202.950 1196.000 203.230 1200.000 ;
    END
  END io[62]
  PIN io[63]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met2 ;
        RECT 219.050 1196.000 219.330 1200.000 ;
    END
  END io[63]
  PIN io[64]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1009.840 4.000 1010.440 ;
    END
  END io[64]
  PIN io[65]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.953500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met2 ;
        RECT 312.430 1196.000 312.710 1200.000 ;
    END
  END io[65]
  PIN io[66]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met2 ;
        RECT 309.210 1196.000 309.490 1200.000 ;
    END
  END io[66]
  PIN io[67]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met2 ;
        RECT 173.970 1196.000 174.250 1200.000 ;
    END
  END io[67]
  PIN io[68]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1003.040 4.000 1003.640 ;
    END
  END io[68]
  PIN io[69]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 928.240 4.000 928.840 ;
    END
  END io[69]
  PIN io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 972.440 4.000 973.040 ;
    END
  END io[6]
  PIN io[70]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 921.440 4.000 922.040 ;
    END
  END io[70]
  PIN io[71]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.953500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 771.840 4.000 772.440 ;
    END
  END io[71]
  PIN io[72]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 986.040 4.000 986.640 ;
    END
  END io[72]
  PIN io[73]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 958.840 4.000 959.440 ;
    END
  END io[73]
  PIN io[74]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 941.840 4.000 942.440 ;
    END
  END io[74]
  PIN io[75]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1122.040 4.000 1122.640 ;
    END
  END io[75]
  PIN io[76]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.953500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 924.840 4.000 925.440 ;
    END
  END io[76]
  PIN io[77]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1128.840 4.000 1129.440 ;
    END
  END io[77]
  PIN io[78]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1030.240 4.000 1030.840 ;
    END
  END io[78]
  PIN io[79]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1013.240 4.000 1013.840 ;
    END
  END io[79]
  PIN io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1057.440 4.000 1058.040 ;
    END
  END io[7]
  PIN io[80]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 816.040 4.000 816.640 ;
    END
  END io[80]
  PIN io[81]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 863.640 4.000 864.240 ;
    END
  END io[81]
  PIN io[82]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 999.640 4.000 1000.240 ;
    END
  END io[82]
  PIN io[83]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1033.640 4.000 1034.240 ;
    END
  END io[83]
  PIN io[84]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.953500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 931.640 4.000 932.240 ;
    END
  END io[84]
  PIN io[85]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.953500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 880.640 4.000 881.240 ;
    END
  END io[85]
  PIN io[86]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 812.640 4.000 813.240 ;
    END
  END io[86]
  PIN io[87]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.953500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 765.040 4.000 765.640 ;
    END
  END io[87]
  PIN io[88]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 737.840 4.000 738.440 ;
    END
  END io[88]
  PIN io[89]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 622.240 4.000 622.840 ;
    END
  END io[89]
  PIN io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met2 ;
        RECT 164.310 1196.000 164.590 1200.000 ;
    END
  END io[8]
  PIN io[90]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 680.040 4.000 680.640 ;
    END
  END io[90]
  PIN io[91]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 564.440 4.000 565.040 ;
    END
  END io[91]
  PIN io[92]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.953500 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 632.440 4.000 633.040 ;
    END
  END io[92]
  PIN io[93]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 605.240 4.000 605.840 ;
    END
  END io[93]
  PIN io[94]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 683.440 4.000 684.040 ;
    END
  END io[94]
  PIN io[95]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 703.840 4.000 704.440 ;
    END
  END io[95]
  PIN io[96]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 727.640 4.000 728.240 ;
    END
  END io[96]
  PIN io[97]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 795.640 4.000 796.240 ;
    END
  END io[97]
  PIN io[98]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 734.440 4.000 735.040 ;
    END
  END io[98]
  PIN io[99]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 5.737500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 843.240 4.000 843.840 ;
    END
  END io[99]
  PIN io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.635600 ;
    ANTENNADIFFAREA 7.041600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 969.040 4.000 969.640 ;
    END
  END io[9]
  PIN nrst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.860700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 17.040 1200.000 17.640 ;
    END
  END nrst
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 1194.350 1188.830 ;
      LAYER li1 ;
        RECT 5.520 10.795 1194.160 1188.725 ;
      LAYER met1 ;
        RECT 0.530 10.640 1194.160 1196.760 ;
      LAYER met2 ;
        RECT 0.550 1195.720 164.030 1196.790 ;
        RECT 164.870 1195.720 167.250 1196.790 ;
        RECT 168.090 1195.720 170.470 1196.790 ;
        RECT 171.310 1195.720 173.690 1196.790 ;
        RECT 174.530 1195.720 176.910 1196.790 ;
        RECT 177.750 1195.720 180.130 1196.790 ;
        RECT 180.970 1195.720 183.350 1196.790 ;
        RECT 184.190 1195.720 186.570 1196.790 ;
        RECT 187.410 1195.720 189.790 1196.790 ;
        RECT 190.630 1195.720 193.010 1196.790 ;
        RECT 193.850 1195.720 196.230 1196.790 ;
        RECT 197.070 1195.720 199.450 1196.790 ;
        RECT 200.290 1195.720 202.670 1196.790 ;
        RECT 203.510 1195.720 205.890 1196.790 ;
        RECT 206.730 1195.720 209.110 1196.790 ;
        RECT 209.950 1195.720 212.330 1196.790 ;
        RECT 213.170 1195.720 215.550 1196.790 ;
        RECT 216.390 1195.720 218.770 1196.790 ;
        RECT 219.610 1195.720 221.990 1196.790 ;
        RECT 222.830 1195.720 225.210 1196.790 ;
        RECT 226.050 1195.720 228.430 1196.790 ;
        RECT 229.270 1195.720 231.650 1196.790 ;
        RECT 232.490 1195.720 234.870 1196.790 ;
        RECT 235.710 1195.720 238.090 1196.790 ;
        RECT 238.930 1195.720 241.310 1196.790 ;
        RECT 242.150 1195.720 244.530 1196.790 ;
        RECT 245.370 1195.720 247.750 1196.790 ;
        RECT 248.590 1195.720 250.970 1196.790 ;
        RECT 251.810 1195.720 254.190 1196.790 ;
        RECT 255.030 1195.720 257.410 1196.790 ;
        RECT 258.250 1195.720 260.630 1196.790 ;
        RECT 261.470 1195.720 263.850 1196.790 ;
        RECT 264.690 1195.720 267.070 1196.790 ;
        RECT 267.910 1195.720 270.290 1196.790 ;
        RECT 271.130 1195.720 273.510 1196.790 ;
        RECT 274.350 1195.720 276.730 1196.790 ;
        RECT 277.570 1195.720 279.950 1196.790 ;
        RECT 280.790 1195.720 283.170 1196.790 ;
        RECT 284.010 1195.720 286.390 1196.790 ;
        RECT 287.230 1195.720 289.610 1196.790 ;
        RECT 290.450 1195.720 292.830 1196.790 ;
        RECT 293.670 1195.720 296.050 1196.790 ;
        RECT 296.890 1195.720 299.270 1196.790 ;
        RECT 300.110 1195.720 302.490 1196.790 ;
        RECT 303.330 1195.720 305.710 1196.790 ;
        RECT 306.550 1195.720 308.930 1196.790 ;
        RECT 309.770 1195.720 312.150 1196.790 ;
        RECT 312.990 1195.720 315.370 1196.790 ;
        RECT 316.210 1195.720 318.590 1196.790 ;
        RECT 319.430 1195.720 321.810 1196.790 ;
        RECT 322.650 1195.720 325.030 1196.790 ;
        RECT 325.870 1195.720 328.250 1196.790 ;
        RECT 329.090 1195.720 331.470 1196.790 ;
        RECT 332.310 1195.720 334.690 1196.790 ;
        RECT 335.530 1195.720 337.910 1196.790 ;
        RECT 338.750 1195.720 341.130 1196.790 ;
        RECT 341.970 1195.720 344.350 1196.790 ;
        RECT 345.190 1195.720 347.570 1196.790 ;
        RECT 348.410 1195.720 350.790 1196.790 ;
        RECT 351.630 1195.720 354.010 1196.790 ;
        RECT 354.850 1195.720 357.230 1196.790 ;
        RECT 358.070 1195.720 360.450 1196.790 ;
        RECT 361.290 1195.720 363.670 1196.790 ;
        RECT 364.510 1195.720 366.890 1196.790 ;
        RECT 367.730 1195.720 370.110 1196.790 ;
        RECT 370.950 1195.720 373.330 1196.790 ;
        RECT 374.170 1195.720 386.210 1196.790 ;
        RECT 387.050 1195.720 389.430 1196.790 ;
        RECT 390.270 1195.720 399.090 1196.790 ;
        RECT 399.930 1195.720 402.310 1196.790 ;
        RECT 403.150 1195.720 405.530 1196.790 ;
        RECT 406.370 1195.720 408.750 1196.790 ;
        RECT 409.590 1195.720 411.970 1196.790 ;
        RECT 412.810 1195.720 415.190 1196.790 ;
        RECT 416.030 1195.720 418.410 1196.790 ;
        RECT 419.250 1195.720 421.630 1196.790 ;
        RECT 422.470 1195.720 424.850 1196.790 ;
        RECT 425.690 1195.720 428.070 1196.790 ;
        RECT 428.910 1195.720 431.290 1196.790 ;
        RECT 432.130 1195.720 434.510 1196.790 ;
        RECT 435.350 1195.720 1193.150 1196.790 ;
        RECT 0.550 10.695 1193.150 1195.720 ;
      LAYER met3 ;
        RECT 0.270 1157.040 1196.000 1196.625 ;
        RECT 4.400 1155.640 1196.000 1157.040 ;
        RECT 0.270 1153.640 1196.000 1155.640 ;
        RECT 4.400 1152.240 1196.000 1153.640 ;
        RECT 0.270 1150.240 1196.000 1152.240 ;
        RECT 4.400 1148.840 1196.000 1150.240 ;
        RECT 0.270 1146.840 1196.000 1148.840 ;
        RECT 4.400 1145.440 1196.000 1146.840 ;
        RECT 0.270 1143.440 1196.000 1145.440 ;
        RECT 4.400 1142.040 1196.000 1143.440 ;
        RECT 0.270 1140.040 1196.000 1142.040 ;
        RECT 4.400 1138.640 1196.000 1140.040 ;
        RECT 0.270 1136.640 1196.000 1138.640 ;
        RECT 4.400 1135.240 1196.000 1136.640 ;
        RECT 0.270 1133.240 1196.000 1135.240 ;
        RECT 4.400 1131.840 1196.000 1133.240 ;
        RECT 0.270 1129.840 1196.000 1131.840 ;
        RECT 4.400 1128.440 1196.000 1129.840 ;
        RECT 0.270 1126.440 1196.000 1128.440 ;
        RECT 4.400 1125.040 1196.000 1126.440 ;
        RECT 0.270 1123.040 1196.000 1125.040 ;
        RECT 4.400 1121.640 1196.000 1123.040 ;
        RECT 0.270 1119.640 1196.000 1121.640 ;
        RECT 4.400 1118.240 1196.000 1119.640 ;
        RECT 0.270 1116.240 1196.000 1118.240 ;
        RECT 4.400 1114.840 1196.000 1116.240 ;
        RECT 0.270 1112.840 1196.000 1114.840 ;
        RECT 4.400 1111.440 1196.000 1112.840 ;
        RECT 0.270 1109.440 1196.000 1111.440 ;
        RECT 4.400 1108.040 1196.000 1109.440 ;
        RECT 0.270 1106.040 1196.000 1108.040 ;
        RECT 4.400 1104.640 1196.000 1106.040 ;
        RECT 0.270 1102.640 1196.000 1104.640 ;
        RECT 4.400 1101.240 1196.000 1102.640 ;
        RECT 0.270 1099.240 1196.000 1101.240 ;
        RECT 4.400 1097.840 1196.000 1099.240 ;
        RECT 0.270 1095.840 1196.000 1097.840 ;
        RECT 4.400 1094.440 1196.000 1095.840 ;
        RECT 0.270 1092.440 1196.000 1094.440 ;
        RECT 4.400 1091.040 1196.000 1092.440 ;
        RECT 0.270 1089.040 1196.000 1091.040 ;
        RECT 4.400 1087.640 1196.000 1089.040 ;
        RECT 0.270 1085.640 1196.000 1087.640 ;
        RECT 4.400 1084.240 1196.000 1085.640 ;
        RECT 0.270 1082.240 1196.000 1084.240 ;
        RECT 4.400 1080.840 1196.000 1082.240 ;
        RECT 0.270 1078.840 1196.000 1080.840 ;
        RECT 4.400 1077.440 1196.000 1078.840 ;
        RECT 0.270 1075.440 1196.000 1077.440 ;
        RECT 4.400 1074.040 1196.000 1075.440 ;
        RECT 0.270 1072.040 1196.000 1074.040 ;
        RECT 4.400 1070.640 1196.000 1072.040 ;
        RECT 0.270 1068.640 1196.000 1070.640 ;
        RECT 4.400 1067.240 1196.000 1068.640 ;
        RECT 0.270 1065.240 1196.000 1067.240 ;
        RECT 4.400 1063.840 1196.000 1065.240 ;
        RECT 0.270 1061.840 1196.000 1063.840 ;
        RECT 4.400 1060.440 1196.000 1061.840 ;
        RECT 0.270 1058.440 1196.000 1060.440 ;
        RECT 4.400 1057.040 1196.000 1058.440 ;
        RECT 0.270 1055.040 1196.000 1057.040 ;
        RECT 4.400 1053.640 1196.000 1055.040 ;
        RECT 0.270 1051.640 1196.000 1053.640 ;
        RECT 4.400 1050.240 1196.000 1051.640 ;
        RECT 0.270 1048.240 1196.000 1050.240 ;
        RECT 4.400 1046.840 1196.000 1048.240 ;
        RECT 0.270 1044.840 1196.000 1046.840 ;
        RECT 4.400 1043.440 1196.000 1044.840 ;
        RECT 0.270 1041.440 1196.000 1043.440 ;
        RECT 4.400 1040.040 1196.000 1041.440 ;
        RECT 0.270 1038.040 1196.000 1040.040 ;
        RECT 4.400 1036.640 1196.000 1038.040 ;
        RECT 0.270 1034.640 1196.000 1036.640 ;
        RECT 4.400 1033.240 1196.000 1034.640 ;
        RECT 0.270 1031.240 1196.000 1033.240 ;
        RECT 4.400 1029.840 1196.000 1031.240 ;
        RECT 0.270 1027.840 1196.000 1029.840 ;
        RECT 4.400 1026.440 1196.000 1027.840 ;
        RECT 0.270 1024.440 1196.000 1026.440 ;
        RECT 4.400 1023.040 1196.000 1024.440 ;
        RECT 0.270 1021.040 1196.000 1023.040 ;
        RECT 4.400 1019.640 1196.000 1021.040 ;
        RECT 0.270 1017.640 1196.000 1019.640 ;
        RECT 4.400 1016.240 1196.000 1017.640 ;
        RECT 0.270 1014.240 1196.000 1016.240 ;
        RECT 4.400 1012.840 1196.000 1014.240 ;
        RECT 0.270 1010.840 1196.000 1012.840 ;
        RECT 4.400 1009.440 1196.000 1010.840 ;
        RECT 0.270 1007.440 1196.000 1009.440 ;
        RECT 4.400 1006.040 1196.000 1007.440 ;
        RECT 0.270 1004.040 1196.000 1006.040 ;
        RECT 4.400 1002.640 1196.000 1004.040 ;
        RECT 0.270 1000.640 1196.000 1002.640 ;
        RECT 4.400 999.240 1196.000 1000.640 ;
        RECT 0.270 997.240 1196.000 999.240 ;
        RECT 4.400 995.840 1196.000 997.240 ;
        RECT 0.270 993.840 1196.000 995.840 ;
        RECT 4.400 992.440 1196.000 993.840 ;
        RECT 0.270 990.440 1196.000 992.440 ;
        RECT 4.400 989.040 1196.000 990.440 ;
        RECT 0.270 987.040 1196.000 989.040 ;
        RECT 4.400 985.640 1196.000 987.040 ;
        RECT 0.270 983.640 1196.000 985.640 ;
        RECT 4.400 982.240 1196.000 983.640 ;
        RECT 0.270 980.240 1196.000 982.240 ;
        RECT 4.400 978.840 1196.000 980.240 ;
        RECT 0.270 976.840 1196.000 978.840 ;
        RECT 4.400 975.440 1196.000 976.840 ;
        RECT 0.270 973.440 1196.000 975.440 ;
        RECT 4.400 972.040 1196.000 973.440 ;
        RECT 0.270 970.040 1196.000 972.040 ;
        RECT 4.400 968.640 1196.000 970.040 ;
        RECT 0.270 966.640 1196.000 968.640 ;
        RECT 4.400 965.240 1196.000 966.640 ;
        RECT 0.270 963.240 1196.000 965.240 ;
        RECT 4.400 961.840 1196.000 963.240 ;
        RECT 0.270 959.840 1196.000 961.840 ;
        RECT 4.400 958.440 1196.000 959.840 ;
        RECT 0.270 956.440 1196.000 958.440 ;
        RECT 4.400 955.040 1196.000 956.440 ;
        RECT 0.270 953.040 1196.000 955.040 ;
        RECT 4.400 951.640 1196.000 953.040 ;
        RECT 0.270 949.640 1196.000 951.640 ;
        RECT 4.400 948.240 1196.000 949.640 ;
        RECT 0.270 946.240 1196.000 948.240 ;
        RECT 4.400 944.840 1196.000 946.240 ;
        RECT 0.270 942.840 1196.000 944.840 ;
        RECT 4.400 941.440 1196.000 942.840 ;
        RECT 0.270 939.440 1196.000 941.440 ;
        RECT 4.400 938.040 1196.000 939.440 ;
        RECT 0.270 936.040 1196.000 938.040 ;
        RECT 4.400 934.640 1196.000 936.040 ;
        RECT 0.270 932.640 1196.000 934.640 ;
        RECT 4.400 931.240 1196.000 932.640 ;
        RECT 0.270 929.240 1196.000 931.240 ;
        RECT 4.400 927.840 1196.000 929.240 ;
        RECT 0.270 925.840 1196.000 927.840 ;
        RECT 4.400 924.440 1196.000 925.840 ;
        RECT 0.270 922.440 1196.000 924.440 ;
        RECT 4.400 921.040 1196.000 922.440 ;
        RECT 0.270 919.040 1196.000 921.040 ;
        RECT 4.400 917.640 1196.000 919.040 ;
        RECT 0.270 915.640 1196.000 917.640 ;
        RECT 4.400 914.240 1196.000 915.640 ;
        RECT 0.270 912.240 1196.000 914.240 ;
        RECT 4.400 910.840 1196.000 912.240 ;
        RECT 0.270 908.840 1196.000 910.840 ;
        RECT 4.400 907.440 1196.000 908.840 ;
        RECT 0.270 905.440 1196.000 907.440 ;
        RECT 4.400 904.040 1196.000 905.440 ;
        RECT 0.270 902.040 1196.000 904.040 ;
        RECT 4.400 900.640 1196.000 902.040 ;
        RECT 0.270 898.640 1196.000 900.640 ;
        RECT 4.400 897.240 1196.000 898.640 ;
        RECT 0.270 895.240 1196.000 897.240 ;
        RECT 4.400 893.840 1196.000 895.240 ;
        RECT 0.270 891.840 1196.000 893.840 ;
        RECT 4.400 890.440 1196.000 891.840 ;
        RECT 0.270 888.440 1196.000 890.440 ;
        RECT 4.400 887.040 1196.000 888.440 ;
        RECT 0.270 885.040 1196.000 887.040 ;
        RECT 4.400 883.640 1196.000 885.040 ;
        RECT 0.270 881.640 1196.000 883.640 ;
        RECT 4.400 880.240 1196.000 881.640 ;
        RECT 0.270 878.240 1196.000 880.240 ;
        RECT 4.400 876.840 1196.000 878.240 ;
        RECT 0.270 874.840 1196.000 876.840 ;
        RECT 4.400 873.440 1196.000 874.840 ;
        RECT 0.270 871.440 1196.000 873.440 ;
        RECT 4.400 870.040 1196.000 871.440 ;
        RECT 0.270 868.040 1196.000 870.040 ;
        RECT 4.400 866.640 1196.000 868.040 ;
        RECT 0.270 864.640 1196.000 866.640 ;
        RECT 4.400 863.240 1196.000 864.640 ;
        RECT 0.270 861.240 1196.000 863.240 ;
        RECT 4.400 859.840 1196.000 861.240 ;
        RECT 0.270 857.840 1196.000 859.840 ;
        RECT 4.400 856.440 1196.000 857.840 ;
        RECT 0.270 854.440 1196.000 856.440 ;
        RECT 4.400 853.040 1196.000 854.440 ;
        RECT 0.270 851.040 1196.000 853.040 ;
        RECT 4.400 849.640 1196.000 851.040 ;
        RECT 0.270 847.640 1196.000 849.640 ;
        RECT 4.400 846.240 1196.000 847.640 ;
        RECT 0.270 844.240 1196.000 846.240 ;
        RECT 4.400 842.840 1196.000 844.240 ;
        RECT 0.270 840.840 1196.000 842.840 ;
        RECT 4.400 839.440 1196.000 840.840 ;
        RECT 0.270 837.440 1196.000 839.440 ;
        RECT 4.400 836.040 1196.000 837.440 ;
        RECT 0.270 834.040 1196.000 836.040 ;
        RECT 4.400 832.640 1196.000 834.040 ;
        RECT 0.270 830.640 1196.000 832.640 ;
        RECT 4.400 829.240 1196.000 830.640 ;
        RECT 0.270 827.240 1196.000 829.240 ;
        RECT 4.400 825.840 1196.000 827.240 ;
        RECT 0.270 823.840 1196.000 825.840 ;
        RECT 4.400 822.440 1196.000 823.840 ;
        RECT 0.270 820.440 1196.000 822.440 ;
        RECT 4.400 819.040 1196.000 820.440 ;
        RECT 0.270 817.040 1196.000 819.040 ;
        RECT 4.400 815.640 1196.000 817.040 ;
        RECT 0.270 813.640 1196.000 815.640 ;
        RECT 4.400 812.240 1196.000 813.640 ;
        RECT 0.270 810.240 1196.000 812.240 ;
        RECT 4.400 808.840 1196.000 810.240 ;
        RECT 0.270 806.840 1196.000 808.840 ;
        RECT 4.400 805.440 1196.000 806.840 ;
        RECT 0.270 803.440 1196.000 805.440 ;
        RECT 4.400 802.040 1196.000 803.440 ;
        RECT 0.270 800.040 1196.000 802.040 ;
        RECT 4.400 798.640 1196.000 800.040 ;
        RECT 0.270 796.640 1196.000 798.640 ;
        RECT 4.400 795.240 1196.000 796.640 ;
        RECT 0.270 793.240 1196.000 795.240 ;
        RECT 4.400 791.840 1196.000 793.240 ;
        RECT 0.270 789.840 1196.000 791.840 ;
        RECT 4.400 788.440 1196.000 789.840 ;
        RECT 0.270 786.440 1196.000 788.440 ;
        RECT 4.400 785.040 1196.000 786.440 ;
        RECT 0.270 783.040 1196.000 785.040 ;
        RECT 4.400 781.640 1196.000 783.040 ;
        RECT 0.270 779.640 1196.000 781.640 ;
        RECT 4.400 778.240 1196.000 779.640 ;
        RECT 0.270 776.240 1196.000 778.240 ;
        RECT 4.400 774.840 1196.000 776.240 ;
        RECT 0.270 772.840 1196.000 774.840 ;
        RECT 4.400 771.440 1196.000 772.840 ;
        RECT 0.270 769.440 1196.000 771.440 ;
        RECT 4.400 768.040 1196.000 769.440 ;
        RECT 0.270 766.040 1196.000 768.040 ;
        RECT 4.400 764.640 1196.000 766.040 ;
        RECT 0.270 762.640 1196.000 764.640 ;
        RECT 4.400 761.240 1196.000 762.640 ;
        RECT 0.270 759.240 1196.000 761.240 ;
        RECT 4.400 757.840 1196.000 759.240 ;
        RECT 0.270 755.840 1196.000 757.840 ;
        RECT 4.400 754.440 1196.000 755.840 ;
        RECT 0.270 752.440 1196.000 754.440 ;
        RECT 4.400 751.040 1196.000 752.440 ;
        RECT 0.270 749.040 1196.000 751.040 ;
        RECT 4.400 747.640 1196.000 749.040 ;
        RECT 0.270 745.640 1196.000 747.640 ;
        RECT 4.400 744.240 1196.000 745.640 ;
        RECT 0.270 742.240 1196.000 744.240 ;
        RECT 4.400 740.840 1196.000 742.240 ;
        RECT 0.270 738.840 1196.000 740.840 ;
        RECT 4.400 737.440 1196.000 738.840 ;
        RECT 0.270 735.440 1196.000 737.440 ;
        RECT 4.400 734.040 1196.000 735.440 ;
        RECT 0.270 732.040 1196.000 734.040 ;
        RECT 4.400 730.640 1196.000 732.040 ;
        RECT 0.270 728.640 1196.000 730.640 ;
        RECT 4.400 727.240 1196.000 728.640 ;
        RECT 0.270 725.240 1196.000 727.240 ;
        RECT 4.400 723.840 1196.000 725.240 ;
        RECT 0.270 721.840 1196.000 723.840 ;
        RECT 4.400 720.440 1196.000 721.840 ;
        RECT 0.270 718.440 1196.000 720.440 ;
        RECT 4.400 717.040 1196.000 718.440 ;
        RECT 0.270 715.040 1196.000 717.040 ;
        RECT 4.400 713.640 1196.000 715.040 ;
        RECT 0.270 711.640 1196.000 713.640 ;
        RECT 4.400 710.240 1196.000 711.640 ;
        RECT 0.270 708.240 1196.000 710.240 ;
        RECT 4.400 706.840 1196.000 708.240 ;
        RECT 0.270 704.840 1196.000 706.840 ;
        RECT 4.400 703.440 1196.000 704.840 ;
        RECT 0.270 701.440 1196.000 703.440 ;
        RECT 4.400 700.040 1196.000 701.440 ;
        RECT 0.270 698.040 1196.000 700.040 ;
        RECT 4.400 696.640 1196.000 698.040 ;
        RECT 0.270 694.640 1196.000 696.640 ;
        RECT 4.400 693.240 1196.000 694.640 ;
        RECT 0.270 691.240 1196.000 693.240 ;
        RECT 4.400 689.840 1196.000 691.240 ;
        RECT 0.270 687.840 1196.000 689.840 ;
        RECT 4.400 686.440 1196.000 687.840 ;
        RECT 0.270 684.440 1196.000 686.440 ;
        RECT 4.400 683.040 1196.000 684.440 ;
        RECT 0.270 681.040 1196.000 683.040 ;
        RECT 4.400 679.640 1196.000 681.040 ;
        RECT 0.270 677.640 1196.000 679.640 ;
        RECT 4.400 676.240 1196.000 677.640 ;
        RECT 0.270 674.240 1196.000 676.240 ;
        RECT 4.400 672.840 1196.000 674.240 ;
        RECT 0.270 670.840 1196.000 672.840 ;
        RECT 4.400 669.440 1196.000 670.840 ;
        RECT 0.270 667.440 1196.000 669.440 ;
        RECT 4.400 666.040 1196.000 667.440 ;
        RECT 0.270 664.040 1196.000 666.040 ;
        RECT 4.400 662.640 1196.000 664.040 ;
        RECT 0.270 660.640 1196.000 662.640 ;
        RECT 4.400 659.240 1196.000 660.640 ;
        RECT 0.270 657.240 1196.000 659.240 ;
        RECT 4.400 655.840 1196.000 657.240 ;
        RECT 0.270 653.840 1196.000 655.840 ;
        RECT 4.400 652.440 1196.000 653.840 ;
        RECT 0.270 650.440 1196.000 652.440 ;
        RECT 4.400 649.040 1196.000 650.440 ;
        RECT 0.270 647.040 1196.000 649.040 ;
        RECT 4.400 645.640 1196.000 647.040 ;
        RECT 0.270 643.640 1196.000 645.640 ;
        RECT 4.400 642.240 1196.000 643.640 ;
        RECT 0.270 640.240 1196.000 642.240 ;
        RECT 4.400 638.840 1196.000 640.240 ;
        RECT 0.270 636.840 1196.000 638.840 ;
        RECT 4.400 635.440 1196.000 636.840 ;
        RECT 0.270 633.440 1196.000 635.440 ;
        RECT 4.400 632.040 1196.000 633.440 ;
        RECT 0.270 630.040 1196.000 632.040 ;
        RECT 4.400 628.640 1196.000 630.040 ;
        RECT 0.270 626.640 1196.000 628.640 ;
        RECT 4.400 625.240 1196.000 626.640 ;
        RECT 0.270 623.240 1196.000 625.240 ;
        RECT 4.400 621.840 1196.000 623.240 ;
        RECT 0.270 619.840 1196.000 621.840 ;
        RECT 4.400 618.440 1196.000 619.840 ;
        RECT 0.270 616.440 1196.000 618.440 ;
        RECT 4.400 615.040 1196.000 616.440 ;
        RECT 0.270 613.040 1196.000 615.040 ;
        RECT 4.400 611.640 1196.000 613.040 ;
        RECT 0.270 609.640 1196.000 611.640 ;
        RECT 4.400 608.240 1196.000 609.640 ;
        RECT 0.270 606.240 1196.000 608.240 ;
        RECT 4.400 604.840 1196.000 606.240 ;
        RECT 0.270 602.840 1196.000 604.840 ;
        RECT 4.400 601.440 1196.000 602.840 ;
        RECT 0.270 599.440 1196.000 601.440 ;
        RECT 4.400 598.040 1196.000 599.440 ;
        RECT 0.270 596.040 1196.000 598.040 ;
        RECT 4.400 594.640 1196.000 596.040 ;
        RECT 0.270 592.640 1196.000 594.640 ;
        RECT 4.400 591.240 1196.000 592.640 ;
        RECT 0.270 589.240 1196.000 591.240 ;
        RECT 4.400 587.840 1196.000 589.240 ;
        RECT 0.270 585.840 1196.000 587.840 ;
        RECT 4.400 584.440 1196.000 585.840 ;
        RECT 0.270 582.440 1196.000 584.440 ;
        RECT 4.400 581.040 1196.000 582.440 ;
        RECT 0.270 579.040 1196.000 581.040 ;
        RECT 4.400 577.640 1196.000 579.040 ;
        RECT 0.270 575.640 1196.000 577.640 ;
        RECT 4.400 574.240 1196.000 575.640 ;
        RECT 0.270 572.240 1196.000 574.240 ;
        RECT 4.400 570.840 1196.000 572.240 ;
        RECT 0.270 568.840 1196.000 570.840 ;
        RECT 4.400 567.440 1196.000 568.840 ;
        RECT 0.270 565.440 1196.000 567.440 ;
        RECT 4.400 564.040 1196.000 565.440 ;
        RECT 0.270 562.040 1196.000 564.040 ;
        RECT 4.400 560.640 1196.000 562.040 ;
        RECT 0.270 558.640 1196.000 560.640 ;
        RECT 4.400 557.240 1196.000 558.640 ;
        RECT 0.270 555.240 1196.000 557.240 ;
        RECT 4.400 553.840 1196.000 555.240 ;
        RECT 0.270 551.840 1196.000 553.840 ;
        RECT 4.400 550.440 1196.000 551.840 ;
        RECT 0.270 18.040 1196.000 550.440 ;
        RECT 0.270 16.640 1195.600 18.040 ;
        RECT 0.270 10.715 1196.000 16.640 ;
      LAYER met4 ;
        RECT 0.295 1189.280 1180.065 1196.625 ;
        RECT 0.295 15.815 20.640 1189.280 ;
        RECT 23.040 15.815 23.940 1189.280 ;
        RECT 26.340 15.815 174.240 1189.280 ;
        RECT 176.640 15.815 177.540 1189.280 ;
        RECT 179.940 15.815 327.840 1189.280 ;
        RECT 330.240 15.815 331.140 1189.280 ;
        RECT 333.540 15.815 481.440 1189.280 ;
        RECT 483.840 15.815 484.740 1189.280 ;
        RECT 487.140 15.815 635.040 1189.280 ;
        RECT 637.440 15.815 638.340 1189.280 ;
        RECT 640.740 15.815 788.640 1189.280 ;
        RECT 791.040 15.815 791.940 1189.280 ;
        RECT 794.340 15.815 942.240 1189.280 ;
        RECT 944.640 15.815 945.540 1189.280 ;
        RECT 947.940 15.815 1095.840 1189.280 ;
        RECT 1098.240 15.815 1099.140 1189.280 ;
        RECT 1101.540 15.815 1180.065 1189.280 ;
  END
END fpga
END LIBRARY

