magic
tech sky130A
magscale 1 2
timestamp 1752639015
<< viali >>
rect 8677 95625 8711 95659
rect 14749 95625 14783 95659
rect 16681 95625 16715 95659
rect 17969 95625 18003 95659
rect 19349 95625 19383 95659
rect 20453 95625 20487 95659
rect 21189 95625 21223 95659
rect 22477 95625 22511 95659
rect 23121 95625 23155 95659
rect 24409 95625 24443 95659
rect 25697 95625 25731 95659
rect 26985 95625 27019 95659
rect 27629 95625 27663 95659
rect 29009 95625 29043 95659
rect 30573 95625 30607 95659
rect 31125 95625 31159 95659
rect 32505 95625 32539 95659
rect 33793 95625 33827 95659
rect 35081 95625 35115 95659
rect 35633 95625 35667 95659
rect 37013 95625 37047 95659
rect 38301 95625 38335 95659
rect 38853 95625 38887 95659
rect 40233 95625 40267 95659
rect 41521 95625 41555 95659
rect 42809 95625 42843 95659
rect 43361 95625 43395 95659
rect 44741 95625 44775 95659
rect 50813 95625 50847 95659
rect 56517 95625 56551 95659
rect 57161 95625 57195 95659
rect 57989 95625 58023 95659
rect 59185 95625 59219 95659
rect 61117 95625 61151 95659
rect 62405 95625 62439 95659
rect 63693 95625 63727 95659
rect 65165 95625 65199 95659
rect 65625 95625 65659 95659
rect 66913 95625 66947 95659
rect 67649 95625 67683 95659
rect 68845 95625 68879 95659
rect 70501 95625 70535 95659
rect 71789 95625 71823 95659
rect 72433 95625 72467 95659
rect 73721 95625 73755 95659
rect 75009 95625 75043 95659
rect 75561 95625 75595 95659
rect 76941 95625 76975 95659
rect 78229 95625 78263 95659
rect 79517 95625 79551 95659
rect 80161 95625 80195 95659
rect 81449 95625 81483 95659
rect 82737 95625 82771 95659
rect 15025 95557 15059 95591
rect 22845 95557 22879 95591
rect 26065 95557 26099 95591
rect 27353 95557 27387 95591
rect 55689 95557 55723 95591
rect 55873 95557 55907 95591
rect 62773 95557 62807 95591
rect 65993 95557 66027 95591
rect 67281 95557 67315 95591
rect 8493 95489 8527 95523
rect 15577 95489 15611 95523
rect 15945 95489 15979 95523
rect 16865 95489 16899 95523
rect 18153 95489 18187 95523
rect 19441 95489 19475 95523
rect 20361 95489 20395 95523
rect 21373 95489 21407 95523
rect 23305 95489 23339 95523
rect 24593 95489 24627 95523
rect 27813 95489 27847 95523
rect 29285 95489 29319 95523
rect 30389 95489 30423 95523
rect 31309 95489 31343 95523
rect 32321 95489 32355 95523
rect 33609 95489 33643 95523
rect 34897 95489 34931 95523
rect 35817 95489 35851 95523
rect 36829 95489 36863 95523
rect 38117 95489 38151 95523
rect 39037 95489 39071 95523
rect 40049 95489 40083 95523
rect 41337 95489 41371 95523
rect 42625 95489 42659 95523
rect 43545 95489 43579 95523
rect 44557 95489 44591 95523
rect 50997 95489 51031 95523
rect 52745 95489 52779 95523
rect 56425 95489 56459 95523
rect 57069 95489 57103 95523
rect 58081 95489 58115 95523
rect 59369 95489 59403 95523
rect 60013 95489 60047 95523
rect 60473 95489 60507 95523
rect 61301 95489 61335 95523
rect 63877 95489 63911 95523
rect 65073 95489 65107 95523
rect 67741 95489 67775 95523
rect 69213 95489 69247 95523
rect 70317 95489 70351 95523
rect 71605 95489 71639 95523
rect 72249 95489 72283 95523
rect 73537 95489 73571 95523
rect 74825 95489 74859 95523
rect 75745 95489 75779 95523
rect 76757 95489 76791 95523
rect 78045 95489 78079 95523
rect 79333 95489 79367 95523
rect 79977 95489 80011 95523
rect 81265 95489 81299 95523
rect 82553 95489 82587 95523
rect 19625 95421 19659 95455
rect 23581 95421 23615 95455
rect 52193 95421 52227 95455
rect 52469 95421 52503 95455
rect 53757 95421 53791 95455
rect 54217 95421 54251 95455
rect 59553 95421 59587 95455
rect 64153 95421 64187 95455
rect 22661 95353 22695 95387
rect 25881 95353 25915 95387
rect 27169 95353 27203 95387
rect 62589 95353 62623 95387
rect 65809 95353 65843 95387
rect 67097 95353 67131 95387
rect 15117 95285 15151 95319
rect 15761 95285 15795 95319
rect 17049 95285 17083 95319
rect 18337 95285 18371 95319
rect 20177 95285 20211 95319
rect 21557 95285 21591 95319
rect 24777 95285 24811 95319
rect 27997 95285 28031 95319
rect 29101 95285 29135 95319
rect 55413 95285 55447 95319
rect 56241 95285 56275 95319
rect 56885 95285 56919 95319
rect 58265 95285 58299 95319
rect 60197 95285 60231 95319
rect 61485 95285 61519 95319
rect 64889 95285 64923 95319
rect 67925 95285 67959 95319
rect 69029 95285 69063 95319
rect 52561 95081 52595 95115
rect 88441 94197 88475 94231
rect 87889 93925 87923 93959
rect 88349 93857 88383 93891
rect 88533 93857 88567 93891
rect 88073 93653 88107 93687
rect 88073 93177 88107 93211
rect 88349 93177 88383 93211
rect 87337 93109 87371 93143
rect 87705 93109 87739 93143
rect 87889 93109 87923 93143
rect 88441 93109 88475 93143
rect 87705 92837 87739 92871
rect 86785 92769 86819 92803
rect 86509 92701 86543 92735
rect 87521 92701 87555 92735
rect 87889 92701 87923 92735
rect 87981 92701 88015 92735
rect 88257 92701 88291 92735
rect 87153 92633 87187 92667
rect 87429 92633 87463 92667
rect 86601 92565 86635 92599
rect 87061 92565 87095 92599
rect 88165 92565 88199 92599
rect 88441 92565 88475 92599
rect 31953 92225 31987 92259
rect 53113 92225 53147 92259
rect 87245 92225 87279 92259
rect 87521 92225 87555 92259
rect 87797 92225 87831 92259
rect 88165 92225 88199 92259
rect 88441 92225 88475 92259
rect 51917 92157 51951 92191
rect 52929 92157 52963 92191
rect 86233 92157 86267 92191
rect 32413 92089 32447 92123
rect 52745 92089 52779 92123
rect 87981 92089 88015 92123
rect 88257 92089 88291 92123
rect 30481 92021 30515 92055
rect 32229 92021 32263 92055
rect 52561 92021 52595 92055
rect 85681 92021 85715 92055
rect 85957 92021 85991 92055
rect 86049 92021 86083 92055
rect 86509 92021 86543 92055
rect 86693 92021 86727 92055
rect 86785 92021 86819 92055
rect 87061 92021 87095 92055
rect 87337 92021 87371 92055
rect 87613 92021 87647 92055
rect 50261 91817 50295 91851
rect 86049 91817 86083 91851
rect 86969 91749 87003 91783
rect 32229 91613 32263 91647
rect 51181 91613 51215 91647
rect 52745 91613 52779 91647
rect 54401 91613 54435 91647
rect 85681 91613 85715 91647
rect 86693 91613 86727 91647
rect 86785 91613 86819 91647
rect 88073 91613 88107 91647
rect 10333 91545 10367 91579
rect 30389 91545 30423 91579
rect 31953 91545 31987 91579
rect 32505 91545 32539 91579
rect 50813 91545 50847 91579
rect 52377 91545 52411 91579
rect 53849 91545 53883 91579
rect 54585 91545 54619 91579
rect 85221 91545 85255 91579
rect 87153 91545 87187 91579
rect 87337 91545 87371 91579
rect 87521 91545 87555 91579
rect 87705 91545 87739 91579
rect 88257 91545 88291 91579
rect 88441 91545 88475 91579
rect 11621 91477 11655 91511
rect 12541 91477 12575 91511
rect 13553 91477 13587 91511
rect 49709 91477 49743 91511
rect 51089 91477 51123 91511
rect 54217 91477 54251 91511
rect 85037 91477 85071 91511
rect 85405 91477 85439 91511
rect 85773 91477 85807 91511
rect 86325 91477 86359 91511
rect 86509 91477 86543 91511
rect 87981 91477 88015 91511
rect 1685 86785 1719 86819
rect 1501 86581 1535 86615
rect 1501 85221 1535 85255
rect 1685 85085 1719 85119
rect 1685 83997 1719 84031
rect 1501 83861 1535 83895
rect 1685 82433 1719 82467
rect 1501 82229 1535 82263
rect 1685 81345 1719 81379
rect 1501 81141 1535 81175
rect 1685 79645 1719 79679
rect 1501 79509 1535 79543
rect 1685 78557 1719 78591
rect 1501 78421 1535 78455
rect 1685 76993 1719 77027
rect 1501 76789 1535 76823
rect 1501 76041 1535 76075
rect 1685 75905 1719 75939
rect 1685 74205 1719 74239
rect 1501 74069 1535 74103
rect 1685 73117 1719 73151
rect 1501 72981 1535 73015
rect 1685 71553 1719 71587
rect 5181 71553 5215 71587
rect 5641 71553 5675 71587
rect 5273 71417 5307 71451
rect 5457 71417 5491 71451
rect 1501 71349 1535 71383
rect 1501 70601 1535 70635
rect 5273 70601 5307 70635
rect 5457 70601 5491 70635
rect 1685 70465 1719 70499
rect 5641 70465 5675 70499
rect 5181 70397 5215 70431
rect 1593 68901 1627 68935
rect 1409 68765 1443 68799
rect 1685 68765 1719 68799
rect 5365 68765 5399 68799
rect 5273 68697 5307 68731
rect 5549 68629 5583 68663
rect 1593 67881 1627 67915
rect 5273 67813 5307 67847
rect 5549 67813 5583 67847
rect 1409 67677 1443 67711
rect 1685 67677 1719 67711
rect 5365 67677 5399 67711
rect 1409 66113 1443 66147
rect 1685 66113 1719 66147
rect 5365 66113 5399 66147
rect 1593 65977 1627 66011
rect 5181 65909 5215 65943
rect 5549 65909 5583 65943
rect 5273 65161 5307 65195
rect 1409 65025 1443 65059
rect 1685 65025 1719 65059
rect 5365 65025 5399 65059
rect 1593 64889 1627 64923
rect 5549 64889 5583 64923
rect 1593 63461 1627 63495
rect 1409 63325 1443 63359
rect 1685 63325 1719 63359
rect 5365 63325 5399 63359
rect 5181 63189 5215 63223
rect 5549 63189 5583 63223
rect 5273 62441 5307 62475
rect 1593 62373 1627 62407
rect 1409 62237 1443 62271
rect 1685 62237 1719 62271
rect 5365 62237 5399 62271
rect 5549 62101 5583 62135
rect 1409 61761 1443 61795
rect 1685 61761 1719 61795
rect 1593 61625 1627 61659
rect 5181 60673 5215 60707
rect 5365 60673 5399 60707
rect 1409 60469 1443 60503
rect 5549 60469 5583 60503
rect 1409 60061 1443 60095
rect 1685 60061 1719 60095
rect 1593 59925 1627 59959
rect 5365 59585 5399 59619
rect 1409 59381 1443 59415
rect 5273 59381 5307 59415
rect 5549 59381 5583 59415
rect 1593 59109 1627 59143
rect 1409 58973 1443 59007
rect 1685 58973 1719 59007
rect 1409 57953 1443 57987
rect 5365 57885 5399 57919
rect 5273 57749 5307 57783
rect 5549 57749 5583 57783
rect 5457 57545 5491 57579
rect 1409 57409 1443 57443
rect 1685 57409 1719 57443
rect 1593 57273 1627 57307
rect 5549 57205 5583 57239
rect 1409 56797 1443 56831
rect 5641 56797 5675 56831
rect 4353 56661 4387 56695
rect 1409 56321 1443 56355
rect 1685 56321 1719 56355
rect 5365 56321 5399 56355
rect 1593 56185 1627 56219
rect 5181 56117 5215 56151
rect 5549 56117 5583 56151
rect 5181 55369 5215 55403
rect 5549 55369 5583 55403
rect 5365 55233 5399 55267
rect 1409 55029 1443 55063
rect 1409 54621 1443 54655
rect 1685 54621 1719 54655
rect 1593 54485 1627 54519
rect 5365 54145 5399 54179
rect 1409 53941 1443 53975
rect 5181 53941 5215 53975
rect 5549 53941 5583 53975
rect 1593 53669 1627 53703
rect 1409 53533 1443 53567
rect 1685 53533 1719 53567
rect 5549 52581 5583 52615
rect 1409 52445 1443 52479
rect 5181 52445 5215 52479
rect 5365 52445 5399 52479
rect 1409 51901 1443 51935
rect 1409 51357 1443 51391
rect 5365 51357 5399 51391
rect 5273 51221 5307 51255
rect 5549 51221 5583 51255
rect 4905 50881 4939 50915
rect 5365 50881 5399 50915
rect 5089 50813 5123 50847
rect 5273 50745 5307 50779
rect 1409 50677 1443 50711
rect 5549 50677 5583 50711
rect 5457 50269 5491 50303
rect 5641 50133 5675 50167
rect 1409 49589 1443 49623
rect 1409 49317 1443 49351
rect 1593 48841 1627 48875
rect 1409 48705 1443 48739
rect 1685 48705 1719 48739
rect 1409 48093 1443 48127
rect 5549 47209 5583 47243
rect 1409 47005 1443 47039
rect 5273 47005 5307 47039
rect 5457 46937 5491 46971
rect 1409 46325 1443 46359
rect 5273 46053 5307 46087
rect 5641 46053 5675 46087
rect 1685 45917 1719 45951
rect 5089 45849 5123 45883
rect 5457 45849 5491 45883
rect 1501 45781 1535 45815
rect 1409 45237 1443 45271
rect 5273 44489 5307 44523
rect 5457 44489 5491 44523
rect 1685 44353 1719 44387
rect 5089 44353 5123 44387
rect 5641 44353 5675 44387
rect 1501 44217 1535 44251
rect 1777 43945 1811 43979
rect 1501 43673 1535 43707
rect 1961 43673 1995 43707
rect 5273 43401 5307 43435
rect 5457 43401 5491 43435
rect 1685 43265 1719 43299
rect 5089 43265 5123 43299
rect 5549 43265 5583 43299
rect 1501 43061 1535 43095
rect 5089 41769 5123 41803
rect 5273 41701 5307 41735
rect 5641 41701 5675 41735
rect 1685 41565 1719 41599
rect 5457 41497 5491 41531
rect 1501 41429 1535 41463
rect 4997 40681 5031 40715
rect 5273 40681 5307 40715
rect 5549 40681 5583 40715
rect 1685 40477 1719 40511
rect 5457 40409 5491 40443
rect 1501 40341 1535 40375
rect 5273 39049 5307 39083
rect 5457 39049 5491 39083
rect 1685 38913 1719 38947
rect 5181 38913 5215 38947
rect 5641 38913 5675 38947
rect 1501 38709 1535 38743
rect 5273 37961 5307 37995
rect 5457 37961 5491 37995
rect 1685 37825 1719 37859
rect 5089 37825 5123 37859
rect 5549 37825 5583 37859
rect 1501 37621 1535 37655
rect 5273 36329 5307 36363
rect 5641 36329 5675 36363
rect 1501 36261 1535 36295
rect 1685 36125 1719 36159
rect 5181 36125 5215 36159
rect 5457 36125 5491 36159
rect 1685 35037 1719 35071
rect 5181 35037 5215 35071
rect 5457 35037 5491 35071
rect 1501 34901 1535 34935
rect 5273 34901 5307 34935
rect 5641 34901 5675 34935
rect 1685 33473 1719 33507
rect 5181 33473 5215 33507
rect 5641 33473 5675 33507
rect 1501 33269 1535 33303
rect 5365 33269 5399 33303
rect 5457 33269 5491 33303
rect 5089 32521 5123 32555
rect 1685 32385 1719 32419
rect 5641 32385 5675 32419
rect 1501 32181 1535 32215
rect 5365 32181 5399 32215
rect 5457 32181 5491 32215
rect 5273 30889 5307 30923
rect 5457 30889 5491 30923
rect 1501 30821 1535 30855
rect 1685 30685 1719 30719
rect 5181 30685 5215 30719
rect 5641 30685 5675 30719
rect 1685 29597 1719 29631
rect 5181 29597 5215 29631
rect 5457 29597 5491 29631
rect 1501 29461 1535 29495
rect 5365 29461 5399 29495
rect 5641 29461 5675 29495
rect 5089 28169 5123 28203
rect 5273 28169 5307 28203
rect 5457 28169 5491 28203
rect 1685 28033 1719 28067
rect 5641 28033 5675 28067
rect 1501 27829 1535 27863
rect 1593 27081 1627 27115
rect 5273 27013 5307 27047
rect 1409 26945 1443 26979
rect 1685 26945 1719 26979
rect 5365 26945 5399 26979
rect 5549 26741 5583 26775
rect 5549 25449 5583 25483
rect 1593 25381 1627 25415
rect 1409 25245 1443 25279
rect 1685 25245 1719 25279
rect 5365 25245 5399 25279
rect 5273 25109 5307 25143
rect 1593 24293 1627 24327
rect 1409 24157 1443 24191
rect 1685 24157 1719 24191
rect 1409 22593 1443 22627
rect 1685 22593 1719 22627
rect 1593 22457 1627 22491
rect 1593 21641 1627 21675
rect 1409 21505 1443 21539
rect 1685 21505 1719 21539
rect 1593 20009 1627 20043
rect 1409 19805 1443 19839
rect 1685 19805 1719 19839
rect 1593 18853 1627 18887
rect 1409 18717 1443 18751
rect 1685 18717 1719 18751
rect 1409 17153 1443 17187
rect 1685 17153 1719 17187
rect 1593 17017 1627 17051
rect 1593 16201 1627 16235
rect 1409 16065 1443 16099
rect 1685 16065 1719 16099
rect 1593 14569 1627 14603
rect 1409 14365 1443 14399
rect 1685 14365 1719 14399
rect 1593 13413 1627 13447
rect 1409 13277 1443 13311
rect 1685 13277 1719 13311
rect 1409 11713 1443 11747
rect 1685 11713 1719 11747
rect 1593 11577 1627 11611
rect 10885 5865 10919 5899
rect 13001 5865 13035 5899
rect 49709 5865 49743 5899
rect 50261 5865 50295 5899
rect 50813 5865 50847 5899
rect 84761 5865 84795 5899
rect 85313 5865 85347 5899
rect 86325 5865 86359 5899
rect 86601 5865 86635 5899
rect 88073 5865 88107 5899
rect 88441 5865 88475 5899
rect 53573 5797 53607 5831
rect 85129 5797 85163 5831
rect 85865 5797 85899 5831
rect 86969 5797 87003 5831
rect 87705 5797 87739 5831
rect 51365 5729 51399 5763
rect 85773 5729 85807 5763
rect 9781 5661 9815 5695
rect 52469 5661 52503 5695
rect 86049 5661 86083 5695
rect 86417 5661 86451 5695
rect 86785 5661 86819 5695
rect 87153 5661 87187 5695
rect 87521 5661 87555 5695
rect 87889 5661 87923 5695
rect 88257 5661 88291 5695
rect 11989 5593 12023 5627
rect 51917 5593 51951 5627
rect 85589 5593 85623 5627
rect 53021 5525 53055 5559
rect 85037 5525 85071 5559
rect 87337 5525 87371 5559
rect 85865 5321 85899 5355
rect 86049 5321 86083 5355
rect 86509 5321 86543 5355
rect 86693 5321 86727 5355
rect 87705 5321 87739 5355
rect 88441 5321 88475 5355
rect 86325 5253 86359 5287
rect 86969 5185 87003 5219
rect 87153 5185 87187 5219
rect 87521 5185 87555 5219
rect 87889 5185 87923 5219
rect 88257 5185 88291 5219
rect 86785 5117 86819 5151
rect 85681 5049 85715 5083
rect 88073 5049 88107 5083
rect 87337 4981 87371 5015
rect 86785 4777 86819 4811
rect 87245 4777 87279 4811
rect 87429 4777 87463 4811
rect 88441 4777 88475 4811
rect 87705 4709 87739 4743
rect 88073 4709 88107 4743
rect 87613 4641 87647 4675
rect 87889 4573 87923 4607
rect 88257 4573 88291 4607
rect 86601 4505 86635 4539
rect 86969 4505 87003 4539
rect 86417 4437 86451 4471
rect 88165 4233 88199 4267
rect 8033 2601 8067 2635
rect 11621 2601 11655 2635
rect 13369 2601 13403 2635
rect 15117 2601 15151 2635
rect 31033 2601 31067 2635
rect 31861 2601 31895 2635
rect 32965 2601 32999 2635
rect 34253 2601 34287 2635
rect 35081 2601 35115 2635
rect 36185 2601 36219 2635
rect 37473 2601 37507 2635
rect 42809 2601 42843 2635
rect 45201 2601 45235 2635
rect 70961 2601 70995 2635
rect 71789 2601 71823 2635
rect 72893 2601 72927 2635
rect 74181 2601 74215 2635
rect 75469 2601 75503 2635
rect 76297 2601 76331 2635
rect 77401 2601 77435 2635
rect 8493 2533 8527 2567
rect 39865 2533 39899 2567
rect 40693 2533 40727 2567
rect 41981 2533 42015 2567
rect 43913 2533 43947 2567
rect 79609 2533 79643 2567
rect 80621 2533 80655 2567
rect 81909 2533 81943 2567
rect 83197 2533 83231 2567
rect 10609 2465 10643 2499
rect 13185 2465 13219 2499
rect 14933 2465 14967 2499
rect 39037 2465 39071 2499
rect 78965 2465 78999 2499
rect 7849 2397 7883 2431
rect 8677 2397 8711 2431
rect 15577 2397 15611 2431
rect 16497 2397 16531 2431
rect 17509 2397 17543 2431
rect 18797 2397 18831 2431
rect 19717 2397 19751 2431
rect 20729 2397 20763 2431
rect 22017 2397 22051 2431
rect 23305 2397 23339 2431
rect 24225 2397 24259 2431
rect 25237 2397 25271 2431
rect 26525 2397 26559 2431
rect 27445 2397 27479 2431
rect 28457 2397 28491 2431
rect 29745 2397 29779 2431
rect 31217 2397 31251 2431
rect 31677 2397 31711 2431
rect 33149 2397 33183 2431
rect 34437 2397 34471 2431
rect 34897 2397 34931 2431
rect 36369 2397 36403 2431
rect 37657 2397 37691 2431
rect 38761 2397 38795 2431
rect 45385 2397 45419 2431
rect 55505 2397 55539 2431
rect 56425 2397 56459 2431
rect 57437 2397 57471 2431
rect 58725 2397 58759 2431
rect 60013 2397 60047 2431
rect 60657 2397 60691 2431
rect 61945 2397 61979 2431
rect 63233 2397 63267 2431
rect 64153 2397 64187 2431
rect 65165 2397 65199 2431
rect 66453 2397 66487 2431
rect 67741 2397 67775 2431
rect 68385 2397 68419 2431
rect 69673 2397 69707 2431
rect 71145 2397 71179 2431
rect 71605 2397 71639 2431
rect 73077 2397 73111 2431
rect 74365 2397 74399 2431
rect 75653 2397 75687 2431
rect 76113 2397 76147 2431
rect 77585 2397 77619 2431
rect 78689 2397 78723 2431
rect 11345 2329 11379 2363
rect 11805 2329 11839 2363
rect 12357 2329 12391 2363
rect 14105 2329 14139 2363
rect 40049 2329 40083 2363
rect 40233 2329 40267 2363
rect 40877 2329 40911 2363
rect 42165 2329 42199 2363
rect 42717 2329 42751 2363
rect 44097 2329 44131 2363
rect 79793 2329 79827 2363
rect 79977 2329 80011 2363
rect 80805 2329 80839 2363
rect 82093 2329 82127 2363
rect 83381 2329 83415 2363
rect 7757 2261 7791 2295
rect 8401 2261 8435 2295
rect 12265 2261 12299 2295
rect 13829 2261 13863 2295
rect 15761 2261 15795 2295
rect 16313 2261 16347 2295
rect 17693 2261 17727 2295
rect 18981 2261 19015 2295
rect 19533 2261 19567 2295
rect 20913 2261 20947 2295
rect 22201 2261 22235 2295
rect 23489 2261 23523 2295
rect 24041 2261 24075 2295
rect 25421 2261 25455 2295
rect 26709 2261 26743 2295
rect 27261 2261 27295 2295
rect 28641 2261 28675 2295
rect 29929 2261 29963 2295
rect 30941 2261 30975 2295
rect 31585 2261 31619 2295
rect 32873 2261 32907 2295
rect 34161 2261 34195 2295
rect 34805 2261 34839 2295
rect 36093 2261 36127 2295
rect 37381 2261 37415 2295
rect 38669 2261 38703 2295
rect 40601 2261 40635 2295
rect 41889 2261 41923 2295
rect 42533 2261 42567 2295
rect 43821 2261 43855 2295
rect 45109 2261 45143 2295
rect 55689 2261 55723 2295
rect 56241 2261 56275 2295
rect 57621 2261 57655 2295
rect 58909 2261 58943 2295
rect 60197 2261 60231 2295
rect 60841 2261 60875 2295
rect 62129 2261 62163 2295
rect 63417 2261 63451 2295
rect 63969 2261 64003 2295
rect 65349 2261 65383 2295
rect 66637 2261 66671 2295
rect 67925 2261 67959 2295
rect 68569 2261 68603 2295
rect 69857 2261 69891 2295
rect 70869 2261 70903 2295
rect 71513 2261 71547 2295
rect 72801 2261 72835 2295
rect 74089 2261 74123 2295
rect 75377 2261 75411 2295
rect 76021 2261 76055 2295
rect 77309 2261 77343 2295
rect 78597 2261 78631 2295
rect 80529 2261 80563 2295
rect 81817 2261 81851 2295
rect 83105 2261 83139 2295
<< metal1 >>
rect 1104 95770 88872 95792
rect 1104 95718 37610 95770
rect 37662 95718 37674 95770
rect 37726 95718 37738 95770
rect 37790 95718 37802 95770
rect 37854 95718 37866 95770
rect 37918 95718 73610 95770
rect 73662 95718 73674 95770
rect 73726 95718 73738 95770
rect 73790 95718 73802 95770
rect 73854 95718 73866 95770
rect 73918 95718 88872 95770
rect 1104 95696 88872 95718
rect 8662 95616 8668 95668
rect 8720 95616 8726 95668
rect 14734 95616 14740 95668
rect 14792 95656 14798 95668
rect 14792 95628 15056 95656
rect 14792 95616 14798 95628
rect 15028 95597 15056 95628
rect 16666 95616 16672 95668
rect 16724 95616 16730 95668
rect 17954 95616 17960 95668
rect 18012 95616 18018 95668
rect 19337 95659 19395 95665
rect 19337 95625 19349 95659
rect 19383 95656 19395 95659
rect 19426 95656 19432 95668
rect 19383 95628 19432 95656
rect 19383 95625 19395 95628
rect 19337 95619 19395 95625
rect 19426 95616 19432 95628
rect 19484 95616 19490 95668
rect 20346 95616 20352 95668
rect 20404 95656 20410 95668
rect 20441 95659 20499 95665
rect 20441 95656 20453 95659
rect 20404 95628 20453 95656
rect 20404 95616 20410 95628
rect 20441 95625 20453 95628
rect 20487 95625 20499 95659
rect 20441 95619 20499 95625
rect 21174 95616 21180 95668
rect 21232 95616 21238 95668
rect 22462 95616 22468 95668
rect 22520 95656 22526 95668
rect 22520 95628 22876 95656
rect 22520 95616 22526 95628
rect 15013 95591 15071 95597
rect 15013 95557 15025 95591
rect 15059 95557 15071 95591
rect 15013 95551 15071 95557
rect 8478 95480 8484 95532
rect 8536 95480 8542 95532
rect 15562 95480 15568 95532
rect 15620 95520 15626 95532
rect 15933 95523 15991 95529
rect 15933 95520 15945 95523
rect 15620 95492 15945 95520
rect 15620 95480 15626 95492
rect 15933 95489 15945 95492
rect 15979 95489 15991 95523
rect 16684 95520 16712 95616
rect 16853 95523 16911 95529
rect 16853 95520 16865 95523
rect 16684 95492 16865 95520
rect 15933 95483 15991 95489
rect 16853 95489 16865 95492
rect 16899 95489 16911 95523
rect 17972 95520 18000 95616
rect 19444 95529 19472 95616
rect 20364 95529 20392 95616
rect 18141 95523 18199 95529
rect 18141 95520 18153 95523
rect 17972 95492 18153 95520
rect 16853 95483 16911 95489
rect 18141 95489 18153 95492
rect 18187 95489 18199 95523
rect 18141 95483 18199 95489
rect 19429 95523 19487 95529
rect 19429 95489 19441 95523
rect 19475 95489 19487 95523
rect 19429 95483 19487 95489
rect 20349 95523 20407 95529
rect 20349 95489 20361 95523
rect 20395 95489 20407 95523
rect 21192 95520 21220 95616
rect 22848 95597 22876 95628
rect 23106 95616 23112 95668
rect 23164 95616 23170 95668
rect 24394 95616 24400 95668
rect 24452 95616 24458 95668
rect 25682 95616 25688 95668
rect 25740 95656 25746 95668
rect 25740 95628 26096 95656
rect 25740 95616 25746 95628
rect 22833 95591 22891 95597
rect 22833 95557 22845 95591
rect 22879 95557 22891 95591
rect 22833 95551 22891 95557
rect 21361 95523 21419 95529
rect 21361 95520 21373 95523
rect 21192 95492 21373 95520
rect 20349 95483 20407 95489
rect 21361 95489 21373 95492
rect 21407 95489 21419 95523
rect 23124 95520 23152 95616
rect 23293 95523 23351 95529
rect 23293 95520 23305 95523
rect 23124 95492 23305 95520
rect 21361 95483 21419 95489
rect 23293 95489 23305 95492
rect 23339 95489 23351 95523
rect 24412 95520 24440 95616
rect 26068 95597 26096 95628
rect 26970 95616 26976 95668
rect 27028 95656 27034 95668
rect 27028 95628 27384 95656
rect 27028 95616 27034 95628
rect 27356 95597 27384 95628
rect 27614 95616 27620 95668
rect 27672 95616 27678 95668
rect 28997 95659 29055 95665
rect 28997 95625 29009 95659
rect 29043 95656 29055 95659
rect 29086 95656 29092 95668
rect 29043 95628 29092 95656
rect 29043 95625 29055 95628
rect 28997 95619 29055 95625
rect 29086 95616 29092 95628
rect 29144 95616 29150 95668
rect 30190 95616 30196 95668
rect 30248 95656 30254 95668
rect 30561 95659 30619 95665
rect 30561 95656 30573 95659
rect 30248 95628 30573 95656
rect 30248 95616 30254 95628
rect 30561 95625 30573 95628
rect 30607 95625 30619 95659
rect 30561 95619 30619 95625
rect 31110 95616 31116 95668
rect 31168 95616 31174 95668
rect 32490 95616 32496 95668
rect 32548 95616 32554 95668
rect 33778 95616 33784 95668
rect 33836 95616 33842 95668
rect 35066 95616 35072 95668
rect 35124 95616 35130 95668
rect 35618 95616 35624 95668
rect 35676 95616 35682 95668
rect 36998 95616 37004 95668
rect 37056 95616 37062 95668
rect 38286 95616 38292 95668
rect 38344 95616 38350 95668
rect 38838 95616 38844 95668
rect 38896 95616 38902 95668
rect 39850 95616 39856 95668
rect 39908 95656 39914 95668
rect 40221 95659 40279 95665
rect 40221 95656 40233 95659
rect 39908 95628 40233 95656
rect 39908 95616 39914 95628
rect 40221 95625 40233 95628
rect 40267 95625 40279 95659
rect 40221 95619 40279 95625
rect 41322 95616 41328 95668
rect 41380 95656 41386 95668
rect 41509 95659 41567 95665
rect 41509 95656 41521 95659
rect 41380 95628 41521 95656
rect 41380 95616 41386 95628
rect 41509 95625 41521 95628
rect 41555 95625 41567 95659
rect 41509 95619 41567 95625
rect 42702 95616 42708 95668
rect 42760 95656 42766 95668
rect 42797 95659 42855 95665
rect 42797 95656 42809 95659
rect 42760 95628 42809 95656
rect 42760 95616 42766 95628
rect 42797 95625 42809 95628
rect 42843 95625 42855 95659
rect 42797 95619 42855 95625
rect 43346 95616 43352 95668
rect 43404 95616 43410 95668
rect 44726 95616 44732 95668
rect 44784 95616 44790 95668
rect 50798 95616 50804 95668
rect 50856 95616 50862 95668
rect 56410 95616 56416 95668
rect 56468 95656 56474 95668
rect 56505 95659 56563 95665
rect 56505 95656 56517 95659
rect 56468 95628 56517 95656
rect 56468 95616 56474 95628
rect 56505 95625 56517 95628
rect 56551 95625 56563 95659
rect 56505 95619 56563 95625
rect 56962 95616 56968 95668
rect 57020 95656 57026 95668
rect 57149 95659 57207 95665
rect 57149 95656 57161 95659
rect 57020 95628 57161 95656
rect 57020 95616 57026 95628
rect 26053 95591 26111 95597
rect 26053 95557 26065 95591
rect 26099 95557 26111 95591
rect 26053 95551 26111 95557
rect 27341 95591 27399 95597
rect 27341 95557 27353 95591
rect 27387 95557 27399 95591
rect 27341 95551 27399 95557
rect 24581 95523 24639 95529
rect 24581 95520 24593 95523
rect 24412 95492 24593 95520
rect 23293 95483 23351 95489
rect 24581 95489 24593 95492
rect 24627 95489 24639 95523
rect 27632 95520 27660 95616
rect 27801 95523 27859 95529
rect 27801 95520 27813 95523
rect 27632 95492 27813 95520
rect 24581 95483 24639 95489
rect 27801 95489 27813 95492
rect 27847 95489 27859 95523
rect 29104 95520 29132 95616
rect 29273 95523 29331 95529
rect 29273 95520 29285 95523
rect 29104 95492 29285 95520
rect 27801 95483 27859 95489
rect 29273 95489 29285 95492
rect 29319 95489 29331 95523
rect 29273 95483 29331 95489
rect 30098 95480 30104 95532
rect 30156 95520 30162 95532
rect 30377 95523 30435 95529
rect 30377 95520 30389 95523
rect 30156 95492 30389 95520
rect 30156 95480 30162 95492
rect 30377 95489 30389 95492
rect 30423 95489 30435 95523
rect 30377 95483 30435 95489
rect 31294 95480 31300 95532
rect 31352 95480 31358 95532
rect 32306 95480 32312 95532
rect 32364 95480 32370 95532
rect 33594 95480 33600 95532
rect 33652 95480 33658 95532
rect 34882 95480 34888 95532
rect 34940 95480 34946 95532
rect 35802 95480 35808 95532
rect 35860 95480 35866 95532
rect 36814 95480 36820 95532
rect 36872 95480 36878 95532
rect 38102 95480 38108 95532
rect 38160 95480 38166 95532
rect 39022 95480 39028 95532
rect 39080 95480 39086 95532
rect 40034 95480 40040 95532
rect 40092 95480 40098 95532
rect 41322 95480 41328 95532
rect 41380 95480 41386 95532
rect 42610 95480 42616 95532
rect 42668 95480 42674 95532
rect 43530 95480 43536 95532
rect 43588 95480 43594 95532
rect 44542 95480 44548 95532
rect 44600 95480 44606 95532
rect 50816 95520 50844 95616
rect 54938 95548 54944 95600
rect 54996 95588 55002 95600
rect 55677 95591 55735 95597
rect 55677 95588 55689 95591
rect 54996 95560 55689 95588
rect 54996 95548 55002 95560
rect 55677 95557 55689 95560
rect 55723 95588 55735 95591
rect 55861 95591 55919 95597
rect 55861 95588 55873 95591
rect 55723 95560 55873 95588
rect 55723 95557 55735 95560
rect 55677 95551 55735 95557
rect 55861 95557 55873 95560
rect 55907 95557 55919 95591
rect 55861 95551 55919 95557
rect 50985 95523 51043 95529
rect 50985 95520 50997 95523
rect 50816 95492 50997 95520
rect 50985 95489 50997 95492
rect 51031 95489 51043 95523
rect 50985 95483 51043 95489
rect 52270 95480 52276 95532
rect 52328 95520 52334 95532
rect 56428 95529 56456 95616
rect 57072 95529 57100 95628
rect 57149 95625 57161 95628
rect 57195 95625 57207 95659
rect 57149 95619 57207 95625
rect 57977 95659 58035 95665
rect 57977 95625 57989 95659
rect 58023 95656 58035 95659
rect 58066 95656 58072 95668
rect 58023 95628 58072 95656
rect 58023 95625 58035 95628
rect 57977 95619 58035 95625
rect 58066 95616 58072 95628
rect 58124 95616 58130 95668
rect 59170 95616 59176 95668
rect 59228 95616 59234 95668
rect 61102 95616 61108 95668
rect 61160 95616 61166 95668
rect 62390 95616 62396 95668
rect 62448 95656 62454 95668
rect 62448 95628 62804 95656
rect 62448 95616 62454 95628
rect 58084 95529 58112 95616
rect 52733 95523 52791 95529
rect 52733 95520 52745 95523
rect 52328 95492 52745 95520
rect 52328 95480 52334 95492
rect 52733 95489 52745 95492
rect 52779 95489 52791 95523
rect 52733 95483 52791 95489
rect 56413 95523 56471 95529
rect 56413 95489 56425 95523
rect 56459 95489 56471 95523
rect 56413 95483 56471 95489
rect 57057 95523 57115 95529
rect 57057 95489 57069 95523
rect 57103 95489 57115 95523
rect 57057 95483 57115 95489
rect 58069 95523 58127 95529
rect 58069 95489 58081 95523
rect 58115 95489 58127 95523
rect 59188 95520 59216 95616
rect 59357 95523 59415 95529
rect 59357 95520 59369 95523
rect 59188 95492 59369 95520
rect 58069 95483 58127 95489
rect 59357 95489 59369 95492
rect 59403 95489 59415 95523
rect 59357 95483 59415 95489
rect 59998 95480 60004 95532
rect 60056 95520 60062 95532
rect 60461 95523 60519 95529
rect 60461 95520 60473 95523
rect 60056 95492 60473 95520
rect 60056 95480 60062 95492
rect 60461 95489 60473 95492
rect 60507 95489 60519 95523
rect 61120 95520 61148 95616
rect 62776 95597 62804 95628
rect 63678 95616 63684 95668
rect 63736 95616 63742 95668
rect 64598 95616 64604 95668
rect 64656 95656 64662 95668
rect 65153 95659 65211 95665
rect 65153 95656 65165 95659
rect 64656 95628 65165 95656
rect 64656 95616 64662 95628
rect 62761 95591 62819 95597
rect 62761 95557 62773 95591
rect 62807 95557 62819 95591
rect 62761 95551 62819 95557
rect 61289 95523 61347 95529
rect 61289 95520 61301 95523
rect 61120 95492 61301 95520
rect 60461 95483 60519 95489
rect 61289 95489 61301 95492
rect 61335 95489 61347 95523
rect 63696 95520 63724 95616
rect 65076 95529 65104 95628
rect 65153 95625 65165 95628
rect 65199 95625 65211 95659
rect 65153 95619 65211 95625
rect 65610 95616 65616 95668
rect 65668 95656 65674 95668
rect 65668 95628 66024 95656
rect 65668 95616 65674 95628
rect 65996 95597 66024 95628
rect 66898 95616 66904 95668
rect 66956 95656 66962 95668
rect 67637 95659 67695 95665
rect 66956 95628 67312 95656
rect 66956 95616 66962 95628
rect 67284 95597 67312 95628
rect 67637 95625 67649 95659
rect 67683 95656 67695 95659
rect 67726 95656 67732 95668
rect 67683 95628 67732 95656
rect 67683 95625 67695 95628
rect 67637 95619 67695 95625
rect 67726 95616 67732 95628
rect 67784 95616 67790 95668
rect 68830 95616 68836 95668
rect 68888 95616 68894 95668
rect 70302 95616 70308 95668
rect 70360 95656 70366 95668
rect 70489 95659 70547 95665
rect 70489 95656 70501 95659
rect 70360 95628 70501 95656
rect 70360 95616 70366 95628
rect 70489 95625 70501 95628
rect 70535 95625 70547 95659
rect 70489 95619 70547 95625
rect 71682 95616 71688 95668
rect 71740 95656 71746 95668
rect 71777 95659 71835 95665
rect 71777 95656 71789 95659
rect 71740 95628 71789 95656
rect 71740 95616 71746 95628
rect 71777 95625 71789 95628
rect 71823 95625 71835 95659
rect 71777 95619 71835 95625
rect 72418 95616 72424 95668
rect 72476 95616 72482 95668
rect 73522 95616 73528 95668
rect 73580 95656 73586 95668
rect 73709 95659 73767 95665
rect 73709 95656 73721 95659
rect 73580 95628 73721 95656
rect 73580 95616 73586 95628
rect 73709 95625 73721 95628
rect 73755 95625 73767 95659
rect 73709 95619 73767 95625
rect 74994 95616 75000 95668
rect 75052 95616 75058 95668
rect 75546 95616 75552 95668
rect 75604 95616 75610 95668
rect 76926 95616 76932 95668
rect 76984 95616 76990 95668
rect 78214 95616 78220 95668
rect 78272 95616 78278 95668
rect 79502 95616 79508 95668
rect 79560 95616 79566 95668
rect 79962 95616 79968 95668
rect 80020 95656 80026 95668
rect 80149 95659 80207 95665
rect 80149 95656 80161 95659
rect 80020 95628 80161 95656
rect 80020 95616 80026 95628
rect 80149 95625 80161 95628
rect 80195 95625 80207 95659
rect 80149 95619 80207 95625
rect 81342 95616 81348 95668
rect 81400 95656 81406 95668
rect 81437 95659 81495 95665
rect 81437 95656 81449 95659
rect 81400 95628 81449 95656
rect 81400 95616 81406 95628
rect 81437 95625 81449 95628
rect 81483 95625 81495 95659
rect 81437 95619 81495 95625
rect 82722 95616 82728 95668
rect 82780 95616 82786 95668
rect 65981 95591 66039 95597
rect 65981 95557 65993 95591
rect 66027 95557 66039 95591
rect 65981 95551 66039 95557
rect 67269 95591 67327 95597
rect 67269 95557 67281 95591
rect 67315 95557 67327 95591
rect 67269 95551 67327 95557
rect 67744 95529 67772 95616
rect 63865 95523 63923 95529
rect 63865 95520 63877 95523
rect 63696 95492 63877 95520
rect 61289 95483 61347 95489
rect 63865 95489 63877 95492
rect 63911 95489 63923 95523
rect 63865 95483 63923 95489
rect 65061 95523 65119 95529
rect 65061 95489 65073 95523
rect 65107 95489 65119 95523
rect 65061 95483 65119 95489
rect 67729 95523 67787 95529
rect 67729 95489 67741 95523
rect 67775 95489 67787 95523
rect 68848 95520 68876 95616
rect 69201 95523 69259 95529
rect 69201 95520 69213 95523
rect 68848 95492 69213 95520
rect 67729 95483 67787 95489
rect 69201 95489 69213 95492
rect 69247 95489 69259 95523
rect 69201 95483 69259 95489
rect 70302 95480 70308 95532
rect 70360 95480 70366 95532
rect 71222 95480 71228 95532
rect 71280 95520 71286 95532
rect 71593 95523 71651 95529
rect 71593 95520 71605 95523
rect 71280 95492 71605 95520
rect 71280 95480 71286 95492
rect 71593 95489 71605 95492
rect 71639 95489 71651 95523
rect 71593 95483 71651 95489
rect 72234 95480 72240 95532
rect 72292 95480 72298 95532
rect 73522 95480 73528 95532
rect 73580 95480 73586 95532
rect 74810 95480 74816 95532
rect 74868 95480 74874 95532
rect 75730 95480 75736 95532
rect 75788 95480 75794 95532
rect 76742 95480 76748 95532
rect 76800 95480 76806 95532
rect 78030 95480 78036 95532
rect 78088 95480 78094 95532
rect 78950 95480 78956 95532
rect 79008 95520 79014 95532
rect 79321 95523 79379 95529
rect 79321 95520 79333 95523
rect 79008 95492 79333 95520
rect 79008 95480 79014 95492
rect 79321 95489 79333 95492
rect 79367 95489 79379 95523
rect 79321 95483 79379 95489
rect 79965 95523 80023 95529
rect 79965 95489 79977 95523
rect 80011 95520 80023 95523
rect 80054 95520 80060 95532
rect 80011 95492 80060 95520
rect 80011 95489 80023 95492
rect 79965 95483 80023 95489
rect 80054 95480 80060 95492
rect 80112 95480 80118 95532
rect 81250 95480 81256 95532
rect 81308 95480 81314 95532
rect 82538 95480 82544 95532
rect 82596 95480 82602 95532
rect 19058 95412 19064 95464
rect 19116 95452 19122 95464
rect 19613 95455 19671 95461
rect 19613 95452 19625 95455
rect 19116 95424 19625 95452
rect 19116 95412 19122 95424
rect 19613 95421 19625 95424
rect 19659 95421 19671 95455
rect 19613 95415 19671 95421
rect 23566 95412 23572 95464
rect 23624 95412 23630 95464
rect 52181 95455 52239 95461
rect 52181 95421 52193 95455
rect 52227 95452 52239 95455
rect 52362 95452 52368 95464
rect 52227 95424 52368 95452
rect 52227 95421 52239 95424
rect 52181 95415 52239 95421
rect 52362 95412 52368 95424
rect 52420 95452 52426 95464
rect 52457 95455 52515 95461
rect 52457 95452 52469 95455
rect 52420 95424 52469 95452
rect 52420 95412 52426 95424
rect 52457 95421 52469 95424
rect 52503 95421 52515 95455
rect 52457 95415 52515 95421
rect 53742 95412 53748 95464
rect 53800 95452 53806 95464
rect 54205 95455 54263 95461
rect 54205 95452 54217 95455
rect 53800 95424 54217 95452
rect 53800 95412 53806 95424
rect 54205 95421 54217 95424
rect 54251 95421 54263 95455
rect 54205 95415 54263 95421
rect 59078 95412 59084 95464
rect 59136 95452 59142 95464
rect 59541 95455 59599 95461
rect 59541 95452 59553 95455
rect 59136 95424 59553 95452
rect 59136 95412 59142 95424
rect 59541 95421 59553 95424
rect 59587 95421 59599 95455
rect 59541 95415 59599 95421
rect 63494 95412 63500 95464
rect 63552 95452 63558 95464
rect 64141 95455 64199 95461
rect 64141 95452 64153 95455
rect 63552 95424 64153 95452
rect 63552 95412 63558 95424
rect 64141 95421 64153 95424
rect 64187 95421 64199 95455
rect 64141 95415 64199 95421
rect 22646 95344 22652 95396
rect 22704 95344 22710 95396
rect 25866 95344 25872 95396
rect 25924 95344 25930 95396
rect 27154 95344 27160 95396
rect 27212 95344 27218 95396
rect 62574 95344 62580 95396
rect 62632 95344 62638 95396
rect 65794 95344 65800 95396
rect 65852 95344 65858 95396
rect 67082 95344 67088 95396
rect 67140 95344 67146 95396
rect 14642 95276 14648 95328
rect 14700 95316 14706 95328
rect 15105 95319 15163 95325
rect 15105 95316 15117 95319
rect 14700 95288 15117 95316
rect 14700 95276 14706 95288
rect 15105 95285 15117 95288
rect 15151 95285 15163 95319
rect 15105 95279 15163 95285
rect 15746 95276 15752 95328
rect 15804 95276 15810 95328
rect 17034 95276 17040 95328
rect 17092 95276 17098 95328
rect 18322 95276 18328 95328
rect 18380 95276 18386 95328
rect 20162 95276 20168 95328
rect 20220 95276 20226 95328
rect 21542 95276 21548 95328
rect 21600 95276 21606 95328
rect 24762 95276 24768 95328
rect 24820 95276 24826 95328
rect 27982 95276 27988 95328
rect 28040 95276 28046 95328
rect 29086 95276 29092 95328
rect 29144 95276 29150 95328
rect 54662 95276 54668 95328
rect 54720 95316 54726 95328
rect 55401 95319 55459 95325
rect 55401 95316 55413 95319
rect 54720 95288 55413 95316
rect 54720 95276 54726 95288
rect 55401 95285 55413 95288
rect 55447 95285 55459 95319
rect 55401 95279 55459 95285
rect 55950 95276 55956 95328
rect 56008 95316 56014 95328
rect 56229 95319 56287 95325
rect 56229 95316 56241 95319
rect 56008 95288 56241 95316
rect 56008 95276 56014 95288
rect 56229 95285 56241 95288
rect 56275 95285 56287 95319
rect 56229 95279 56287 95285
rect 56870 95276 56876 95328
rect 56928 95276 56934 95328
rect 58250 95276 58256 95328
rect 58308 95276 58314 95328
rect 60182 95276 60188 95328
rect 60240 95276 60246 95328
rect 61470 95276 61476 95328
rect 61528 95276 61534 95328
rect 64598 95276 64604 95328
rect 64656 95316 64662 95328
rect 64877 95319 64935 95325
rect 64877 95316 64889 95319
rect 64656 95288 64889 95316
rect 64656 95276 64662 95288
rect 64877 95285 64889 95288
rect 64923 95285 64935 95319
rect 64877 95279 64935 95285
rect 67910 95276 67916 95328
rect 67968 95276 67974 95328
rect 69014 95276 69020 95328
rect 69072 95276 69078 95328
rect 1104 95226 88872 95248
rect 1104 95174 36950 95226
rect 37002 95174 37014 95226
rect 37066 95174 37078 95226
rect 37130 95174 37142 95226
rect 37194 95174 37206 95226
rect 37258 95174 72950 95226
rect 73002 95174 73014 95226
rect 73066 95174 73078 95226
rect 73130 95174 73142 95226
rect 73194 95174 73206 95226
rect 73258 95174 88872 95226
rect 1104 95152 88872 95174
rect 52270 95072 52276 95124
rect 52328 95112 52334 95124
rect 52549 95115 52607 95121
rect 52549 95112 52561 95115
rect 52328 95084 52561 95112
rect 52328 95072 52334 95084
rect 52549 95081 52561 95084
rect 52595 95081 52607 95115
rect 52549 95075 52607 95081
rect 1104 94682 88872 94704
rect 1104 94630 37610 94682
rect 37662 94630 37674 94682
rect 37726 94630 37738 94682
rect 37790 94630 37802 94682
rect 37854 94630 37866 94682
rect 37918 94630 73610 94682
rect 73662 94630 73674 94682
rect 73726 94630 73738 94682
rect 73790 94630 73802 94682
rect 73854 94630 73866 94682
rect 73918 94630 88872 94682
rect 1104 94608 88872 94630
rect 88150 94188 88156 94240
rect 88208 94228 88214 94240
rect 88429 94231 88487 94237
rect 88429 94228 88441 94231
rect 88208 94200 88441 94228
rect 88208 94188 88214 94200
rect 88429 94197 88441 94200
rect 88475 94197 88487 94231
rect 88429 94191 88487 94197
rect 1104 94138 88872 94160
rect 1104 94086 36950 94138
rect 37002 94086 37014 94138
rect 37066 94086 37078 94138
rect 37130 94086 37142 94138
rect 37194 94086 37206 94138
rect 37258 94086 72950 94138
rect 73002 94086 73014 94138
rect 73066 94086 73078 94138
rect 73130 94086 73142 94138
rect 73194 94086 73206 94138
rect 73258 94086 88872 94138
rect 1104 94064 88872 94086
rect 87877 93959 87935 93965
rect 87877 93925 87889 93959
rect 87923 93956 87935 93959
rect 88610 93956 88616 93968
rect 87923 93928 88616 93956
rect 87923 93925 87935 93928
rect 87877 93919 87935 93925
rect 88610 93916 88616 93928
rect 88668 93916 88674 93968
rect 88334 93848 88340 93900
rect 88392 93848 88398 93900
rect 88518 93848 88524 93900
rect 88576 93848 88582 93900
rect 88058 93644 88064 93696
rect 88116 93644 88122 93696
rect 1104 93594 88872 93616
rect 1104 93542 37610 93594
rect 37662 93542 37674 93594
rect 37726 93542 37738 93594
rect 37790 93542 37802 93594
rect 37854 93542 37866 93594
rect 37918 93542 73610 93594
rect 73662 93542 73674 93594
rect 73726 93542 73738 93594
rect 73790 93542 73802 93594
rect 73854 93542 73866 93594
rect 73918 93542 88872 93594
rect 1104 93520 88872 93542
rect 87782 93168 87788 93220
rect 87840 93208 87846 93220
rect 88061 93211 88119 93217
rect 88061 93208 88073 93211
rect 87840 93180 88073 93208
rect 87840 93168 87846 93180
rect 88061 93177 88073 93180
rect 88107 93177 88119 93211
rect 88061 93171 88119 93177
rect 88337 93211 88395 93217
rect 88337 93177 88349 93211
rect 88383 93208 88395 93211
rect 88518 93208 88524 93220
rect 88383 93180 88524 93208
rect 88383 93177 88395 93180
rect 88337 93171 88395 93177
rect 88518 93168 88524 93180
rect 88576 93168 88582 93220
rect 87230 93100 87236 93152
rect 87288 93140 87294 93152
rect 87325 93143 87383 93149
rect 87325 93140 87337 93143
rect 87288 93112 87337 93140
rect 87288 93100 87294 93112
rect 87325 93109 87337 93112
rect 87371 93109 87383 93143
rect 87325 93103 87383 93109
rect 87690 93100 87696 93152
rect 87748 93100 87754 93152
rect 87874 93100 87880 93152
rect 87932 93100 87938 93152
rect 88429 93143 88487 93149
rect 88429 93109 88441 93143
rect 88475 93140 88487 93143
rect 88794 93140 88800 93152
rect 88475 93112 88800 93140
rect 88475 93109 88487 93112
rect 88429 93103 88487 93109
rect 88794 93100 88800 93112
rect 88852 93100 88858 93152
rect 1104 93050 88872 93072
rect 1104 92998 36950 93050
rect 37002 92998 37014 93050
rect 37066 92998 37078 93050
rect 37130 92998 37142 93050
rect 37194 92998 37206 93050
rect 37258 92998 72950 93050
rect 73002 92998 73014 93050
rect 73066 92998 73078 93050
rect 73130 92998 73142 93050
rect 73194 92998 73206 93050
rect 73258 92998 88872 93050
rect 1104 92976 88872 92998
rect 83366 92896 83372 92948
rect 83424 92936 83430 92948
rect 83424 92908 88288 92936
rect 83424 92896 83430 92908
rect 86402 92828 86408 92880
rect 86460 92868 86466 92880
rect 87693 92871 87751 92877
rect 87693 92868 87705 92871
rect 86460 92840 87705 92868
rect 86460 92828 86466 92840
rect 87693 92837 87705 92840
rect 87739 92837 87751 92871
rect 87693 92831 87751 92837
rect 86770 92760 86776 92812
rect 86828 92760 86834 92812
rect 87248 92772 88012 92800
rect 86497 92735 86555 92741
rect 86497 92701 86509 92735
rect 86543 92732 86555 92735
rect 87248 92732 87276 92772
rect 87984 92744 88012 92772
rect 86543 92704 87276 92732
rect 86543 92701 86555 92704
rect 86497 92695 86555 92701
rect 87322 92692 87328 92744
rect 87380 92732 87386 92744
rect 87509 92735 87567 92741
rect 87509 92732 87521 92735
rect 87380 92704 87521 92732
rect 87380 92692 87386 92704
rect 87509 92701 87521 92704
rect 87555 92701 87567 92735
rect 87509 92695 87567 92701
rect 87877 92735 87935 92741
rect 87877 92701 87889 92735
rect 87923 92701 87935 92735
rect 87877 92695 87935 92701
rect 87138 92624 87144 92676
rect 87196 92624 87202 92676
rect 87417 92667 87475 92673
rect 87417 92633 87429 92667
rect 87463 92664 87475 92667
rect 87598 92664 87604 92676
rect 87463 92636 87604 92664
rect 87463 92633 87475 92636
rect 87417 92627 87475 92633
rect 87598 92624 87604 92636
rect 87656 92624 87662 92676
rect 87892 92664 87920 92695
rect 87966 92692 87972 92744
rect 88024 92692 88030 92744
rect 88260 92741 88288 92908
rect 88245 92735 88303 92741
rect 88245 92701 88257 92735
rect 88291 92701 88303 92735
rect 88245 92695 88303 92701
rect 88058 92664 88064 92676
rect 87892 92636 88064 92664
rect 88058 92624 88064 92636
rect 88116 92664 88122 92676
rect 89346 92664 89352 92676
rect 88116 92636 89352 92664
rect 88116 92624 88122 92636
rect 89346 92624 89352 92636
rect 89404 92624 89410 92676
rect 86586 92556 86592 92608
rect 86644 92556 86650 92608
rect 87046 92556 87052 92608
rect 87104 92556 87110 92608
rect 87506 92556 87512 92608
rect 87564 92596 87570 92608
rect 88150 92596 88156 92608
rect 87564 92568 88156 92596
rect 87564 92556 87570 92568
rect 88150 92556 88156 92568
rect 88208 92556 88214 92608
rect 88426 92556 88432 92608
rect 88484 92556 88490 92608
rect 1104 92506 88872 92528
rect 1104 92454 37610 92506
rect 37662 92454 37674 92506
rect 37726 92454 37738 92506
rect 37790 92454 37802 92506
rect 37854 92454 37866 92506
rect 37918 92454 73610 92506
rect 73662 92454 73674 92506
rect 73726 92454 73738 92506
rect 73790 92454 73802 92506
rect 73854 92454 73866 92506
rect 73918 92454 88872 92506
rect 1104 92432 88872 92454
rect 87690 92392 87696 92404
rect 87524 92364 87696 92392
rect 31941 92259 31999 92265
rect 31941 92225 31953 92259
rect 31987 92256 31999 92259
rect 31987 92228 32444 92256
rect 31987 92225 31999 92228
rect 31941 92219 31999 92225
rect 32416 92132 32444 92228
rect 47486 92216 47492 92268
rect 47544 92256 47550 92268
rect 53101 92259 53159 92265
rect 53101 92256 53113 92259
rect 47544 92228 53113 92256
rect 47544 92216 47550 92228
rect 53101 92225 53113 92228
rect 53147 92225 53159 92259
rect 53101 92219 53159 92225
rect 87230 92216 87236 92268
rect 87288 92216 87294 92268
rect 87524 92265 87552 92364
rect 87690 92352 87696 92364
rect 87748 92392 87754 92404
rect 89254 92392 89260 92404
rect 87748 92364 89260 92392
rect 87748 92352 87754 92364
rect 89254 92352 89260 92364
rect 89312 92352 89318 92404
rect 88702 92284 88708 92336
rect 88760 92284 88766 92336
rect 87509 92259 87567 92265
rect 87509 92225 87521 92259
rect 87555 92225 87567 92259
rect 87509 92219 87567 92225
rect 87782 92216 87788 92268
rect 87840 92216 87846 92268
rect 88153 92259 88211 92265
rect 88153 92225 88165 92259
rect 88199 92225 88211 92259
rect 88153 92219 88211 92225
rect 88429 92259 88487 92265
rect 88429 92225 88441 92259
rect 88475 92256 88487 92259
rect 88720 92256 88748 92284
rect 89530 92256 89536 92268
rect 88475 92228 89536 92256
rect 88475 92225 88487 92228
rect 88429 92219 88487 92225
rect 47394 92148 47400 92200
rect 47452 92188 47458 92200
rect 51905 92191 51963 92197
rect 51905 92188 51917 92191
rect 47452 92160 51917 92188
rect 47452 92148 47458 92160
rect 51905 92157 51917 92160
rect 51951 92157 51963 92191
rect 51905 92151 51963 92157
rect 52454 92148 52460 92200
rect 52512 92188 52518 92200
rect 52917 92191 52975 92197
rect 52917 92188 52929 92191
rect 52512 92160 52929 92188
rect 52512 92148 52518 92160
rect 52917 92157 52929 92160
rect 52963 92157 52975 92191
rect 52917 92151 52975 92157
rect 86218 92148 86224 92200
rect 86276 92148 86282 92200
rect 86310 92148 86316 92200
rect 86368 92188 86374 92200
rect 88168 92188 88196 92219
rect 89530 92216 89536 92228
rect 89588 92216 89594 92268
rect 88334 92188 88340 92200
rect 86368 92160 87644 92188
rect 88168 92160 88340 92188
rect 86368 92148 86374 92160
rect 32398 92080 32404 92132
rect 32456 92080 32462 92132
rect 51074 92080 51080 92132
rect 51132 92120 51138 92132
rect 52362 92120 52368 92132
rect 51132 92092 52368 92120
rect 51132 92080 51138 92092
rect 52362 92080 52368 92092
rect 52420 92120 52426 92132
rect 52733 92123 52791 92129
rect 52733 92120 52745 92123
rect 52420 92092 52745 92120
rect 52420 92080 52426 92092
rect 52733 92089 52745 92092
rect 52779 92089 52791 92123
rect 87506 92120 87512 92132
rect 52733 92083 52791 92089
rect 86788 92092 87512 92120
rect 86788 92064 86816 92092
rect 87506 92080 87512 92092
rect 87564 92080 87570 92132
rect 30466 92012 30472 92064
rect 30524 92052 30530 92064
rect 32217 92055 32275 92061
rect 32217 92052 32229 92055
rect 30524 92024 32229 92052
rect 30524 92012 30530 92024
rect 32217 92021 32229 92024
rect 32263 92052 32275 92055
rect 50246 92052 50252 92064
rect 32263 92024 50252 92052
rect 32263 92021 32275 92024
rect 32217 92015 32275 92021
rect 50246 92012 50252 92024
rect 50304 92012 50310 92064
rect 52549 92055 52607 92061
rect 52549 92021 52561 92055
rect 52595 92052 52607 92055
rect 52638 92052 52644 92064
rect 52595 92024 52644 92052
rect 52595 92021 52607 92024
rect 52549 92015 52607 92021
rect 52638 92012 52644 92024
rect 52696 92012 52702 92064
rect 85666 92012 85672 92064
rect 85724 92012 85730 92064
rect 85942 92012 85948 92064
rect 86000 92012 86006 92064
rect 86034 92012 86040 92064
rect 86092 92012 86098 92064
rect 86494 92012 86500 92064
rect 86552 92012 86558 92064
rect 86678 92012 86684 92064
rect 86736 92012 86742 92064
rect 86770 92012 86776 92064
rect 86828 92012 86834 92064
rect 87046 92012 87052 92064
rect 87104 92012 87110 92064
rect 87325 92055 87383 92061
rect 87325 92021 87337 92055
rect 87371 92052 87383 92055
rect 87414 92052 87420 92064
rect 87371 92024 87420 92052
rect 87371 92021 87383 92024
rect 87325 92015 87383 92021
rect 87414 92012 87420 92024
rect 87472 92012 87478 92064
rect 87616 92061 87644 92160
rect 88334 92148 88340 92160
rect 88392 92188 88398 92200
rect 88702 92188 88708 92200
rect 88392 92160 88708 92188
rect 88392 92148 88398 92160
rect 88702 92148 88708 92160
rect 88760 92148 88766 92200
rect 87690 92080 87696 92132
rect 87748 92120 87754 92132
rect 87969 92123 88027 92129
rect 87969 92120 87981 92123
rect 87748 92092 87981 92120
rect 87748 92080 87754 92092
rect 87969 92089 87981 92092
rect 88015 92089 88027 92123
rect 87969 92083 88027 92089
rect 88058 92080 88064 92132
rect 88116 92120 88122 92132
rect 88245 92123 88303 92129
rect 88245 92120 88257 92123
rect 88116 92092 88257 92120
rect 88116 92080 88122 92092
rect 88245 92089 88257 92092
rect 88291 92089 88303 92123
rect 88245 92083 88303 92089
rect 87601 92055 87659 92061
rect 87601 92021 87613 92055
rect 87647 92052 87659 92055
rect 88794 92052 88800 92064
rect 87647 92024 88800 92052
rect 87647 92021 87659 92024
rect 87601 92015 87659 92021
rect 88794 92012 88800 92024
rect 88852 92012 88858 92064
rect 1104 91962 88872 91984
rect 1104 91910 3066 91962
rect 3118 91910 3130 91962
rect 3182 91910 3194 91962
rect 3246 91910 3258 91962
rect 3310 91910 3322 91962
rect 3374 91910 36950 91962
rect 37002 91910 37014 91962
rect 37066 91910 37078 91962
rect 37130 91910 37142 91962
rect 37194 91910 37206 91962
rect 37258 91910 72950 91962
rect 73002 91910 73014 91962
rect 73066 91910 73078 91962
rect 73130 91910 73142 91962
rect 73194 91910 73206 91962
rect 73258 91910 88872 91962
rect 1104 91888 88872 91910
rect 50246 91808 50252 91860
rect 50304 91808 50310 91860
rect 86037 91851 86095 91857
rect 86037 91817 86049 91851
rect 86083 91848 86095 91851
rect 86310 91848 86316 91860
rect 86083 91820 86316 91848
rect 86083 91817 86095 91820
rect 86037 91811 86095 91817
rect 86310 91808 86316 91820
rect 86368 91808 86374 91860
rect 87230 91808 87236 91860
rect 87288 91848 87294 91860
rect 89162 91848 89168 91860
rect 87288 91820 89168 91848
rect 87288 91808 87294 91820
rect 89162 91808 89168 91820
rect 89220 91808 89226 91860
rect 86957 91783 87015 91789
rect 86957 91749 86969 91783
rect 87003 91780 87015 91783
rect 88334 91780 88340 91792
rect 87003 91752 88340 91780
rect 87003 91749 87015 91752
rect 86957 91743 87015 91749
rect 88334 91740 88340 91752
rect 88392 91740 88398 91792
rect 9646 91684 19334 91712
rect 5626 91536 5632 91588
rect 5684 91576 5690 91588
rect 9646 91576 9674 91684
rect 5684 91548 9674 91576
rect 5684 91536 5690 91548
rect 10318 91536 10324 91588
rect 10376 91576 10382 91588
rect 19306 91576 19334 91684
rect 47946 91672 47952 91724
rect 48004 91712 48010 91724
rect 86034 91712 86040 91724
rect 48004 91684 86040 91712
rect 48004 91672 48010 91684
rect 86034 91672 86040 91684
rect 86092 91672 86098 91724
rect 87598 91712 87604 91724
rect 86696 91684 87604 91712
rect 32217 91647 32275 91653
rect 32217 91644 32229 91647
rect 30392 91616 32229 91644
rect 30392 91585 30420 91616
rect 32217 91613 32229 91616
rect 32263 91644 32275 91647
rect 32398 91644 32404 91656
rect 32263 91616 32404 91644
rect 32263 91613 32275 91616
rect 32217 91607 32275 91613
rect 32398 91604 32404 91616
rect 32456 91604 32462 91656
rect 51169 91647 51227 91653
rect 51169 91644 51181 91647
rect 51092 91616 51181 91644
rect 30377 91579 30435 91585
rect 30377 91576 30389 91579
rect 10376 91548 13676 91576
rect 19306 91548 30389 91576
rect 10376 91536 10382 91548
rect 11606 91468 11612 91520
rect 11664 91468 11670 91520
rect 12526 91468 12532 91520
rect 12584 91468 12590 91520
rect 13538 91468 13544 91520
rect 13596 91468 13602 91520
rect 13648 91508 13676 91548
rect 30377 91545 30389 91548
rect 30423 91545 30435 91579
rect 30377 91539 30435 91545
rect 31941 91579 31999 91585
rect 31941 91545 31953 91579
rect 31987 91576 31999 91579
rect 32493 91579 32551 91585
rect 32493 91576 32505 91579
rect 31987 91548 32505 91576
rect 31987 91545 31999 91548
rect 31941 91539 31999 91545
rect 32493 91545 32505 91548
rect 32539 91576 32551 91579
rect 43438 91576 43444 91588
rect 32539 91548 43444 91576
rect 32539 91545 32551 91548
rect 32493 91539 32551 91545
rect 43438 91536 43444 91548
rect 43496 91536 43502 91588
rect 47762 91536 47768 91588
rect 47820 91576 47826 91588
rect 50801 91579 50859 91585
rect 50801 91576 50813 91579
rect 47820 91548 50813 91576
rect 47820 91536 47826 91548
rect 50801 91545 50813 91548
rect 50847 91545 50859 91579
rect 50801 91539 50859 91545
rect 51092 91520 51120 91616
rect 51169 91613 51181 91616
rect 51215 91613 51227 91647
rect 51169 91607 51227 91613
rect 52730 91604 52736 91656
rect 52788 91644 52794 91656
rect 53742 91644 53748 91656
rect 52788 91616 53748 91644
rect 52788 91604 52794 91616
rect 53742 91604 53748 91616
rect 53800 91644 53806 91656
rect 54389 91647 54447 91653
rect 54389 91644 54401 91647
rect 53800 91616 54401 91644
rect 53800 91604 53806 91616
rect 54389 91613 54401 91616
rect 54435 91613 54447 91647
rect 54389 91607 54447 91613
rect 84470 91604 84476 91656
rect 84528 91644 84534 91656
rect 85669 91647 85727 91653
rect 84528 91616 85344 91644
rect 84528 91604 84534 91616
rect 52365 91579 52423 91585
rect 52365 91545 52377 91579
rect 52411 91576 52423 91579
rect 52454 91576 52460 91588
rect 52411 91548 52460 91576
rect 52411 91545 52423 91548
rect 52365 91539 52423 91545
rect 52454 91536 52460 91548
rect 52512 91536 52518 91588
rect 53834 91536 53840 91588
rect 53892 91576 53898 91588
rect 54573 91579 54631 91585
rect 54573 91576 54585 91579
rect 53892 91548 54585 91576
rect 53892 91536 53898 91548
rect 54573 91545 54585 91548
rect 54619 91545 54631 91579
rect 54573 91539 54631 91545
rect 85206 91536 85212 91588
rect 85264 91536 85270 91588
rect 85316 91576 85344 91616
rect 85669 91613 85681 91647
rect 85715 91644 85727 91647
rect 85850 91644 85856 91656
rect 85715 91616 85856 91644
rect 85715 91613 85727 91616
rect 85669 91607 85727 91613
rect 85850 91604 85856 91616
rect 85908 91604 85914 91656
rect 86696 91653 86724 91684
rect 87598 91672 87604 91684
rect 87656 91712 87662 91724
rect 89070 91712 89076 91724
rect 87656 91684 89076 91712
rect 87656 91672 87662 91684
rect 89070 91672 89076 91684
rect 89128 91672 89134 91724
rect 86681 91647 86739 91653
rect 86681 91613 86693 91647
rect 86727 91613 86739 91647
rect 86681 91607 86739 91613
rect 86773 91647 86831 91653
rect 86773 91613 86785 91647
rect 86819 91613 86831 91647
rect 86773 91607 86831 91613
rect 88061 91647 88119 91653
rect 88061 91613 88073 91647
rect 88107 91644 88119 91647
rect 88518 91644 88524 91656
rect 88107 91616 88524 91644
rect 88107 91613 88119 91616
rect 88061 91607 88119 91613
rect 86788 91576 86816 91607
rect 88518 91604 88524 91616
rect 88576 91644 88582 91656
rect 88978 91644 88984 91656
rect 88576 91616 88984 91644
rect 88576 91604 88582 91616
rect 88978 91604 88984 91616
rect 89036 91604 89042 91656
rect 85316 91548 86816 91576
rect 87138 91536 87144 91588
rect 87196 91536 87202 91588
rect 87322 91536 87328 91588
rect 87380 91536 87386 91588
rect 87506 91536 87512 91588
rect 87564 91536 87570 91588
rect 87693 91579 87751 91585
rect 87693 91545 87705 91579
rect 87739 91576 87751 91579
rect 87874 91576 87880 91588
rect 87739 91548 87880 91576
rect 87739 91545 87751 91548
rect 87693 91539 87751 91545
rect 87874 91536 87880 91548
rect 87932 91576 87938 91588
rect 87932 91548 88196 91576
rect 87932 91536 87938 91548
rect 30466 91508 30472 91520
rect 13648 91480 30472 91508
rect 30466 91468 30472 91480
rect 30524 91468 30530 91520
rect 47670 91468 47676 91520
rect 47728 91508 47734 91520
rect 49697 91511 49755 91517
rect 49697 91508 49709 91511
rect 47728 91480 49709 91508
rect 47728 91468 47734 91480
rect 49697 91477 49709 91480
rect 49743 91477 49755 91511
rect 49697 91471 49755 91477
rect 51074 91468 51080 91520
rect 51132 91468 51138 91520
rect 53742 91468 53748 91520
rect 53800 91508 53806 91520
rect 54205 91511 54263 91517
rect 54205 91508 54217 91511
rect 53800 91480 54217 91508
rect 53800 91468 53806 91480
rect 54205 91477 54217 91480
rect 54251 91477 54263 91511
rect 54205 91471 54263 91477
rect 85022 91468 85028 91520
rect 85080 91468 85086 91520
rect 85390 91468 85396 91520
rect 85448 91468 85454 91520
rect 85758 91468 85764 91520
rect 85816 91468 85822 91520
rect 86310 91468 86316 91520
rect 86368 91468 86374 91520
rect 86497 91511 86555 91517
rect 86497 91477 86509 91511
rect 86543 91508 86555 91511
rect 86678 91508 86684 91520
rect 86543 91480 86684 91508
rect 86543 91477 86555 91480
rect 86497 91471 86555 91477
rect 86678 91468 86684 91480
rect 86736 91468 86742 91520
rect 87966 91468 87972 91520
rect 88024 91468 88030 91520
rect 88168 91508 88196 91548
rect 88242 91536 88248 91588
rect 88300 91536 88306 91588
rect 88429 91579 88487 91585
rect 88429 91545 88441 91579
rect 88475 91576 88487 91579
rect 88610 91576 88616 91588
rect 88475 91548 88616 91576
rect 88475 91545 88487 91548
rect 88429 91539 88487 91545
rect 88610 91536 88616 91548
rect 88668 91576 88674 91588
rect 89438 91576 89444 91588
rect 88668 91548 89444 91576
rect 88668 91536 88674 91548
rect 89438 91536 89444 91548
rect 89496 91536 89502 91588
rect 88518 91508 88524 91520
rect 88168 91480 88524 91508
rect 88518 91468 88524 91480
rect 88576 91468 88582 91520
rect 1104 91418 88872 91440
rect 1104 91366 3802 91418
rect 3854 91366 3866 91418
rect 3918 91366 3930 91418
rect 3982 91366 3994 91418
rect 4046 91366 4058 91418
rect 4110 91366 37610 91418
rect 37662 91366 37674 91418
rect 37726 91366 37738 91418
rect 37790 91366 37802 91418
rect 37854 91366 37866 91418
rect 37918 91366 73610 91418
rect 73662 91366 73674 91418
rect 73726 91366 73738 91418
rect 73790 91366 73802 91418
rect 73854 91366 73866 91418
rect 73918 91366 88872 91418
rect 1104 91344 88872 91366
rect 12526 91264 12532 91316
rect 12584 91304 12590 91316
rect 52730 91304 52736 91316
rect 12584 91276 52736 91304
rect 12584 91264 12590 91276
rect 52730 91264 52736 91276
rect 52788 91264 52794 91316
rect 11606 91196 11612 91248
rect 11664 91236 11670 91248
rect 51074 91236 51080 91248
rect 11664 91208 51080 91236
rect 11664 91196 11670 91208
rect 51074 91196 51080 91208
rect 51132 91196 51138 91248
rect 47854 91128 47860 91180
rect 47912 91168 47918 91180
rect 85390 91168 85396 91180
rect 47912 91140 85396 91168
rect 47912 91128 47918 91140
rect 85390 91128 85396 91140
rect 85448 91128 85454 91180
rect 48130 91060 48136 91112
rect 48188 91100 48194 91112
rect 85758 91100 85764 91112
rect 48188 91072 85764 91100
rect 48188 91060 48194 91072
rect 85758 91060 85764 91072
rect 85816 91060 85822 91112
rect 48222 90992 48228 91044
rect 48280 91032 48286 91044
rect 52454 91032 52460 91044
rect 48280 91004 52460 91032
rect 48280 90992 48286 91004
rect 52454 90992 52460 91004
rect 52512 90992 52518 91044
rect 48038 90924 48044 90976
rect 48096 90964 48102 90976
rect 53834 90964 53840 90976
rect 48096 90936 53840 90964
rect 48096 90924 48102 90936
rect 53834 90924 53840 90936
rect 53892 90924 53898 90976
rect 1104 90874 5980 90896
rect 1104 90822 3066 90874
rect 3118 90822 3130 90874
rect 3182 90822 3194 90874
rect 3246 90822 3258 90874
rect 3310 90822 3322 90874
rect 3374 90822 5980 90874
rect 1104 90800 5980 90822
rect 1104 90330 5980 90352
rect 1104 90278 3802 90330
rect 3854 90278 3866 90330
rect 3918 90278 3930 90330
rect 3982 90278 3994 90330
rect 4046 90278 4058 90330
rect 4110 90278 5980 90330
rect 1104 90256 5980 90278
rect 1104 89786 5980 89808
rect 1104 89734 3066 89786
rect 3118 89734 3130 89786
rect 3182 89734 3194 89786
rect 3246 89734 3258 89786
rect 3310 89734 3322 89786
rect 3374 89734 5980 89786
rect 1104 89712 5980 89734
rect 47302 89632 47308 89684
rect 47360 89672 47366 89684
rect 85022 89672 85028 89684
rect 47360 89644 85028 89672
rect 47360 89632 47366 89644
rect 85022 89632 85028 89644
rect 85080 89632 85086 89684
rect 5166 89292 5172 89344
rect 5224 89332 5230 89344
rect 85666 89332 85672 89344
rect 5224 89304 85672 89332
rect 5224 89292 5230 89304
rect 85666 89292 85672 89304
rect 85724 89292 85730 89344
rect 1104 89242 5980 89264
rect 1104 89190 3802 89242
rect 3854 89190 3866 89242
rect 3918 89190 3930 89242
rect 3982 89190 3994 89242
rect 4046 89190 4058 89242
rect 4110 89190 5980 89242
rect 1104 89168 5980 89190
rect 5350 89088 5356 89140
rect 5408 89128 5414 89140
rect 86494 89128 86500 89140
rect 5408 89100 86500 89128
rect 5408 89088 5414 89100
rect 86494 89088 86500 89100
rect 86552 89088 86558 89140
rect 5442 89020 5448 89072
rect 5500 89060 5506 89072
rect 86034 89060 86040 89072
rect 5500 89032 86040 89060
rect 5500 89020 5506 89032
rect 86034 89020 86040 89032
rect 86092 89020 86098 89072
rect 5074 88952 5080 89004
rect 5132 88992 5138 89004
rect 86310 88992 86316 89004
rect 5132 88964 86316 88992
rect 5132 88952 5138 88964
rect 86310 88952 86316 88964
rect 86368 88952 86374 89004
rect 1104 88698 5980 88720
rect 1104 88646 3066 88698
rect 3118 88646 3130 88698
rect 3182 88646 3194 88698
rect 3246 88646 3258 88698
rect 3310 88646 3322 88698
rect 3374 88646 5980 88698
rect 1104 88624 5980 88646
rect 6730 88476 6736 88528
rect 6788 88516 6794 88528
rect 53190 88516 53196 88528
rect 6788 88488 53196 88516
rect 6788 88476 6794 88488
rect 53190 88476 53196 88488
rect 53248 88476 53254 88528
rect 86310 88476 86316 88528
rect 86368 88516 86374 88528
rect 88610 88516 88616 88528
rect 86368 88488 88616 88516
rect 86368 88476 86374 88488
rect 88610 88476 88616 88488
rect 88668 88476 88674 88528
rect 13722 88408 13728 88460
rect 13780 88448 13786 88460
rect 47578 88448 47584 88460
rect 13780 88420 47584 88448
rect 13780 88408 13786 88420
rect 47578 88408 47584 88420
rect 47636 88408 47642 88460
rect 85666 88408 85672 88460
rect 85724 88448 85730 88460
rect 86862 88448 86868 88460
rect 85724 88420 86868 88448
rect 85724 88408 85730 88420
rect 86862 88408 86868 88420
rect 86920 88408 86926 88460
rect 5258 88340 5264 88392
rect 5316 88380 5322 88392
rect 47302 88380 47308 88392
rect 5316 88352 47308 88380
rect 5316 88340 5322 88352
rect 47302 88340 47308 88352
rect 47360 88340 47366 88392
rect 1104 88154 5980 88176
rect 1104 88102 3802 88154
rect 3854 88102 3866 88154
rect 3918 88102 3930 88154
rect 3982 88102 3994 88154
rect 4046 88102 4058 88154
rect 4110 88102 5980 88154
rect 1104 88080 5980 88102
rect 1104 87610 5980 87632
rect 1104 87558 3066 87610
rect 3118 87558 3130 87610
rect 3182 87558 3194 87610
rect 3246 87558 3258 87610
rect 3310 87558 3322 87610
rect 3374 87558 5980 87610
rect 1104 87536 5980 87558
rect 1104 87066 5980 87088
rect 1104 87014 3802 87066
rect 3854 87014 3866 87066
rect 3918 87014 3930 87066
rect 3982 87014 3994 87066
rect 4046 87014 4058 87066
rect 4110 87014 5980 87066
rect 1104 86992 5980 87014
rect 1673 86819 1731 86825
rect 1673 86785 1685 86819
rect 1719 86816 1731 86819
rect 8294 86816 8300 86828
rect 1719 86788 8300 86816
rect 1719 86785 1731 86788
rect 1673 86779 1731 86785
rect 8294 86776 8300 86788
rect 8352 86776 8358 86828
rect 842 86572 848 86624
rect 900 86612 906 86624
rect 1489 86615 1547 86621
rect 1489 86612 1501 86615
rect 900 86584 1501 86612
rect 900 86572 906 86584
rect 1489 86581 1501 86584
rect 1535 86581 1547 86615
rect 1489 86575 1547 86581
rect 1104 86522 5980 86544
rect 1104 86470 3066 86522
rect 3118 86470 3130 86522
rect 3182 86470 3194 86522
rect 3246 86470 3258 86522
rect 3310 86470 3322 86522
rect 3374 86470 5980 86522
rect 1104 86448 5980 86470
rect 1104 85978 5980 86000
rect 1104 85926 3802 85978
rect 3854 85926 3866 85978
rect 3918 85926 3930 85978
rect 3982 85926 3994 85978
rect 4046 85926 4058 85978
rect 4110 85926 5980 85978
rect 1104 85904 5980 85926
rect 1104 85434 5980 85456
rect 1104 85382 3066 85434
rect 3118 85382 3130 85434
rect 3182 85382 3194 85434
rect 3246 85382 3258 85434
rect 3310 85382 3322 85434
rect 3374 85382 5980 85434
rect 1104 85360 5980 85382
rect 842 85212 848 85264
rect 900 85252 906 85264
rect 1489 85255 1547 85261
rect 1489 85252 1501 85255
rect 900 85224 1501 85252
rect 900 85212 906 85224
rect 1489 85221 1501 85224
rect 1535 85221 1547 85255
rect 1489 85215 1547 85221
rect 1673 85119 1731 85125
rect 1673 85085 1685 85119
rect 1719 85116 1731 85119
rect 8294 85116 8300 85128
rect 1719 85088 8300 85116
rect 1719 85085 1731 85088
rect 1673 85079 1731 85085
rect 8294 85076 8300 85088
rect 8352 85076 8358 85128
rect 1104 84890 5980 84912
rect 1104 84838 3802 84890
rect 3854 84838 3866 84890
rect 3918 84838 3930 84890
rect 3982 84838 3994 84890
rect 4046 84838 4058 84890
rect 4110 84838 5980 84890
rect 1104 84816 5980 84838
rect 1104 84346 5980 84368
rect 1104 84294 3066 84346
rect 3118 84294 3130 84346
rect 3182 84294 3194 84346
rect 3246 84294 3258 84346
rect 3310 84294 3322 84346
rect 3374 84294 5980 84346
rect 1104 84272 5980 84294
rect 1673 84031 1731 84037
rect 1673 83997 1685 84031
rect 1719 84028 1731 84031
rect 8294 84028 8300 84040
rect 1719 84000 8300 84028
rect 1719 83997 1731 84000
rect 1673 83991 1731 83997
rect 8294 83988 8300 84000
rect 8352 83988 8358 84040
rect 842 83852 848 83904
rect 900 83892 906 83904
rect 1489 83895 1547 83901
rect 1489 83892 1501 83895
rect 900 83864 1501 83892
rect 900 83852 906 83864
rect 1489 83861 1501 83864
rect 1535 83861 1547 83895
rect 1489 83855 1547 83861
rect 1104 83802 5980 83824
rect 1104 83750 3802 83802
rect 3854 83750 3866 83802
rect 3918 83750 3930 83802
rect 3982 83750 3994 83802
rect 4046 83750 4058 83802
rect 4110 83750 5980 83802
rect 1104 83728 5980 83750
rect 1104 83258 5980 83280
rect 1104 83206 3066 83258
rect 3118 83206 3130 83258
rect 3182 83206 3194 83258
rect 3246 83206 3258 83258
rect 3310 83206 3322 83258
rect 3374 83206 5980 83258
rect 1104 83184 5980 83206
rect 1104 82714 5980 82736
rect 1104 82662 3802 82714
rect 3854 82662 3866 82714
rect 3918 82662 3930 82714
rect 3982 82662 3994 82714
rect 4046 82662 4058 82714
rect 4110 82662 5980 82714
rect 1104 82640 5980 82662
rect 1673 82467 1731 82473
rect 1673 82433 1685 82467
rect 1719 82464 1731 82467
rect 8294 82464 8300 82476
rect 1719 82436 8300 82464
rect 1719 82433 1731 82436
rect 1673 82427 1731 82433
rect 8294 82424 8300 82436
rect 8352 82424 8358 82476
rect 842 82220 848 82272
rect 900 82260 906 82272
rect 1489 82263 1547 82269
rect 1489 82260 1501 82263
rect 900 82232 1501 82260
rect 900 82220 906 82232
rect 1489 82229 1501 82232
rect 1535 82229 1547 82263
rect 1489 82223 1547 82229
rect 1104 82170 5980 82192
rect 1104 82118 3066 82170
rect 3118 82118 3130 82170
rect 3182 82118 3194 82170
rect 3246 82118 3258 82170
rect 3310 82118 3322 82170
rect 3374 82118 5980 82170
rect 1104 82096 5980 82118
rect 88426 81744 88432 81796
rect 88484 81784 88490 81796
rect 88794 81784 88800 81796
rect 88484 81756 88800 81784
rect 88484 81744 88490 81756
rect 88794 81744 88800 81756
rect 88852 81744 88858 81796
rect 1104 81626 5980 81648
rect 1104 81574 3802 81626
rect 3854 81574 3866 81626
rect 3918 81574 3930 81626
rect 3982 81574 3994 81626
rect 4046 81574 4058 81626
rect 4110 81574 5980 81626
rect 1104 81552 5980 81574
rect 1673 81379 1731 81385
rect 1673 81345 1685 81379
rect 1719 81376 1731 81379
rect 8294 81376 8300 81388
rect 1719 81348 8300 81376
rect 1719 81345 1731 81348
rect 1673 81339 1731 81345
rect 8294 81336 8300 81348
rect 8352 81336 8358 81388
rect 842 81132 848 81184
rect 900 81172 906 81184
rect 1489 81175 1547 81181
rect 1489 81172 1501 81175
rect 900 81144 1501 81172
rect 900 81132 906 81144
rect 1489 81141 1501 81144
rect 1535 81141 1547 81175
rect 1489 81135 1547 81141
rect 1104 81082 5980 81104
rect 1104 81030 3066 81082
rect 3118 81030 3130 81082
rect 3182 81030 3194 81082
rect 3246 81030 3258 81082
rect 3310 81030 3322 81082
rect 3374 81030 5980 81082
rect 1104 81008 5980 81030
rect 1104 80538 5980 80560
rect 1104 80486 3802 80538
rect 3854 80486 3866 80538
rect 3918 80486 3930 80538
rect 3982 80486 3994 80538
rect 4046 80486 4058 80538
rect 4110 80486 5980 80538
rect 1104 80464 5980 80486
rect 1104 79994 5980 80016
rect 1104 79942 3066 79994
rect 3118 79942 3130 79994
rect 3182 79942 3194 79994
rect 3246 79942 3258 79994
rect 3310 79942 3322 79994
rect 3374 79942 5980 79994
rect 1104 79920 5980 79942
rect 1673 79679 1731 79685
rect 1673 79645 1685 79679
rect 1719 79676 1731 79679
rect 8294 79676 8300 79688
rect 1719 79648 8300 79676
rect 1719 79645 1731 79648
rect 1673 79639 1731 79645
rect 8294 79636 8300 79648
rect 8352 79636 8358 79688
rect 842 79500 848 79552
rect 900 79540 906 79552
rect 1489 79543 1547 79549
rect 1489 79540 1501 79543
rect 900 79512 1501 79540
rect 900 79500 906 79512
rect 1489 79509 1501 79512
rect 1535 79509 1547 79543
rect 1489 79503 1547 79509
rect 1104 79450 5980 79472
rect 1104 79398 3802 79450
rect 3854 79398 3866 79450
rect 3918 79398 3930 79450
rect 3982 79398 3994 79450
rect 4046 79398 4058 79450
rect 4110 79398 5980 79450
rect 1104 79376 5980 79398
rect 1104 78906 5980 78928
rect 1104 78854 3066 78906
rect 3118 78854 3130 78906
rect 3182 78854 3194 78906
rect 3246 78854 3258 78906
rect 3310 78854 3322 78906
rect 3374 78854 5980 78906
rect 1104 78832 5980 78854
rect 1673 78591 1731 78597
rect 1673 78557 1685 78591
rect 1719 78588 1731 78591
rect 8294 78588 8300 78600
rect 1719 78560 8300 78588
rect 1719 78557 1731 78560
rect 1673 78551 1731 78557
rect 8294 78548 8300 78560
rect 8352 78548 8358 78600
rect 842 78412 848 78464
rect 900 78452 906 78464
rect 1489 78455 1547 78461
rect 1489 78452 1501 78455
rect 900 78424 1501 78452
rect 900 78412 906 78424
rect 1489 78421 1501 78424
rect 1535 78421 1547 78455
rect 1489 78415 1547 78421
rect 1104 78362 5980 78384
rect 1104 78310 3802 78362
rect 3854 78310 3866 78362
rect 3918 78310 3930 78362
rect 3982 78310 3994 78362
rect 4046 78310 4058 78362
rect 4110 78310 5980 78362
rect 1104 78288 5980 78310
rect 1104 77818 5980 77840
rect 1104 77766 3066 77818
rect 3118 77766 3130 77818
rect 3182 77766 3194 77818
rect 3246 77766 3258 77818
rect 3310 77766 3322 77818
rect 3374 77766 5980 77818
rect 1104 77744 5980 77766
rect 1104 77274 5980 77296
rect 1104 77222 3802 77274
rect 3854 77222 3866 77274
rect 3918 77222 3930 77274
rect 3982 77222 3994 77274
rect 4046 77222 4058 77274
rect 4110 77222 5980 77274
rect 1104 77200 5980 77222
rect 89162 77052 89168 77104
rect 89220 77092 89226 77104
rect 89346 77092 89352 77104
rect 89220 77064 89352 77092
rect 89220 77052 89226 77064
rect 89346 77052 89352 77064
rect 89404 77052 89410 77104
rect 1673 77027 1731 77033
rect 1673 76993 1685 77027
rect 1719 77024 1731 77027
rect 8294 77024 8300 77036
rect 1719 76996 8300 77024
rect 1719 76993 1731 76996
rect 1673 76987 1731 76993
rect 8294 76984 8300 76996
rect 8352 76984 8358 77036
rect 842 76780 848 76832
rect 900 76820 906 76832
rect 1489 76823 1547 76829
rect 1489 76820 1501 76823
rect 900 76792 1501 76820
rect 900 76780 906 76792
rect 1489 76789 1501 76792
rect 1535 76789 1547 76823
rect 1489 76783 1547 76789
rect 1104 76730 5980 76752
rect 1104 76678 3066 76730
rect 3118 76678 3130 76730
rect 3182 76678 3194 76730
rect 3246 76678 3258 76730
rect 3310 76678 3322 76730
rect 3374 76678 5980 76730
rect 1104 76656 5980 76678
rect 1104 76186 5980 76208
rect 1104 76134 3802 76186
rect 3854 76134 3866 76186
rect 3918 76134 3930 76186
rect 3982 76134 3994 76186
rect 4046 76134 4058 76186
rect 4110 76134 5980 76186
rect 1104 76112 5980 76134
rect 842 76032 848 76084
rect 900 76072 906 76084
rect 1489 76075 1547 76081
rect 1489 76072 1501 76075
rect 900 76044 1501 76072
rect 900 76032 906 76044
rect 1489 76041 1501 76044
rect 1535 76041 1547 76075
rect 1489 76035 1547 76041
rect 1673 75939 1731 75945
rect 1673 75905 1685 75939
rect 1719 75936 1731 75939
rect 5534 75936 5540 75948
rect 1719 75908 5540 75936
rect 1719 75905 1731 75908
rect 1673 75899 1731 75905
rect 5534 75896 5540 75908
rect 5592 75896 5598 75948
rect 1104 75642 5980 75664
rect 1104 75590 3066 75642
rect 3118 75590 3130 75642
rect 3182 75590 3194 75642
rect 3246 75590 3258 75642
rect 3310 75590 3322 75642
rect 3374 75590 5980 75642
rect 1104 75568 5980 75590
rect 1104 75098 5980 75120
rect 1104 75046 3802 75098
rect 3854 75046 3866 75098
rect 3918 75046 3930 75098
rect 3982 75046 3994 75098
rect 4046 75046 4058 75098
rect 4110 75046 5980 75098
rect 1104 75024 5980 75046
rect 1104 74554 5980 74576
rect 1104 74502 3066 74554
rect 3118 74502 3130 74554
rect 3182 74502 3194 74554
rect 3246 74502 3258 74554
rect 3310 74502 3322 74554
rect 3374 74502 5980 74554
rect 1104 74480 5980 74502
rect 1673 74239 1731 74245
rect 1673 74205 1685 74239
rect 1719 74236 1731 74239
rect 8294 74236 8300 74248
rect 1719 74208 8300 74236
rect 1719 74205 1731 74208
rect 1673 74199 1731 74205
rect 8294 74196 8300 74208
rect 8352 74196 8358 74248
rect 842 74060 848 74112
rect 900 74100 906 74112
rect 1489 74103 1547 74109
rect 1489 74100 1501 74103
rect 900 74072 1501 74100
rect 900 74060 906 74072
rect 1489 74069 1501 74072
rect 1535 74069 1547 74103
rect 1489 74063 1547 74069
rect 1104 74010 5980 74032
rect 1104 73958 3802 74010
rect 3854 73958 3866 74010
rect 3918 73958 3930 74010
rect 3982 73958 3994 74010
rect 4046 73958 4058 74010
rect 4110 73958 5980 74010
rect 1104 73936 5980 73958
rect 1104 73466 5980 73488
rect 1104 73414 3066 73466
rect 3118 73414 3130 73466
rect 3182 73414 3194 73466
rect 3246 73414 3258 73466
rect 3310 73414 3322 73466
rect 3374 73414 5980 73466
rect 1104 73392 5980 73414
rect 1673 73151 1731 73157
rect 1673 73117 1685 73151
rect 1719 73148 1731 73151
rect 8294 73148 8300 73160
rect 1719 73120 8300 73148
rect 1719 73117 1731 73120
rect 1673 73111 1731 73117
rect 8294 73108 8300 73120
rect 8352 73108 8358 73160
rect 842 72972 848 73024
rect 900 73012 906 73024
rect 1489 73015 1547 73021
rect 1489 73012 1501 73015
rect 900 72984 1501 73012
rect 900 72972 906 72984
rect 1489 72981 1501 72984
rect 1535 72981 1547 73015
rect 1489 72975 1547 72981
rect 1104 72922 5980 72944
rect 1104 72870 3802 72922
rect 3854 72870 3866 72922
rect 3918 72870 3930 72922
rect 3982 72870 3994 72922
rect 4046 72870 4058 72922
rect 4110 72870 5980 72922
rect 1104 72848 5980 72870
rect 1104 72378 5980 72400
rect 1104 72326 3066 72378
rect 3118 72326 3130 72378
rect 3182 72326 3194 72378
rect 3246 72326 3258 72378
rect 3310 72326 3322 72378
rect 3374 72326 5980 72378
rect 1104 72304 5980 72326
rect 1104 71834 5980 71856
rect 1104 71782 3802 71834
rect 3854 71782 3866 71834
rect 3918 71782 3930 71834
rect 3982 71782 3994 71834
rect 4046 71782 4058 71834
rect 4110 71782 5980 71834
rect 1104 71760 5980 71782
rect 8294 71652 8300 71664
rect 1688 71624 8300 71652
rect 1688 71593 1716 71624
rect 8294 71612 8300 71624
rect 8352 71612 8358 71664
rect 1673 71587 1731 71593
rect 1673 71553 1685 71587
rect 1719 71553 1731 71587
rect 1673 71547 1731 71553
rect 5169 71587 5227 71593
rect 5169 71553 5181 71587
rect 5215 71584 5227 71587
rect 5629 71587 5687 71593
rect 5629 71584 5641 71587
rect 5215 71556 5641 71584
rect 5215 71553 5227 71556
rect 5169 71547 5227 71553
rect 5629 71553 5641 71556
rect 5675 71584 5687 71587
rect 5902 71584 5908 71596
rect 5675 71556 5908 71584
rect 5675 71553 5687 71556
rect 5629 71547 5687 71553
rect 5902 71544 5908 71556
rect 5960 71544 5966 71596
rect 4614 71408 4620 71460
rect 4672 71448 4678 71460
rect 5261 71451 5319 71457
rect 5261 71448 5273 71451
rect 4672 71420 5273 71448
rect 4672 71408 4678 71420
rect 5261 71417 5273 71420
rect 5307 71448 5319 71451
rect 5445 71451 5503 71457
rect 5445 71448 5457 71451
rect 5307 71420 5457 71448
rect 5307 71417 5319 71420
rect 5261 71411 5319 71417
rect 5445 71417 5457 71420
rect 5491 71417 5503 71451
rect 5445 71411 5503 71417
rect 842 71340 848 71392
rect 900 71380 906 71392
rect 1489 71383 1547 71389
rect 1489 71380 1501 71383
rect 900 71352 1501 71380
rect 900 71340 906 71352
rect 1489 71349 1501 71352
rect 1535 71349 1547 71383
rect 1489 71343 1547 71349
rect 1104 71290 5980 71312
rect 1104 71238 3066 71290
rect 3118 71238 3130 71290
rect 3182 71238 3194 71290
rect 3246 71238 3258 71290
rect 3310 71238 3322 71290
rect 3374 71238 5980 71290
rect 1104 71216 5980 71238
rect 1104 70746 5980 70768
rect 1104 70694 3802 70746
rect 3854 70694 3866 70746
rect 3918 70694 3930 70746
rect 3982 70694 3994 70746
rect 4046 70694 4058 70746
rect 4110 70694 5980 70746
rect 1104 70672 5980 70694
rect 842 70592 848 70644
rect 900 70632 906 70644
rect 1489 70635 1547 70641
rect 1489 70632 1501 70635
rect 900 70604 1501 70632
rect 900 70592 906 70604
rect 1489 70601 1501 70604
rect 1535 70601 1547 70635
rect 1489 70595 1547 70601
rect 5074 70592 5080 70644
rect 5132 70632 5138 70644
rect 5261 70635 5319 70641
rect 5261 70632 5273 70635
rect 5132 70604 5273 70632
rect 5132 70592 5138 70604
rect 5261 70601 5273 70604
rect 5307 70632 5319 70635
rect 5445 70635 5503 70641
rect 5445 70632 5457 70635
rect 5307 70604 5457 70632
rect 5307 70601 5319 70604
rect 5261 70595 5319 70601
rect 5445 70601 5457 70604
rect 5491 70601 5503 70635
rect 5445 70595 5503 70601
rect 1673 70499 1731 70505
rect 1673 70465 1685 70499
rect 1719 70496 1731 70499
rect 5534 70496 5540 70508
rect 1719 70468 5540 70496
rect 1719 70465 1731 70468
rect 1673 70459 1731 70465
rect 5534 70456 5540 70468
rect 5592 70456 5598 70508
rect 5629 70499 5687 70505
rect 5629 70465 5641 70499
rect 5675 70496 5687 70499
rect 5810 70496 5816 70508
rect 5675 70468 5816 70496
rect 5675 70465 5687 70468
rect 5629 70459 5687 70465
rect 5169 70431 5227 70437
rect 5169 70397 5181 70431
rect 5215 70428 5227 70431
rect 5644 70428 5672 70459
rect 5810 70456 5816 70468
rect 5868 70456 5874 70508
rect 5215 70400 5672 70428
rect 5215 70397 5227 70400
rect 5169 70391 5227 70397
rect 1104 70202 5980 70224
rect 1104 70150 3066 70202
rect 3118 70150 3130 70202
rect 3182 70150 3194 70202
rect 3246 70150 3258 70202
rect 3310 70150 3322 70202
rect 3374 70150 5980 70202
rect 1104 70128 5980 70150
rect 1104 69658 5980 69680
rect 1104 69606 3802 69658
rect 3854 69606 3866 69658
rect 3918 69606 3930 69658
rect 3982 69606 3994 69658
rect 4046 69606 4058 69658
rect 4110 69606 5980 69658
rect 1104 69584 5980 69606
rect 1104 69114 5980 69136
rect 1104 69062 3066 69114
rect 3118 69062 3130 69114
rect 3182 69062 3194 69114
rect 3246 69062 3258 69114
rect 3310 69062 3322 69114
rect 3374 69062 5980 69114
rect 1104 69040 5980 69062
rect 1581 68935 1639 68941
rect 1581 68901 1593 68935
rect 1627 68932 1639 68935
rect 8294 68932 8300 68944
rect 1627 68904 8300 68932
rect 1627 68901 1639 68904
rect 1581 68895 1639 68901
rect 8294 68892 8300 68904
rect 8352 68892 8358 68944
rect 1210 68756 1216 68808
rect 1268 68796 1274 68808
rect 1397 68799 1455 68805
rect 1397 68796 1409 68799
rect 1268 68768 1409 68796
rect 1268 68756 1274 68768
rect 1397 68765 1409 68768
rect 1443 68796 1455 68799
rect 1673 68799 1731 68805
rect 1673 68796 1685 68799
rect 1443 68768 1685 68796
rect 1443 68765 1455 68768
rect 1397 68759 1455 68765
rect 1673 68765 1685 68768
rect 1719 68765 1731 68799
rect 1673 68759 1731 68765
rect 5353 68799 5411 68805
rect 5353 68765 5365 68799
rect 5399 68796 5411 68799
rect 5399 68768 5433 68796
rect 5399 68765 5411 68768
rect 5353 68759 5411 68765
rect 5261 68731 5319 68737
rect 5261 68697 5273 68731
rect 5307 68728 5319 68731
rect 5368 68728 5396 68759
rect 6178 68728 6184 68740
rect 5307 68700 6184 68728
rect 5307 68697 5319 68700
rect 5261 68691 5319 68697
rect 6178 68688 6184 68700
rect 6236 68688 6242 68740
rect 5537 68663 5595 68669
rect 5537 68629 5549 68663
rect 5583 68660 5595 68663
rect 6086 68660 6092 68672
rect 5583 68632 6092 68660
rect 5583 68629 5595 68632
rect 5537 68623 5595 68629
rect 6086 68620 6092 68632
rect 6144 68620 6150 68672
rect 1104 68570 5980 68592
rect 1104 68518 3802 68570
rect 3854 68518 3866 68570
rect 3918 68518 3930 68570
rect 3982 68518 3994 68570
rect 4046 68518 4058 68570
rect 4110 68518 5980 68570
rect 1104 68496 5980 68518
rect 1104 68026 5980 68048
rect 1104 67974 3066 68026
rect 3118 67974 3130 68026
rect 3182 67974 3194 68026
rect 3246 67974 3258 68026
rect 3310 67974 3322 68026
rect 3374 67974 5980 68026
rect 1104 67952 5980 67974
rect 1581 67915 1639 67921
rect 1581 67881 1593 67915
rect 1627 67912 1639 67915
rect 5718 67912 5724 67924
rect 1627 67884 5724 67912
rect 1627 67881 1639 67884
rect 1581 67875 1639 67881
rect 5718 67872 5724 67884
rect 5776 67872 5782 67924
rect 5261 67847 5319 67853
rect 5261 67813 5273 67847
rect 5307 67844 5319 67847
rect 5442 67844 5448 67856
rect 5307 67816 5448 67844
rect 5307 67813 5319 67816
rect 5261 67807 5319 67813
rect 1302 67668 1308 67720
rect 1360 67708 1366 67720
rect 5368 67717 5396 67816
rect 5442 67804 5448 67816
rect 5500 67804 5506 67856
rect 5534 67804 5540 67856
rect 5592 67804 5598 67856
rect 1397 67711 1455 67717
rect 1397 67708 1409 67711
rect 1360 67680 1409 67708
rect 1360 67668 1366 67680
rect 1397 67677 1409 67680
rect 1443 67708 1455 67711
rect 1673 67711 1731 67717
rect 1673 67708 1685 67711
rect 1443 67680 1685 67708
rect 1443 67677 1455 67680
rect 1397 67671 1455 67677
rect 1673 67677 1685 67680
rect 1719 67677 1731 67711
rect 1673 67671 1731 67677
rect 5353 67711 5411 67717
rect 5353 67677 5365 67711
rect 5399 67677 5411 67711
rect 5353 67671 5411 67677
rect 1104 67482 5980 67504
rect 1104 67430 3802 67482
rect 3854 67430 3866 67482
rect 3918 67430 3930 67482
rect 3982 67430 3994 67482
rect 4046 67430 4058 67482
rect 4110 67430 5980 67482
rect 1104 67408 5980 67430
rect 1104 66938 5980 66960
rect 1104 66886 3066 66938
rect 3118 66886 3130 66938
rect 3182 66886 3194 66938
rect 3246 66886 3258 66938
rect 3310 66886 3322 66938
rect 3374 66886 5980 66938
rect 1104 66864 5980 66886
rect 1104 66394 5980 66416
rect 1104 66342 3802 66394
rect 3854 66342 3866 66394
rect 3918 66342 3930 66394
rect 3982 66342 3994 66394
rect 4046 66342 4058 66394
rect 4110 66342 5980 66394
rect 1104 66320 5980 66342
rect 1302 66104 1308 66156
rect 1360 66144 1366 66156
rect 1397 66147 1455 66153
rect 1397 66144 1409 66147
rect 1360 66116 1409 66144
rect 1360 66104 1366 66116
rect 1397 66113 1409 66116
rect 1443 66144 1455 66147
rect 1673 66147 1731 66153
rect 1673 66144 1685 66147
rect 1443 66116 1685 66144
rect 1443 66113 1455 66116
rect 1397 66107 1455 66113
rect 1673 66113 1685 66116
rect 1719 66113 1731 66147
rect 1673 66107 1731 66113
rect 4890 66104 4896 66156
rect 4948 66144 4954 66156
rect 5353 66147 5411 66153
rect 5353 66144 5365 66147
rect 4948 66116 5365 66144
rect 4948 66104 4954 66116
rect 5353 66113 5365 66116
rect 5399 66113 5411 66147
rect 5353 66107 5411 66113
rect 1581 66011 1639 66017
rect 1581 65977 1593 66011
rect 1627 66008 1639 66011
rect 8294 66008 8300 66020
rect 1627 65980 8300 66008
rect 1627 65977 1639 65980
rect 1581 65971 1639 65977
rect 8294 65968 8300 65980
rect 8352 65968 8358 66020
rect 4890 65900 4896 65952
rect 4948 65940 4954 65952
rect 5169 65943 5227 65949
rect 5169 65940 5181 65943
rect 4948 65912 5181 65940
rect 4948 65900 4954 65912
rect 5169 65909 5181 65912
rect 5215 65909 5227 65943
rect 5169 65903 5227 65909
rect 5537 65943 5595 65949
rect 5537 65909 5549 65943
rect 5583 65940 5595 65943
rect 7558 65940 7564 65952
rect 5583 65912 7564 65940
rect 5583 65909 5595 65912
rect 5537 65903 5595 65909
rect 7558 65900 7564 65912
rect 7616 65900 7622 65952
rect 1104 65850 5980 65872
rect 1104 65798 3066 65850
rect 3118 65798 3130 65850
rect 3182 65798 3194 65850
rect 3246 65798 3258 65850
rect 3310 65798 3322 65850
rect 3374 65798 5980 65850
rect 1104 65776 5980 65798
rect 1104 65306 5980 65328
rect 1104 65254 3802 65306
rect 3854 65254 3866 65306
rect 3918 65254 3930 65306
rect 3982 65254 3994 65306
rect 4046 65254 4058 65306
rect 4110 65254 5980 65306
rect 1104 65232 5980 65254
rect 5261 65195 5319 65201
rect 5261 65161 5273 65195
rect 5307 65192 5319 65195
rect 5350 65192 5356 65204
rect 5307 65164 5356 65192
rect 5307 65161 5319 65164
rect 5261 65155 5319 65161
rect 5350 65152 5356 65164
rect 5408 65152 5414 65204
rect 1302 65016 1308 65068
rect 1360 65056 1366 65068
rect 5368 65065 5396 65152
rect 1397 65059 1455 65065
rect 1397 65056 1409 65059
rect 1360 65028 1409 65056
rect 1360 65016 1366 65028
rect 1397 65025 1409 65028
rect 1443 65056 1455 65059
rect 1673 65059 1731 65065
rect 1673 65056 1685 65059
rect 1443 65028 1685 65056
rect 1443 65025 1455 65028
rect 1397 65019 1455 65025
rect 1673 65025 1685 65028
rect 1719 65025 1731 65059
rect 1673 65019 1731 65025
rect 5353 65059 5411 65065
rect 5353 65025 5365 65059
rect 5399 65025 5411 65059
rect 5353 65019 5411 65025
rect 5902 64988 5908 65000
rect 1596 64960 5908 64988
rect 1596 64929 1624 64960
rect 5902 64948 5908 64960
rect 5960 64948 5966 65000
rect 1581 64923 1639 64929
rect 1581 64889 1593 64923
rect 1627 64889 1639 64923
rect 1581 64883 1639 64889
rect 5534 64880 5540 64932
rect 5592 64880 5598 64932
rect 1104 64762 5980 64784
rect 1104 64710 3066 64762
rect 3118 64710 3130 64762
rect 3182 64710 3194 64762
rect 3246 64710 3258 64762
rect 3310 64710 3322 64762
rect 3374 64710 5980 64762
rect 1104 64688 5980 64710
rect 1104 64218 5980 64240
rect 1104 64166 3802 64218
rect 3854 64166 3866 64218
rect 3918 64166 3930 64218
rect 3982 64166 3994 64218
rect 4046 64166 4058 64218
rect 4110 64166 5980 64218
rect 1104 64144 5980 64166
rect 1104 63674 5980 63696
rect 1104 63622 3066 63674
rect 3118 63622 3130 63674
rect 3182 63622 3194 63674
rect 3246 63622 3258 63674
rect 3310 63622 3322 63674
rect 3374 63622 5980 63674
rect 1104 63600 5980 63622
rect 1581 63495 1639 63501
rect 1581 63461 1593 63495
rect 1627 63492 1639 63495
rect 8294 63492 8300 63504
rect 1627 63464 8300 63492
rect 1627 63461 1639 63464
rect 1581 63455 1639 63461
rect 8294 63452 8300 63464
rect 8352 63452 8358 63504
rect 1210 63316 1216 63368
rect 1268 63356 1274 63368
rect 1397 63359 1455 63365
rect 1397 63356 1409 63359
rect 1268 63328 1409 63356
rect 1268 63316 1274 63328
rect 1397 63325 1409 63328
rect 1443 63356 1455 63359
rect 1673 63359 1731 63365
rect 1673 63356 1685 63359
rect 1443 63328 1685 63356
rect 1443 63325 1455 63328
rect 1397 63319 1455 63325
rect 1673 63325 1685 63328
rect 1719 63325 1731 63359
rect 5353 63359 5411 63365
rect 5353 63356 5365 63359
rect 1673 63319 1731 63325
rect 5184 63328 5365 63356
rect 4522 63180 4528 63232
rect 4580 63220 4586 63232
rect 5184 63229 5212 63328
rect 5353 63325 5365 63328
rect 5399 63325 5411 63359
rect 5353 63319 5411 63325
rect 5169 63223 5227 63229
rect 5169 63220 5181 63223
rect 4580 63192 5181 63220
rect 4580 63180 4586 63192
rect 5169 63189 5181 63192
rect 5215 63189 5227 63223
rect 5169 63183 5227 63189
rect 5537 63223 5595 63229
rect 5537 63189 5549 63223
rect 5583 63220 5595 63223
rect 7650 63220 7656 63232
rect 5583 63192 7656 63220
rect 5583 63189 5595 63192
rect 5537 63183 5595 63189
rect 7650 63180 7656 63192
rect 7708 63180 7714 63232
rect 1104 63130 5980 63152
rect 1104 63078 3802 63130
rect 3854 63078 3866 63130
rect 3918 63078 3930 63130
rect 3982 63078 3994 63130
rect 4046 63078 4058 63130
rect 4110 63078 5980 63130
rect 1104 63056 5980 63078
rect 1104 62586 5980 62608
rect 1104 62534 3066 62586
rect 3118 62534 3130 62586
rect 3182 62534 3194 62586
rect 3246 62534 3258 62586
rect 3310 62534 3322 62586
rect 3374 62534 5980 62586
rect 1104 62512 5980 62534
rect 5258 62432 5264 62484
rect 5316 62432 5322 62484
rect 1581 62407 1639 62413
rect 1581 62373 1593 62407
rect 1627 62404 1639 62407
rect 5534 62404 5540 62416
rect 1627 62376 5540 62404
rect 1627 62373 1639 62376
rect 1581 62367 1639 62373
rect 5534 62364 5540 62376
rect 5592 62364 5598 62416
rect 1302 62228 1308 62280
rect 1360 62268 1366 62280
rect 1397 62271 1455 62277
rect 1397 62268 1409 62271
rect 1360 62240 1409 62268
rect 1360 62228 1366 62240
rect 1397 62237 1409 62240
rect 1443 62268 1455 62271
rect 1673 62271 1731 62277
rect 1673 62268 1685 62271
rect 1443 62240 1685 62268
rect 1443 62237 1455 62240
rect 1397 62231 1455 62237
rect 1673 62237 1685 62240
rect 1719 62237 1731 62271
rect 1673 62231 1731 62237
rect 5258 62228 5264 62280
rect 5316 62268 5322 62280
rect 5353 62271 5411 62277
rect 5353 62268 5365 62271
rect 5316 62240 5365 62268
rect 5316 62228 5322 62240
rect 5353 62237 5365 62240
rect 5399 62237 5411 62271
rect 5353 62231 5411 62237
rect 5537 62135 5595 62141
rect 5537 62101 5549 62135
rect 5583 62132 5595 62135
rect 5902 62132 5908 62144
rect 5583 62104 5908 62132
rect 5583 62101 5595 62104
rect 5537 62095 5595 62101
rect 5902 62092 5908 62104
rect 5960 62092 5966 62144
rect 1104 62042 5980 62064
rect 1104 61990 3802 62042
rect 3854 61990 3866 62042
rect 3918 61990 3930 62042
rect 3982 61990 3994 62042
rect 4046 61990 4058 62042
rect 4110 61990 5980 62042
rect 1104 61968 5980 61990
rect 1302 61752 1308 61804
rect 1360 61792 1366 61804
rect 1397 61795 1455 61801
rect 1397 61792 1409 61795
rect 1360 61764 1409 61792
rect 1360 61752 1366 61764
rect 1397 61761 1409 61764
rect 1443 61792 1455 61795
rect 1673 61795 1731 61801
rect 1673 61792 1685 61795
rect 1443 61764 1685 61792
rect 1443 61761 1455 61764
rect 1397 61755 1455 61761
rect 1673 61761 1685 61764
rect 1719 61761 1731 61795
rect 1673 61755 1731 61761
rect 1581 61659 1639 61665
rect 1581 61625 1593 61659
rect 1627 61656 1639 61659
rect 8294 61656 8300 61668
rect 1627 61628 8300 61656
rect 1627 61625 1639 61628
rect 1581 61619 1639 61625
rect 8294 61616 8300 61628
rect 8352 61616 8358 61668
rect 1104 61498 5980 61520
rect 1104 61446 3066 61498
rect 3118 61446 3130 61498
rect 3182 61446 3194 61498
rect 3246 61446 3258 61498
rect 3310 61446 3322 61498
rect 3374 61446 5980 61498
rect 1104 61424 5980 61446
rect 1104 60954 5980 60976
rect 1104 60902 3802 60954
rect 3854 60902 3866 60954
rect 3918 60902 3930 60954
rect 3982 60902 3994 60954
rect 4046 60902 4058 60954
rect 4110 60902 5980 60954
rect 1104 60880 5980 60902
rect 5166 60664 5172 60716
rect 5224 60704 5230 60716
rect 5353 60707 5411 60713
rect 5353 60704 5365 60707
rect 5224 60676 5365 60704
rect 5224 60664 5230 60676
rect 5353 60673 5365 60676
rect 5399 60673 5411 60707
rect 5353 60667 5411 60673
rect 842 60460 848 60512
rect 900 60500 906 60512
rect 1397 60503 1455 60509
rect 1397 60500 1409 60503
rect 900 60472 1409 60500
rect 900 60460 906 60472
rect 1397 60469 1409 60472
rect 1443 60469 1455 60503
rect 1397 60463 1455 60469
rect 5537 60503 5595 60509
rect 5537 60469 5549 60503
rect 5583 60500 5595 60503
rect 7834 60500 7840 60512
rect 5583 60472 7840 60500
rect 5583 60469 5595 60472
rect 5537 60463 5595 60469
rect 7834 60460 7840 60472
rect 7892 60460 7898 60512
rect 1104 60410 5980 60432
rect 1104 60358 3066 60410
rect 3118 60358 3130 60410
rect 3182 60358 3194 60410
rect 3246 60358 3258 60410
rect 3310 60358 3322 60410
rect 3374 60358 5980 60410
rect 1104 60336 5980 60358
rect 1210 60052 1216 60104
rect 1268 60092 1274 60104
rect 1397 60095 1455 60101
rect 1397 60092 1409 60095
rect 1268 60064 1409 60092
rect 1268 60052 1274 60064
rect 1397 60061 1409 60064
rect 1443 60092 1455 60095
rect 1673 60095 1731 60101
rect 1673 60092 1685 60095
rect 1443 60064 1685 60092
rect 1443 60061 1455 60064
rect 1397 60055 1455 60061
rect 1673 60061 1685 60064
rect 1719 60061 1731 60095
rect 1673 60055 1731 60061
rect 8294 60024 8300 60036
rect 1596 59996 8300 60024
rect 1596 59965 1624 59996
rect 8294 59984 8300 59996
rect 8352 59984 8358 60036
rect 1581 59959 1639 59965
rect 1581 59925 1593 59959
rect 1627 59925 1639 59959
rect 1581 59919 1639 59925
rect 1104 59866 5980 59888
rect 1104 59814 3802 59866
rect 3854 59814 3866 59866
rect 3918 59814 3930 59866
rect 3982 59814 3994 59866
rect 4046 59814 4058 59866
rect 4110 59814 5980 59866
rect 1104 59792 5980 59814
rect 5258 59576 5264 59628
rect 5316 59616 5322 59628
rect 5353 59619 5411 59625
rect 5353 59616 5365 59619
rect 5316 59588 5365 59616
rect 5316 59576 5322 59588
rect 5353 59585 5365 59588
rect 5399 59585 5411 59619
rect 5353 59579 5411 59585
rect 842 59372 848 59424
rect 900 59412 906 59424
rect 1397 59415 1455 59421
rect 1397 59412 1409 59415
rect 900 59384 1409 59412
rect 900 59372 906 59384
rect 1397 59381 1409 59384
rect 1443 59381 1455 59415
rect 1397 59375 1455 59381
rect 5258 59372 5264 59424
rect 5316 59372 5322 59424
rect 5537 59415 5595 59421
rect 5537 59381 5549 59415
rect 5583 59412 5595 59415
rect 5902 59412 5908 59424
rect 5583 59384 5908 59412
rect 5583 59381 5595 59384
rect 5537 59375 5595 59381
rect 5902 59372 5908 59384
rect 5960 59372 5966 59424
rect 1104 59322 5980 59344
rect 1104 59270 3066 59322
rect 3118 59270 3130 59322
rect 3182 59270 3194 59322
rect 3246 59270 3258 59322
rect 3310 59270 3322 59322
rect 3374 59270 5980 59322
rect 1104 59248 5980 59270
rect 1581 59143 1639 59149
rect 1581 59109 1593 59143
rect 1627 59140 1639 59143
rect 8294 59140 8300 59152
rect 1627 59112 8300 59140
rect 1627 59109 1639 59112
rect 1581 59103 1639 59109
rect 8294 59100 8300 59112
rect 8352 59100 8358 59152
rect 1302 58964 1308 59016
rect 1360 59004 1366 59016
rect 1397 59007 1455 59013
rect 1397 59004 1409 59007
rect 1360 58976 1409 59004
rect 1360 58964 1366 58976
rect 1397 58973 1409 58976
rect 1443 59004 1455 59007
rect 1673 59007 1731 59013
rect 1673 59004 1685 59007
rect 1443 58976 1685 59004
rect 1443 58973 1455 58976
rect 1397 58967 1455 58973
rect 1673 58973 1685 58976
rect 1719 58973 1731 59007
rect 1673 58967 1731 58973
rect 1104 58778 5980 58800
rect 1104 58726 3802 58778
rect 3854 58726 3866 58778
rect 3918 58726 3930 58778
rect 3982 58726 3994 58778
rect 4046 58726 4058 58778
rect 4110 58726 5980 58778
rect 1104 58704 5980 58726
rect 1104 58234 5980 58256
rect 1104 58182 3066 58234
rect 3118 58182 3130 58234
rect 3182 58182 3194 58234
rect 3246 58182 3258 58234
rect 3310 58182 3322 58234
rect 3374 58182 5980 58234
rect 1104 58160 5980 58182
rect 842 57944 848 57996
rect 900 57984 906 57996
rect 1397 57987 1455 57993
rect 1397 57984 1409 57987
rect 900 57956 1409 57984
rect 900 57944 906 57956
rect 1397 57953 1409 57956
rect 1443 57953 1455 57987
rect 1397 57947 1455 57953
rect 5353 57919 5411 57925
rect 5353 57885 5365 57919
rect 5399 57885 5411 57919
rect 5353 57879 5411 57885
rect 5261 57783 5319 57789
rect 5261 57749 5273 57783
rect 5307 57780 5319 57783
rect 5368 57780 5396 57879
rect 5442 57780 5448 57792
rect 5307 57752 5448 57780
rect 5307 57749 5319 57752
rect 5261 57743 5319 57749
rect 5442 57740 5448 57752
rect 5500 57740 5506 57792
rect 5537 57783 5595 57789
rect 5537 57749 5549 57783
rect 5583 57780 5595 57783
rect 7190 57780 7196 57792
rect 5583 57752 7196 57780
rect 5583 57749 5595 57752
rect 5537 57743 5595 57749
rect 7190 57740 7196 57752
rect 7248 57740 7254 57792
rect 1104 57690 5980 57712
rect 1104 57638 3802 57690
rect 3854 57638 3866 57690
rect 3918 57638 3930 57690
rect 3982 57638 3994 57690
rect 4046 57638 4058 57690
rect 4110 57638 5980 57690
rect 1104 57616 5980 57638
rect 5445 57579 5503 57585
rect 5445 57545 5457 57579
rect 5491 57576 5503 57579
rect 5626 57576 5632 57588
rect 5491 57548 5632 57576
rect 5491 57545 5503 57548
rect 5445 57539 5503 57545
rect 5626 57536 5632 57548
rect 5684 57536 5690 57588
rect 1302 57400 1308 57452
rect 1360 57440 1366 57452
rect 1397 57443 1455 57449
rect 1397 57440 1409 57443
rect 1360 57412 1409 57440
rect 1360 57400 1366 57412
rect 1397 57409 1409 57412
rect 1443 57440 1455 57443
rect 1673 57443 1731 57449
rect 1673 57440 1685 57443
rect 1443 57412 1685 57440
rect 1443 57409 1455 57412
rect 1397 57403 1455 57409
rect 1673 57409 1685 57412
rect 1719 57409 1731 57443
rect 1673 57403 1731 57409
rect 1581 57307 1639 57313
rect 1581 57273 1593 57307
rect 1627 57304 1639 57307
rect 8294 57304 8300 57316
rect 1627 57276 8300 57304
rect 1627 57273 1639 57276
rect 1581 57267 1639 57273
rect 8294 57264 8300 57276
rect 8352 57264 8358 57316
rect 5534 57196 5540 57248
rect 5592 57196 5598 57248
rect 1104 57146 5980 57168
rect 1104 57094 3066 57146
rect 3118 57094 3130 57146
rect 3182 57094 3194 57146
rect 3246 57094 3258 57146
rect 3310 57094 3322 57146
rect 3374 57094 5980 57146
rect 1104 57072 5980 57094
rect 842 56788 848 56840
rect 900 56828 906 56840
rect 1397 56831 1455 56837
rect 1397 56828 1409 56831
rect 900 56800 1409 56828
rect 900 56788 906 56800
rect 1397 56797 1409 56800
rect 1443 56797 1455 56831
rect 1397 56791 1455 56797
rect 5626 56788 5632 56840
rect 5684 56788 5690 56840
rect 4341 56695 4399 56701
rect 4341 56661 4353 56695
rect 4387 56692 4399 56695
rect 5534 56692 5540 56704
rect 4387 56664 5540 56692
rect 4387 56661 4399 56664
rect 4341 56655 4399 56661
rect 5534 56652 5540 56664
rect 5592 56652 5598 56704
rect 1104 56602 5980 56624
rect 1104 56550 3802 56602
rect 3854 56550 3866 56602
rect 3918 56550 3930 56602
rect 3982 56550 3994 56602
rect 4046 56550 4058 56602
rect 4110 56550 5980 56602
rect 1104 56528 5980 56550
rect 1302 56312 1308 56364
rect 1360 56352 1366 56364
rect 1397 56355 1455 56361
rect 1397 56352 1409 56355
rect 1360 56324 1409 56352
rect 1360 56312 1366 56324
rect 1397 56321 1409 56324
rect 1443 56352 1455 56355
rect 1673 56355 1731 56361
rect 1673 56352 1685 56355
rect 1443 56324 1685 56352
rect 1443 56321 1455 56324
rect 1397 56315 1455 56321
rect 1673 56321 1685 56324
rect 1719 56321 1731 56355
rect 1673 56315 1731 56321
rect 5074 56312 5080 56364
rect 5132 56352 5138 56364
rect 5353 56355 5411 56361
rect 5353 56352 5365 56355
rect 5132 56324 5365 56352
rect 5132 56312 5138 56324
rect 5353 56321 5365 56324
rect 5399 56321 5411 56355
rect 5353 56315 5411 56321
rect 1581 56219 1639 56225
rect 1581 56185 1593 56219
rect 1627 56216 1639 56219
rect 8294 56216 8300 56228
rect 1627 56188 8300 56216
rect 1627 56185 1639 56188
rect 1581 56179 1639 56185
rect 8294 56176 8300 56188
rect 8352 56176 8358 56228
rect 5074 56108 5080 56160
rect 5132 56148 5138 56160
rect 5169 56151 5227 56157
rect 5169 56148 5181 56151
rect 5132 56120 5181 56148
rect 5132 56108 5138 56120
rect 5169 56117 5181 56120
rect 5215 56117 5227 56151
rect 5169 56111 5227 56117
rect 5537 56151 5595 56157
rect 5537 56117 5549 56151
rect 5583 56148 5595 56151
rect 6730 56148 6736 56160
rect 5583 56120 6736 56148
rect 5583 56117 5595 56120
rect 5537 56111 5595 56117
rect 6730 56108 6736 56120
rect 6788 56108 6794 56160
rect 1104 56058 5980 56080
rect 1104 56006 3066 56058
rect 3118 56006 3130 56058
rect 3182 56006 3194 56058
rect 3246 56006 3258 56058
rect 3310 56006 3322 56058
rect 3374 56006 5980 56058
rect 1104 55984 5980 56006
rect 1104 55514 5980 55536
rect 1104 55462 3802 55514
rect 3854 55462 3866 55514
rect 3918 55462 3930 55514
rect 3982 55462 3994 55514
rect 4046 55462 4058 55514
rect 4110 55462 5980 55514
rect 1104 55440 5980 55462
rect 4890 55360 4896 55412
rect 4948 55400 4954 55412
rect 5169 55403 5227 55409
rect 5169 55400 5181 55403
rect 4948 55372 5181 55400
rect 4948 55360 4954 55372
rect 5169 55369 5181 55372
rect 5215 55369 5227 55403
rect 5169 55363 5227 55369
rect 5537 55403 5595 55409
rect 5537 55369 5549 55403
rect 5583 55400 5595 55403
rect 6822 55400 6828 55412
rect 5583 55372 6828 55400
rect 5583 55369 5595 55372
rect 5537 55363 5595 55369
rect 5184 55264 5212 55363
rect 6822 55360 6828 55372
rect 6880 55360 6886 55412
rect 5353 55267 5411 55273
rect 5353 55264 5365 55267
rect 5184 55236 5365 55264
rect 5353 55233 5365 55236
rect 5399 55233 5411 55267
rect 5353 55227 5411 55233
rect 842 55020 848 55072
rect 900 55060 906 55072
rect 1397 55063 1455 55069
rect 1397 55060 1409 55063
rect 900 55032 1409 55060
rect 900 55020 906 55032
rect 1397 55029 1409 55032
rect 1443 55029 1455 55063
rect 1397 55023 1455 55029
rect 1104 54970 5980 54992
rect 1104 54918 3066 54970
rect 3118 54918 3130 54970
rect 3182 54918 3194 54970
rect 3246 54918 3258 54970
rect 3310 54918 3322 54970
rect 3374 54918 5980 54970
rect 1104 54896 5980 54918
rect 1210 54612 1216 54664
rect 1268 54652 1274 54664
rect 1397 54655 1455 54661
rect 1397 54652 1409 54655
rect 1268 54624 1409 54652
rect 1268 54612 1274 54624
rect 1397 54621 1409 54624
rect 1443 54652 1455 54655
rect 1673 54655 1731 54661
rect 1673 54652 1685 54655
rect 1443 54624 1685 54652
rect 1443 54621 1455 54624
rect 1397 54615 1455 54621
rect 1673 54621 1685 54624
rect 1719 54621 1731 54655
rect 1673 54615 1731 54621
rect 8294 54584 8300 54596
rect 1596 54556 8300 54584
rect 1596 54525 1624 54556
rect 8294 54544 8300 54556
rect 8352 54544 8358 54596
rect 1581 54519 1639 54525
rect 1581 54485 1593 54519
rect 1627 54485 1639 54519
rect 1581 54479 1639 54485
rect 1104 54426 5980 54448
rect 1104 54374 3802 54426
rect 3854 54374 3866 54426
rect 3918 54374 3930 54426
rect 3982 54374 3994 54426
rect 4046 54374 4058 54426
rect 4110 54374 5980 54426
rect 1104 54352 5980 54374
rect 4706 54272 4712 54324
rect 4764 54312 4770 54324
rect 4890 54312 4896 54324
rect 4764 54284 4896 54312
rect 4764 54272 4770 54284
rect 4890 54272 4896 54284
rect 4948 54272 4954 54324
rect 5353 54179 5411 54185
rect 5353 54176 5365 54179
rect 5184 54148 5365 54176
rect 842 53932 848 53984
rect 900 53972 906 53984
rect 1397 53975 1455 53981
rect 1397 53972 1409 53975
rect 900 53944 1409 53972
rect 900 53932 906 53944
rect 1397 53941 1409 53944
rect 1443 53941 1455 53975
rect 1397 53935 1455 53941
rect 5074 53932 5080 53984
rect 5132 53972 5138 53984
rect 5184 53981 5212 54148
rect 5353 54145 5365 54148
rect 5399 54145 5411 54179
rect 5353 54139 5411 54145
rect 5169 53975 5227 53981
rect 5169 53972 5181 53975
rect 5132 53944 5181 53972
rect 5132 53932 5138 53944
rect 5169 53941 5181 53944
rect 5215 53941 5227 53975
rect 5169 53935 5227 53941
rect 5537 53975 5595 53981
rect 5537 53941 5549 53975
rect 5583 53972 5595 53975
rect 7926 53972 7932 53984
rect 5583 53944 7932 53972
rect 5583 53941 5595 53944
rect 5537 53935 5595 53941
rect 7926 53932 7932 53944
rect 7984 53932 7990 53984
rect 1104 53882 5980 53904
rect 1104 53830 3066 53882
rect 3118 53830 3130 53882
rect 3182 53830 3194 53882
rect 3246 53830 3258 53882
rect 3310 53830 3322 53882
rect 3374 53830 5980 53882
rect 1104 53808 5980 53830
rect 1581 53703 1639 53709
rect 1581 53669 1593 53703
rect 1627 53700 1639 53703
rect 8294 53700 8300 53712
rect 1627 53672 8300 53700
rect 1627 53669 1639 53672
rect 1581 53663 1639 53669
rect 8294 53660 8300 53672
rect 8352 53660 8358 53712
rect 1302 53524 1308 53576
rect 1360 53564 1366 53576
rect 1397 53567 1455 53573
rect 1397 53564 1409 53567
rect 1360 53536 1409 53564
rect 1360 53524 1366 53536
rect 1397 53533 1409 53536
rect 1443 53564 1455 53567
rect 1673 53567 1731 53573
rect 1673 53564 1685 53567
rect 1443 53536 1685 53564
rect 1443 53533 1455 53536
rect 1397 53527 1455 53533
rect 1673 53533 1685 53536
rect 1719 53533 1731 53567
rect 1673 53527 1731 53533
rect 1104 53338 5980 53360
rect 1104 53286 3802 53338
rect 3854 53286 3866 53338
rect 3918 53286 3930 53338
rect 3982 53286 3994 53338
rect 4046 53286 4058 53338
rect 4110 53286 5980 53338
rect 1104 53264 5980 53286
rect 1104 52794 5980 52816
rect 1104 52742 3066 52794
rect 3118 52742 3130 52794
rect 3182 52742 3194 52794
rect 3246 52742 3258 52794
rect 3310 52742 3322 52794
rect 3374 52742 5980 52794
rect 1104 52720 5980 52742
rect 5537 52615 5595 52621
rect 5537 52581 5549 52615
rect 5583 52612 5595 52615
rect 8202 52612 8208 52624
rect 5583 52584 8208 52612
rect 5583 52581 5595 52584
rect 5537 52575 5595 52581
rect 8202 52572 8208 52584
rect 8260 52572 8266 52624
rect 842 52436 848 52488
rect 900 52476 906 52488
rect 1397 52479 1455 52485
rect 1397 52476 1409 52479
rect 900 52448 1409 52476
rect 900 52436 906 52448
rect 1397 52445 1409 52448
rect 1443 52445 1455 52479
rect 1397 52439 1455 52445
rect 5166 52436 5172 52488
rect 5224 52476 5230 52488
rect 5353 52479 5411 52485
rect 5353 52476 5365 52479
rect 5224 52448 5365 52476
rect 5224 52436 5230 52448
rect 5353 52445 5365 52448
rect 5399 52445 5411 52479
rect 5353 52439 5411 52445
rect 1104 52250 5980 52272
rect 1104 52198 3802 52250
rect 3854 52198 3866 52250
rect 3918 52198 3930 52250
rect 3982 52198 3994 52250
rect 4046 52198 4058 52250
rect 4110 52198 5980 52250
rect 1104 52176 5980 52198
rect 842 51892 848 51944
rect 900 51932 906 51944
rect 1397 51935 1455 51941
rect 1397 51932 1409 51935
rect 900 51904 1409 51932
rect 900 51892 906 51904
rect 1397 51901 1409 51904
rect 1443 51901 1455 51935
rect 1397 51895 1455 51901
rect 1104 51706 5980 51728
rect 1104 51654 3066 51706
rect 3118 51654 3130 51706
rect 3182 51654 3194 51706
rect 3246 51654 3258 51706
rect 3310 51654 3322 51706
rect 3374 51654 5980 51706
rect 1104 51632 5980 51654
rect 1026 51348 1032 51400
rect 1084 51388 1090 51400
rect 1397 51391 1455 51397
rect 1397 51388 1409 51391
rect 1084 51360 1409 51388
rect 1084 51348 1090 51360
rect 1397 51357 1409 51360
rect 1443 51357 1455 51391
rect 5353 51391 5411 51397
rect 5353 51388 5365 51391
rect 1397 51351 1455 51357
rect 5276 51360 5365 51388
rect 5276 51264 5304 51360
rect 5353 51357 5365 51360
rect 5399 51357 5411 51391
rect 5353 51351 5411 51357
rect 5258 51212 5264 51264
rect 5316 51212 5322 51264
rect 5537 51255 5595 51261
rect 5537 51221 5549 51255
rect 5583 51252 5595 51255
rect 5583 51224 6914 51252
rect 5583 51221 5595 51224
rect 5537 51215 5595 51221
rect 1104 51162 5980 51184
rect 1104 51110 3802 51162
rect 3854 51110 3866 51162
rect 3918 51110 3930 51162
rect 3982 51110 3994 51162
rect 4046 51110 4058 51162
rect 4110 51110 5980 51162
rect 1104 51088 5980 51110
rect 6886 51048 6914 51224
rect 87138 51048 87144 51060
rect 6886 51020 87144 51048
rect 87138 51008 87144 51020
rect 87196 51008 87202 51060
rect 6546 50940 6552 50992
rect 6604 50980 6610 50992
rect 6730 50980 6736 50992
rect 6604 50952 6736 50980
rect 6604 50940 6610 50952
rect 6730 50940 6736 50952
rect 6788 50940 6794 50992
rect 7558 50940 7564 50992
rect 7616 50980 7622 50992
rect 89070 50980 89076 50992
rect 7616 50952 89076 50980
rect 7616 50940 7622 50952
rect 89070 50940 89076 50952
rect 89128 50940 89134 50992
rect 4893 50915 4951 50921
rect 4893 50881 4905 50915
rect 4939 50912 4951 50915
rect 5350 50912 5356 50924
rect 4939 50884 5356 50912
rect 4939 50881 4951 50884
rect 4893 50875 4951 50881
rect 5350 50872 5356 50884
rect 5408 50872 5414 50924
rect 5077 50847 5135 50853
rect 5077 50813 5089 50847
rect 5123 50844 5135 50847
rect 5626 50844 5632 50856
rect 5123 50816 5632 50844
rect 5123 50813 5135 50816
rect 5077 50807 5135 50813
rect 5626 50804 5632 50816
rect 5684 50804 5690 50856
rect 7926 50804 7932 50856
rect 7984 50844 7990 50856
rect 88334 50844 88340 50856
rect 7984 50816 88340 50844
rect 7984 50804 7990 50816
rect 88334 50804 88340 50816
rect 88392 50804 88398 50856
rect 5261 50779 5319 50785
rect 5261 50745 5273 50779
rect 5307 50776 5319 50779
rect 6638 50776 6644 50788
rect 5307 50748 6644 50776
rect 5307 50745 5319 50748
rect 5261 50739 5319 50745
rect 6638 50736 6644 50748
rect 6696 50736 6702 50788
rect 1394 50668 1400 50720
rect 1452 50668 1458 50720
rect 5537 50711 5595 50717
rect 5537 50677 5549 50711
rect 5583 50708 5595 50711
rect 6730 50708 6736 50720
rect 5583 50680 6736 50708
rect 5583 50677 5595 50680
rect 5537 50671 5595 50677
rect 6730 50668 6736 50680
rect 6788 50668 6794 50720
rect 1104 50618 5980 50640
rect 1104 50566 3066 50618
rect 3118 50566 3130 50618
rect 3182 50566 3194 50618
rect 3246 50566 3258 50618
rect 3310 50566 3322 50618
rect 3374 50566 5980 50618
rect 6638 50600 6644 50652
rect 6696 50640 6702 50652
rect 9582 50640 9588 50652
rect 6696 50612 9588 50640
rect 6696 50600 6702 50612
rect 9582 50600 9588 50612
rect 9640 50600 9646 50652
rect 46842 50600 46848 50652
rect 46900 50640 46906 50652
rect 85574 50640 85580 50652
rect 46900 50612 85580 50640
rect 46900 50600 46906 50612
rect 85574 50600 85580 50612
rect 85632 50600 85638 50652
rect 1104 50544 5980 50566
rect 8202 50532 8208 50584
rect 8260 50572 8266 50584
rect 88426 50572 88432 50584
rect 8260 50544 88432 50572
rect 8260 50532 8266 50544
rect 88426 50532 88432 50544
rect 88484 50532 88490 50584
rect 5626 50464 5632 50516
rect 5684 50504 5690 50516
rect 6638 50504 6644 50516
rect 5684 50476 6644 50504
rect 5684 50464 5690 50476
rect 6638 50464 6644 50476
rect 6696 50504 6702 50516
rect 11606 50504 11612 50516
rect 6696 50476 11612 50504
rect 6696 50464 6702 50476
rect 11606 50464 11612 50476
rect 11664 50464 11670 50516
rect 47486 50436 47492 50448
rect 26206 50408 47492 50436
rect 5445 50303 5503 50309
rect 5445 50269 5457 50303
rect 5491 50300 5503 50303
rect 8202 50300 8208 50312
rect 5491 50272 8208 50300
rect 5491 50269 5503 50272
rect 5445 50263 5503 50269
rect 8202 50260 8208 50272
rect 8260 50300 8266 50312
rect 13078 50300 13084 50312
rect 8260 50272 13084 50300
rect 8260 50260 8266 50272
rect 13078 50260 13084 50272
rect 13136 50300 13142 50312
rect 26206 50300 26234 50408
rect 47486 50396 47492 50408
rect 47544 50436 47550 50448
rect 52638 50436 52644 50448
rect 47544 50408 52644 50436
rect 47544 50396 47550 50408
rect 52638 50396 52644 50408
rect 52696 50396 52702 50448
rect 13136 50272 26234 50300
rect 13136 50260 13142 50272
rect 12250 50192 12256 50244
rect 12308 50232 12314 50244
rect 47394 50232 47400 50244
rect 12308 50204 47400 50232
rect 12308 50192 12314 50204
rect 47394 50192 47400 50204
rect 47452 50232 47458 50244
rect 51534 50232 51540 50244
rect 47452 50204 51540 50232
rect 47452 50192 47458 50204
rect 51534 50192 51540 50204
rect 51592 50192 51598 50244
rect 5629 50167 5687 50173
rect 5629 50133 5641 50167
rect 5675 50164 5687 50167
rect 8018 50164 8024 50176
rect 5675 50136 8024 50164
rect 5675 50133 5687 50136
rect 5629 50127 5687 50133
rect 8018 50124 8024 50136
rect 8076 50124 8082 50176
rect 10870 50124 10876 50176
rect 10928 50164 10934 50176
rect 47762 50164 47768 50176
rect 10928 50136 47768 50164
rect 10928 50124 10934 50136
rect 47762 50124 47768 50136
rect 47820 50164 47826 50176
rect 50430 50164 50436 50176
rect 47820 50136 50436 50164
rect 47820 50124 47826 50136
rect 50430 50124 50436 50136
rect 50488 50124 50494 50176
rect 1104 50074 5980 50096
rect 1104 50022 3802 50074
rect 3854 50022 3866 50074
rect 3918 50022 3930 50074
rect 3982 50022 3994 50074
rect 4046 50022 4058 50074
rect 4110 50022 5980 50074
rect 1104 50000 5980 50022
rect 8018 49920 8024 49972
rect 8076 49960 8082 49972
rect 10502 49960 10508 49972
rect 8076 49932 10508 49960
rect 8076 49920 8082 49932
rect 10502 49920 10508 49932
rect 10560 49920 10566 49972
rect 4614 49852 4620 49904
rect 4672 49892 4678 49904
rect 86678 49892 86684 49904
rect 4672 49864 86684 49892
rect 4672 49852 4678 49864
rect 86678 49852 86684 49864
rect 86736 49852 86742 49904
rect 6454 49784 6460 49836
rect 6512 49824 6518 49836
rect 6512 49796 12434 49824
rect 6512 49784 6518 49796
rect 6086 49716 6092 49768
rect 6144 49756 6150 49768
rect 9674 49756 9680 49768
rect 6144 49728 9680 49756
rect 6144 49716 6150 49728
rect 9674 49716 9680 49728
rect 9732 49716 9738 49768
rect 12406 49756 12434 49796
rect 46842 49784 46848 49836
rect 46900 49824 46906 49836
rect 47670 49824 47676 49836
rect 46900 49796 47676 49824
rect 46900 49784 46906 49796
rect 47670 49784 47676 49796
rect 47728 49824 47734 49836
rect 49694 49824 49700 49836
rect 47728 49796 49700 49824
rect 47728 49784 47734 49796
rect 49694 49784 49700 49796
rect 49752 49784 49758 49836
rect 86862 49756 86868 49768
rect 12406 49728 86868 49756
rect 86862 49716 86868 49728
rect 86920 49716 86926 49768
rect 5810 49648 5816 49700
rect 5868 49688 5874 49700
rect 89162 49688 89168 49700
rect 5868 49660 89168 49688
rect 5868 49648 5874 49660
rect 89162 49648 89168 49660
rect 89220 49648 89226 49700
rect 1394 49580 1400 49632
rect 1452 49580 1458 49632
rect 6822 49580 6828 49632
rect 6880 49620 6886 49632
rect 88518 49620 88524 49632
rect 6880 49592 88524 49620
rect 6880 49580 6886 49592
rect 88518 49580 88524 49592
rect 88576 49580 88582 49632
rect 1104 49530 5980 49552
rect 1104 49478 3066 49530
rect 3118 49478 3130 49530
rect 3182 49478 3194 49530
rect 3246 49478 3258 49530
rect 3310 49478 3322 49530
rect 3374 49478 5980 49530
rect 1104 49456 5980 49478
rect 47762 49444 47768 49496
rect 47820 49484 47826 49496
rect 48222 49484 48228 49496
rect 47820 49456 48228 49484
rect 47820 49444 47826 49456
rect 48222 49444 48228 49456
rect 48280 49444 48286 49496
rect 4890 49376 4896 49428
rect 4948 49416 4954 49428
rect 87414 49416 87420 49428
rect 4948 49388 87420 49416
rect 4948 49376 4954 49388
rect 87414 49376 87420 49388
rect 87472 49376 87478 49428
rect 1394 49308 1400 49360
rect 1452 49308 1458 49360
rect 7650 49308 7656 49360
rect 7708 49348 7714 49360
rect 88886 49348 88892 49360
rect 7708 49320 88892 49348
rect 7708 49308 7714 49320
rect 88886 49308 88892 49320
rect 88944 49308 88950 49360
rect 7834 49240 7840 49292
rect 7892 49280 7898 49292
rect 88794 49280 88800 49292
rect 7892 49252 88800 49280
rect 7892 49240 7898 49252
rect 88794 49240 88800 49252
rect 88852 49240 88858 49292
rect 7190 49172 7196 49224
rect 7248 49212 7254 49224
rect 88610 49212 88616 49224
rect 7248 49184 88616 49212
rect 7248 49172 7254 49184
rect 88610 49172 88616 49184
rect 88668 49172 88674 49224
rect 5258 49104 5264 49156
rect 5316 49144 5322 49156
rect 48130 49144 48136 49156
rect 5316 49116 48136 49144
rect 5316 49104 5322 49116
rect 48130 49104 48136 49116
rect 48188 49144 48194 49156
rect 87138 49144 87144 49156
rect 48188 49116 87144 49144
rect 48188 49104 48194 49116
rect 87138 49104 87144 49116
rect 87196 49104 87202 49156
rect 5166 49036 5172 49088
rect 5224 49076 5230 49088
rect 47946 49076 47952 49088
rect 5224 49048 47952 49076
rect 5224 49036 5230 49048
rect 47946 49036 47952 49048
rect 48004 49076 48010 49088
rect 48222 49076 48228 49088
rect 48004 49048 48228 49076
rect 48004 49036 48010 49048
rect 48222 49036 48228 49048
rect 48280 49036 48286 49088
rect 1104 48986 5980 49008
rect 1104 48934 3802 48986
rect 3854 48934 3866 48986
rect 3918 48934 3930 48986
rect 3982 48934 3994 48986
rect 4046 48934 4058 48986
rect 4110 48934 5980 48986
rect 1104 48912 5980 48934
rect 1578 48832 1584 48884
rect 1636 48832 1642 48884
rect 5350 48832 5356 48884
rect 5408 48872 5414 48884
rect 46842 48872 46848 48884
rect 5408 48844 46848 48872
rect 5408 48832 5414 48844
rect 46842 48832 46848 48844
rect 46900 48832 46906 48884
rect 5902 48764 5908 48816
rect 5960 48804 5966 48816
rect 87782 48804 87788 48816
rect 5960 48776 87788 48804
rect 5960 48764 5966 48776
rect 87782 48764 87788 48776
rect 87840 48764 87846 48816
rect 1302 48696 1308 48748
rect 1360 48736 1366 48748
rect 1397 48739 1455 48745
rect 1397 48736 1409 48739
rect 1360 48708 1409 48736
rect 1360 48696 1366 48708
rect 1397 48705 1409 48708
rect 1443 48736 1455 48739
rect 1673 48739 1731 48745
rect 1673 48736 1685 48739
rect 1443 48708 1685 48736
rect 1443 48705 1455 48708
rect 1397 48699 1455 48705
rect 1673 48705 1685 48708
rect 1719 48705 1731 48739
rect 1673 48699 1731 48705
rect 6546 48696 6552 48748
rect 6604 48736 6610 48748
rect 88702 48736 88708 48748
rect 6604 48708 88708 48736
rect 6604 48696 6610 48708
rect 88702 48696 88708 48708
rect 88760 48696 88766 48748
rect 6178 48628 6184 48680
rect 6236 48668 6242 48680
rect 89346 48668 89352 48680
rect 6236 48640 89352 48668
rect 6236 48628 6242 48640
rect 89346 48628 89352 48640
rect 89404 48628 89410 48680
rect 5166 48560 5172 48612
rect 5224 48600 5230 48612
rect 89070 48600 89076 48612
rect 5224 48572 89076 48600
rect 5224 48560 5230 48572
rect 89070 48560 89076 48572
rect 89128 48560 89134 48612
rect 47946 48492 47952 48544
rect 48004 48532 48010 48544
rect 87322 48532 87328 48544
rect 48004 48504 87328 48532
rect 48004 48492 48010 48504
rect 87322 48492 87328 48504
rect 87380 48492 87386 48544
rect 1104 48442 5980 48464
rect 1104 48390 3066 48442
rect 3118 48390 3130 48442
rect 3182 48390 3194 48442
rect 3246 48390 3258 48442
rect 3310 48390 3322 48442
rect 3374 48390 5980 48442
rect 7006 48424 7012 48476
rect 7064 48464 7070 48476
rect 86678 48464 86684 48476
rect 7064 48436 86684 48464
rect 7064 48424 7070 48436
rect 86678 48424 86684 48436
rect 86736 48424 86742 48476
rect 1104 48368 5980 48390
rect 5718 48220 5724 48272
rect 5776 48260 5782 48272
rect 89254 48260 89260 48272
rect 5776 48232 89260 48260
rect 5776 48220 5782 48232
rect 89254 48220 89260 48232
rect 89312 48220 89318 48272
rect 6270 48152 6276 48204
rect 6328 48192 6334 48204
rect 86770 48192 86776 48204
rect 6328 48164 86776 48192
rect 6328 48152 6334 48164
rect 86770 48152 86776 48164
rect 86828 48152 86834 48204
rect 1394 48084 1400 48136
rect 1452 48084 1458 48136
rect 9674 48084 9680 48136
rect 9732 48124 9738 48136
rect 88978 48124 88984 48136
rect 9732 48096 88984 48124
rect 9732 48084 9738 48096
rect 88978 48084 88984 48096
rect 89036 48084 89042 48136
rect 6730 48016 6736 48068
rect 6788 48056 6794 48068
rect 46750 48056 46756 48068
rect 6788 48028 46756 48056
rect 6788 48016 6794 48028
rect 46750 48016 46756 48028
rect 46808 48016 46814 48068
rect 1104 47898 5980 47920
rect 1104 47846 3802 47898
rect 3854 47846 3866 47898
rect 3918 47846 3930 47898
rect 3982 47846 3994 47898
rect 4046 47846 4058 47898
rect 4110 47846 5980 47898
rect 1104 47824 5980 47846
rect 5626 47676 5632 47728
rect 5684 47716 5690 47728
rect 51166 47716 51172 47728
rect 5684 47688 51172 47716
rect 5684 47676 5690 47688
rect 51166 47676 51172 47688
rect 51224 47676 51230 47728
rect 5074 47608 5080 47660
rect 5132 47648 5138 47660
rect 88702 47648 88708 47660
rect 5132 47620 88708 47648
rect 5132 47608 5138 47620
rect 88702 47608 88708 47620
rect 88760 47608 88766 47660
rect 6914 47540 6920 47592
rect 6972 47580 6978 47592
rect 10502 47580 10508 47592
rect 6972 47552 10508 47580
rect 6972 47540 6978 47552
rect 10502 47540 10508 47552
rect 10560 47540 10566 47592
rect 11238 47540 11244 47592
rect 11296 47580 11302 47592
rect 46842 47580 46848 47592
rect 11296 47552 46848 47580
rect 11296 47540 11302 47552
rect 46842 47540 46848 47552
rect 46900 47540 46906 47592
rect 47486 47540 47492 47592
rect 47544 47580 47550 47592
rect 89438 47580 89444 47592
rect 47544 47552 89444 47580
rect 47544 47540 47550 47552
rect 89438 47540 89444 47552
rect 89496 47540 89502 47592
rect 11422 47472 11428 47524
rect 11480 47512 11486 47524
rect 11480 47484 12434 47512
rect 11480 47472 11486 47484
rect 5442 47404 5448 47456
rect 5500 47444 5506 47456
rect 11146 47444 11152 47456
rect 5500 47416 11152 47444
rect 5500 47404 5506 47416
rect 11146 47404 11152 47416
rect 11204 47404 11210 47456
rect 12406 47444 12434 47484
rect 48130 47472 48136 47524
rect 48188 47512 48194 47524
rect 89162 47512 89168 47524
rect 48188 47484 89168 47512
rect 48188 47472 48194 47484
rect 89162 47472 89168 47484
rect 89220 47472 89226 47524
rect 88334 47444 88340 47456
rect 12406 47416 88340 47444
rect 88334 47404 88340 47416
rect 88392 47404 88398 47456
rect 1104 47354 5980 47376
rect 1104 47302 3066 47354
rect 3118 47302 3130 47354
rect 3182 47302 3194 47354
rect 3246 47302 3258 47354
rect 3310 47302 3322 47354
rect 3374 47302 5980 47354
rect 6546 47336 6552 47388
rect 6604 47376 6610 47388
rect 86954 47376 86960 47388
rect 6604 47348 86960 47376
rect 6604 47336 6610 47348
rect 86954 47336 86960 47348
rect 87012 47336 87018 47388
rect 1104 47280 5980 47302
rect 6086 47268 6092 47320
rect 6144 47308 6150 47320
rect 10410 47308 10416 47320
rect 6144 47280 10416 47308
rect 6144 47268 6150 47280
rect 10410 47268 10416 47280
rect 10468 47268 10474 47320
rect 10502 47268 10508 47320
rect 10560 47308 10566 47320
rect 88518 47308 88524 47320
rect 10560 47280 88524 47308
rect 10560 47268 10566 47280
rect 88518 47268 88524 47280
rect 88576 47268 88582 47320
rect 5534 47200 5540 47252
rect 5592 47240 5598 47252
rect 10226 47240 10232 47252
rect 5592 47212 10232 47240
rect 5592 47200 5598 47212
rect 10226 47200 10232 47212
rect 10284 47200 10290 47252
rect 88610 47240 88616 47252
rect 10336 47212 88616 47240
rect 7834 47132 7840 47184
rect 7892 47172 7898 47184
rect 10336 47172 10364 47212
rect 88610 47200 88616 47212
rect 88668 47200 88674 47252
rect 7892 47144 10364 47172
rect 7892 47132 7898 47144
rect 10410 47132 10416 47184
rect 10468 47172 10474 47184
rect 87690 47172 87696 47184
rect 10468 47144 87696 47172
rect 10468 47132 10474 47144
rect 87690 47132 87696 47144
rect 87748 47132 87754 47184
rect 6270 47064 6276 47116
rect 6328 47104 6334 47116
rect 88794 47104 88800 47116
rect 6328 47076 88800 47104
rect 6328 47064 6334 47076
rect 88794 47064 88800 47076
rect 88852 47064 88858 47116
rect 1394 46996 1400 47048
rect 1452 46996 1458 47048
rect 5261 47039 5319 47045
rect 5261 47005 5273 47039
rect 5307 47036 5319 47039
rect 11054 47036 11060 47048
rect 5307 47008 11060 47036
rect 5307 47005 5319 47008
rect 5261 46999 5319 47005
rect 11054 46996 11060 47008
rect 11112 46996 11118 47048
rect 11146 46996 11152 47048
rect 11204 47036 11210 47048
rect 88426 47036 88432 47048
rect 11204 47008 88432 47036
rect 11204 46996 11210 47008
rect 88426 46996 88432 47008
rect 88484 46996 88490 47048
rect 5445 46971 5503 46977
rect 5445 46937 5457 46971
rect 5491 46968 5503 46971
rect 5491 46940 8248 46968
rect 5491 46937 5503 46940
rect 5445 46931 5503 46937
rect 8220 46900 8248 46940
rect 9674 46928 9680 46980
rect 9732 46968 9738 46980
rect 11422 46968 11428 46980
rect 9732 46940 11428 46968
rect 9732 46928 9738 46940
rect 11422 46928 11428 46940
rect 11480 46928 11486 46980
rect 12526 46900 12532 46912
rect 8220 46872 12532 46900
rect 12526 46860 12532 46872
rect 12584 46860 12590 46912
rect 1104 46810 5980 46832
rect 1104 46758 3802 46810
rect 3854 46758 3866 46810
rect 3918 46758 3930 46810
rect 3982 46758 3994 46810
rect 4046 46758 4058 46810
rect 4110 46758 5980 46810
rect 48038 46792 48044 46844
rect 48096 46832 48102 46844
rect 52546 46832 52552 46844
rect 48096 46804 52552 46832
rect 48096 46792 48102 46804
rect 52546 46792 52552 46804
rect 52604 46792 52610 46844
rect 51442 46764 51448 46776
rect 1104 46736 5980 46758
rect 47780 46736 51448 46764
rect 47780 46708 47808 46736
rect 51442 46724 51448 46736
rect 51500 46724 51506 46776
rect 6822 46656 6828 46708
rect 6880 46696 6886 46708
rect 13262 46696 13268 46708
rect 6880 46668 13268 46696
rect 6880 46656 6886 46668
rect 13262 46656 13268 46668
rect 13320 46656 13326 46708
rect 47762 46696 47768 46708
rect 45526 46668 47768 46696
rect 11698 46588 11704 46640
rect 11756 46628 11762 46640
rect 45526 46628 45554 46668
rect 47762 46656 47768 46668
rect 47820 46656 47826 46708
rect 51074 46656 51080 46708
rect 51132 46696 51138 46708
rect 51132 46668 55214 46696
rect 51132 46656 51138 46668
rect 11756 46600 45554 46628
rect 11756 46588 11762 46600
rect 47670 46588 47676 46640
rect 47728 46628 47734 46640
rect 55186 46628 55214 46668
rect 89254 46628 89260 46640
rect 47728 46600 53328 46628
rect 55186 46600 89260 46628
rect 47728 46588 47734 46600
rect 47854 46520 47860 46572
rect 47912 46560 47918 46572
rect 53190 46560 53196 46572
rect 47912 46532 53196 46560
rect 47912 46520 47918 46532
rect 53190 46520 53196 46532
rect 53248 46520 53254 46572
rect 53300 46560 53328 46600
rect 89254 46588 89260 46600
rect 89312 46588 89318 46640
rect 87598 46560 87604 46572
rect 53300 46532 87604 46560
rect 87598 46520 87604 46532
rect 87656 46520 87662 46572
rect 4798 46452 4804 46504
rect 4856 46492 4862 46504
rect 4856 46464 9812 46492
rect 4856 46452 4862 46464
rect 9674 46384 9680 46436
rect 9732 46384 9738 46436
rect 1394 46316 1400 46368
rect 1452 46316 1458 46368
rect 1104 46266 5980 46288
rect 1104 46214 3066 46266
rect 3118 46214 3130 46266
rect 3182 46214 3194 46266
rect 3246 46214 3258 46266
rect 3310 46214 3322 46266
rect 3374 46214 5980 46266
rect 1104 46192 5980 46214
rect 5261 46087 5319 46093
rect 5261 46053 5273 46087
rect 5307 46084 5319 46087
rect 5629 46087 5687 46093
rect 5629 46084 5641 46087
rect 5307 46056 5641 46084
rect 5307 46053 5319 46056
rect 5261 46047 5319 46053
rect 5629 46053 5641 46056
rect 5675 46084 5687 46087
rect 8386 46084 8392 46096
rect 5675 46056 8392 46084
rect 5675 46053 5687 46056
rect 5629 46047 5687 46053
rect 8386 46044 8392 46056
rect 8444 46044 8450 46096
rect 1673 45951 1731 45957
rect 1673 45917 1685 45951
rect 1719 45948 1731 45951
rect 8294 45948 8300 45960
rect 1719 45920 8300 45948
rect 1719 45917 1731 45920
rect 1673 45911 1731 45917
rect 8294 45908 8300 45920
rect 8352 45908 8358 45960
rect 5077 45883 5135 45889
rect 5077 45849 5089 45883
rect 5123 45880 5135 45883
rect 5445 45883 5503 45889
rect 5445 45880 5457 45883
rect 5123 45852 5457 45880
rect 5123 45849 5135 45852
rect 5077 45843 5135 45849
rect 5445 45849 5457 45852
rect 5491 45880 5503 45883
rect 9692 45880 9720 46384
rect 9784 46356 9812 46464
rect 10318 46452 10324 46504
rect 10376 46492 10382 46504
rect 10376 46464 48268 46492
rect 10376 46452 10382 46464
rect 48240 46436 48268 46464
rect 51166 46452 51172 46504
rect 51224 46492 51230 46504
rect 88978 46492 88984 46504
rect 51224 46464 88984 46492
rect 51224 46452 51230 46464
rect 88978 46452 88984 46464
rect 89036 46452 89042 46504
rect 12526 46384 12532 46436
rect 12584 46424 12590 46436
rect 48038 46424 48044 46436
rect 12584 46396 48044 46424
rect 12584 46384 12590 46396
rect 48038 46384 48044 46396
rect 48096 46384 48102 46436
rect 48222 46384 48228 46436
rect 48280 46424 48286 46436
rect 49878 46424 49884 46436
rect 48280 46396 49884 46424
rect 48280 46384 48286 46396
rect 49878 46384 49884 46396
rect 49936 46384 49942 46436
rect 48130 46356 48136 46368
rect 9784 46328 48136 46356
rect 48130 46316 48136 46328
rect 48188 46316 48194 46368
rect 5491 45852 9720 45880
rect 5491 45849 5503 45852
rect 5445 45843 5503 45849
rect 1486 45772 1492 45824
rect 1544 45772 1550 45824
rect 1104 45722 5980 45744
rect 1104 45670 3802 45722
rect 3854 45670 3866 45722
rect 3918 45670 3930 45722
rect 3982 45670 3994 45722
rect 4046 45670 4058 45722
rect 4110 45670 5980 45722
rect 1104 45648 5980 45670
rect 1394 45228 1400 45280
rect 1452 45228 1458 45280
rect 1104 45178 5980 45200
rect 1104 45126 3066 45178
rect 3118 45126 3130 45178
rect 3182 45126 3194 45178
rect 3246 45126 3258 45178
rect 3310 45126 3322 45178
rect 3374 45126 5980 45178
rect 1104 45104 5980 45126
rect 1104 44634 5980 44656
rect 1104 44582 3802 44634
rect 3854 44582 3866 44634
rect 3918 44582 3930 44634
rect 3982 44582 3994 44634
rect 4046 44582 4058 44634
rect 4110 44582 5980 44634
rect 1104 44560 5980 44582
rect 5261 44523 5319 44529
rect 5261 44489 5273 44523
rect 5307 44520 5319 44523
rect 5445 44523 5503 44529
rect 5445 44520 5457 44523
rect 5307 44492 5457 44520
rect 5307 44489 5319 44492
rect 5261 44483 5319 44489
rect 5445 44489 5457 44492
rect 5491 44520 5503 44523
rect 6546 44520 6552 44532
rect 5491 44492 6552 44520
rect 5491 44489 5503 44492
rect 5445 44483 5503 44489
rect 6546 44480 6552 44492
rect 6604 44480 6610 44532
rect 1673 44387 1731 44393
rect 1673 44353 1685 44387
rect 1719 44384 1731 44387
rect 5077 44387 5135 44393
rect 1719 44356 2774 44384
rect 1719 44353 1731 44356
rect 1673 44347 1731 44353
rect 2746 44316 2774 44356
rect 5077 44353 5089 44387
rect 5123 44384 5135 44387
rect 5442 44384 5448 44396
rect 5123 44356 5448 44384
rect 5123 44353 5135 44356
rect 5077 44347 5135 44353
rect 5442 44344 5448 44356
rect 5500 44384 5506 44396
rect 5629 44387 5687 44393
rect 5629 44384 5641 44387
rect 5500 44356 5641 44384
rect 5500 44344 5506 44356
rect 5629 44353 5641 44356
rect 5675 44353 5687 44387
rect 5629 44347 5687 44353
rect 8294 44316 8300 44328
rect 2746 44288 8300 44316
rect 8294 44276 8300 44288
rect 8352 44276 8358 44328
rect 1486 44208 1492 44260
rect 1544 44208 1550 44260
rect 1104 44090 5980 44112
rect 1104 44038 3066 44090
rect 3118 44038 3130 44090
rect 3182 44038 3194 44090
rect 3246 44038 3258 44090
rect 3310 44038 3322 44090
rect 3374 44038 5980 44090
rect 1104 44016 5980 44038
rect 1765 43979 1823 43985
rect 1765 43945 1777 43979
rect 1811 43976 1823 43979
rect 6822 43976 6828 43988
rect 1811 43948 6828 43976
rect 1811 43945 1823 43948
rect 1765 43939 1823 43945
rect 6822 43936 6828 43948
rect 6880 43936 6886 43988
rect 1210 43664 1216 43716
rect 1268 43704 1274 43716
rect 1489 43707 1547 43713
rect 1489 43704 1501 43707
rect 1268 43676 1501 43704
rect 1268 43664 1274 43676
rect 1489 43673 1501 43676
rect 1535 43704 1547 43707
rect 1949 43707 2007 43713
rect 1949 43704 1961 43707
rect 1535 43676 1961 43704
rect 1535 43673 1547 43676
rect 1489 43667 1547 43673
rect 1949 43673 1961 43676
rect 1995 43673 2007 43707
rect 1949 43667 2007 43673
rect 1104 43546 5980 43568
rect 1104 43494 3802 43546
rect 3854 43494 3866 43546
rect 3918 43494 3930 43546
rect 3982 43494 3994 43546
rect 4046 43494 4058 43546
rect 4110 43494 5980 43546
rect 1104 43472 5980 43494
rect 5261 43435 5319 43441
rect 5261 43401 5273 43435
rect 5307 43432 5319 43435
rect 5445 43435 5503 43441
rect 5445 43432 5457 43435
rect 5307 43404 5457 43432
rect 5307 43401 5319 43404
rect 5261 43395 5319 43401
rect 5445 43401 5457 43404
rect 5491 43432 5503 43435
rect 7006 43432 7012 43444
rect 5491 43404 7012 43432
rect 5491 43401 5503 43404
rect 5445 43395 5503 43401
rect 7006 43392 7012 43404
rect 7064 43392 7070 43444
rect 8294 43364 8300 43376
rect 2746 43336 8300 43364
rect 1673 43299 1731 43305
rect 1673 43265 1685 43299
rect 1719 43296 1731 43299
rect 2746 43296 2774 43336
rect 8294 43324 8300 43336
rect 8352 43324 8358 43376
rect 1719 43268 2774 43296
rect 5077 43299 5135 43305
rect 1719 43265 1731 43268
rect 1673 43259 1731 43265
rect 5077 43265 5089 43299
rect 5123 43296 5135 43299
rect 5537 43299 5595 43305
rect 5537 43296 5549 43299
rect 5123 43268 5549 43296
rect 5123 43265 5135 43268
rect 5077 43259 5135 43265
rect 5537 43265 5549 43268
rect 5583 43296 5595 43299
rect 6914 43296 6920 43308
rect 5583 43268 6920 43296
rect 5583 43265 5595 43268
rect 5537 43259 5595 43265
rect 6914 43256 6920 43268
rect 6972 43256 6978 43308
rect 1486 43052 1492 43104
rect 1544 43052 1550 43104
rect 1104 43002 5980 43024
rect 1104 42950 3066 43002
rect 3118 42950 3130 43002
rect 3182 42950 3194 43002
rect 3246 42950 3258 43002
rect 3310 42950 3322 43002
rect 3374 42950 5980 43002
rect 1104 42928 5980 42950
rect 1104 42458 5980 42480
rect 1104 42406 3802 42458
rect 3854 42406 3866 42458
rect 3918 42406 3930 42458
rect 3982 42406 3994 42458
rect 4046 42406 4058 42458
rect 4110 42406 5980 42458
rect 1104 42384 5980 42406
rect 1104 41914 5980 41936
rect 1104 41862 3066 41914
rect 3118 41862 3130 41914
rect 3182 41862 3194 41914
rect 3246 41862 3258 41914
rect 3310 41862 3322 41914
rect 3374 41862 5980 41914
rect 1104 41840 5980 41862
rect 5074 41760 5080 41812
rect 5132 41760 5138 41812
rect 5261 41735 5319 41741
rect 5261 41701 5273 41735
rect 5307 41732 5319 41735
rect 5629 41735 5687 41741
rect 5629 41732 5641 41735
rect 5307 41704 5641 41732
rect 5307 41701 5319 41704
rect 5261 41695 5319 41701
rect 5629 41701 5641 41704
rect 5675 41732 5687 41735
rect 6454 41732 6460 41744
rect 5675 41704 6460 41732
rect 5675 41701 5687 41704
rect 5629 41695 5687 41701
rect 6454 41692 6460 41704
rect 6512 41692 6518 41744
rect 1673 41599 1731 41605
rect 1673 41565 1685 41599
rect 1719 41596 1731 41599
rect 8294 41596 8300 41608
rect 1719 41568 8300 41596
rect 1719 41565 1731 41568
rect 1673 41559 1731 41565
rect 8294 41556 8300 41568
rect 8352 41556 8358 41608
rect 5074 41488 5080 41540
rect 5132 41528 5138 41540
rect 5445 41531 5503 41537
rect 5445 41528 5457 41531
rect 5132 41500 5457 41528
rect 5132 41488 5138 41500
rect 5445 41497 5457 41500
rect 5491 41497 5503 41531
rect 5445 41491 5503 41497
rect 1486 41420 1492 41472
rect 1544 41420 1550 41472
rect 1104 41370 5980 41392
rect 1104 41318 3802 41370
rect 3854 41318 3866 41370
rect 3918 41318 3930 41370
rect 3982 41318 3994 41370
rect 4046 41318 4058 41370
rect 4110 41318 5980 41370
rect 1104 41296 5980 41318
rect 88794 41080 88800 41132
rect 88852 41080 88858 41132
rect 88812 40860 88840 41080
rect 1104 40826 5980 40848
rect 1104 40774 3066 40826
rect 3118 40774 3130 40826
rect 3182 40774 3194 40826
rect 3246 40774 3258 40826
rect 3310 40774 3322 40826
rect 3374 40774 5980 40826
rect 88794 40808 88800 40860
rect 88852 40808 88858 40860
rect 1104 40752 5980 40774
rect 4890 40672 4896 40724
rect 4948 40712 4954 40724
rect 4985 40715 5043 40721
rect 4985 40712 4997 40715
rect 4948 40684 4997 40712
rect 4948 40672 4954 40684
rect 4985 40681 4997 40684
rect 5031 40681 5043 40715
rect 4985 40675 5043 40681
rect 5261 40715 5319 40721
rect 5261 40681 5273 40715
rect 5307 40712 5319 40715
rect 5350 40712 5356 40724
rect 5307 40684 5356 40712
rect 5307 40681 5319 40684
rect 5261 40675 5319 40681
rect 5350 40672 5356 40684
rect 5408 40712 5414 40724
rect 5537 40715 5595 40721
rect 5537 40712 5549 40715
rect 5408 40684 5549 40712
rect 5408 40672 5414 40684
rect 5537 40681 5549 40684
rect 5583 40681 5595 40715
rect 5537 40675 5595 40681
rect 88886 40672 88892 40724
rect 88944 40712 88950 40724
rect 89162 40712 89168 40724
rect 88944 40684 89168 40712
rect 88944 40672 88950 40684
rect 89162 40672 89168 40684
rect 89220 40672 89226 40724
rect 89162 40536 89168 40588
rect 89220 40576 89226 40588
rect 89438 40576 89444 40588
rect 89220 40548 89444 40576
rect 89220 40536 89226 40548
rect 89438 40536 89444 40548
rect 89496 40536 89502 40588
rect 1673 40511 1731 40517
rect 1673 40477 1685 40511
rect 1719 40508 1731 40511
rect 8294 40508 8300 40520
rect 1719 40480 8300 40508
rect 1719 40477 1731 40480
rect 1673 40471 1731 40477
rect 8294 40468 8300 40480
rect 8352 40468 8358 40520
rect 4890 40400 4896 40452
rect 4948 40440 4954 40452
rect 5445 40443 5503 40449
rect 5445 40440 5457 40443
rect 4948 40412 5457 40440
rect 4948 40400 4954 40412
rect 5445 40409 5457 40412
rect 5491 40409 5503 40443
rect 5445 40403 5503 40409
rect 842 40332 848 40384
rect 900 40372 906 40384
rect 1489 40375 1547 40381
rect 1489 40372 1501 40375
rect 900 40344 1501 40372
rect 900 40332 906 40344
rect 1489 40341 1501 40344
rect 1535 40341 1547 40375
rect 1489 40335 1547 40341
rect 1104 40282 5980 40304
rect 1104 40230 3802 40282
rect 3854 40230 3866 40282
rect 3918 40230 3930 40282
rect 3982 40230 3994 40282
rect 4046 40230 4058 40282
rect 4110 40230 5980 40282
rect 1104 40208 5980 40230
rect 1104 39738 5980 39760
rect 1104 39686 3066 39738
rect 3118 39686 3130 39738
rect 3182 39686 3194 39738
rect 3246 39686 3258 39738
rect 3310 39686 3322 39738
rect 3374 39686 5980 39738
rect 1104 39664 5980 39686
rect 1104 39194 5980 39216
rect 1104 39142 3802 39194
rect 3854 39142 3866 39194
rect 3918 39142 3930 39194
rect 3982 39142 3994 39194
rect 4046 39142 4058 39194
rect 4110 39142 5980 39194
rect 1104 39120 5980 39142
rect 4982 39040 4988 39092
rect 5040 39080 5046 39092
rect 5261 39083 5319 39089
rect 5261 39080 5273 39083
rect 5040 39052 5273 39080
rect 5040 39040 5046 39052
rect 5261 39049 5273 39052
rect 5307 39080 5319 39083
rect 5445 39083 5503 39089
rect 5445 39080 5457 39083
rect 5307 39052 5457 39080
rect 5307 39049 5319 39052
rect 5261 39043 5319 39049
rect 5445 39049 5457 39052
rect 5491 39049 5503 39083
rect 5445 39043 5503 39049
rect 1673 38947 1731 38953
rect 1673 38913 1685 38947
rect 1719 38913 1731 38947
rect 1673 38907 1731 38913
rect 5169 38947 5227 38953
rect 5169 38913 5181 38947
rect 5215 38944 5227 38947
rect 5629 38947 5687 38953
rect 5629 38944 5641 38947
rect 5215 38916 5641 38944
rect 5215 38913 5227 38916
rect 5169 38907 5227 38913
rect 5629 38913 5641 38916
rect 5675 38944 5687 38947
rect 7834 38944 7840 38956
rect 5675 38916 7840 38944
rect 5675 38913 5687 38916
rect 5629 38907 5687 38913
rect 1688 38876 1716 38907
rect 7834 38904 7840 38916
rect 7892 38904 7898 38956
rect 8294 38876 8300 38888
rect 1688 38848 8300 38876
rect 8294 38836 8300 38848
rect 8352 38836 8358 38888
rect 842 38700 848 38752
rect 900 38740 906 38752
rect 1489 38743 1547 38749
rect 1489 38740 1501 38743
rect 900 38712 1501 38740
rect 900 38700 906 38712
rect 1489 38709 1501 38712
rect 1535 38709 1547 38743
rect 1489 38703 1547 38709
rect 1104 38650 5980 38672
rect 1104 38598 3066 38650
rect 3118 38598 3130 38650
rect 3182 38598 3194 38650
rect 3246 38598 3258 38650
rect 3310 38598 3322 38650
rect 3374 38598 5980 38650
rect 1104 38576 5980 38598
rect 1104 38106 5980 38128
rect 1104 38054 3802 38106
rect 3854 38054 3866 38106
rect 3918 38054 3930 38106
rect 3982 38054 3994 38106
rect 4046 38054 4058 38106
rect 4110 38054 5980 38106
rect 1104 38032 5980 38054
rect 5261 37995 5319 38001
rect 5261 37961 5273 37995
rect 5307 37992 5319 37995
rect 5445 37995 5503 38001
rect 5445 37992 5457 37995
rect 5307 37964 5457 37992
rect 5307 37961 5319 37964
rect 5261 37955 5319 37961
rect 5445 37961 5457 37964
rect 5491 37992 5503 37995
rect 6362 37992 6368 38004
rect 5491 37964 6368 37992
rect 5491 37961 5503 37964
rect 5445 37955 5503 37961
rect 6362 37952 6368 37964
rect 6420 37952 6426 38004
rect 8294 37924 8300 37936
rect 1688 37896 8300 37924
rect 1688 37865 1716 37896
rect 8294 37884 8300 37896
rect 8352 37884 8358 37936
rect 1673 37859 1731 37865
rect 1673 37825 1685 37859
rect 1719 37825 1731 37859
rect 1673 37819 1731 37825
rect 5077 37859 5135 37865
rect 5077 37825 5089 37859
rect 5123 37856 5135 37859
rect 5537 37859 5595 37865
rect 5537 37856 5549 37859
rect 5123 37828 5549 37856
rect 5123 37825 5135 37828
rect 5077 37819 5135 37825
rect 5537 37825 5549 37828
rect 5583 37856 5595 37859
rect 5718 37856 5724 37868
rect 5583 37828 5724 37856
rect 5583 37825 5595 37828
rect 5537 37819 5595 37825
rect 5718 37816 5724 37828
rect 5776 37816 5782 37868
rect 842 37612 848 37664
rect 900 37652 906 37664
rect 1489 37655 1547 37661
rect 1489 37652 1501 37655
rect 900 37624 1501 37652
rect 900 37612 906 37624
rect 1489 37621 1501 37624
rect 1535 37621 1547 37655
rect 1489 37615 1547 37621
rect 1104 37562 5980 37584
rect 1104 37510 3066 37562
rect 3118 37510 3130 37562
rect 3182 37510 3194 37562
rect 3246 37510 3258 37562
rect 3310 37510 3322 37562
rect 3374 37510 5980 37562
rect 1104 37488 5980 37510
rect 1104 37018 5980 37040
rect 1104 36966 3802 37018
rect 3854 36966 3866 37018
rect 3918 36966 3930 37018
rect 3982 36966 3994 37018
rect 4046 36966 4058 37018
rect 4110 36966 5980 37018
rect 1104 36944 5980 36966
rect 1104 36474 5980 36496
rect 1104 36422 3066 36474
rect 3118 36422 3130 36474
rect 3182 36422 3194 36474
rect 3246 36422 3258 36474
rect 3310 36422 3322 36474
rect 3374 36422 5980 36474
rect 1104 36400 5980 36422
rect 4614 36320 4620 36372
rect 4672 36360 4678 36372
rect 5261 36363 5319 36369
rect 5261 36360 5273 36363
rect 4672 36332 5273 36360
rect 4672 36320 4678 36332
rect 5261 36329 5273 36332
rect 5307 36360 5319 36363
rect 5629 36363 5687 36369
rect 5629 36360 5641 36363
rect 5307 36332 5641 36360
rect 5307 36329 5319 36332
rect 5261 36323 5319 36329
rect 5629 36329 5641 36332
rect 5675 36329 5687 36363
rect 5629 36323 5687 36329
rect 842 36252 848 36304
rect 900 36292 906 36304
rect 1489 36295 1547 36301
rect 1489 36292 1501 36295
rect 900 36264 1501 36292
rect 900 36252 906 36264
rect 1489 36261 1501 36264
rect 1535 36261 1547 36295
rect 1489 36255 1547 36261
rect 1673 36159 1731 36165
rect 1673 36125 1685 36159
rect 1719 36125 1731 36159
rect 1673 36119 1731 36125
rect 5169 36159 5227 36165
rect 5169 36125 5181 36159
rect 5215 36156 5227 36159
rect 5445 36159 5503 36165
rect 5445 36156 5457 36159
rect 5215 36128 5457 36156
rect 5215 36125 5227 36128
rect 5169 36119 5227 36125
rect 5445 36125 5457 36128
rect 5491 36156 5503 36159
rect 7558 36156 7564 36168
rect 5491 36128 7564 36156
rect 5491 36125 5503 36128
rect 5445 36119 5503 36125
rect 1688 36088 1716 36119
rect 7558 36116 7564 36128
rect 7616 36116 7622 36168
rect 8294 36088 8300 36100
rect 1688 36060 8300 36088
rect 8294 36048 8300 36060
rect 8352 36048 8358 36100
rect 1104 35930 5980 35952
rect 1104 35878 3802 35930
rect 3854 35878 3866 35930
rect 3918 35878 3930 35930
rect 3982 35878 3994 35930
rect 4046 35878 4058 35930
rect 4110 35878 5980 35930
rect 1104 35856 5980 35878
rect 1104 35386 5980 35408
rect 1104 35334 3066 35386
rect 3118 35334 3130 35386
rect 3182 35334 3194 35386
rect 3246 35334 3258 35386
rect 3310 35334 3322 35386
rect 3374 35334 5980 35386
rect 1104 35312 5980 35334
rect 8294 35136 8300 35148
rect 1688 35108 8300 35136
rect 1688 35077 1716 35108
rect 8294 35096 8300 35108
rect 8352 35096 8358 35148
rect 1673 35071 1731 35077
rect 1673 35037 1685 35071
rect 1719 35037 1731 35071
rect 1673 35031 1731 35037
rect 5169 35071 5227 35077
rect 5169 35037 5181 35071
rect 5215 35068 5227 35071
rect 5445 35071 5503 35077
rect 5445 35068 5457 35071
rect 5215 35040 5457 35068
rect 5215 35037 5227 35040
rect 5169 35031 5227 35037
rect 5445 35037 5457 35040
rect 5491 35068 5503 35071
rect 6270 35068 6276 35080
rect 5491 35040 6276 35068
rect 5491 35037 5503 35040
rect 5445 35031 5503 35037
rect 6270 35028 6276 35040
rect 6328 35028 6334 35080
rect 842 34892 848 34944
rect 900 34932 906 34944
rect 1489 34935 1547 34941
rect 1489 34932 1501 34935
rect 900 34904 1501 34932
rect 900 34892 906 34904
rect 1489 34901 1501 34904
rect 1535 34901 1547 34935
rect 1489 34895 1547 34901
rect 4982 34892 4988 34944
rect 5040 34932 5046 34944
rect 5261 34935 5319 34941
rect 5261 34932 5273 34935
rect 5040 34904 5273 34932
rect 5040 34892 5046 34904
rect 5261 34901 5273 34904
rect 5307 34932 5319 34935
rect 5629 34935 5687 34941
rect 5629 34932 5641 34935
rect 5307 34904 5641 34932
rect 5307 34901 5319 34904
rect 5261 34895 5319 34901
rect 5629 34901 5641 34904
rect 5675 34901 5687 34935
rect 5629 34895 5687 34901
rect 1104 34842 5980 34864
rect 1104 34790 3802 34842
rect 3854 34790 3866 34842
rect 3918 34790 3930 34842
rect 3982 34790 3994 34842
rect 4046 34790 4058 34842
rect 4110 34790 5980 34842
rect 1104 34768 5980 34790
rect 1104 34298 5980 34320
rect 1104 34246 3066 34298
rect 3118 34246 3130 34298
rect 3182 34246 3194 34298
rect 3246 34246 3258 34298
rect 3310 34246 3322 34298
rect 3374 34246 5980 34298
rect 1104 34224 5980 34246
rect 1104 33754 5980 33776
rect 1104 33702 3802 33754
rect 3854 33702 3866 33754
rect 3918 33702 3930 33754
rect 3982 33702 3994 33754
rect 4046 33702 4058 33754
rect 4110 33702 5980 33754
rect 1104 33680 5980 33702
rect 1673 33507 1731 33513
rect 1673 33473 1685 33507
rect 1719 33473 1731 33507
rect 1673 33467 1731 33473
rect 5169 33507 5227 33513
rect 5169 33473 5181 33507
rect 5215 33504 5227 33507
rect 5626 33504 5632 33516
rect 5215 33476 5632 33504
rect 5215 33473 5227 33476
rect 5169 33467 5227 33473
rect 1688 33436 1716 33467
rect 5626 33464 5632 33476
rect 5684 33464 5690 33516
rect 8294 33436 8300 33448
rect 1688 33408 8300 33436
rect 8294 33396 8300 33408
rect 8352 33396 8358 33448
rect 842 33260 848 33312
rect 900 33300 906 33312
rect 1489 33303 1547 33309
rect 1489 33300 1501 33303
rect 900 33272 1501 33300
rect 900 33260 906 33272
rect 1489 33269 1501 33272
rect 1535 33269 1547 33303
rect 1489 33263 1547 33269
rect 5353 33303 5411 33309
rect 5353 33269 5365 33303
rect 5399 33300 5411 33303
rect 5445 33303 5503 33309
rect 5445 33300 5457 33303
rect 5399 33272 5457 33300
rect 5399 33269 5411 33272
rect 5353 33263 5411 33269
rect 5445 33269 5457 33272
rect 5491 33300 5503 33303
rect 6178 33300 6184 33312
rect 5491 33272 6184 33300
rect 5491 33269 5503 33272
rect 5445 33263 5503 33269
rect 6178 33260 6184 33272
rect 6236 33260 6242 33312
rect 1104 33210 5980 33232
rect 1104 33158 3066 33210
rect 3118 33158 3130 33210
rect 3182 33158 3194 33210
rect 3246 33158 3258 33210
rect 3310 33158 3322 33210
rect 3374 33158 5980 33210
rect 1104 33136 5980 33158
rect 1104 32666 5980 32688
rect 1104 32614 3802 32666
rect 3854 32614 3866 32666
rect 3918 32614 3930 32666
rect 3982 32614 3994 32666
rect 4046 32614 4058 32666
rect 4110 32614 5980 32666
rect 1104 32592 5980 32614
rect 4798 32512 4804 32564
rect 4856 32552 4862 32564
rect 5077 32555 5135 32561
rect 5077 32552 5089 32555
rect 4856 32524 5089 32552
rect 4856 32512 4862 32524
rect 5077 32521 5089 32524
rect 5123 32521 5135 32555
rect 5077 32515 5135 32521
rect 8294 32484 8300 32496
rect 1688 32456 8300 32484
rect 1688 32425 1716 32456
rect 8294 32444 8300 32456
rect 8352 32444 8358 32496
rect 1673 32419 1731 32425
rect 1673 32385 1685 32419
rect 1719 32385 1731 32419
rect 1673 32379 1731 32385
rect 4798 32376 4804 32428
rect 4856 32416 4862 32428
rect 5629 32419 5687 32425
rect 5629 32416 5641 32419
rect 4856 32388 5641 32416
rect 4856 32376 4862 32388
rect 5629 32385 5641 32388
rect 5675 32385 5687 32419
rect 5629 32379 5687 32385
rect 842 32172 848 32224
rect 900 32212 906 32224
rect 1489 32215 1547 32221
rect 1489 32212 1501 32215
rect 900 32184 1501 32212
rect 900 32172 906 32184
rect 1489 32181 1501 32184
rect 1535 32181 1547 32215
rect 1489 32175 1547 32181
rect 5353 32215 5411 32221
rect 5353 32181 5365 32215
rect 5399 32212 5411 32215
rect 5445 32215 5503 32221
rect 5445 32212 5457 32215
rect 5399 32184 5457 32212
rect 5399 32181 5411 32184
rect 5353 32175 5411 32181
rect 5445 32181 5457 32184
rect 5491 32212 5503 32215
rect 6270 32212 6276 32224
rect 5491 32184 6276 32212
rect 5491 32181 5503 32184
rect 5445 32175 5503 32181
rect 6270 32172 6276 32184
rect 6328 32172 6334 32224
rect 1104 32122 5980 32144
rect 1104 32070 3066 32122
rect 3118 32070 3130 32122
rect 3182 32070 3194 32122
rect 3246 32070 3258 32122
rect 3310 32070 3322 32122
rect 3374 32070 5980 32122
rect 1104 32048 5980 32070
rect 1104 31578 5980 31600
rect 1104 31526 3802 31578
rect 3854 31526 3866 31578
rect 3918 31526 3930 31578
rect 3982 31526 3994 31578
rect 4046 31526 4058 31578
rect 4110 31526 5980 31578
rect 1104 31504 5980 31526
rect 1104 31034 5980 31056
rect 1104 30982 3066 31034
rect 3118 30982 3130 31034
rect 3182 30982 3194 31034
rect 3246 30982 3258 31034
rect 3310 30982 3322 31034
rect 3374 30982 5980 31034
rect 1104 30960 5980 30982
rect 4706 30880 4712 30932
rect 4764 30920 4770 30932
rect 5261 30923 5319 30929
rect 5261 30920 5273 30923
rect 4764 30892 5273 30920
rect 4764 30880 4770 30892
rect 5261 30889 5273 30892
rect 5307 30920 5319 30923
rect 5445 30923 5503 30929
rect 5445 30920 5457 30923
rect 5307 30892 5457 30920
rect 5307 30889 5319 30892
rect 5261 30883 5319 30889
rect 5445 30889 5457 30892
rect 5491 30889 5503 30923
rect 5445 30883 5503 30889
rect 842 30812 848 30864
rect 900 30852 906 30864
rect 1489 30855 1547 30861
rect 1489 30852 1501 30855
rect 900 30824 1501 30852
rect 900 30812 906 30824
rect 1489 30821 1501 30824
rect 1535 30821 1547 30855
rect 1489 30815 1547 30821
rect 1673 30719 1731 30725
rect 1673 30685 1685 30719
rect 1719 30685 1731 30719
rect 1673 30679 1731 30685
rect 5169 30719 5227 30725
rect 5169 30685 5181 30719
rect 5215 30716 5227 30719
rect 5626 30716 5632 30728
rect 5215 30688 5632 30716
rect 5215 30685 5227 30688
rect 5169 30679 5227 30685
rect 1688 30648 1716 30679
rect 5626 30676 5632 30688
rect 5684 30676 5690 30728
rect 8294 30648 8300 30660
rect 1688 30620 8300 30648
rect 8294 30608 8300 30620
rect 8352 30608 8358 30660
rect 1104 30490 5980 30512
rect 1104 30438 3802 30490
rect 3854 30438 3866 30490
rect 3918 30438 3930 30490
rect 3982 30438 3994 30490
rect 4046 30438 4058 30490
rect 4110 30438 5980 30490
rect 1104 30416 5980 30438
rect 1104 29946 5980 29968
rect 1104 29894 3066 29946
rect 3118 29894 3130 29946
rect 3182 29894 3194 29946
rect 3246 29894 3258 29946
rect 3310 29894 3322 29946
rect 3374 29894 5980 29946
rect 1104 29872 5980 29894
rect 8294 29696 8300 29708
rect 1688 29668 8300 29696
rect 1688 29637 1716 29668
rect 8294 29656 8300 29668
rect 8352 29656 8358 29708
rect 1673 29631 1731 29637
rect 1673 29597 1685 29631
rect 1719 29597 1731 29631
rect 1673 29591 1731 29597
rect 5169 29631 5227 29637
rect 5169 29597 5181 29631
rect 5215 29628 5227 29631
rect 5442 29628 5448 29640
rect 5215 29600 5448 29628
rect 5215 29597 5227 29600
rect 5169 29591 5227 29597
rect 5442 29588 5448 29600
rect 5500 29588 5506 29640
rect 842 29452 848 29504
rect 900 29492 906 29504
rect 1489 29495 1547 29501
rect 1489 29492 1501 29495
rect 900 29464 1501 29492
rect 900 29452 906 29464
rect 1489 29461 1501 29464
rect 1535 29461 1547 29495
rect 1489 29455 1547 29461
rect 5350 29452 5356 29504
rect 5408 29492 5414 29504
rect 5629 29495 5687 29501
rect 5629 29492 5641 29495
rect 5408 29464 5641 29492
rect 5408 29452 5414 29464
rect 5629 29461 5641 29464
rect 5675 29461 5687 29495
rect 5629 29455 5687 29461
rect 1104 29402 5980 29424
rect 1104 29350 3802 29402
rect 3854 29350 3866 29402
rect 3918 29350 3930 29402
rect 3982 29350 3994 29402
rect 4046 29350 4058 29402
rect 4110 29350 5980 29402
rect 1104 29328 5980 29350
rect 1104 28858 5980 28880
rect 1104 28806 3066 28858
rect 3118 28806 3130 28858
rect 3182 28806 3194 28858
rect 3246 28806 3258 28858
rect 3310 28806 3322 28858
rect 3374 28806 5980 28858
rect 1104 28784 5980 28806
rect 1104 28314 5980 28336
rect 1104 28262 3802 28314
rect 3854 28262 3866 28314
rect 3918 28262 3930 28314
rect 3982 28262 3994 28314
rect 4046 28262 4058 28314
rect 4110 28262 5980 28314
rect 1104 28240 5980 28262
rect 5074 28160 5080 28212
rect 5132 28160 5138 28212
rect 5258 28160 5264 28212
rect 5316 28200 5322 28212
rect 5445 28203 5503 28209
rect 5445 28200 5457 28203
rect 5316 28172 5457 28200
rect 5316 28160 5322 28172
rect 5445 28169 5457 28172
rect 5491 28169 5503 28203
rect 5445 28163 5503 28169
rect 1673 28067 1731 28073
rect 1673 28033 1685 28067
rect 1719 28033 1731 28067
rect 5092 28064 5120 28160
rect 5629 28067 5687 28073
rect 5629 28064 5641 28067
rect 5092 28036 5641 28064
rect 1673 28027 1731 28033
rect 5629 28033 5641 28036
rect 5675 28033 5687 28067
rect 5629 28027 5687 28033
rect 1688 27996 1716 28027
rect 8294 27996 8300 28008
rect 1688 27968 8300 27996
rect 8294 27956 8300 27968
rect 8352 27956 8358 28008
rect 842 27820 848 27872
rect 900 27860 906 27872
rect 1489 27863 1547 27869
rect 1489 27860 1501 27863
rect 900 27832 1501 27860
rect 900 27820 906 27832
rect 1489 27829 1501 27832
rect 1535 27829 1547 27863
rect 1489 27823 1547 27829
rect 1104 27770 5980 27792
rect 1104 27718 3066 27770
rect 3118 27718 3130 27770
rect 3182 27718 3194 27770
rect 3246 27718 3258 27770
rect 3310 27718 3322 27770
rect 3374 27718 5980 27770
rect 1104 27696 5980 27718
rect 1104 27226 5980 27248
rect 1104 27174 3802 27226
rect 3854 27174 3866 27226
rect 3918 27174 3930 27226
rect 3982 27174 3994 27226
rect 4046 27174 4058 27226
rect 4110 27174 5980 27226
rect 1104 27152 5980 27174
rect 1581 27115 1639 27121
rect 1581 27081 1593 27115
rect 1627 27112 1639 27115
rect 8294 27112 8300 27124
rect 1627 27084 8300 27112
rect 1627 27081 1639 27084
rect 1581 27075 1639 27081
rect 8294 27072 8300 27084
rect 8352 27072 8358 27124
rect 5258 27004 5264 27056
rect 5316 27004 5322 27056
rect 1302 26936 1308 26988
rect 1360 26976 1366 26988
rect 1397 26979 1455 26985
rect 1397 26976 1409 26979
rect 1360 26948 1409 26976
rect 1360 26936 1366 26948
rect 1397 26945 1409 26948
rect 1443 26976 1455 26979
rect 1673 26979 1731 26985
rect 1673 26976 1685 26979
rect 1443 26948 1685 26976
rect 1443 26945 1455 26948
rect 1397 26939 1455 26945
rect 1673 26945 1685 26948
rect 1719 26945 1731 26979
rect 5276 26976 5304 27004
rect 5353 26979 5411 26985
rect 5353 26976 5365 26979
rect 5276 26948 5365 26976
rect 1673 26939 1731 26945
rect 5353 26945 5365 26948
rect 5399 26945 5411 26979
rect 5353 26939 5411 26945
rect 5534 26732 5540 26784
rect 5592 26732 5598 26784
rect 1104 26682 5980 26704
rect 1104 26630 3066 26682
rect 3118 26630 3130 26682
rect 3182 26630 3194 26682
rect 3246 26630 3258 26682
rect 3310 26630 3322 26682
rect 3374 26630 5980 26682
rect 1104 26608 5980 26630
rect 1104 26138 5980 26160
rect 1104 26086 3802 26138
rect 3854 26086 3866 26138
rect 3918 26086 3930 26138
rect 3982 26086 3994 26138
rect 4046 26086 4058 26138
rect 4110 26086 5980 26138
rect 1104 26064 5980 26086
rect 1104 25594 5980 25616
rect 1104 25542 3066 25594
rect 3118 25542 3130 25594
rect 3182 25542 3194 25594
rect 3246 25542 3258 25594
rect 3310 25542 3322 25594
rect 3374 25542 5980 25594
rect 1104 25520 5980 25542
rect 5537 25483 5595 25489
rect 5537 25449 5549 25483
rect 5583 25480 5595 25483
rect 5810 25480 5816 25492
rect 5583 25452 5816 25480
rect 5583 25449 5595 25452
rect 5537 25443 5595 25449
rect 5810 25440 5816 25452
rect 5868 25440 5874 25492
rect 1581 25415 1639 25421
rect 1581 25381 1593 25415
rect 1627 25412 1639 25415
rect 8294 25412 8300 25424
rect 1627 25384 8300 25412
rect 1627 25381 1639 25384
rect 1581 25375 1639 25381
rect 8294 25372 8300 25384
rect 8352 25372 8358 25424
rect 1210 25236 1216 25288
rect 1268 25276 1274 25288
rect 1397 25279 1455 25285
rect 1397 25276 1409 25279
rect 1268 25248 1409 25276
rect 1268 25236 1274 25248
rect 1397 25245 1409 25248
rect 1443 25276 1455 25279
rect 1673 25279 1731 25285
rect 1673 25276 1685 25279
rect 1443 25248 1685 25276
rect 1443 25245 1455 25248
rect 1397 25239 1455 25245
rect 1673 25245 1685 25248
rect 1719 25245 1731 25279
rect 1673 25239 1731 25245
rect 5353 25279 5411 25285
rect 5353 25245 5365 25279
rect 5399 25245 5411 25279
rect 5353 25239 5411 25245
rect 5261 25143 5319 25149
rect 5261 25109 5273 25143
rect 5307 25140 5319 25143
rect 5368 25140 5396 25239
rect 6362 25140 6368 25152
rect 5307 25112 6368 25140
rect 5307 25109 5319 25112
rect 5261 25103 5319 25109
rect 6362 25100 6368 25112
rect 6420 25100 6426 25152
rect 1104 25050 5980 25072
rect 1104 24998 3802 25050
rect 3854 24998 3866 25050
rect 3918 24998 3930 25050
rect 3982 24998 3994 25050
rect 4046 24998 4058 25050
rect 4110 24998 5980 25050
rect 1104 24976 5980 24998
rect 1104 24506 5980 24528
rect 1104 24454 3066 24506
rect 3118 24454 3130 24506
rect 3182 24454 3194 24506
rect 3246 24454 3258 24506
rect 3310 24454 3322 24506
rect 3374 24454 5980 24506
rect 1104 24432 5980 24454
rect 1581 24327 1639 24333
rect 1581 24293 1593 24327
rect 1627 24324 1639 24327
rect 8294 24324 8300 24336
rect 1627 24296 8300 24324
rect 1627 24293 1639 24296
rect 1581 24287 1639 24293
rect 8294 24284 8300 24296
rect 8352 24284 8358 24336
rect 1302 24148 1308 24200
rect 1360 24188 1366 24200
rect 1397 24191 1455 24197
rect 1397 24188 1409 24191
rect 1360 24160 1409 24188
rect 1360 24148 1366 24160
rect 1397 24157 1409 24160
rect 1443 24188 1455 24191
rect 1673 24191 1731 24197
rect 1673 24188 1685 24191
rect 1443 24160 1685 24188
rect 1443 24157 1455 24160
rect 1397 24151 1455 24157
rect 1673 24157 1685 24160
rect 1719 24157 1731 24191
rect 1673 24151 1731 24157
rect 1104 23962 5980 23984
rect 1104 23910 3802 23962
rect 3854 23910 3866 23962
rect 3918 23910 3930 23962
rect 3982 23910 3994 23962
rect 4046 23910 4058 23962
rect 4110 23910 5980 23962
rect 1104 23888 5980 23910
rect 1104 23418 5980 23440
rect 1104 23366 3066 23418
rect 3118 23366 3130 23418
rect 3182 23366 3194 23418
rect 3246 23366 3258 23418
rect 3310 23366 3322 23418
rect 3374 23366 5980 23418
rect 1104 23344 5980 23366
rect 1104 22874 5980 22896
rect 1104 22822 3802 22874
rect 3854 22822 3866 22874
rect 3918 22822 3930 22874
rect 3982 22822 3994 22874
rect 4046 22822 4058 22874
rect 4110 22822 5980 22874
rect 1104 22800 5980 22822
rect 1302 22584 1308 22636
rect 1360 22624 1366 22636
rect 1397 22627 1455 22633
rect 1397 22624 1409 22627
rect 1360 22596 1409 22624
rect 1360 22584 1366 22596
rect 1397 22593 1409 22596
rect 1443 22624 1455 22627
rect 1673 22627 1731 22633
rect 1673 22624 1685 22627
rect 1443 22596 1685 22624
rect 1443 22593 1455 22596
rect 1397 22587 1455 22593
rect 1673 22593 1685 22596
rect 1719 22593 1731 22627
rect 1673 22587 1731 22593
rect 1581 22491 1639 22497
rect 1581 22457 1593 22491
rect 1627 22488 1639 22491
rect 8294 22488 8300 22500
rect 1627 22460 8300 22488
rect 1627 22457 1639 22460
rect 1581 22451 1639 22457
rect 8294 22448 8300 22460
rect 8352 22448 8358 22500
rect 1104 22330 5980 22352
rect 1104 22278 3066 22330
rect 3118 22278 3130 22330
rect 3182 22278 3194 22330
rect 3246 22278 3258 22330
rect 3310 22278 3322 22330
rect 3374 22278 5980 22330
rect 1104 22256 5980 22278
rect 1104 21786 5980 21808
rect 1104 21734 3802 21786
rect 3854 21734 3866 21786
rect 3918 21734 3930 21786
rect 3982 21734 3994 21786
rect 4046 21734 4058 21786
rect 4110 21734 5980 21786
rect 1104 21712 5980 21734
rect 1581 21675 1639 21681
rect 1581 21641 1593 21675
rect 1627 21672 1639 21675
rect 8294 21672 8300 21684
rect 1627 21644 8300 21672
rect 1627 21641 1639 21644
rect 1581 21635 1639 21641
rect 8294 21632 8300 21644
rect 8352 21632 8358 21684
rect 1302 21496 1308 21548
rect 1360 21536 1366 21548
rect 1397 21539 1455 21545
rect 1397 21536 1409 21539
rect 1360 21508 1409 21536
rect 1360 21496 1366 21508
rect 1397 21505 1409 21508
rect 1443 21536 1455 21539
rect 1673 21539 1731 21545
rect 1673 21536 1685 21539
rect 1443 21508 1685 21536
rect 1443 21505 1455 21508
rect 1397 21499 1455 21505
rect 1673 21505 1685 21508
rect 1719 21505 1731 21539
rect 1673 21499 1731 21505
rect 1104 21242 5980 21264
rect 1104 21190 3066 21242
rect 3118 21190 3130 21242
rect 3182 21190 3194 21242
rect 3246 21190 3258 21242
rect 3310 21190 3322 21242
rect 3374 21190 5980 21242
rect 1104 21168 5980 21190
rect 1104 20698 5980 20720
rect 1104 20646 3802 20698
rect 3854 20646 3866 20698
rect 3918 20646 3930 20698
rect 3982 20646 3994 20698
rect 4046 20646 4058 20698
rect 4110 20646 5980 20698
rect 1104 20624 5980 20646
rect 1104 20154 5980 20176
rect 1104 20102 3066 20154
rect 3118 20102 3130 20154
rect 3182 20102 3194 20154
rect 3246 20102 3258 20154
rect 3310 20102 3322 20154
rect 3374 20102 5980 20154
rect 1104 20080 5980 20102
rect 1581 20043 1639 20049
rect 1581 20009 1593 20043
rect 1627 20040 1639 20043
rect 8294 20040 8300 20052
rect 1627 20012 8300 20040
rect 1627 20009 1639 20012
rect 1581 20003 1639 20009
rect 8294 20000 8300 20012
rect 8352 20000 8358 20052
rect 1210 19796 1216 19848
rect 1268 19836 1274 19848
rect 1397 19839 1455 19845
rect 1397 19836 1409 19839
rect 1268 19808 1409 19836
rect 1268 19796 1274 19808
rect 1397 19805 1409 19808
rect 1443 19836 1455 19839
rect 1673 19839 1731 19845
rect 1673 19836 1685 19839
rect 1443 19808 1685 19836
rect 1443 19805 1455 19808
rect 1397 19799 1455 19805
rect 1673 19805 1685 19808
rect 1719 19805 1731 19839
rect 1673 19799 1731 19805
rect 1104 19610 5980 19632
rect 1104 19558 3802 19610
rect 3854 19558 3866 19610
rect 3918 19558 3930 19610
rect 3982 19558 3994 19610
rect 4046 19558 4058 19610
rect 4110 19558 5980 19610
rect 1104 19536 5980 19558
rect 1104 19066 5980 19088
rect 1104 19014 3066 19066
rect 3118 19014 3130 19066
rect 3182 19014 3194 19066
rect 3246 19014 3258 19066
rect 3310 19014 3322 19066
rect 3374 19014 5980 19066
rect 1104 18992 5980 19014
rect 1581 18887 1639 18893
rect 1581 18853 1593 18887
rect 1627 18884 1639 18887
rect 8294 18884 8300 18896
rect 1627 18856 8300 18884
rect 1627 18853 1639 18856
rect 1581 18847 1639 18853
rect 8294 18844 8300 18856
rect 8352 18844 8358 18896
rect 1302 18708 1308 18760
rect 1360 18748 1366 18760
rect 1397 18751 1455 18757
rect 1397 18748 1409 18751
rect 1360 18720 1409 18748
rect 1360 18708 1366 18720
rect 1397 18717 1409 18720
rect 1443 18748 1455 18751
rect 1673 18751 1731 18757
rect 1673 18748 1685 18751
rect 1443 18720 1685 18748
rect 1443 18717 1455 18720
rect 1397 18711 1455 18717
rect 1673 18717 1685 18720
rect 1719 18717 1731 18751
rect 1673 18711 1731 18717
rect 1104 18522 5980 18544
rect 1104 18470 3802 18522
rect 3854 18470 3866 18522
rect 3918 18470 3930 18522
rect 3982 18470 3994 18522
rect 4046 18470 4058 18522
rect 4110 18470 5980 18522
rect 1104 18448 5980 18470
rect 1104 17978 5980 18000
rect 1104 17926 3066 17978
rect 3118 17926 3130 17978
rect 3182 17926 3194 17978
rect 3246 17926 3258 17978
rect 3310 17926 3322 17978
rect 3374 17926 5980 17978
rect 1104 17904 5980 17926
rect 1104 17434 5980 17456
rect 1104 17382 3802 17434
rect 3854 17382 3866 17434
rect 3918 17382 3930 17434
rect 3982 17382 3994 17434
rect 4046 17382 4058 17434
rect 4110 17382 5980 17434
rect 1104 17360 5980 17382
rect 1302 17144 1308 17196
rect 1360 17184 1366 17196
rect 1397 17187 1455 17193
rect 1397 17184 1409 17187
rect 1360 17156 1409 17184
rect 1360 17144 1366 17156
rect 1397 17153 1409 17156
rect 1443 17184 1455 17187
rect 1673 17187 1731 17193
rect 1673 17184 1685 17187
rect 1443 17156 1685 17184
rect 1443 17153 1455 17156
rect 1397 17147 1455 17153
rect 1673 17153 1685 17156
rect 1719 17153 1731 17187
rect 1673 17147 1731 17153
rect 1581 17051 1639 17057
rect 1581 17017 1593 17051
rect 1627 17048 1639 17051
rect 8294 17048 8300 17060
rect 1627 17020 8300 17048
rect 1627 17017 1639 17020
rect 1581 17011 1639 17017
rect 8294 17008 8300 17020
rect 8352 17008 8358 17060
rect 1104 16890 5980 16912
rect 1104 16838 3066 16890
rect 3118 16838 3130 16890
rect 3182 16838 3194 16890
rect 3246 16838 3258 16890
rect 3310 16838 3322 16890
rect 3374 16838 5980 16890
rect 1104 16816 5980 16838
rect 1104 16346 5980 16368
rect 1104 16294 3802 16346
rect 3854 16294 3866 16346
rect 3918 16294 3930 16346
rect 3982 16294 3994 16346
rect 4046 16294 4058 16346
rect 4110 16294 5980 16346
rect 1104 16272 5980 16294
rect 1581 16235 1639 16241
rect 1581 16201 1593 16235
rect 1627 16232 1639 16235
rect 8294 16232 8300 16244
rect 1627 16204 8300 16232
rect 1627 16201 1639 16204
rect 1581 16195 1639 16201
rect 8294 16192 8300 16204
rect 8352 16192 8358 16244
rect 1302 16056 1308 16108
rect 1360 16096 1366 16108
rect 1397 16099 1455 16105
rect 1397 16096 1409 16099
rect 1360 16068 1409 16096
rect 1360 16056 1366 16068
rect 1397 16065 1409 16068
rect 1443 16096 1455 16099
rect 1673 16099 1731 16105
rect 1673 16096 1685 16099
rect 1443 16068 1685 16096
rect 1443 16065 1455 16068
rect 1397 16059 1455 16065
rect 1673 16065 1685 16068
rect 1719 16065 1731 16099
rect 1673 16059 1731 16065
rect 1104 15802 5980 15824
rect 1104 15750 3066 15802
rect 3118 15750 3130 15802
rect 3182 15750 3194 15802
rect 3246 15750 3258 15802
rect 3310 15750 3322 15802
rect 3374 15750 5980 15802
rect 1104 15728 5980 15750
rect 1104 15258 5980 15280
rect 1104 15206 3802 15258
rect 3854 15206 3866 15258
rect 3918 15206 3930 15258
rect 3982 15206 3994 15258
rect 4046 15206 4058 15258
rect 4110 15206 5980 15258
rect 1104 15184 5980 15206
rect 1104 14714 5980 14736
rect 1104 14662 3066 14714
rect 3118 14662 3130 14714
rect 3182 14662 3194 14714
rect 3246 14662 3258 14714
rect 3310 14662 3322 14714
rect 3374 14662 5980 14714
rect 1104 14640 5980 14662
rect 1581 14603 1639 14609
rect 1581 14569 1593 14603
rect 1627 14600 1639 14603
rect 8294 14600 8300 14612
rect 1627 14572 8300 14600
rect 1627 14569 1639 14572
rect 1581 14563 1639 14569
rect 8294 14560 8300 14572
rect 8352 14560 8358 14612
rect 1210 14356 1216 14408
rect 1268 14396 1274 14408
rect 1397 14399 1455 14405
rect 1397 14396 1409 14399
rect 1268 14368 1409 14396
rect 1268 14356 1274 14368
rect 1397 14365 1409 14368
rect 1443 14396 1455 14399
rect 1673 14399 1731 14405
rect 1673 14396 1685 14399
rect 1443 14368 1685 14396
rect 1443 14365 1455 14368
rect 1397 14359 1455 14365
rect 1673 14365 1685 14368
rect 1719 14365 1731 14399
rect 1673 14359 1731 14365
rect 1104 14170 5980 14192
rect 1104 14118 3802 14170
rect 3854 14118 3866 14170
rect 3918 14118 3930 14170
rect 3982 14118 3994 14170
rect 4046 14118 4058 14170
rect 4110 14118 5980 14170
rect 1104 14096 5980 14118
rect 1104 13626 5980 13648
rect 1104 13574 3066 13626
rect 3118 13574 3130 13626
rect 3182 13574 3194 13626
rect 3246 13574 3258 13626
rect 3310 13574 3322 13626
rect 3374 13574 5980 13626
rect 1104 13552 5980 13574
rect 1581 13447 1639 13453
rect 1581 13413 1593 13447
rect 1627 13444 1639 13447
rect 8294 13444 8300 13456
rect 1627 13416 8300 13444
rect 1627 13413 1639 13416
rect 1581 13407 1639 13413
rect 8294 13404 8300 13416
rect 8352 13404 8358 13456
rect 1302 13268 1308 13320
rect 1360 13308 1366 13320
rect 1397 13311 1455 13317
rect 1397 13308 1409 13311
rect 1360 13280 1409 13308
rect 1360 13268 1366 13280
rect 1397 13277 1409 13280
rect 1443 13308 1455 13311
rect 1673 13311 1731 13317
rect 1673 13308 1685 13311
rect 1443 13280 1685 13308
rect 1443 13277 1455 13280
rect 1397 13271 1455 13277
rect 1673 13277 1685 13280
rect 1719 13277 1731 13311
rect 1673 13271 1731 13277
rect 1104 13082 5980 13104
rect 1104 13030 3802 13082
rect 3854 13030 3866 13082
rect 3918 13030 3930 13082
rect 3982 13030 3994 13082
rect 4046 13030 4058 13082
rect 4110 13030 5980 13082
rect 1104 13008 5980 13030
rect 1104 12538 5980 12560
rect 1104 12486 3066 12538
rect 3118 12486 3130 12538
rect 3182 12486 3194 12538
rect 3246 12486 3258 12538
rect 3310 12486 3322 12538
rect 3374 12486 5980 12538
rect 1104 12464 5980 12486
rect 1104 11994 5980 12016
rect 1104 11942 3802 11994
rect 3854 11942 3866 11994
rect 3918 11942 3930 11994
rect 3982 11942 3994 11994
rect 4046 11942 4058 11994
rect 4110 11942 5980 11994
rect 1104 11920 5980 11942
rect 1302 11704 1308 11756
rect 1360 11744 1366 11756
rect 1397 11747 1455 11753
rect 1397 11744 1409 11747
rect 1360 11716 1409 11744
rect 1360 11704 1366 11716
rect 1397 11713 1409 11716
rect 1443 11744 1455 11747
rect 1673 11747 1731 11753
rect 1673 11744 1685 11747
rect 1443 11716 1685 11744
rect 1443 11713 1455 11716
rect 1397 11707 1455 11713
rect 1673 11713 1685 11716
rect 1719 11713 1731 11747
rect 1673 11707 1731 11713
rect 1581 11611 1639 11617
rect 1581 11577 1593 11611
rect 1627 11608 1639 11611
rect 8294 11608 8300 11620
rect 1627 11580 8300 11608
rect 1627 11577 1639 11580
rect 1581 11571 1639 11577
rect 8294 11568 8300 11580
rect 8352 11568 8358 11620
rect 1104 11450 5980 11472
rect 1104 11398 3066 11450
rect 3118 11398 3130 11450
rect 3182 11398 3194 11450
rect 3246 11398 3258 11450
rect 3310 11398 3322 11450
rect 3374 11398 5980 11450
rect 1104 11376 5980 11398
rect 1104 10906 5980 10928
rect 1104 10854 3802 10906
rect 3854 10854 3866 10906
rect 3918 10854 3930 10906
rect 3982 10854 3994 10906
rect 4046 10854 4058 10906
rect 4110 10854 5980 10906
rect 1104 10832 5980 10854
rect 1104 10362 5980 10384
rect 1104 10310 3066 10362
rect 3118 10310 3130 10362
rect 3182 10310 3194 10362
rect 3246 10310 3258 10362
rect 3310 10310 3322 10362
rect 3374 10310 5980 10362
rect 1104 10288 5980 10310
rect 1104 9818 5980 9840
rect 1104 9766 3802 9818
rect 3854 9766 3866 9818
rect 3918 9766 3930 9818
rect 3982 9766 3994 9818
rect 4046 9766 4058 9818
rect 4110 9766 5980 9818
rect 1104 9744 5980 9766
rect 46750 9596 46756 9648
rect 46808 9636 46814 9648
rect 48682 9636 48688 9648
rect 46808 9608 48688 9636
rect 46808 9596 46814 9608
rect 48682 9596 48688 9608
rect 48740 9596 48746 9648
rect 86862 9460 86868 9512
rect 86920 9500 86926 9512
rect 88150 9500 88156 9512
rect 86920 9472 88156 9500
rect 86920 9460 86926 9472
rect 88150 9460 88156 9472
rect 88208 9460 88214 9512
rect 1104 9274 5980 9296
rect 1104 9222 3066 9274
rect 3118 9222 3130 9274
rect 3182 9222 3194 9274
rect 3246 9222 3258 9274
rect 3310 9222 3322 9274
rect 3374 9222 5980 9274
rect 1104 9200 5980 9222
rect 88058 8780 88064 8832
rect 88116 8820 88122 8832
rect 89162 8820 89168 8832
rect 88116 8792 89168 8820
rect 88116 8780 88122 8792
rect 89162 8780 89168 8792
rect 89220 8780 89226 8832
rect 1104 8730 5980 8752
rect 1104 8678 3802 8730
rect 3854 8678 3866 8730
rect 3918 8678 3930 8730
rect 3982 8678 3994 8730
rect 4046 8678 4058 8730
rect 4110 8678 5980 8730
rect 1104 8656 5980 8678
rect 47578 8576 47584 8628
rect 47636 8616 47642 8628
rect 49326 8616 49332 8628
rect 47636 8588 49332 8616
rect 47636 8576 47642 8588
rect 49326 8576 49332 8588
rect 49384 8576 49390 8628
rect 5350 8236 5356 8288
rect 5408 8276 5414 8288
rect 5408 8248 84194 8276
rect 5408 8236 5414 8248
rect 1104 8186 5980 8208
rect 1104 8134 3066 8186
rect 3118 8134 3130 8186
rect 3182 8134 3194 8186
rect 3246 8134 3258 8186
rect 3310 8134 3322 8186
rect 3374 8134 5980 8186
rect 8202 8168 8208 8220
rect 8260 8208 8266 8220
rect 12710 8208 12716 8220
rect 8260 8180 12716 8208
rect 8260 8168 8266 8180
rect 12710 8168 12716 8180
rect 12768 8168 12774 8220
rect 48682 8168 48688 8220
rect 48740 8208 48746 8220
rect 53834 8208 53840 8220
rect 48740 8180 53840 8208
rect 48740 8168 48746 8180
rect 53834 8168 53840 8180
rect 53892 8168 53898 8220
rect 84166 8208 84194 8248
rect 84746 8236 84752 8288
rect 84804 8276 84810 8288
rect 87230 8276 87236 8288
rect 84804 8248 87236 8276
rect 84804 8236 84810 8248
rect 87230 8236 87236 8248
rect 87288 8236 87294 8288
rect 86034 8208 86040 8220
rect 84166 8180 86040 8208
rect 86034 8168 86040 8180
rect 86092 8168 86098 8220
rect 1104 8112 5980 8134
rect 6822 8100 6828 8152
rect 6880 8140 6886 8152
rect 6880 8100 6914 8140
rect 8018 8100 8024 8152
rect 8076 8140 8082 8152
rect 10502 8140 10508 8152
rect 8076 8112 10508 8140
rect 8076 8100 8082 8112
rect 10502 8100 10508 8112
rect 10560 8100 10566 8152
rect 6886 8072 6914 8100
rect 11606 8072 11612 8084
rect 6886 8044 11612 8072
rect 11606 8032 11612 8044
rect 11664 8032 11670 8084
rect 5442 7964 5448 8016
rect 5500 8004 5506 8016
rect 47394 8004 47400 8016
rect 5500 7976 47400 8004
rect 5500 7964 5506 7976
rect 47394 7964 47400 7976
rect 47452 7964 47458 8016
rect 5534 7896 5540 7948
rect 5592 7936 5598 7948
rect 47670 7936 47676 7948
rect 5592 7908 47676 7936
rect 5592 7896 5598 7908
rect 47670 7896 47676 7908
rect 47728 7896 47734 7948
rect 4982 7828 4988 7880
rect 5040 7868 5046 7880
rect 47946 7868 47952 7880
rect 5040 7840 47952 7868
rect 5040 7828 5046 7840
rect 47946 7828 47952 7840
rect 48004 7868 48010 7880
rect 48004 7840 55214 7868
rect 48004 7828 48010 7840
rect 5626 7760 5632 7812
rect 5684 7800 5690 7812
rect 47486 7800 47492 7812
rect 5684 7772 47492 7800
rect 5684 7760 5690 7772
rect 47486 7760 47492 7772
rect 47544 7760 47550 7812
rect 55186 7800 55214 7840
rect 85298 7800 85304 7812
rect 55186 7772 85304 7800
rect 85298 7760 85304 7772
rect 85356 7760 85362 7812
rect 6362 7692 6368 7744
rect 6420 7732 6426 7744
rect 84746 7732 84752 7744
rect 6420 7704 84752 7732
rect 6420 7692 6426 7704
rect 84746 7692 84752 7704
rect 84804 7692 84810 7744
rect 1104 7642 5980 7664
rect 1104 7590 3802 7642
rect 3854 7590 3866 7642
rect 3918 7590 3930 7642
rect 3982 7590 3994 7642
rect 4046 7590 4058 7642
rect 4110 7590 5980 7642
rect 6178 7624 6184 7676
rect 6236 7664 6242 7676
rect 85666 7664 85672 7676
rect 6236 7636 85672 7664
rect 6236 7624 6242 7636
rect 85666 7624 85672 7636
rect 85724 7624 85730 7676
rect 1104 7568 5980 7590
rect 6270 7556 6276 7608
rect 6328 7596 6334 7608
rect 85758 7596 85764 7608
rect 6328 7568 85764 7596
rect 6328 7556 6334 7568
rect 85758 7556 85764 7568
rect 85816 7556 85822 7608
rect 1104 7098 5980 7120
rect 1104 7046 3066 7098
rect 3118 7046 3130 7098
rect 3182 7046 3194 7098
rect 3246 7046 3258 7098
rect 3310 7046 3322 7098
rect 3374 7046 5980 7098
rect 1104 7024 5980 7046
rect 1104 6554 5980 6576
rect 1104 6502 3802 6554
rect 3854 6502 3866 6554
rect 3918 6502 3930 6554
rect 3982 6502 3994 6554
rect 4046 6502 4058 6554
rect 4110 6502 5980 6554
rect 1104 6480 5980 6502
rect 48222 6196 48228 6248
rect 48280 6236 48286 6248
rect 50246 6236 50252 6248
rect 48280 6208 50252 6236
rect 48280 6196 48286 6208
rect 50246 6196 50252 6208
rect 50304 6196 50310 6248
rect 10870 6128 10876 6180
rect 10928 6168 10934 6180
rect 50798 6168 50804 6180
rect 10928 6140 50804 6168
rect 10928 6128 10934 6140
rect 50798 6128 50804 6140
rect 50856 6128 50862 6180
rect 1104 6010 88872 6032
rect 1104 5958 3066 6010
rect 3118 5958 3130 6010
rect 3182 5958 3194 6010
rect 3246 5958 3258 6010
rect 3310 5958 3322 6010
rect 3374 5958 72950 6010
rect 73002 5958 73014 6010
rect 73066 5958 73078 6010
rect 73130 5958 73142 6010
rect 73194 5958 73206 6010
rect 73258 5958 88872 6010
rect 1104 5936 88872 5958
rect 10870 5856 10876 5908
rect 10928 5856 10934 5908
rect 12986 5856 12992 5908
rect 13044 5896 13050 5908
rect 15102 5896 15108 5908
rect 13044 5868 15108 5896
rect 13044 5856 13050 5868
rect 15102 5856 15108 5868
rect 15160 5896 15166 5908
rect 15160 5868 16574 5896
rect 15160 5856 15166 5868
rect 16546 5760 16574 5868
rect 49694 5856 49700 5908
rect 49752 5856 49758 5908
rect 50246 5856 50252 5908
rect 50304 5856 50310 5908
rect 50798 5856 50804 5908
rect 50856 5856 50862 5908
rect 50908 5868 51074 5896
rect 46934 5788 46940 5840
rect 46992 5828 46998 5840
rect 47854 5828 47860 5840
rect 46992 5800 47860 5828
rect 46992 5788 46998 5800
rect 47854 5788 47860 5800
rect 47912 5828 47918 5840
rect 50908 5828 50936 5868
rect 47912 5800 50936 5828
rect 51046 5828 51074 5868
rect 84746 5856 84752 5908
rect 84804 5856 84810 5908
rect 85022 5856 85028 5908
rect 85080 5896 85086 5908
rect 85080 5868 85252 5896
rect 85080 5856 85086 5868
rect 53561 5831 53619 5837
rect 53561 5828 53573 5831
rect 51046 5800 53573 5828
rect 47912 5788 47918 5800
rect 53561 5797 53573 5800
rect 53607 5797 53619 5831
rect 53561 5791 53619 5797
rect 85114 5788 85120 5840
rect 85172 5788 85178 5840
rect 85224 5828 85252 5868
rect 85298 5856 85304 5908
rect 85356 5856 85362 5908
rect 86310 5856 86316 5908
rect 86368 5856 86374 5908
rect 86586 5856 86592 5908
rect 86644 5856 86650 5908
rect 88058 5856 88064 5908
rect 88116 5856 88122 5908
rect 88429 5899 88487 5905
rect 88429 5865 88441 5899
rect 88475 5896 88487 5899
rect 88518 5896 88524 5908
rect 88475 5868 88524 5896
rect 88475 5865 88487 5868
rect 88429 5859 88487 5865
rect 88518 5856 88524 5868
rect 88576 5856 88582 5908
rect 85853 5831 85911 5837
rect 85853 5828 85865 5831
rect 85224 5800 85865 5828
rect 85853 5797 85865 5800
rect 85899 5797 85911 5831
rect 85853 5791 85911 5797
rect 86957 5831 87015 5837
rect 86957 5797 86969 5831
rect 87003 5797 87015 5831
rect 86957 5791 87015 5797
rect 87693 5831 87751 5837
rect 87693 5797 87705 5831
rect 87739 5828 87751 5831
rect 89254 5828 89260 5840
rect 87739 5800 89260 5828
rect 87739 5797 87751 5800
rect 87693 5791 87751 5797
rect 43438 5760 43444 5772
rect 16546 5732 43444 5760
rect 43438 5720 43444 5732
rect 43496 5720 43502 5772
rect 47762 5720 47768 5772
rect 47820 5760 47826 5772
rect 51353 5763 51411 5769
rect 51353 5760 51365 5763
rect 47820 5732 51365 5760
rect 47820 5720 47826 5732
rect 51353 5729 51365 5732
rect 51399 5729 51411 5763
rect 51353 5723 51411 5729
rect 85761 5763 85819 5769
rect 85761 5729 85773 5763
rect 85807 5760 85819 5763
rect 86862 5760 86868 5772
rect 85807 5732 86868 5760
rect 85807 5729 85819 5732
rect 85761 5723 85819 5729
rect 86862 5720 86868 5732
rect 86920 5720 86926 5772
rect 86972 5760 87000 5791
rect 89254 5788 89260 5800
rect 89312 5788 89318 5840
rect 88978 5760 88984 5772
rect 86972 5732 88984 5760
rect 88978 5720 88984 5732
rect 89036 5720 89042 5772
rect 9766 5652 9772 5704
rect 9824 5692 9830 5704
rect 46934 5692 46940 5704
rect 9824 5664 46940 5692
rect 9824 5652 9830 5664
rect 46934 5652 46940 5664
rect 46992 5652 46998 5704
rect 47044 5664 47348 5692
rect 11974 5584 11980 5636
rect 12032 5624 12038 5636
rect 13354 5624 13360 5636
rect 12032 5596 13360 5624
rect 12032 5584 12038 5596
rect 13354 5584 13360 5596
rect 13412 5624 13418 5636
rect 47044 5624 47072 5664
rect 13412 5596 47072 5624
rect 47320 5624 47348 5664
rect 48038 5652 48044 5704
rect 48096 5692 48102 5704
rect 52457 5695 52515 5701
rect 52457 5692 52469 5695
rect 48096 5664 52469 5692
rect 48096 5652 48102 5664
rect 52457 5661 52469 5664
rect 52503 5661 52515 5695
rect 52457 5655 52515 5661
rect 86037 5695 86095 5701
rect 86037 5661 86049 5695
rect 86083 5692 86095 5695
rect 86310 5692 86316 5704
rect 86083 5664 86316 5692
rect 86083 5661 86095 5664
rect 86037 5655 86095 5661
rect 86310 5652 86316 5664
rect 86368 5652 86374 5704
rect 86402 5652 86408 5704
rect 86460 5652 86466 5704
rect 86773 5695 86831 5701
rect 86773 5661 86785 5695
rect 86819 5692 86831 5695
rect 87046 5692 87052 5704
rect 86819 5664 87052 5692
rect 86819 5661 86831 5664
rect 86773 5655 86831 5661
rect 87046 5652 87052 5664
rect 87104 5652 87110 5704
rect 87138 5652 87144 5704
rect 87196 5652 87202 5704
rect 87506 5652 87512 5704
rect 87564 5652 87570 5704
rect 87690 5652 87696 5704
rect 87748 5692 87754 5704
rect 87877 5695 87935 5701
rect 87877 5692 87889 5695
rect 87748 5664 87889 5692
rect 87748 5652 87754 5664
rect 87877 5661 87889 5664
rect 87923 5661 87935 5695
rect 87877 5655 87935 5661
rect 88242 5652 88248 5704
rect 88300 5652 88306 5704
rect 51902 5624 51908 5636
rect 47320 5596 51908 5624
rect 13412 5584 13418 5596
rect 51902 5584 51908 5596
rect 51960 5584 51966 5636
rect 85574 5584 85580 5636
rect 85632 5584 85638 5636
rect 86494 5584 86500 5636
rect 86552 5624 86558 5636
rect 87708 5624 87736 5652
rect 86552 5596 87736 5624
rect 86552 5584 86558 5596
rect 43438 5516 43444 5568
rect 43496 5556 43502 5568
rect 53006 5556 53012 5568
rect 43496 5528 53012 5556
rect 43496 5516 43502 5528
rect 53006 5516 53012 5528
rect 53064 5516 53070 5568
rect 85025 5559 85083 5565
rect 85025 5525 85037 5559
rect 85071 5556 85083 5559
rect 86512 5556 86540 5584
rect 85071 5528 86540 5556
rect 87325 5559 87383 5565
rect 85071 5525 85083 5528
rect 85025 5519 85083 5525
rect 87325 5525 87337 5559
rect 87371 5556 87383 5559
rect 89070 5556 89076 5568
rect 87371 5528 89076 5556
rect 87371 5525 87383 5528
rect 87325 5519 87383 5525
rect 89070 5516 89076 5528
rect 89128 5516 89134 5568
rect 1104 5466 88872 5488
rect 1104 5414 3802 5466
rect 3854 5414 3866 5466
rect 3918 5414 3930 5466
rect 3982 5414 3994 5466
rect 4046 5414 4058 5466
rect 4110 5414 37610 5466
rect 37662 5414 37674 5466
rect 37726 5414 37738 5466
rect 37790 5414 37802 5466
rect 37854 5414 37866 5466
rect 37918 5414 73610 5466
rect 73662 5414 73674 5466
rect 73726 5414 73738 5466
rect 73790 5414 73802 5466
rect 73854 5414 73866 5466
rect 73918 5414 88872 5466
rect 1104 5392 88872 5414
rect 85666 5312 85672 5364
rect 85724 5352 85730 5364
rect 85853 5355 85911 5361
rect 85853 5352 85865 5355
rect 85724 5324 85865 5352
rect 85724 5312 85730 5324
rect 85853 5321 85865 5324
rect 85899 5321 85911 5355
rect 85853 5315 85911 5321
rect 86034 5312 86040 5364
rect 86092 5312 86098 5364
rect 86494 5312 86500 5364
rect 86552 5312 86558 5364
rect 86678 5312 86684 5364
rect 86736 5312 86742 5364
rect 87693 5355 87751 5361
rect 87693 5321 87705 5355
rect 87739 5352 87751 5355
rect 87739 5324 88288 5352
rect 87739 5321 87751 5324
rect 87693 5315 87751 5321
rect 86313 5287 86371 5293
rect 86313 5253 86325 5287
rect 86359 5284 86371 5287
rect 86770 5284 86776 5296
rect 86359 5256 86776 5284
rect 86359 5253 86371 5256
rect 86313 5247 86371 5253
rect 86770 5244 86776 5256
rect 86828 5244 86834 5296
rect 87966 5284 87972 5296
rect 87156 5256 87972 5284
rect 87156 5225 87184 5256
rect 87966 5244 87972 5256
rect 88024 5244 88030 5296
rect 88260 5284 88288 5324
rect 88426 5312 88432 5364
rect 88484 5312 88490 5364
rect 88886 5284 88892 5296
rect 88260 5256 88892 5284
rect 88886 5244 88892 5256
rect 88944 5244 88950 5296
rect 86957 5219 87015 5225
rect 86957 5185 86969 5219
rect 87003 5185 87015 5219
rect 86957 5179 87015 5185
rect 87141 5219 87199 5225
rect 87141 5185 87153 5219
rect 87187 5185 87199 5219
rect 87141 5179 87199 5185
rect 83918 5108 83924 5160
rect 83976 5148 83982 5160
rect 86773 5151 86831 5157
rect 86773 5148 86785 5151
rect 83976 5120 86785 5148
rect 83976 5108 83982 5120
rect 86773 5117 86785 5120
rect 86819 5117 86831 5151
rect 86972 5148 87000 5179
rect 87414 5176 87420 5228
rect 87472 5216 87478 5228
rect 87509 5219 87567 5225
rect 87509 5216 87521 5219
rect 87472 5188 87521 5216
rect 87472 5176 87478 5188
rect 87509 5185 87521 5188
rect 87555 5185 87567 5219
rect 87509 5179 87567 5185
rect 87874 5176 87880 5228
rect 87932 5176 87938 5228
rect 88242 5176 88248 5228
rect 88300 5176 88306 5228
rect 88334 5148 88340 5160
rect 86972 5120 88340 5148
rect 86773 5111 86831 5117
rect 88334 5108 88340 5120
rect 88392 5108 88398 5160
rect 53834 5040 53840 5092
rect 53892 5080 53898 5092
rect 85669 5083 85727 5089
rect 85669 5080 85681 5083
rect 53892 5052 85681 5080
rect 53892 5040 53898 5052
rect 85669 5049 85681 5052
rect 85715 5049 85727 5083
rect 85669 5043 85727 5049
rect 88061 5083 88119 5089
rect 88061 5049 88073 5083
rect 88107 5080 88119 5083
rect 89346 5080 89352 5092
rect 88107 5052 89352 5080
rect 88107 5049 88119 5052
rect 88061 5043 88119 5049
rect 89346 5040 89352 5052
rect 89404 5040 89410 5092
rect 87325 5015 87383 5021
rect 87325 4981 87337 5015
rect 87371 5012 87383 5015
rect 88702 5012 88708 5024
rect 87371 4984 88708 5012
rect 87371 4981 87383 4984
rect 87325 4975 87383 4981
rect 88702 4972 88708 4984
rect 88760 4972 88766 5024
rect 1104 4922 88872 4944
rect 1104 4870 36950 4922
rect 37002 4870 37014 4922
rect 37066 4870 37078 4922
rect 37130 4870 37142 4922
rect 37194 4870 37206 4922
rect 37258 4870 72950 4922
rect 73002 4870 73014 4922
rect 73066 4870 73078 4922
rect 73130 4870 73142 4922
rect 73194 4870 73206 4922
rect 73258 4870 88872 4922
rect 1104 4848 88872 4870
rect 85758 4768 85764 4820
rect 85816 4808 85822 4820
rect 86773 4811 86831 4817
rect 86773 4808 86785 4811
rect 85816 4780 86785 4808
rect 85816 4768 85822 4780
rect 86773 4777 86785 4780
rect 86819 4777 86831 4811
rect 86773 4771 86831 4777
rect 87230 4768 87236 4820
rect 87288 4768 87294 4820
rect 87417 4811 87475 4817
rect 87417 4777 87429 4811
rect 87463 4808 87475 4811
rect 88150 4808 88156 4820
rect 87463 4780 88156 4808
rect 87463 4777 87475 4780
rect 87417 4771 87475 4777
rect 88150 4768 88156 4780
rect 88208 4768 88214 4820
rect 88429 4811 88487 4817
rect 88429 4777 88441 4811
rect 88475 4808 88487 4811
rect 89438 4808 89444 4820
rect 88475 4780 89444 4808
rect 88475 4777 88487 4780
rect 88429 4771 88487 4777
rect 89438 4768 89444 4780
rect 89496 4768 89502 4820
rect 87690 4700 87696 4752
rect 87748 4700 87754 4752
rect 88061 4743 88119 4749
rect 88061 4709 88073 4743
rect 88107 4740 88119 4743
rect 88794 4740 88800 4752
rect 88107 4712 88800 4740
rect 88107 4709 88119 4712
rect 88061 4703 88119 4709
rect 88794 4700 88800 4712
rect 88852 4700 88858 4752
rect 87601 4675 87659 4681
rect 87601 4641 87613 4675
rect 87647 4672 87659 4675
rect 88334 4672 88340 4684
rect 87647 4644 88340 4672
rect 87647 4641 87659 4644
rect 87601 4635 87659 4641
rect 88334 4632 88340 4644
rect 88392 4632 88398 4684
rect 87782 4564 87788 4616
rect 87840 4604 87846 4616
rect 87877 4607 87935 4613
rect 87877 4604 87889 4607
rect 87840 4576 87889 4604
rect 87840 4564 87846 4576
rect 87877 4573 87889 4576
rect 87923 4573 87935 4607
rect 87877 4567 87935 4573
rect 88245 4607 88303 4613
rect 88245 4573 88257 4607
rect 88291 4604 88303 4607
rect 88610 4604 88616 4616
rect 88291 4576 88616 4604
rect 88291 4573 88303 4576
rect 88245 4567 88303 4573
rect 88610 4564 88616 4576
rect 88668 4564 88674 4616
rect 47210 4496 47216 4548
rect 47268 4536 47274 4548
rect 86589 4539 86647 4545
rect 86589 4536 86601 4539
rect 47268 4508 86601 4536
rect 47268 4496 47274 4508
rect 86589 4505 86601 4508
rect 86635 4505 86647 4539
rect 86589 4499 86647 4505
rect 86954 4496 86960 4548
rect 87012 4496 87018 4548
rect 46842 4428 46848 4480
rect 46900 4468 46906 4480
rect 86405 4471 86463 4477
rect 86405 4468 86417 4471
rect 46900 4440 86417 4468
rect 46900 4428 46906 4440
rect 86405 4437 86417 4440
rect 86451 4437 86463 4471
rect 86405 4431 86463 4437
rect 1104 4378 88872 4400
rect 1104 4326 37610 4378
rect 37662 4326 37674 4378
rect 37726 4326 37738 4378
rect 37790 4326 37802 4378
rect 37854 4326 37866 4378
rect 37918 4326 73610 4378
rect 73662 4326 73674 4378
rect 73726 4326 73738 4378
rect 73790 4326 73802 4378
rect 73854 4326 73866 4378
rect 73918 4326 88872 4378
rect 1104 4304 88872 4326
rect 88150 4224 88156 4276
rect 88208 4224 88214 4276
rect 1104 3834 88872 3856
rect 1104 3782 36950 3834
rect 37002 3782 37014 3834
rect 37066 3782 37078 3834
rect 37130 3782 37142 3834
rect 37194 3782 37206 3834
rect 37258 3782 72950 3834
rect 73002 3782 73014 3834
rect 73066 3782 73078 3834
rect 73130 3782 73142 3834
rect 73194 3782 73206 3834
rect 73258 3782 88872 3834
rect 1104 3760 88872 3782
rect 1104 3290 88872 3312
rect 1104 3238 37610 3290
rect 37662 3238 37674 3290
rect 37726 3238 37738 3290
rect 37790 3238 37802 3290
rect 37854 3238 37866 3290
rect 37918 3238 73610 3290
rect 73662 3238 73674 3290
rect 73726 3238 73738 3290
rect 73790 3238 73802 3290
rect 73854 3238 73866 3290
rect 73918 3238 88872 3290
rect 1104 3216 88872 3238
rect 1104 2746 88872 2768
rect 1104 2694 36950 2746
rect 37002 2694 37014 2746
rect 37066 2694 37078 2746
rect 37130 2694 37142 2746
rect 37194 2694 37206 2746
rect 37258 2694 72950 2746
rect 73002 2694 73014 2746
rect 73066 2694 73078 2746
rect 73130 2694 73142 2746
rect 73194 2694 73206 2746
rect 73258 2694 88872 2746
rect 1104 2672 88872 2694
rect 8021 2635 8079 2641
rect 8021 2601 8033 2635
rect 8067 2632 8079 2635
rect 8294 2632 8300 2644
rect 8067 2604 8300 2632
rect 8067 2601 8079 2604
rect 8021 2595 8079 2601
rect 8294 2592 8300 2604
rect 8352 2592 8358 2644
rect 10870 2592 10876 2644
rect 10928 2632 10934 2644
rect 11609 2635 11667 2641
rect 11609 2632 11621 2635
rect 10928 2604 11621 2632
rect 10928 2592 10934 2604
rect 11609 2601 11621 2604
rect 11655 2601 11667 2635
rect 11609 2595 11667 2601
rect 13354 2592 13360 2644
rect 13412 2592 13418 2644
rect 15102 2632 15108 2644
rect 14936 2604 15108 2632
rect 8110 2524 8116 2576
rect 8168 2564 8174 2576
rect 8481 2567 8539 2573
rect 8481 2564 8493 2567
rect 8168 2536 8493 2564
rect 8168 2524 8174 2536
rect 8481 2533 8493 2536
rect 8527 2533 8539 2567
rect 8481 2527 8539 2533
rect 10597 2499 10655 2505
rect 10597 2465 10609 2499
rect 10643 2496 10655 2499
rect 10888 2496 10916 2592
rect 10643 2468 10916 2496
rect 13173 2499 13231 2505
rect 10643 2465 10655 2468
rect 10597 2459 10655 2465
rect 13173 2465 13185 2499
rect 13219 2496 13231 2499
rect 13372 2496 13400 2592
rect 14936 2505 14964 2604
rect 15102 2592 15108 2604
rect 15160 2592 15166 2644
rect 31018 2592 31024 2644
rect 31076 2592 31082 2644
rect 31846 2592 31852 2644
rect 31904 2592 31910 2644
rect 32950 2592 32956 2644
rect 33008 2592 33014 2644
rect 34238 2592 34244 2644
rect 34296 2592 34302 2644
rect 35066 2592 35072 2644
rect 35124 2592 35130 2644
rect 36170 2592 36176 2644
rect 36228 2592 36234 2644
rect 37458 2592 37464 2644
rect 37516 2592 37522 2644
rect 42794 2592 42800 2644
rect 42852 2592 42858 2644
rect 45186 2592 45192 2644
rect 45244 2592 45250 2644
rect 70946 2592 70952 2644
rect 71004 2592 71010 2644
rect 71774 2592 71780 2644
rect 71832 2592 71838 2644
rect 72786 2592 72792 2644
rect 72844 2632 72850 2644
rect 72881 2635 72939 2641
rect 72881 2632 72893 2635
rect 72844 2604 72893 2632
rect 72844 2592 72850 2604
rect 72881 2601 72893 2604
rect 72927 2601 72939 2635
rect 72881 2595 72939 2601
rect 74166 2592 74172 2644
rect 74224 2592 74230 2644
rect 75086 2592 75092 2644
rect 75144 2632 75150 2644
rect 75457 2635 75515 2641
rect 75457 2632 75469 2635
rect 75144 2604 75469 2632
rect 75144 2592 75150 2604
rect 75457 2601 75469 2604
rect 75503 2601 75515 2635
rect 75457 2595 75515 2601
rect 76282 2592 76288 2644
rect 76340 2592 76346 2644
rect 77386 2592 77392 2644
rect 77444 2592 77450 2644
rect 39850 2524 39856 2576
rect 39908 2524 39914 2576
rect 40678 2524 40684 2576
rect 40736 2524 40742 2576
rect 41966 2524 41972 2576
rect 42024 2524 42030 2576
rect 43898 2524 43904 2576
rect 43956 2524 43962 2576
rect 79594 2524 79600 2576
rect 79652 2524 79658 2576
rect 80606 2524 80612 2576
rect 80664 2524 80670 2576
rect 81894 2524 81900 2576
rect 81952 2524 81958 2576
rect 82814 2524 82820 2576
rect 82872 2564 82878 2576
rect 83185 2567 83243 2573
rect 83185 2564 83197 2567
rect 82872 2536 83197 2564
rect 82872 2524 82878 2536
rect 83185 2533 83197 2536
rect 83231 2533 83243 2567
rect 83185 2527 83243 2533
rect 13219 2468 13400 2496
rect 14921 2499 14979 2505
rect 13219 2465 13231 2468
rect 13173 2459 13231 2465
rect 14921 2465 14933 2499
rect 14967 2465 14979 2499
rect 14921 2459 14979 2465
rect 38378 2456 38384 2508
rect 38436 2496 38442 2508
rect 39025 2499 39083 2505
rect 39025 2496 39037 2499
rect 38436 2468 39037 2496
rect 38436 2456 38442 2468
rect 39025 2465 39037 2468
rect 39071 2465 39083 2499
rect 39025 2459 39083 2465
rect 78398 2456 78404 2508
rect 78456 2496 78462 2508
rect 78953 2499 79011 2505
rect 78953 2496 78965 2499
rect 78456 2468 78965 2496
rect 78456 2456 78462 2468
rect 78953 2465 78965 2468
rect 78999 2465 79011 2499
rect 78953 2459 79011 2465
rect 7837 2431 7895 2437
rect 7837 2428 7849 2431
rect 7760 2400 7849 2428
rect 7760 2304 7788 2400
rect 7837 2397 7849 2400
rect 7883 2397 7895 2431
rect 8665 2431 8723 2437
rect 8665 2428 8677 2431
rect 7837 2391 7895 2397
rect 8404 2400 8677 2428
rect 8404 2304 8432 2400
rect 8665 2397 8677 2400
rect 8711 2397 8723 2431
rect 8665 2391 8723 2397
rect 15562 2388 15568 2440
rect 15620 2388 15626 2440
rect 16482 2388 16488 2440
rect 16540 2388 16546 2440
rect 17494 2388 17500 2440
rect 17552 2388 17558 2440
rect 18782 2388 18788 2440
rect 18840 2388 18846 2440
rect 19702 2388 19708 2440
rect 19760 2388 19766 2440
rect 20714 2388 20720 2440
rect 20772 2388 20778 2440
rect 22002 2388 22008 2440
rect 22060 2388 22066 2440
rect 23290 2388 23296 2440
rect 23348 2388 23354 2440
rect 24210 2388 24216 2440
rect 24268 2388 24274 2440
rect 25222 2388 25228 2440
rect 25280 2388 25286 2440
rect 26510 2388 26516 2440
rect 26568 2388 26574 2440
rect 27430 2388 27436 2440
rect 27488 2388 27494 2440
rect 28442 2388 28448 2440
rect 28500 2388 28506 2440
rect 29730 2388 29736 2440
rect 29788 2388 29794 2440
rect 31205 2431 31263 2437
rect 31205 2428 31217 2431
rect 30944 2400 31217 2428
rect 10962 2320 10968 2372
rect 11020 2360 11026 2372
rect 11333 2363 11391 2369
rect 11333 2360 11345 2363
rect 11020 2332 11345 2360
rect 11020 2320 11026 2332
rect 11333 2329 11345 2332
rect 11379 2360 11391 2363
rect 11793 2363 11851 2369
rect 11793 2360 11805 2363
rect 11379 2332 11805 2360
rect 11379 2329 11391 2332
rect 11333 2323 11391 2329
rect 11793 2329 11805 2332
rect 11839 2329 11851 2363
rect 11793 2323 11851 2329
rect 12345 2363 12403 2369
rect 12345 2329 12357 2363
rect 12391 2329 12403 2363
rect 12345 2323 12403 2329
rect 14093 2363 14151 2369
rect 14093 2329 14105 2363
rect 14139 2329 14151 2363
rect 14093 2323 14151 2329
rect 7742 2252 7748 2304
rect 7800 2252 7806 2304
rect 8386 2252 8392 2304
rect 8444 2252 8450 2304
rect 12250 2252 12256 2304
rect 12308 2292 12314 2304
rect 12360 2292 12388 2323
rect 12308 2264 12388 2292
rect 12308 2252 12314 2264
rect 13538 2252 13544 2304
rect 13596 2292 13602 2304
rect 13817 2295 13875 2301
rect 13817 2292 13829 2295
rect 13596 2264 13829 2292
rect 13596 2252 13602 2264
rect 13817 2261 13829 2264
rect 13863 2292 13875 2295
rect 14108 2292 14136 2323
rect 30944 2304 30972 2400
rect 31205 2397 31217 2400
rect 31251 2397 31263 2431
rect 31665 2431 31723 2437
rect 31665 2428 31677 2431
rect 31205 2391 31263 2397
rect 31588 2400 31677 2428
rect 31588 2304 31616 2400
rect 31665 2397 31677 2400
rect 31711 2397 31723 2431
rect 33137 2431 33195 2437
rect 33137 2428 33149 2431
rect 31665 2391 31723 2397
rect 32876 2400 33149 2428
rect 32876 2304 32904 2400
rect 33137 2397 33149 2400
rect 33183 2397 33195 2431
rect 34425 2431 34483 2437
rect 34425 2428 34437 2431
rect 33137 2391 33195 2397
rect 34164 2400 34437 2428
rect 34164 2304 34192 2400
rect 34425 2397 34437 2400
rect 34471 2397 34483 2431
rect 34885 2431 34943 2437
rect 34885 2428 34897 2431
rect 34425 2391 34483 2397
rect 34808 2400 34897 2428
rect 34808 2304 34836 2400
rect 34885 2397 34897 2400
rect 34931 2397 34943 2431
rect 36357 2431 36415 2437
rect 36357 2428 36369 2431
rect 34885 2391 34943 2397
rect 36096 2400 36369 2428
rect 36096 2304 36124 2400
rect 36357 2397 36369 2400
rect 36403 2397 36415 2431
rect 37645 2431 37703 2437
rect 37645 2428 37657 2431
rect 36357 2391 36415 2397
rect 37384 2400 37657 2428
rect 37384 2304 37412 2400
rect 37645 2397 37657 2400
rect 37691 2397 37703 2431
rect 38749 2431 38807 2437
rect 38749 2428 38761 2431
rect 37645 2391 37703 2397
rect 38672 2400 38761 2428
rect 38672 2304 38700 2400
rect 38749 2397 38761 2400
rect 38795 2397 38807 2431
rect 45373 2431 45431 2437
rect 45373 2428 45385 2431
rect 38749 2391 38807 2397
rect 45112 2400 45385 2428
rect 39298 2320 39304 2372
rect 39356 2360 39362 2372
rect 40037 2363 40095 2369
rect 40037 2360 40049 2363
rect 39356 2332 40049 2360
rect 39356 2320 39362 2332
rect 40037 2329 40049 2332
rect 40083 2360 40095 2363
rect 40221 2363 40279 2369
rect 40221 2360 40233 2363
rect 40083 2332 40233 2360
rect 40083 2329 40095 2332
rect 40037 2323 40095 2329
rect 40221 2329 40233 2332
rect 40267 2329 40279 2363
rect 40221 2323 40279 2329
rect 40865 2363 40923 2369
rect 40865 2329 40877 2363
rect 40911 2329 40923 2363
rect 40865 2323 40923 2329
rect 42153 2363 42211 2369
rect 42153 2329 42165 2363
rect 42199 2329 42211 2363
rect 42153 2323 42211 2329
rect 42705 2363 42763 2369
rect 42705 2329 42717 2363
rect 42751 2329 42763 2363
rect 42705 2323 42763 2329
rect 44085 2363 44143 2369
rect 44085 2329 44097 2363
rect 44131 2329 44143 2363
rect 44085 2323 44143 2329
rect 13863 2264 14136 2292
rect 13863 2261 13875 2264
rect 13817 2255 13875 2261
rect 15470 2252 15476 2304
rect 15528 2292 15534 2304
rect 15749 2295 15807 2301
rect 15749 2292 15761 2295
rect 15528 2264 15761 2292
rect 15528 2252 15534 2264
rect 15749 2261 15761 2264
rect 15795 2261 15807 2295
rect 15749 2255 15807 2261
rect 16114 2252 16120 2304
rect 16172 2292 16178 2304
rect 16301 2295 16359 2301
rect 16301 2292 16313 2295
rect 16172 2264 16313 2292
rect 16172 2252 16178 2264
rect 16301 2261 16313 2264
rect 16347 2261 16359 2295
rect 16301 2255 16359 2261
rect 17402 2252 17408 2304
rect 17460 2292 17466 2304
rect 17681 2295 17739 2301
rect 17681 2292 17693 2295
rect 17460 2264 17693 2292
rect 17460 2252 17466 2264
rect 17681 2261 17693 2264
rect 17727 2261 17739 2295
rect 17681 2255 17739 2261
rect 18690 2252 18696 2304
rect 18748 2292 18754 2304
rect 18969 2295 19027 2301
rect 18969 2292 18981 2295
rect 18748 2264 18981 2292
rect 18748 2252 18754 2264
rect 18969 2261 18981 2264
rect 19015 2261 19027 2295
rect 18969 2255 19027 2261
rect 19334 2252 19340 2304
rect 19392 2292 19398 2304
rect 19521 2295 19579 2301
rect 19521 2292 19533 2295
rect 19392 2264 19533 2292
rect 19392 2252 19398 2264
rect 19521 2261 19533 2264
rect 19567 2261 19579 2295
rect 19521 2255 19579 2261
rect 20622 2252 20628 2304
rect 20680 2292 20686 2304
rect 20901 2295 20959 2301
rect 20901 2292 20913 2295
rect 20680 2264 20913 2292
rect 20680 2252 20686 2264
rect 20901 2261 20913 2264
rect 20947 2261 20959 2295
rect 20901 2255 20959 2261
rect 21910 2252 21916 2304
rect 21968 2292 21974 2304
rect 22189 2295 22247 2301
rect 22189 2292 22201 2295
rect 21968 2264 22201 2292
rect 21968 2252 21974 2264
rect 22189 2261 22201 2264
rect 22235 2261 22247 2295
rect 22189 2255 22247 2261
rect 23198 2252 23204 2304
rect 23256 2292 23262 2304
rect 23477 2295 23535 2301
rect 23477 2292 23489 2295
rect 23256 2264 23489 2292
rect 23256 2252 23262 2264
rect 23477 2261 23489 2264
rect 23523 2261 23535 2295
rect 23477 2255 23535 2261
rect 23842 2252 23848 2304
rect 23900 2292 23906 2304
rect 24029 2295 24087 2301
rect 24029 2292 24041 2295
rect 23900 2264 24041 2292
rect 23900 2252 23906 2264
rect 24029 2261 24041 2264
rect 24075 2261 24087 2295
rect 24029 2255 24087 2261
rect 25130 2252 25136 2304
rect 25188 2292 25194 2304
rect 25409 2295 25467 2301
rect 25409 2292 25421 2295
rect 25188 2264 25421 2292
rect 25188 2252 25194 2264
rect 25409 2261 25421 2264
rect 25455 2261 25467 2295
rect 25409 2255 25467 2261
rect 26418 2252 26424 2304
rect 26476 2292 26482 2304
rect 26697 2295 26755 2301
rect 26697 2292 26709 2295
rect 26476 2264 26709 2292
rect 26476 2252 26482 2264
rect 26697 2261 26709 2264
rect 26743 2261 26755 2295
rect 26697 2255 26755 2261
rect 27062 2252 27068 2304
rect 27120 2292 27126 2304
rect 27249 2295 27307 2301
rect 27249 2292 27261 2295
rect 27120 2264 27261 2292
rect 27120 2252 27126 2264
rect 27249 2261 27261 2264
rect 27295 2261 27307 2295
rect 27249 2255 27307 2261
rect 28350 2252 28356 2304
rect 28408 2292 28414 2304
rect 28629 2295 28687 2301
rect 28629 2292 28641 2295
rect 28408 2264 28641 2292
rect 28408 2252 28414 2264
rect 28629 2261 28641 2264
rect 28675 2261 28687 2295
rect 28629 2255 28687 2261
rect 29638 2252 29644 2304
rect 29696 2292 29702 2304
rect 29917 2295 29975 2301
rect 29917 2292 29929 2295
rect 29696 2264 29929 2292
rect 29696 2252 29702 2264
rect 29917 2261 29929 2264
rect 29963 2261 29975 2295
rect 29917 2255 29975 2261
rect 30926 2252 30932 2304
rect 30984 2252 30990 2304
rect 31570 2252 31576 2304
rect 31628 2252 31634 2304
rect 32858 2252 32864 2304
rect 32916 2252 32922 2304
rect 34146 2252 34152 2304
rect 34204 2252 34210 2304
rect 34790 2252 34796 2304
rect 34848 2252 34854 2304
rect 36078 2252 36084 2304
rect 36136 2252 36142 2304
rect 37366 2252 37372 2304
rect 37424 2252 37430 2304
rect 38654 2252 38660 2304
rect 38712 2252 38718 2304
rect 40586 2252 40592 2304
rect 40644 2292 40650 2304
rect 40880 2292 40908 2323
rect 40644 2264 40908 2292
rect 40644 2252 40650 2264
rect 41874 2252 41880 2304
rect 41932 2292 41938 2304
rect 42168 2292 42196 2323
rect 41932 2264 42196 2292
rect 41932 2252 41938 2264
rect 42518 2252 42524 2304
rect 42576 2292 42582 2304
rect 42720 2292 42748 2323
rect 42576 2264 42748 2292
rect 42576 2252 42582 2264
rect 43806 2252 43812 2304
rect 43864 2292 43870 2304
rect 44100 2292 44128 2323
rect 45112 2304 45140 2400
rect 45373 2397 45385 2400
rect 45419 2397 45431 2431
rect 45373 2391 45431 2397
rect 55490 2388 55496 2440
rect 55548 2388 55554 2440
rect 56410 2388 56416 2440
rect 56468 2388 56474 2440
rect 57422 2388 57428 2440
rect 57480 2388 57486 2440
rect 58710 2388 58716 2440
rect 58768 2388 58774 2440
rect 59630 2388 59636 2440
rect 59688 2428 59694 2440
rect 60001 2431 60059 2437
rect 60001 2428 60013 2431
rect 59688 2400 60013 2428
rect 59688 2388 59694 2400
rect 60001 2397 60013 2400
rect 60047 2397 60059 2431
rect 60001 2391 60059 2397
rect 60645 2431 60703 2437
rect 60645 2397 60657 2431
rect 60691 2428 60703 2431
rect 60734 2428 60740 2440
rect 60691 2400 60740 2428
rect 60691 2397 60703 2400
rect 60645 2391 60703 2397
rect 60734 2388 60740 2400
rect 60792 2388 60798 2440
rect 61930 2388 61936 2440
rect 61988 2388 61994 2440
rect 63218 2388 63224 2440
rect 63276 2388 63282 2440
rect 64138 2388 64144 2440
rect 64196 2388 64202 2440
rect 65150 2388 65156 2440
rect 65208 2388 65214 2440
rect 66438 2388 66444 2440
rect 66496 2388 66502 2440
rect 67358 2388 67364 2440
rect 67416 2428 67422 2440
rect 67729 2431 67787 2437
rect 67729 2428 67741 2431
rect 67416 2400 67741 2428
rect 67416 2388 67422 2400
rect 67729 2397 67741 2400
rect 67775 2397 67787 2431
rect 67729 2391 67787 2397
rect 68370 2388 68376 2440
rect 68428 2388 68434 2440
rect 69658 2388 69664 2440
rect 69716 2388 69722 2440
rect 71133 2431 71191 2437
rect 71133 2428 71145 2431
rect 70872 2400 71145 2428
rect 70872 2304 70900 2400
rect 71133 2397 71145 2400
rect 71179 2397 71191 2431
rect 71593 2431 71651 2437
rect 71593 2428 71605 2431
rect 71133 2391 71191 2397
rect 71516 2400 71605 2428
rect 71516 2304 71544 2400
rect 71593 2397 71605 2400
rect 71639 2397 71651 2431
rect 73065 2431 73123 2437
rect 73065 2428 73077 2431
rect 71593 2391 71651 2397
rect 72804 2400 73077 2428
rect 72804 2304 72832 2400
rect 73065 2397 73077 2400
rect 73111 2397 73123 2431
rect 74353 2431 74411 2437
rect 74353 2428 74365 2431
rect 73065 2391 73123 2397
rect 74092 2400 74365 2428
rect 74092 2304 74120 2400
rect 74353 2397 74365 2400
rect 74399 2397 74411 2431
rect 75641 2431 75699 2437
rect 75641 2428 75653 2431
rect 74353 2391 74411 2397
rect 75380 2400 75653 2428
rect 75380 2304 75408 2400
rect 75641 2397 75653 2400
rect 75687 2397 75699 2431
rect 76101 2431 76159 2437
rect 76101 2428 76113 2431
rect 75641 2391 75699 2397
rect 76024 2400 76113 2428
rect 76024 2304 76052 2400
rect 76101 2397 76113 2400
rect 76147 2397 76159 2431
rect 77573 2431 77631 2437
rect 77573 2428 77585 2431
rect 76101 2391 76159 2397
rect 77312 2400 77585 2428
rect 77312 2304 77340 2400
rect 77573 2397 77585 2400
rect 77619 2397 77631 2431
rect 78677 2431 78735 2437
rect 78677 2428 78689 2431
rect 77573 2391 77631 2397
rect 78600 2400 78689 2428
rect 78600 2304 78628 2400
rect 78677 2397 78689 2400
rect 78723 2397 78735 2431
rect 78677 2391 78735 2397
rect 79226 2320 79232 2372
rect 79284 2360 79290 2372
rect 79781 2363 79839 2369
rect 79781 2360 79793 2363
rect 79284 2332 79793 2360
rect 79284 2320 79290 2332
rect 79781 2329 79793 2332
rect 79827 2360 79839 2363
rect 79965 2363 80023 2369
rect 79965 2360 79977 2363
rect 79827 2332 79977 2360
rect 79827 2329 79839 2332
rect 79781 2323 79839 2329
rect 79965 2329 79977 2332
rect 80011 2329 80023 2363
rect 79965 2323 80023 2329
rect 80793 2363 80851 2369
rect 80793 2329 80805 2363
rect 80839 2329 80851 2363
rect 80793 2323 80851 2329
rect 82081 2363 82139 2369
rect 82081 2329 82093 2363
rect 82127 2329 82139 2363
rect 82081 2323 82139 2329
rect 83369 2363 83427 2369
rect 83369 2329 83381 2363
rect 83415 2329 83427 2363
rect 83369 2323 83427 2329
rect 43864 2264 44128 2292
rect 43864 2252 43870 2264
rect 45094 2252 45100 2304
rect 45152 2252 45158 2304
rect 55398 2252 55404 2304
rect 55456 2292 55462 2304
rect 55677 2295 55735 2301
rect 55677 2292 55689 2295
rect 55456 2264 55689 2292
rect 55456 2252 55462 2264
rect 55677 2261 55689 2264
rect 55723 2261 55735 2295
rect 55677 2255 55735 2261
rect 56042 2252 56048 2304
rect 56100 2292 56106 2304
rect 56229 2295 56287 2301
rect 56229 2292 56241 2295
rect 56100 2264 56241 2292
rect 56100 2252 56106 2264
rect 56229 2261 56241 2264
rect 56275 2261 56287 2295
rect 56229 2255 56287 2261
rect 57330 2252 57336 2304
rect 57388 2292 57394 2304
rect 57609 2295 57667 2301
rect 57609 2292 57621 2295
rect 57388 2264 57621 2292
rect 57388 2252 57394 2264
rect 57609 2261 57621 2264
rect 57655 2261 57667 2295
rect 57609 2255 57667 2261
rect 58618 2252 58624 2304
rect 58676 2292 58682 2304
rect 58897 2295 58955 2301
rect 58897 2292 58909 2295
rect 58676 2264 58909 2292
rect 58676 2252 58682 2264
rect 58897 2261 58909 2264
rect 58943 2261 58955 2295
rect 58897 2255 58955 2261
rect 59906 2252 59912 2304
rect 59964 2292 59970 2304
rect 60185 2295 60243 2301
rect 60185 2292 60197 2295
rect 59964 2264 60197 2292
rect 59964 2252 59970 2264
rect 60185 2261 60197 2264
rect 60231 2261 60243 2295
rect 60185 2255 60243 2261
rect 60550 2252 60556 2304
rect 60608 2292 60614 2304
rect 60829 2295 60887 2301
rect 60829 2292 60841 2295
rect 60608 2264 60841 2292
rect 60608 2252 60614 2264
rect 60829 2261 60841 2264
rect 60875 2261 60887 2295
rect 60829 2255 60887 2261
rect 61838 2252 61844 2304
rect 61896 2292 61902 2304
rect 62117 2295 62175 2301
rect 62117 2292 62129 2295
rect 61896 2264 62129 2292
rect 61896 2252 61902 2264
rect 62117 2261 62129 2264
rect 62163 2261 62175 2295
rect 62117 2255 62175 2261
rect 63126 2252 63132 2304
rect 63184 2292 63190 2304
rect 63405 2295 63463 2301
rect 63405 2292 63417 2295
rect 63184 2264 63417 2292
rect 63184 2252 63190 2264
rect 63405 2261 63417 2264
rect 63451 2261 63463 2295
rect 63405 2255 63463 2261
rect 63770 2252 63776 2304
rect 63828 2292 63834 2304
rect 63957 2295 64015 2301
rect 63957 2292 63969 2295
rect 63828 2264 63969 2292
rect 63828 2252 63834 2264
rect 63957 2261 63969 2264
rect 64003 2261 64015 2295
rect 63957 2255 64015 2261
rect 65058 2252 65064 2304
rect 65116 2292 65122 2304
rect 65337 2295 65395 2301
rect 65337 2292 65349 2295
rect 65116 2264 65349 2292
rect 65116 2252 65122 2264
rect 65337 2261 65349 2264
rect 65383 2261 65395 2295
rect 65337 2255 65395 2261
rect 66346 2252 66352 2304
rect 66404 2292 66410 2304
rect 66625 2295 66683 2301
rect 66625 2292 66637 2295
rect 66404 2264 66637 2292
rect 66404 2252 66410 2264
rect 66625 2261 66637 2264
rect 66671 2261 66683 2295
rect 66625 2255 66683 2261
rect 67634 2252 67640 2304
rect 67692 2292 67698 2304
rect 67913 2295 67971 2301
rect 67913 2292 67925 2295
rect 67692 2264 67925 2292
rect 67692 2252 67698 2264
rect 67913 2261 67925 2264
rect 67959 2261 67971 2295
rect 67913 2255 67971 2261
rect 68278 2252 68284 2304
rect 68336 2292 68342 2304
rect 68557 2295 68615 2301
rect 68557 2292 68569 2295
rect 68336 2264 68569 2292
rect 68336 2252 68342 2264
rect 68557 2261 68569 2264
rect 68603 2261 68615 2295
rect 68557 2255 68615 2261
rect 69566 2252 69572 2304
rect 69624 2292 69630 2304
rect 69845 2295 69903 2301
rect 69845 2292 69857 2295
rect 69624 2264 69857 2292
rect 69624 2252 69630 2264
rect 69845 2261 69857 2264
rect 69891 2261 69903 2295
rect 69845 2255 69903 2261
rect 70854 2252 70860 2304
rect 70912 2252 70918 2304
rect 71498 2252 71504 2304
rect 71556 2252 71562 2304
rect 72786 2252 72792 2304
rect 72844 2252 72850 2304
rect 74074 2252 74080 2304
rect 74132 2252 74138 2304
rect 75362 2252 75368 2304
rect 75420 2252 75426 2304
rect 76006 2252 76012 2304
rect 76064 2252 76070 2304
rect 77294 2252 77300 2304
rect 77352 2252 77358 2304
rect 78582 2252 78588 2304
rect 78640 2252 78646 2304
rect 80514 2252 80520 2304
rect 80572 2292 80578 2304
rect 80808 2292 80836 2323
rect 80572 2264 80836 2292
rect 80572 2252 80578 2264
rect 81802 2252 81808 2304
rect 81860 2292 81866 2304
rect 82096 2292 82124 2323
rect 81860 2264 82124 2292
rect 81860 2252 81866 2264
rect 83090 2252 83096 2304
rect 83148 2292 83154 2304
rect 83384 2292 83412 2323
rect 83148 2264 83412 2292
rect 83148 2252 83154 2264
rect 1104 2202 88872 2224
rect 1104 2150 37610 2202
rect 37662 2150 37674 2202
rect 37726 2150 37738 2202
rect 37790 2150 37802 2202
rect 37854 2150 37866 2202
rect 37918 2150 73610 2202
rect 73662 2150 73674 2202
rect 73726 2150 73738 2202
rect 73790 2150 73802 2202
rect 73854 2150 73866 2202
rect 73918 2150 88872 2202
rect 1104 2128 88872 2150
<< via1 >>
rect 37610 95718 37662 95770
rect 37674 95718 37726 95770
rect 37738 95718 37790 95770
rect 37802 95718 37854 95770
rect 37866 95718 37918 95770
rect 73610 95718 73662 95770
rect 73674 95718 73726 95770
rect 73738 95718 73790 95770
rect 73802 95718 73854 95770
rect 73866 95718 73918 95770
rect 8668 95659 8720 95668
rect 8668 95625 8677 95659
rect 8677 95625 8711 95659
rect 8711 95625 8720 95659
rect 8668 95616 8720 95625
rect 14740 95659 14792 95668
rect 14740 95625 14749 95659
rect 14749 95625 14783 95659
rect 14783 95625 14792 95659
rect 14740 95616 14792 95625
rect 16672 95659 16724 95668
rect 16672 95625 16681 95659
rect 16681 95625 16715 95659
rect 16715 95625 16724 95659
rect 16672 95616 16724 95625
rect 17960 95659 18012 95668
rect 17960 95625 17969 95659
rect 17969 95625 18003 95659
rect 18003 95625 18012 95659
rect 17960 95616 18012 95625
rect 19432 95616 19484 95668
rect 20352 95616 20404 95668
rect 21180 95659 21232 95668
rect 21180 95625 21189 95659
rect 21189 95625 21223 95659
rect 21223 95625 21232 95659
rect 21180 95616 21232 95625
rect 22468 95659 22520 95668
rect 22468 95625 22477 95659
rect 22477 95625 22511 95659
rect 22511 95625 22520 95659
rect 22468 95616 22520 95625
rect 8484 95523 8536 95532
rect 8484 95489 8493 95523
rect 8493 95489 8527 95523
rect 8527 95489 8536 95523
rect 8484 95480 8536 95489
rect 15568 95523 15620 95532
rect 15568 95489 15577 95523
rect 15577 95489 15611 95523
rect 15611 95489 15620 95523
rect 15568 95480 15620 95489
rect 23112 95659 23164 95668
rect 23112 95625 23121 95659
rect 23121 95625 23155 95659
rect 23155 95625 23164 95659
rect 23112 95616 23164 95625
rect 24400 95659 24452 95668
rect 24400 95625 24409 95659
rect 24409 95625 24443 95659
rect 24443 95625 24452 95659
rect 24400 95616 24452 95625
rect 25688 95659 25740 95668
rect 25688 95625 25697 95659
rect 25697 95625 25731 95659
rect 25731 95625 25740 95659
rect 25688 95616 25740 95625
rect 26976 95659 27028 95668
rect 26976 95625 26985 95659
rect 26985 95625 27019 95659
rect 27019 95625 27028 95659
rect 26976 95616 27028 95625
rect 27620 95659 27672 95668
rect 27620 95625 27629 95659
rect 27629 95625 27663 95659
rect 27663 95625 27672 95659
rect 27620 95616 27672 95625
rect 29092 95616 29144 95668
rect 30196 95616 30248 95668
rect 31116 95659 31168 95668
rect 31116 95625 31125 95659
rect 31125 95625 31159 95659
rect 31159 95625 31168 95659
rect 31116 95616 31168 95625
rect 32496 95659 32548 95668
rect 32496 95625 32505 95659
rect 32505 95625 32539 95659
rect 32539 95625 32548 95659
rect 32496 95616 32548 95625
rect 33784 95659 33836 95668
rect 33784 95625 33793 95659
rect 33793 95625 33827 95659
rect 33827 95625 33836 95659
rect 33784 95616 33836 95625
rect 35072 95659 35124 95668
rect 35072 95625 35081 95659
rect 35081 95625 35115 95659
rect 35115 95625 35124 95659
rect 35072 95616 35124 95625
rect 35624 95659 35676 95668
rect 35624 95625 35633 95659
rect 35633 95625 35667 95659
rect 35667 95625 35676 95659
rect 35624 95616 35676 95625
rect 37004 95659 37056 95668
rect 37004 95625 37013 95659
rect 37013 95625 37047 95659
rect 37047 95625 37056 95659
rect 37004 95616 37056 95625
rect 38292 95659 38344 95668
rect 38292 95625 38301 95659
rect 38301 95625 38335 95659
rect 38335 95625 38344 95659
rect 38292 95616 38344 95625
rect 38844 95659 38896 95668
rect 38844 95625 38853 95659
rect 38853 95625 38887 95659
rect 38887 95625 38896 95659
rect 38844 95616 38896 95625
rect 39856 95616 39908 95668
rect 41328 95616 41380 95668
rect 42708 95616 42760 95668
rect 43352 95659 43404 95668
rect 43352 95625 43361 95659
rect 43361 95625 43395 95659
rect 43395 95625 43404 95659
rect 43352 95616 43404 95625
rect 44732 95659 44784 95668
rect 44732 95625 44741 95659
rect 44741 95625 44775 95659
rect 44775 95625 44784 95659
rect 44732 95616 44784 95625
rect 50804 95659 50856 95668
rect 50804 95625 50813 95659
rect 50813 95625 50847 95659
rect 50847 95625 50856 95659
rect 50804 95616 50856 95625
rect 56416 95616 56468 95668
rect 56968 95616 57020 95668
rect 30104 95480 30156 95532
rect 31300 95523 31352 95532
rect 31300 95489 31309 95523
rect 31309 95489 31343 95523
rect 31343 95489 31352 95523
rect 31300 95480 31352 95489
rect 32312 95523 32364 95532
rect 32312 95489 32321 95523
rect 32321 95489 32355 95523
rect 32355 95489 32364 95523
rect 32312 95480 32364 95489
rect 33600 95523 33652 95532
rect 33600 95489 33609 95523
rect 33609 95489 33643 95523
rect 33643 95489 33652 95523
rect 33600 95480 33652 95489
rect 34888 95523 34940 95532
rect 34888 95489 34897 95523
rect 34897 95489 34931 95523
rect 34931 95489 34940 95523
rect 34888 95480 34940 95489
rect 35808 95523 35860 95532
rect 35808 95489 35817 95523
rect 35817 95489 35851 95523
rect 35851 95489 35860 95523
rect 35808 95480 35860 95489
rect 36820 95523 36872 95532
rect 36820 95489 36829 95523
rect 36829 95489 36863 95523
rect 36863 95489 36872 95523
rect 36820 95480 36872 95489
rect 38108 95523 38160 95532
rect 38108 95489 38117 95523
rect 38117 95489 38151 95523
rect 38151 95489 38160 95523
rect 38108 95480 38160 95489
rect 39028 95523 39080 95532
rect 39028 95489 39037 95523
rect 39037 95489 39071 95523
rect 39071 95489 39080 95523
rect 39028 95480 39080 95489
rect 40040 95523 40092 95532
rect 40040 95489 40049 95523
rect 40049 95489 40083 95523
rect 40083 95489 40092 95523
rect 40040 95480 40092 95489
rect 41328 95523 41380 95532
rect 41328 95489 41337 95523
rect 41337 95489 41371 95523
rect 41371 95489 41380 95523
rect 41328 95480 41380 95489
rect 42616 95523 42668 95532
rect 42616 95489 42625 95523
rect 42625 95489 42659 95523
rect 42659 95489 42668 95523
rect 42616 95480 42668 95489
rect 43536 95523 43588 95532
rect 43536 95489 43545 95523
rect 43545 95489 43579 95523
rect 43579 95489 43588 95523
rect 43536 95480 43588 95489
rect 44548 95523 44600 95532
rect 44548 95489 44557 95523
rect 44557 95489 44591 95523
rect 44591 95489 44600 95523
rect 44548 95480 44600 95489
rect 54944 95548 54996 95600
rect 52276 95480 52328 95532
rect 58072 95616 58124 95668
rect 59176 95659 59228 95668
rect 59176 95625 59185 95659
rect 59185 95625 59219 95659
rect 59219 95625 59228 95659
rect 59176 95616 59228 95625
rect 61108 95659 61160 95668
rect 61108 95625 61117 95659
rect 61117 95625 61151 95659
rect 61151 95625 61160 95659
rect 61108 95616 61160 95625
rect 62396 95659 62448 95668
rect 62396 95625 62405 95659
rect 62405 95625 62439 95659
rect 62439 95625 62448 95659
rect 62396 95616 62448 95625
rect 60004 95523 60056 95532
rect 60004 95489 60013 95523
rect 60013 95489 60047 95523
rect 60047 95489 60056 95523
rect 60004 95480 60056 95489
rect 63684 95659 63736 95668
rect 63684 95625 63693 95659
rect 63693 95625 63727 95659
rect 63727 95625 63736 95659
rect 63684 95616 63736 95625
rect 64604 95616 64656 95668
rect 65616 95659 65668 95668
rect 65616 95625 65625 95659
rect 65625 95625 65659 95659
rect 65659 95625 65668 95659
rect 65616 95616 65668 95625
rect 66904 95659 66956 95668
rect 66904 95625 66913 95659
rect 66913 95625 66947 95659
rect 66947 95625 66956 95659
rect 66904 95616 66956 95625
rect 67732 95616 67784 95668
rect 68836 95659 68888 95668
rect 68836 95625 68845 95659
rect 68845 95625 68879 95659
rect 68879 95625 68888 95659
rect 68836 95616 68888 95625
rect 70308 95616 70360 95668
rect 71688 95616 71740 95668
rect 72424 95659 72476 95668
rect 72424 95625 72433 95659
rect 72433 95625 72467 95659
rect 72467 95625 72476 95659
rect 72424 95616 72476 95625
rect 73528 95616 73580 95668
rect 75000 95659 75052 95668
rect 75000 95625 75009 95659
rect 75009 95625 75043 95659
rect 75043 95625 75052 95659
rect 75000 95616 75052 95625
rect 75552 95659 75604 95668
rect 75552 95625 75561 95659
rect 75561 95625 75595 95659
rect 75595 95625 75604 95659
rect 75552 95616 75604 95625
rect 76932 95659 76984 95668
rect 76932 95625 76941 95659
rect 76941 95625 76975 95659
rect 76975 95625 76984 95659
rect 76932 95616 76984 95625
rect 78220 95659 78272 95668
rect 78220 95625 78229 95659
rect 78229 95625 78263 95659
rect 78263 95625 78272 95659
rect 78220 95616 78272 95625
rect 79508 95659 79560 95668
rect 79508 95625 79517 95659
rect 79517 95625 79551 95659
rect 79551 95625 79560 95659
rect 79508 95616 79560 95625
rect 79968 95616 80020 95668
rect 81348 95616 81400 95668
rect 82728 95659 82780 95668
rect 82728 95625 82737 95659
rect 82737 95625 82771 95659
rect 82771 95625 82780 95659
rect 82728 95616 82780 95625
rect 70308 95523 70360 95532
rect 70308 95489 70317 95523
rect 70317 95489 70351 95523
rect 70351 95489 70360 95523
rect 70308 95480 70360 95489
rect 71228 95480 71280 95532
rect 72240 95523 72292 95532
rect 72240 95489 72249 95523
rect 72249 95489 72283 95523
rect 72283 95489 72292 95523
rect 72240 95480 72292 95489
rect 73528 95523 73580 95532
rect 73528 95489 73537 95523
rect 73537 95489 73571 95523
rect 73571 95489 73580 95523
rect 73528 95480 73580 95489
rect 74816 95523 74868 95532
rect 74816 95489 74825 95523
rect 74825 95489 74859 95523
rect 74859 95489 74868 95523
rect 74816 95480 74868 95489
rect 75736 95523 75788 95532
rect 75736 95489 75745 95523
rect 75745 95489 75779 95523
rect 75779 95489 75788 95523
rect 75736 95480 75788 95489
rect 76748 95523 76800 95532
rect 76748 95489 76757 95523
rect 76757 95489 76791 95523
rect 76791 95489 76800 95523
rect 76748 95480 76800 95489
rect 78036 95523 78088 95532
rect 78036 95489 78045 95523
rect 78045 95489 78079 95523
rect 78079 95489 78088 95523
rect 78036 95480 78088 95489
rect 78956 95480 79008 95532
rect 80060 95480 80112 95532
rect 81256 95523 81308 95532
rect 81256 95489 81265 95523
rect 81265 95489 81299 95523
rect 81299 95489 81308 95523
rect 81256 95480 81308 95489
rect 82544 95523 82596 95532
rect 82544 95489 82553 95523
rect 82553 95489 82587 95523
rect 82587 95489 82596 95523
rect 82544 95480 82596 95489
rect 19064 95412 19116 95464
rect 23572 95455 23624 95464
rect 23572 95421 23581 95455
rect 23581 95421 23615 95455
rect 23615 95421 23624 95455
rect 23572 95412 23624 95421
rect 52368 95412 52420 95464
rect 53748 95455 53800 95464
rect 53748 95421 53757 95455
rect 53757 95421 53791 95455
rect 53791 95421 53800 95455
rect 53748 95412 53800 95421
rect 59084 95412 59136 95464
rect 63500 95412 63552 95464
rect 22652 95387 22704 95396
rect 22652 95353 22661 95387
rect 22661 95353 22695 95387
rect 22695 95353 22704 95387
rect 22652 95344 22704 95353
rect 25872 95387 25924 95396
rect 25872 95353 25881 95387
rect 25881 95353 25915 95387
rect 25915 95353 25924 95387
rect 25872 95344 25924 95353
rect 27160 95387 27212 95396
rect 27160 95353 27169 95387
rect 27169 95353 27203 95387
rect 27203 95353 27212 95387
rect 27160 95344 27212 95353
rect 62580 95387 62632 95396
rect 62580 95353 62589 95387
rect 62589 95353 62623 95387
rect 62623 95353 62632 95387
rect 62580 95344 62632 95353
rect 65800 95387 65852 95396
rect 65800 95353 65809 95387
rect 65809 95353 65843 95387
rect 65843 95353 65852 95387
rect 65800 95344 65852 95353
rect 67088 95387 67140 95396
rect 67088 95353 67097 95387
rect 67097 95353 67131 95387
rect 67131 95353 67140 95387
rect 67088 95344 67140 95353
rect 14648 95276 14700 95328
rect 15752 95319 15804 95328
rect 15752 95285 15761 95319
rect 15761 95285 15795 95319
rect 15795 95285 15804 95319
rect 15752 95276 15804 95285
rect 17040 95319 17092 95328
rect 17040 95285 17049 95319
rect 17049 95285 17083 95319
rect 17083 95285 17092 95319
rect 17040 95276 17092 95285
rect 18328 95319 18380 95328
rect 18328 95285 18337 95319
rect 18337 95285 18371 95319
rect 18371 95285 18380 95319
rect 18328 95276 18380 95285
rect 20168 95319 20220 95328
rect 20168 95285 20177 95319
rect 20177 95285 20211 95319
rect 20211 95285 20220 95319
rect 20168 95276 20220 95285
rect 21548 95319 21600 95328
rect 21548 95285 21557 95319
rect 21557 95285 21591 95319
rect 21591 95285 21600 95319
rect 21548 95276 21600 95285
rect 24768 95319 24820 95328
rect 24768 95285 24777 95319
rect 24777 95285 24811 95319
rect 24811 95285 24820 95319
rect 24768 95276 24820 95285
rect 27988 95319 28040 95328
rect 27988 95285 27997 95319
rect 27997 95285 28031 95319
rect 28031 95285 28040 95319
rect 27988 95276 28040 95285
rect 29092 95319 29144 95328
rect 29092 95285 29101 95319
rect 29101 95285 29135 95319
rect 29135 95285 29144 95319
rect 29092 95276 29144 95285
rect 54668 95276 54720 95328
rect 55956 95276 56008 95328
rect 56876 95319 56928 95328
rect 56876 95285 56885 95319
rect 56885 95285 56919 95319
rect 56919 95285 56928 95319
rect 56876 95276 56928 95285
rect 58256 95319 58308 95328
rect 58256 95285 58265 95319
rect 58265 95285 58299 95319
rect 58299 95285 58308 95319
rect 58256 95276 58308 95285
rect 60188 95319 60240 95328
rect 60188 95285 60197 95319
rect 60197 95285 60231 95319
rect 60231 95285 60240 95319
rect 60188 95276 60240 95285
rect 61476 95319 61528 95328
rect 61476 95285 61485 95319
rect 61485 95285 61519 95319
rect 61519 95285 61528 95319
rect 61476 95276 61528 95285
rect 64604 95276 64656 95328
rect 67916 95319 67968 95328
rect 67916 95285 67925 95319
rect 67925 95285 67959 95319
rect 67959 95285 67968 95319
rect 67916 95276 67968 95285
rect 69020 95319 69072 95328
rect 69020 95285 69029 95319
rect 69029 95285 69063 95319
rect 69063 95285 69072 95319
rect 69020 95276 69072 95285
rect 36950 95174 37002 95226
rect 37014 95174 37066 95226
rect 37078 95174 37130 95226
rect 37142 95174 37194 95226
rect 37206 95174 37258 95226
rect 72950 95174 73002 95226
rect 73014 95174 73066 95226
rect 73078 95174 73130 95226
rect 73142 95174 73194 95226
rect 73206 95174 73258 95226
rect 52276 95072 52328 95124
rect 37610 94630 37662 94682
rect 37674 94630 37726 94682
rect 37738 94630 37790 94682
rect 37802 94630 37854 94682
rect 37866 94630 37918 94682
rect 73610 94630 73662 94682
rect 73674 94630 73726 94682
rect 73738 94630 73790 94682
rect 73802 94630 73854 94682
rect 73866 94630 73918 94682
rect 88156 94188 88208 94240
rect 36950 94086 37002 94138
rect 37014 94086 37066 94138
rect 37078 94086 37130 94138
rect 37142 94086 37194 94138
rect 37206 94086 37258 94138
rect 72950 94086 73002 94138
rect 73014 94086 73066 94138
rect 73078 94086 73130 94138
rect 73142 94086 73194 94138
rect 73206 94086 73258 94138
rect 88616 93916 88668 93968
rect 88340 93891 88392 93900
rect 88340 93857 88349 93891
rect 88349 93857 88383 93891
rect 88383 93857 88392 93891
rect 88340 93848 88392 93857
rect 88524 93891 88576 93900
rect 88524 93857 88533 93891
rect 88533 93857 88567 93891
rect 88567 93857 88576 93891
rect 88524 93848 88576 93857
rect 88064 93687 88116 93696
rect 88064 93653 88073 93687
rect 88073 93653 88107 93687
rect 88107 93653 88116 93687
rect 88064 93644 88116 93653
rect 37610 93542 37662 93594
rect 37674 93542 37726 93594
rect 37738 93542 37790 93594
rect 37802 93542 37854 93594
rect 37866 93542 37918 93594
rect 73610 93542 73662 93594
rect 73674 93542 73726 93594
rect 73738 93542 73790 93594
rect 73802 93542 73854 93594
rect 73866 93542 73918 93594
rect 87788 93168 87840 93220
rect 88524 93168 88576 93220
rect 87236 93100 87288 93152
rect 87696 93143 87748 93152
rect 87696 93109 87705 93143
rect 87705 93109 87739 93143
rect 87739 93109 87748 93143
rect 87696 93100 87748 93109
rect 87880 93143 87932 93152
rect 87880 93109 87889 93143
rect 87889 93109 87923 93143
rect 87923 93109 87932 93143
rect 87880 93100 87932 93109
rect 88800 93100 88852 93152
rect 36950 92998 37002 93050
rect 37014 92998 37066 93050
rect 37078 92998 37130 93050
rect 37142 92998 37194 93050
rect 37206 92998 37258 93050
rect 72950 92998 73002 93050
rect 73014 92998 73066 93050
rect 73078 92998 73130 93050
rect 73142 92998 73194 93050
rect 73206 92998 73258 93050
rect 83372 92896 83424 92948
rect 86408 92828 86460 92880
rect 86776 92803 86828 92812
rect 86776 92769 86785 92803
rect 86785 92769 86819 92803
rect 86819 92769 86828 92803
rect 86776 92760 86828 92769
rect 87328 92692 87380 92744
rect 87144 92667 87196 92676
rect 87144 92633 87153 92667
rect 87153 92633 87187 92667
rect 87187 92633 87196 92667
rect 87144 92624 87196 92633
rect 87604 92624 87656 92676
rect 87972 92735 88024 92744
rect 87972 92701 87981 92735
rect 87981 92701 88015 92735
rect 88015 92701 88024 92735
rect 87972 92692 88024 92701
rect 88064 92624 88116 92676
rect 89352 92624 89404 92676
rect 86592 92599 86644 92608
rect 86592 92565 86601 92599
rect 86601 92565 86635 92599
rect 86635 92565 86644 92599
rect 86592 92556 86644 92565
rect 87052 92599 87104 92608
rect 87052 92565 87061 92599
rect 87061 92565 87095 92599
rect 87095 92565 87104 92599
rect 87052 92556 87104 92565
rect 87512 92556 87564 92608
rect 88156 92599 88208 92608
rect 88156 92565 88165 92599
rect 88165 92565 88199 92599
rect 88199 92565 88208 92599
rect 88156 92556 88208 92565
rect 88432 92599 88484 92608
rect 88432 92565 88441 92599
rect 88441 92565 88475 92599
rect 88475 92565 88484 92599
rect 88432 92556 88484 92565
rect 37610 92454 37662 92506
rect 37674 92454 37726 92506
rect 37738 92454 37790 92506
rect 37802 92454 37854 92506
rect 37866 92454 37918 92506
rect 73610 92454 73662 92506
rect 73674 92454 73726 92506
rect 73738 92454 73790 92506
rect 73802 92454 73854 92506
rect 73866 92454 73918 92506
rect 47492 92216 47544 92268
rect 87236 92259 87288 92268
rect 87236 92225 87245 92259
rect 87245 92225 87279 92259
rect 87279 92225 87288 92259
rect 87236 92216 87288 92225
rect 87696 92352 87748 92404
rect 89260 92352 89312 92404
rect 88708 92284 88760 92336
rect 87788 92259 87840 92268
rect 87788 92225 87797 92259
rect 87797 92225 87831 92259
rect 87831 92225 87840 92259
rect 87788 92216 87840 92225
rect 47400 92148 47452 92200
rect 52460 92148 52512 92200
rect 86224 92191 86276 92200
rect 86224 92157 86233 92191
rect 86233 92157 86267 92191
rect 86267 92157 86276 92191
rect 86224 92148 86276 92157
rect 86316 92148 86368 92200
rect 89536 92216 89588 92268
rect 32404 92123 32456 92132
rect 32404 92089 32413 92123
rect 32413 92089 32447 92123
rect 32447 92089 32456 92123
rect 32404 92080 32456 92089
rect 51080 92080 51132 92132
rect 52368 92080 52420 92132
rect 87512 92080 87564 92132
rect 30472 92055 30524 92064
rect 30472 92021 30481 92055
rect 30481 92021 30515 92055
rect 30515 92021 30524 92055
rect 30472 92012 30524 92021
rect 50252 92012 50304 92064
rect 52644 92012 52696 92064
rect 85672 92055 85724 92064
rect 85672 92021 85681 92055
rect 85681 92021 85715 92055
rect 85715 92021 85724 92055
rect 85672 92012 85724 92021
rect 85948 92055 86000 92064
rect 85948 92021 85957 92055
rect 85957 92021 85991 92055
rect 85991 92021 86000 92055
rect 85948 92012 86000 92021
rect 86040 92055 86092 92064
rect 86040 92021 86049 92055
rect 86049 92021 86083 92055
rect 86083 92021 86092 92055
rect 86040 92012 86092 92021
rect 86500 92055 86552 92064
rect 86500 92021 86509 92055
rect 86509 92021 86543 92055
rect 86543 92021 86552 92055
rect 86500 92012 86552 92021
rect 86684 92055 86736 92064
rect 86684 92021 86693 92055
rect 86693 92021 86727 92055
rect 86727 92021 86736 92055
rect 86684 92012 86736 92021
rect 86776 92055 86828 92064
rect 86776 92021 86785 92055
rect 86785 92021 86819 92055
rect 86819 92021 86828 92055
rect 86776 92012 86828 92021
rect 87052 92055 87104 92064
rect 87052 92021 87061 92055
rect 87061 92021 87095 92055
rect 87095 92021 87104 92055
rect 87052 92012 87104 92021
rect 87420 92012 87472 92064
rect 88340 92148 88392 92200
rect 88708 92148 88760 92200
rect 87696 92080 87748 92132
rect 88064 92080 88116 92132
rect 88800 92012 88852 92064
rect 3066 91910 3118 91962
rect 3130 91910 3182 91962
rect 3194 91910 3246 91962
rect 3258 91910 3310 91962
rect 3322 91910 3374 91962
rect 36950 91910 37002 91962
rect 37014 91910 37066 91962
rect 37078 91910 37130 91962
rect 37142 91910 37194 91962
rect 37206 91910 37258 91962
rect 72950 91910 73002 91962
rect 73014 91910 73066 91962
rect 73078 91910 73130 91962
rect 73142 91910 73194 91962
rect 73206 91910 73258 91962
rect 50252 91851 50304 91860
rect 50252 91817 50261 91851
rect 50261 91817 50295 91851
rect 50295 91817 50304 91851
rect 50252 91808 50304 91817
rect 86316 91808 86368 91860
rect 87236 91808 87288 91860
rect 89168 91808 89220 91860
rect 88340 91740 88392 91792
rect 5632 91536 5684 91588
rect 10324 91579 10376 91588
rect 10324 91545 10333 91579
rect 10333 91545 10367 91579
rect 10367 91545 10376 91579
rect 47952 91672 48004 91724
rect 86040 91672 86092 91724
rect 32404 91604 32456 91656
rect 10324 91536 10376 91545
rect 11612 91511 11664 91520
rect 11612 91477 11621 91511
rect 11621 91477 11655 91511
rect 11655 91477 11664 91511
rect 11612 91468 11664 91477
rect 12532 91511 12584 91520
rect 12532 91477 12541 91511
rect 12541 91477 12575 91511
rect 12575 91477 12584 91511
rect 12532 91468 12584 91477
rect 13544 91511 13596 91520
rect 13544 91477 13553 91511
rect 13553 91477 13587 91511
rect 13587 91477 13596 91511
rect 13544 91468 13596 91477
rect 43444 91536 43496 91588
rect 47768 91536 47820 91588
rect 52736 91647 52788 91656
rect 52736 91613 52745 91647
rect 52745 91613 52779 91647
rect 52779 91613 52788 91647
rect 52736 91604 52788 91613
rect 53748 91604 53800 91656
rect 84476 91604 84528 91656
rect 52460 91536 52512 91588
rect 53840 91579 53892 91588
rect 53840 91545 53849 91579
rect 53849 91545 53883 91579
rect 53883 91545 53892 91579
rect 53840 91536 53892 91545
rect 85212 91579 85264 91588
rect 85212 91545 85221 91579
rect 85221 91545 85255 91579
rect 85255 91545 85264 91579
rect 85212 91536 85264 91545
rect 85856 91604 85908 91656
rect 87604 91672 87656 91724
rect 89076 91672 89128 91724
rect 88524 91604 88576 91656
rect 88984 91604 89036 91656
rect 87144 91579 87196 91588
rect 87144 91545 87153 91579
rect 87153 91545 87187 91579
rect 87187 91545 87196 91579
rect 87144 91536 87196 91545
rect 87328 91579 87380 91588
rect 87328 91545 87337 91579
rect 87337 91545 87371 91579
rect 87371 91545 87380 91579
rect 87328 91536 87380 91545
rect 87512 91579 87564 91588
rect 87512 91545 87521 91579
rect 87521 91545 87555 91579
rect 87555 91545 87564 91579
rect 87512 91536 87564 91545
rect 87880 91536 87932 91588
rect 30472 91468 30524 91520
rect 47676 91468 47728 91520
rect 51080 91511 51132 91520
rect 51080 91477 51089 91511
rect 51089 91477 51123 91511
rect 51123 91477 51132 91511
rect 51080 91468 51132 91477
rect 53748 91468 53800 91520
rect 85028 91511 85080 91520
rect 85028 91477 85037 91511
rect 85037 91477 85071 91511
rect 85071 91477 85080 91511
rect 85028 91468 85080 91477
rect 85396 91511 85448 91520
rect 85396 91477 85405 91511
rect 85405 91477 85439 91511
rect 85439 91477 85448 91511
rect 85396 91468 85448 91477
rect 85764 91511 85816 91520
rect 85764 91477 85773 91511
rect 85773 91477 85807 91511
rect 85807 91477 85816 91511
rect 85764 91468 85816 91477
rect 86316 91511 86368 91520
rect 86316 91477 86325 91511
rect 86325 91477 86359 91511
rect 86359 91477 86368 91511
rect 86316 91468 86368 91477
rect 86684 91468 86736 91520
rect 87972 91511 88024 91520
rect 87972 91477 87981 91511
rect 87981 91477 88015 91511
rect 88015 91477 88024 91511
rect 87972 91468 88024 91477
rect 88248 91579 88300 91588
rect 88248 91545 88257 91579
rect 88257 91545 88291 91579
rect 88291 91545 88300 91579
rect 88248 91536 88300 91545
rect 88616 91536 88668 91588
rect 89444 91536 89496 91588
rect 88524 91468 88576 91520
rect 3802 91366 3854 91418
rect 3866 91366 3918 91418
rect 3930 91366 3982 91418
rect 3994 91366 4046 91418
rect 4058 91366 4110 91418
rect 37610 91366 37662 91418
rect 37674 91366 37726 91418
rect 37738 91366 37790 91418
rect 37802 91366 37854 91418
rect 37866 91366 37918 91418
rect 73610 91366 73662 91418
rect 73674 91366 73726 91418
rect 73738 91366 73790 91418
rect 73802 91366 73854 91418
rect 73866 91366 73918 91418
rect 12532 91264 12584 91316
rect 52736 91264 52788 91316
rect 11612 91196 11664 91248
rect 51080 91196 51132 91248
rect 47860 91128 47912 91180
rect 85396 91128 85448 91180
rect 48136 91060 48188 91112
rect 85764 91060 85816 91112
rect 48228 90992 48280 91044
rect 52460 90992 52512 91044
rect 48044 90924 48096 90976
rect 53840 90924 53892 90976
rect 3066 90822 3118 90874
rect 3130 90822 3182 90874
rect 3194 90822 3246 90874
rect 3258 90822 3310 90874
rect 3322 90822 3374 90874
rect 3802 90278 3854 90330
rect 3866 90278 3918 90330
rect 3930 90278 3982 90330
rect 3994 90278 4046 90330
rect 4058 90278 4110 90330
rect 3066 89734 3118 89786
rect 3130 89734 3182 89786
rect 3194 89734 3246 89786
rect 3258 89734 3310 89786
rect 3322 89734 3374 89786
rect 47308 89632 47360 89684
rect 85028 89632 85080 89684
rect 5172 89292 5224 89344
rect 85672 89292 85724 89344
rect 3802 89190 3854 89242
rect 3866 89190 3918 89242
rect 3930 89190 3982 89242
rect 3994 89190 4046 89242
rect 4058 89190 4110 89242
rect 5356 89088 5408 89140
rect 86500 89088 86552 89140
rect 5448 89020 5500 89072
rect 86040 89020 86092 89072
rect 5080 88952 5132 89004
rect 86316 88952 86368 89004
rect 3066 88646 3118 88698
rect 3130 88646 3182 88698
rect 3194 88646 3246 88698
rect 3258 88646 3310 88698
rect 3322 88646 3374 88698
rect 6736 88476 6788 88528
rect 53196 88476 53248 88528
rect 86316 88476 86368 88528
rect 88616 88476 88668 88528
rect 13728 88408 13780 88460
rect 47584 88408 47636 88460
rect 85672 88408 85724 88460
rect 86868 88408 86920 88460
rect 5264 88340 5316 88392
rect 47308 88340 47360 88392
rect 3802 88102 3854 88154
rect 3866 88102 3918 88154
rect 3930 88102 3982 88154
rect 3994 88102 4046 88154
rect 4058 88102 4110 88154
rect 3066 87558 3118 87610
rect 3130 87558 3182 87610
rect 3194 87558 3246 87610
rect 3258 87558 3310 87610
rect 3322 87558 3374 87610
rect 3802 87014 3854 87066
rect 3866 87014 3918 87066
rect 3930 87014 3982 87066
rect 3994 87014 4046 87066
rect 4058 87014 4110 87066
rect 8300 86776 8352 86828
rect 848 86572 900 86624
rect 3066 86470 3118 86522
rect 3130 86470 3182 86522
rect 3194 86470 3246 86522
rect 3258 86470 3310 86522
rect 3322 86470 3374 86522
rect 3802 85926 3854 85978
rect 3866 85926 3918 85978
rect 3930 85926 3982 85978
rect 3994 85926 4046 85978
rect 4058 85926 4110 85978
rect 3066 85382 3118 85434
rect 3130 85382 3182 85434
rect 3194 85382 3246 85434
rect 3258 85382 3310 85434
rect 3322 85382 3374 85434
rect 848 85212 900 85264
rect 8300 85076 8352 85128
rect 3802 84838 3854 84890
rect 3866 84838 3918 84890
rect 3930 84838 3982 84890
rect 3994 84838 4046 84890
rect 4058 84838 4110 84890
rect 3066 84294 3118 84346
rect 3130 84294 3182 84346
rect 3194 84294 3246 84346
rect 3258 84294 3310 84346
rect 3322 84294 3374 84346
rect 8300 83988 8352 84040
rect 848 83852 900 83904
rect 3802 83750 3854 83802
rect 3866 83750 3918 83802
rect 3930 83750 3982 83802
rect 3994 83750 4046 83802
rect 4058 83750 4110 83802
rect 3066 83206 3118 83258
rect 3130 83206 3182 83258
rect 3194 83206 3246 83258
rect 3258 83206 3310 83258
rect 3322 83206 3374 83258
rect 3802 82662 3854 82714
rect 3866 82662 3918 82714
rect 3930 82662 3982 82714
rect 3994 82662 4046 82714
rect 4058 82662 4110 82714
rect 8300 82424 8352 82476
rect 848 82220 900 82272
rect 3066 82118 3118 82170
rect 3130 82118 3182 82170
rect 3194 82118 3246 82170
rect 3258 82118 3310 82170
rect 3322 82118 3374 82170
rect 88432 81744 88484 81796
rect 88800 81744 88852 81796
rect 3802 81574 3854 81626
rect 3866 81574 3918 81626
rect 3930 81574 3982 81626
rect 3994 81574 4046 81626
rect 4058 81574 4110 81626
rect 8300 81336 8352 81388
rect 848 81132 900 81184
rect 3066 81030 3118 81082
rect 3130 81030 3182 81082
rect 3194 81030 3246 81082
rect 3258 81030 3310 81082
rect 3322 81030 3374 81082
rect 3802 80486 3854 80538
rect 3866 80486 3918 80538
rect 3930 80486 3982 80538
rect 3994 80486 4046 80538
rect 4058 80486 4110 80538
rect 3066 79942 3118 79994
rect 3130 79942 3182 79994
rect 3194 79942 3246 79994
rect 3258 79942 3310 79994
rect 3322 79942 3374 79994
rect 8300 79636 8352 79688
rect 848 79500 900 79552
rect 3802 79398 3854 79450
rect 3866 79398 3918 79450
rect 3930 79398 3982 79450
rect 3994 79398 4046 79450
rect 4058 79398 4110 79450
rect 3066 78854 3118 78906
rect 3130 78854 3182 78906
rect 3194 78854 3246 78906
rect 3258 78854 3310 78906
rect 3322 78854 3374 78906
rect 8300 78548 8352 78600
rect 848 78412 900 78464
rect 3802 78310 3854 78362
rect 3866 78310 3918 78362
rect 3930 78310 3982 78362
rect 3994 78310 4046 78362
rect 4058 78310 4110 78362
rect 3066 77766 3118 77818
rect 3130 77766 3182 77818
rect 3194 77766 3246 77818
rect 3258 77766 3310 77818
rect 3322 77766 3374 77818
rect 3802 77222 3854 77274
rect 3866 77222 3918 77274
rect 3930 77222 3982 77274
rect 3994 77222 4046 77274
rect 4058 77222 4110 77274
rect 89168 77052 89220 77104
rect 89352 77052 89404 77104
rect 8300 76984 8352 77036
rect 848 76780 900 76832
rect 3066 76678 3118 76730
rect 3130 76678 3182 76730
rect 3194 76678 3246 76730
rect 3258 76678 3310 76730
rect 3322 76678 3374 76730
rect 3802 76134 3854 76186
rect 3866 76134 3918 76186
rect 3930 76134 3982 76186
rect 3994 76134 4046 76186
rect 4058 76134 4110 76186
rect 848 76032 900 76084
rect 5540 75896 5592 75948
rect 3066 75590 3118 75642
rect 3130 75590 3182 75642
rect 3194 75590 3246 75642
rect 3258 75590 3310 75642
rect 3322 75590 3374 75642
rect 3802 75046 3854 75098
rect 3866 75046 3918 75098
rect 3930 75046 3982 75098
rect 3994 75046 4046 75098
rect 4058 75046 4110 75098
rect 3066 74502 3118 74554
rect 3130 74502 3182 74554
rect 3194 74502 3246 74554
rect 3258 74502 3310 74554
rect 3322 74502 3374 74554
rect 8300 74196 8352 74248
rect 848 74060 900 74112
rect 3802 73958 3854 74010
rect 3866 73958 3918 74010
rect 3930 73958 3982 74010
rect 3994 73958 4046 74010
rect 4058 73958 4110 74010
rect 3066 73414 3118 73466
rect 3130 73414 3182 73466
rect 3194 73414 3246 73466
rect 3258 73414 3310 73466
rect 3322 73414 3374 73466
rect 8300 73108 8352 73160
rect 848 72972 900 73024
rect 3802 72870 3854 72922
rect 3866 72870 3918 72922
rect 3930 72870 3982 72922
rect 3994 72870 4046 72922
rect 4058 72870 4110 72922
rect 3066 72326 3118 72378
rect 3130 72326 3182 72378
rect 3194 72326 3246 72378
rect 3258 72326 3310 72378
rect 3322 72326 3374 72378
rect 3802 71782 3854 71834
rect 3866 71782 3918 71834
rect 3930 71782 3982 71834
rect 3994 71782 4046 71834
rect 4058 71782 4110 71834
rect 8300 71612 8352 71664
rect 5908 71544 5960 71596
rect 4620 71408 4672 71460
rect 848 71340 900 71392
rect 3066 71238 3118 71290
rect 3130 71238 3182 71290
rect 3194 71238 3246 71290
rect 3258 71238 3310 71290
rect 3322 71238 3374 71290
rect 3802 70694 3854 70746
rect 3866 70694 3918 70746
rect 3930 70694 3982 70746
rect 3994 70694 4046 70746
rect 4058 70694 4110 70746
rect 848 70592 900 70644
rect 5080 70592 5132 70644
rect 5540 70456 5592 70508
rect 5816 70456 5868 70508
rect 3066 70150 3118 70202
rect 3130 70150 3182 70202
rect 3194 70150 3246 70202
rect 3258 70150 3310 70202
rect 3322 70150 3374 70202
rect 3802 69606 3854 69658
rect 3866 69606 3918 69658
rect 3930 69606 3982 69658
rect 3994 69606 4046 69658
rect 4058 69606 4110 69658
rect 3066 69062 3118 69114
rect 3130 69062 3182 69114
rect 3194 69062 3246 69114
rect 3258 69062 3310 69114
rect 3322 69062 3374 69114
rect 8300 68892 8352 68944
rect 1216 68756 1268 68808
rect 6184 68688 6236 68740
rect 6092 68620 6144 68672
rect 3802 68518 3854 68570
rect 3866 68518 3918 68570
rect 3930 68518 3982 68570
rect 3994 68518 4046 68570
rect 4058 68518 4110 68570
rect 3066 67974 3118 68026
rect 3130 67974 3182 68026
rect 3194 67974 3246 68026
rect 3258 67974 3310 68026
rect 3322 67974 3374 68026
rect 5724 67872 5776 67924
rect 1308 67668 1360 67720
rect 5448 67804 5500 67856
rect 5540 67847 5592 67856
rect 5540 67813 5549 67847
rect 5549 67813 5583 67847
rect 5583 67813 5592 67847
rect 5540 67804 5592 67813
rect 3802 67430 3854 67482
rect 3866 67430 3918 67482
rect 3930 67430 3982 67482
rect 3994 67430 4046 67482
rect 4058 67430 4110 67482
rect 3066 66886 3118 66938
rect 3130 66886 3182 66938
rect 3194 66886 3246 66938
rect 3258 66886 3310 66938
rect 3322 66886 3374 66938
rect 3802 66342 3854 66394
rect 3866 66342 3918 66394
rect 3930 66342 3982 66394
rect 3994 66342 4046 66394
rect 4058 66342 4110 66394
rect 1308 66104 1360 66156
rect 4896 66104 4948 66156
rect 8300 65968 8352 66020
rect 4896 65900 4948 65952
rect 7564 65900 7616 65952
rect 3066 65798 3118 65850
rect 3130 65798 3182 65850
rect 3194 65798 3246 65850
rect 3258 65798 3310 65850
rect 3322 65798 3374 65850
rect 3802 65254 3854 65306
rect 3866 65254 3918 65306
rect 3930 65254 3982 65306
rect 3994 65254 4046 65306
rect 4058 65254 4110 65306
rect 5356 65152 5408 65204
rect 1308 65016 1360 65068
rect 5908 64948 5960 65000
rect 5540 64923 5592 64932
rect 5540 64889 5549 64923
rect 5549 64889 5583 64923
rect 5583 64889 5592 64923
rect 5540 64880 5592 64889
rect 3066 64710 3118 64762
rect 3130 64710 3182 64762
rect 3194 64710 3246 64762
rect 3258 64710 3310 64762
rect 3322 64710 3374 64762
rect 3802 64166 3854 64218
rect 3866 64166 3918 64218
rect 3930 64166 3982 64218
rect 3994 64166 4046 64218
rect 4058 64166 4110 64218
rect 3066 63622 3118 63674
rect 3130 63622 3182 63674
rect 3194 63622 3246 63674
rect 3258 63622 3310 63674
rect 3322 63622 3374 63674
rect 8300 63452 8352 63504
rect 1216 63316 1268 63368
rect 4528 63180 4580 63232
rect 7656 63180 7708 63232
rect 3802 63078 3854 63130
rect 3866 63078 3918 63130
rect 3930 63078 3982 63130
rect 3994 63078 4046 63130
rect 4058 63078 4110 63130
rect 3066 62534 3118 62586
rect 3130 62534 3182 62586
rect 3194 62534 3246 62586
rect 3258 62534 3310 62586
rect 3322 62534 3374 62586
rect 5264 62475 5316 62484
rect 5264 62441 5273 62475
rect 5273 62441 5307 62475
rect 5307 62441 5316 62475
rect 5264 62432 5316 62441
rect 5540 62364 5592 62416
rect 1308 62228 1360 62280
rect 5264 62228 5316 62280
rect 5908 62092 5960 62144
rect 3802 61990 3854 62042
rect 3866 61990 3918 62042
rect 3930 61990 3982 62042
rect 3994 61990 4046 62042
rect 4058 61990 4110 62042
rect 1308 61752 1360 61804
rect 8300 61616 8352 61668
rect 3066 61446 3118 61498
rect 3130 61446 3182 61498
rect 3194 61446 3246 61498
rect 3258 61446 3310 61498
rect 3322 61446 3374 61498
rect 3802 60902 3854 60954
rect 3866 60902 3918 60954
rect 3930 60902 3982 60954
rect 3994 60902 4046 60954
rect 4058 60902 4110 60954
rect 5172 60707 5224 60716
rect 5172 60673 5181 60707
rect 5181 60673 5215 60707
rect 5215 60673 5224 60707
rect 5172 60664 5224 60673
rect 848 60460 900 60512
rect 7840 60460 7892 60512
rect 3066 60358 3118 60410
rect 3130 60358 3182 60410
rect 3194 60358 3246 60410
rect 3258 60358 3310 60410
rect 3322 60358 3374 60410
rect 1216 60052 1268 60104
rect 8300 59984 8352 60036
rect 3802 59814 3854 59866
rect 3866 59814 3918 59866
rect 3930 59814 3982 59866
rect 3994 59814 4046 59866
rect 4058 59814 4110 59866
rect 5264 59576 5316 59628
rect 848 59372 900 59424
rect 5264 59415 5316 59424
rect 5264 59381 5273 59415
rect 5273 59381 5307 59415
rect 5307 59381 5316 59415
rect 5264 59372 5316 59381
rect 5908 59372 5960 59424
rect 3066 59270 3118 59322
rect 3130 59270 3182 59322
rect 3194 59270 3246 59322
rect 3258 59270 3310 59322
rect 3322 59270 3374 59322
rect 8300 59100 8352 59152
rect 1308 58964 1360 59016
rect 3802 58726 3854 58778
rect 3866 58726 3918 58778
rect 3930 58726 3982 58778
rect 3994 58726 4046 58778
rect 4058 58726 4110 58778
rect 3066 58182 3118 58234
rect 3130 58182 3182 58234
rect 3194 58182 3246 58234
rect 3258 58182 3310 58234
rect 3322 58182 3374 58234
rect 848 57944 900 57996
rect 5448 57740 5500 57792
rect 7196 57740 7248 57792
rect 3802 57638 3854 57690
rect 3866 57638 3918 57690
rect 3930 57638 3982 57690
rect 3994 57638 4046 57690
rect 4058 57638 4110 57690
rect 5632 57536 5684 57588
rect 1308 57400 1360 57452
rect 8300 57264 8352 57316
rect 5540 57239 5592 57248
rect 5540 57205 5549 57239
rect 5549 57205 5583 57239
rect 5583 57205 5592 57239
rect 5540 57196 5592 57205
rect 3066 57094 3118 57146
rect 3130 57094 3182 57146
rect 3194 57094 3246 57146
rect 3258 57094 3310 57146
rect 3322 57094 3374 57146
rect 848 56788 900 56840
rect 5632 56831 5684 56840
rect 5632 56797 5641 56831
rect 5641 56797 5675 56831
rect 5675 56797 5684 56831
rect 5632 56788 5684 56797
rect 5540 56652 5592 56704
rect 3802 56550 3854 56602
rect 3866 56550 3918 56602
rect 3930 56550 3982 56602
rect 3994 56550 4046 56602
rect 4058 56550 4110 56602
rect 1308 56312 1360 56364
rect 5080 56312 5132 56364
rect 8300 56176 8352 56228
rect 5080 56108 5132 56160
rect 6736 56108 6788 56160
rect 3066 56006 3118 56058
rect 3130 56006 3182 56058
rect 3194 56006 3246 56058
rect 3258 56006 3310 56058
rect 3322 56006 3374 56058
rect 3802 55462 3854 55514
rect 3866 55462 3918 55514
rect 3930 55462 3982 55514
rect 3994 55462 4046 55514
rect 4058 55462 4110 55514
rect 4896 55360 4948 55412
rect 6828 55360 6880 55412
rect 848 55020 900 55072
rect 3066 54918 3118 54970
rect 3130 54918 3182 54970
rect 3194 54918 3246 54970
rect 3258 54918 3310 54970
rect 3322 54918 3374 54970
rect 1216 54612 1268 54664
rect 8300 54544 8352 54596
rect 3802 54374 3854 54426
rect 3866 54374 3918 54426
rect 3930 54374 3982 54426
rect 3994 54374 4046 54426
rect 4058 54374 4110 54426
rect 4712 54272 4764 54324
rect 4896 54272 4948 54324
rect 848 53932 900 53984
rect 5080 53932 5132 53984
rect 7932 53932 7984 53984
rect 3066 53830 3118 53882
rect 3130 53830 3182 53882
rect 3194 53830 3246 53882
rect 3258 53830 3310 53882
rect 3322 53830 3374 53882
rect 8300 53660 8352 53712
rect 1308 53524 1360 53576
rect 3802 53286 3854 53338
rect 3866 53286 3918 53338
rect 3930 53286 3982 53338
rect 3994 53286 4046 53338
rect 4058 53286 4110 53338
rect 3066 52742 3118 52794
rect 3130 52742 3182 52794
rect 3194 52742 3246 52794
rect 3258 52742 3310 52794
rect 3322 52742 3374 52794
rect 8208 52572 8260 52624
rect 848 52436 900 52488
rect 5172 52479 5224 52488
rect 5172 52445 5181 52479
rect 5181 52445 5215 52479
rect 5215 52445 5224 52479
rect 5172 52436 5224 52445
rect 3802 52198 3854 52250
rect 3866 52198 3918 52250
rect 3930 52198 3982 52250
rect 3994 52198 4046 52250
rect 4058 52198 4110 52250
rect 848 51892 900 51944
rect 3066 51654 3118 51706
rect 3130 51654 3182 51706
rect 3194 51654 3246 51706
rect 3258 51654 3310 51706
rect 3322 51654 3374 51706
rect 1032 51348 1084 51400
rect 5264 51255 5316 51264
rect 5264 51221 5273 51255
rect 5273 51221 5307 51255
rect 5307 51221 5316 51255
rect 5264 51212 5316 51221
rect 3802 51110 3854 51162
rect 3866 51110 3918 51162
rect 3930 51110 3982 51162
rect 3994 51110 4046 51162
rect 4058 51110 4110 51162
rect 87144 51008 87196 51060
rect 6552 50940 6604 50992
rect 6736 50940 6788 50992
rect 7564 50940 7616 50992
rect 89076 50940 89128 50992
rect 5356 50915 5408 50924
rect 5356 50881 5365 50915
rect 5365 50881 5399 50915
rect 5399 50881 5408 50915
rect 5356 50872 5408 50881
rect 5632 50804 5684 50856
rect 7932 50804 7984 50856
rect 88340 50804 88392 50856
rect 6644 50736 6696 50788
rect 1400 50711 1452 50720
rect 1400 50677 1409 50711
rect 1409 50677 1443 50711
rect 1443 50677 1452 50711
rect 1400 50668 1452 50677
rect 6736 50668 6788 50720
rect 3066 50566 3118 50618
rect 3130 50566 3182 50618
rect 3194 50566 3246 50618
rect 3258 50566 3310 50618
rect 3322 50566 3374 50618
rect 6644 50600 6696 50652
rect 9588 50600 9640 50652
rect 46848 50600 46900 50652
rect 85580 50600 85632 50652
rect 8208 50532 8260 50584
rect 88432 50532 88484 50584
rect 5632 50464 5684 50516
rect 6644 50464 6696 50516
rect 11612 50464 11664 50516
rect 8208 50260 8260 50312
rect 13084 50260 13136 50312
rect 47492 50396 47544 50448
rect 52644 50396 52696 50448
rect 12256 50192 12308 50244
rect 47400 50192 47452 50244
rect 51540 50192 51592 50244
rect 8024 50124 8076 50176
rect 10876 50124 10928 50176
rect 47768 50124 47820 50176
rect 50436 50124 50488 50176
rect 3802 50022 3854 50074
rect 3866 50022 3918 50074
rect 3930 50022 3982 50074
rect 3994 50022 4046 50074
rect 4058 50022 4110 50074
rect 8024 49920 8076 49972
rect 10508 49920 10560 49972
rect 4620 49852 4672 49904
rect 86684 49852 86736 49904
rect 6460 49784 6512 49836
rect 6092 49716 6144 49768
rect 9680 49716 9732 49768
rect 46848 49784 46900 49836
rect 47676 49784 47728 49836
rect 49700 49784 49752 49836
rect 86868 49716 86920 49768
rect 5816 49648 5868 49700
rect 89168 49648 89220 49700
rect 1400 49623 1452 49632
rect 1400 49589 1409 49623
rect 1409 49589 1443 49623
rect 1443 49589 1452 49623
rect 1400 49580 1452 49589
rect 6828 49580 6880 49632
rect 88524 49580 88576 49632
rect 3066 49478 3118 49530
rect 3130 49478 3182 49530
rect 3194 49478 3246 49530
rect 3258 49478 3310 49530
rect 3322 49478 3374 49530
rect 47768 49444 47820 49496
rect 48228 49444 48280 49496
rect 4896 49376 4948 49428
rect 87420 49376 87472 49428
rect 1400 49351 1452 49360
rect 1400 49317 1409 49351
rect 1409 49317 1443 49351
rect 1443 49317 1452 49351
rect 1400 49308 1452 49317
rect 7656 49308 7708 49360
rect 88892 49308 88944 49360
rect 7840 49240 7892 49292
rect 88800 49240 88852 49292
rect 7196 49172 7248 49224
rect 88616 49172 88668 49224
rect 5264 49104 5316 49156
rect 48136 49104 48188 49156
rect 87144 49104 87196 49156
rect 5172 49036 5224 49088
rect 47952 49036 48004 49088
rect 48228 49036 48280 49088
rect 3802 48934 3854 48986
rect 3866 48934 3918 48986
rect 3930 48934 3982 48986
rect 3994 48934 4046 48986
rect 4058 48934 4110 48986
rect 1584 48875 1636 48884
rect 1584 48841 1593 48875
rect 1593 48841 1627 48875
rect 1627 48841 1636 48875
rect 1584 48832 1636 48841
rect 5356 48832 5408 48884
rect 46848 48832 46900 48884
rect 5908 48764 5960 48816
rect 87788 48764 87840 48816
rect 1308 48696 1360 48748
rect 6552 48696 6604 48748
rect 88708 48696 88760 48748
rect 6184 48628 6236 48680
rect 89352 48628 89404 48680
rect 5172 48560 5224 48612
rect 89076 48560 89128 48612
rect 47952 48492 48004 48544
rect 87328 48492 87380 48544
rect 3066 48390 3118 48442
rect 3130 48390 3182 48442
rect 3194 48390 3246 48442
rect 3258 48390 3310 48442
rect 3322 48390 3374 48442
rect 7012 48424 7064 48476
rect 86684 48424 86736 48476
rect 5724 48220 5776 48272
rect 89260 48220 89312 48272
rect 6276 48152 6328 48204
rect 86776 48152 86828 48204
rect 1400 48127 1452 48136
rect 1400 48093 1409 48127
rect 1409 48093 1443 48127
rect 1443 48093 1452 48127
rect 1400 48084 1452 48093
rect 9680 48084 9732 48136
rect 88984 48084 89036 48136
rect 6736 48016 6788 48068
rect 46756 48016 46808 48068
rect 3802 47846 3854 47898
rect 3866 47846 3918 47898
rect 3930 47846 3982 47898
rect 3994 47846 4046 47898
rect 4058 47846 4110 47898
rect 5632 47676 5684 47728
rect 51172 47676 51224 47728
rect 5080 47608 5132 47660
rect 88708 47608 88760 47660
rect 6920 47540 6972 47592
rect 10508 47540 10560 47592
rect 11244 47540 11296 47592
rect 46848 47540 46900 47592
rect 47492 47540 47544 47592
rect 89444 47540 89496 47592
rect 11428 47472 11480 47524
rect 5448 47404 5500 47456
rect 11152 47404 11204 47456
rect 48136 47472 48188 47524
rect 89168 47472 89220 47524
rect 88340 47404 88392 47456
rect 3066 47302 3118 47354
rect 3130 47302 3182 47354
rect 3194 47302 3246 47354
rect 3258 47302 3310 47354
rect 3322 47302 3374 47354
rect 6552 47336 6604 47388
rect 86960 47336 87012 47388
rect 6092 47268 6144 47320
rect 10416 47268 10468 47320
rect 10508 47268 10560 47320
rect 88524 47268 88576 47320
rect 5540 47243 5592 47252
rect 5540 47209 5549 47243
rect 5549 47209 5583 47243
rect 5583 47209 5592 47243
rect 5540 47200 5592 47209
rect 10232 47200 10284 47252
rect 7840 47132 7892 47184
rect 88616 47200 88668 47252
rect 10416 47132 10468 47184
rect 87696 47132 87748 47184
rect 6276 47064 6328 47116
rect 88800 47064 88852 47116
rect 1400 47039 1452 47048
rect 1400 47005 1409 47039
rect 1409 47005 1443 47039
rect 1443 47005 1452 47039
rect 1400 46996 1452 47005
rect 11060 46996 11112 47048
rect 11152 46996 11204 47048
rect 88432 46996 88484 47048
rect 9680 46928 9732 46980
rect 11428 46928 11480 46980
rect 12532 46860 12584 46912
rect 3802 46758 3854 46810
rect 3866 46758 3918 46810
rect 3930 46758 3982 46810
rect 3994 46758 4046 46810
rect 4058 46758 4110 46810
rect 48044 46792 48096 46844
rect 52552 46792 52604 46844
rect 51448 46724 51500 46776
rect 6828 46656 6880 46708
rect 13268 46656 13320 46708
rect 11704 46588 11756 46640
rect 47768 46656 47820 46708
rect 51080 46656 51132 46708
rect 47676 46588 47728 46640
rect 47860 46520 47912 46572
rect 53196 46520 53248 46572
rect 89260 46588 89312 46640
rect 87604 46520 87656 46572
rect 4804 46452 4856 46504
rect 9680 46384 9732 46436
rect 1400 46359 1452 46368
rect 1400 46325 1409 46359
rect 1409 46325 1443 46359
rect 1443 46325 1452 46359
rect 1400 46316 1452 46325
rect 3066 46214 3118 46266
rect 3130 46214 3182 46266
rect 3194 46214 3246 46266
rect 3258 46214 3310 46266
rect 3322 46214 3374 46266
rect 8392 46044 8444 46096
rect 8300 45908 8352 45960
rect 10324 46452 10376 46504
rect 51172 46452 51224 46504
rect 88984 46452 89036 46504
rect 12532 46384 12584 46436
rect 48044 46384 48096 46436
rect 48228 46384 48280 46436
rect 49884 46384 49936 46436
rect 48136 46316 48188 46368
rect 1492 45815 1544 45824
rect 1492 45781 1501 45815
rect 1501 45781 1535 45815
rect 1535 45781 1544 45815
rect 1492 45772 1544 45781
rect 3802 45670 3854 45722
rect 3866 45670 3918 45722
rect 3930 45670 3982 45722
rect 3994 45670 4046 45722
rect 4058 45670 4110 45722
rect 1400 45271 1452 45280
rect 1400 45237 1409 45271
rect 1409 45237 1443 45271
rect 1443 45237 1452 45271
rect 1400 45228 1452 45237
rect 3066 45126 3118 45178
rect 3130 45126 3182 45178
rect 3194 45126 3246 45178
rect 3258 45126 3310 45178
rect 3322 45126 3374 45178
rect 3802 44582 3854 44634
rect 3866 44582 3918 44634
rect 3930 44582 3982 44634
rect 3994 44582 4046 44634
rect 4058 44582 4110 44634
rect 6552 44480 6604 44532
rect 5448 44344 5500 44396
rect 8300 44276 8352 44328
rect 1492 44251 1544 44260
rect 1492 44217 1501 44251
rect 1501 44217 1535 44251
rect 1535 44217 1544 44251
rect 1492 44208 1544 44217
rect 3066 44038 3118 44090
rect 3130 44038 3182 44090
rect 3194 44038 3246 44090
rect 3258 44038 3310 44090
rect 3322 44038 3374 44090
rect 6828 43936 6880 43988
rect 1216 43664 1268 43716
rect 3802 43494 3854 43546
rect 3866 43494 3918 43546
rect 3930 43494 3982 43546
rect 3994 43494 4046 43546
rect 4058 43494 4110 43546
rect 7012 43392 7064 43444
rect 8300 43324 8352 43376
rect 6920 43256 6972 43308
rect 1492 43095 1544 43104
rect 1492 43061 1501 43095
rect 1501 43061 1535 43095
rect 1535 43061 1544 43095
rect 1492 43052 1544 43061
rect 3066 42950 3118 43002
rect 3130 42950 3182 43002
rect 3194 42950 3246 43002
rect 3258 42950 3310 43002
rect 3322 42950 3374 43002
rect 3802 42406 3854 42458
rect 3866 42406 3918 42458
rect 3930 42406 3982 42458
rect 3994 42406 4046 42458
rect 4058 42406 4110 42458
rect 3066 41862 3118 41914
rect 3130 41862 3182 41914
rect 3194 41862 3246 41914
rect 3258 41862 3310 41914
rect 3322 41862 3374 41914
rect 5080 41803 5132 41812
rect 5080 41769 5089 41803
rect 5089 41769 5123 41803
rect 5123 41769 5132 41803
rect 5080 41760 5132 41769
rect 6460 41692 6512 41744
rect 8300 41556 8352 41608
rect 5080 41488 5132 41540
rect 1492 41463 1544 41472
rect 1492 41429 1501 41463
rect 1501 41429 1535 41463
rect 1535 41429 1544 41463
rect 1492 41420 1544 41429
rect 3802 41318 3854 41370
rect 3866 41318 3918 41370
rect 3930 41318 3982 41370
rect 3994 41318 4046 41370
rect 4058 41318 4110 41370
rect 88800 41080 88852 41132
rect 3066 40774 3118 40826
rect 3130 40774 3182 40826
rect 3194 40774 3246 40826
rect 3258 40774 3310 40826
rect 3322 40774 3374 40826
rect 88800 40808 88852 40860
rect 4896 40672 4948 40724
rect 5356 40672 5408 40724
rect 88892 40672 88944 40724
rect 89168 40672 89220 40724
rect 89168 40536 89220 40588
rect 89444 40536 89496 40588
rect 8300 40468 8352 40520
rect 4896 40400 4948 40452
rect 848 40332 900 40384
rect 3802 40230 3854 40282
rect 3866 40230 3918 40282
rect 3930 40230 3982 40282
rect 3994 40230 4046 40282
rect 4058 40230 4110 40282
rect 3066 39686 3118 39738
rect 3130 39686 3182 39738
rect 3194 39686 3246 39738
rect 3258 39686 3310 39738
rect 3322 39686 3374 39738
rect 3802 39142 3854 39194
rect 3866 39142 3918 39194
rect 3930 39142 3982 39194
rect 3994 39142 4046 39194
rect 4058 39142 4110 39194
rect 4988 39040 5040 39092
rect 7840 38904 7892 38956
rect 8300 38836 8352 38888
rect 848 38700 900 38752
rect 3066 38598 3118 38650
rect 3130 38598 3182 38650
rect 3194 38598 3246 38650
rect 3258 38598 3310 38650
rect 3322 38598 3374 38650
rect 3802 38054 3854 38106
rect 3866 38054 3918 38106
rect 3930 38054 3982 38106
rect 3994 38054 4046 38106
rect 4058 38054 4110 38106
rect 6368 37952 6420 38004
rect 8300 37884 8352 37936
rect 5724 37816 5776 37868
rect 848 37612 900 37664
rect 3066 37510 3118 37562
rect 3130 37510 3182 37562
rect 3194 37510 3246 37562
rect 3258 37510 3310 37562
rect 3322 37510 3374 37562
rect 3802 36966 3854 37018
rect 3866 36966 3918 37018
rect 3930 36966 3982 37018
rect 3994 36966 4046 37018
rect 4058 36966 4110 37018
rect 3066 36422 3118 36474
rect 3130 36422 3182 36474
rect 3194 36422 3246 36474
rect 3258 36422 3310 36474
rect 3322 36422 3374 36474
rect 4620 36320 4672 36372
rect 848 36252 900 36304
rect 7564 36116 7616 36168
rect 8300 36048 8352 36100
rect 3802 35878 3854 35930
rect 3866 35878 3918 35930
rect 3930 35878 3982 35930
rect 3994 35878 4046 35930
rect 4058 35878 4110 35930
rect 3066 35334 3118 35386
rect 3130 35334 3182 35386
rect 3194 35334 3246 35386
rect 3258 35334 3310 35386
rect 3322 35334 3374 35386
rect 8300 35096 8352 35148
rect 6276 35028 6328 35080
rect 848 34892 900 34944
rect 4988 34892 5040 34944
rect 3802 34790 3854 34842
rect 3866 34790 3918 34842
rect 3930 34790 3982 34842
rect 3994 34790 4046 34842
rect 4058 34790 4110 34842
rect 3066 34246 3118 34298
rect 3130 34246 3182 34298
rect 3194 34246 3246 34298
rect 3258 34246 3310 34298
rect 3322 34246 3374 34298
rect 3802 33702 3854 33754
rect 3866 33702 3918 33754
rect 3930 33702 3982 33754
rect 3994 33702 4046 33754
rect 4058 33702 4110 33754
rect 5632 33507 5684 33516
rect 5632 33473 5641 33507
rect 5641 33473 5675 33507
rect 5675 33473 5684 33507
rect 5632 33464 5684 33473
rect 8300 33396 8352 33448
rect 848 33260 900 33312
rect 6184 33260 6236 33312
rect 3066 33158 3118 33210
rect 3130 33158 3182 33210
rect 3194 33158 3246 33210
rect 3258 33158 3310 33210
rect 3322 33158 3374 33210
rect 3802 32614 3854 32666
rect 3866 32614 3918 32666
rect 3930 32614 3982 32666
rect 3994 32614 4046 32666
rect 4058 32614 4110 32666
rect 4804 32512 4856 32564
rect 8300 32444 8352 32496
rect 4804 32376 4856 32428
rect 848 32172 900 32224
rect 6276 32172 6328 32224
rect 3066 32070 3118 32122
rect 3130 32070 3182 32122
rect 3194 32070 3246 32122
rect 3258 32070 3310 32122
rect 3322 32070 3374 32122
rect 3802 31526 3854 31578
rect 3866 31526 3918 31578
rect 3930 31526 3982 31578
rect 3994 31526 4046 31578
rect 4058 31526 4110 31578
rect 3066 30982 3118 31034
rect 3130 30982 3182 31034
rect 3194 30982 3246 31034
rect 3258 30982 3310 31034
rect 3322 30982 3374 31034
rect 4712 30880 4764 30932
rect 848 30812 900 30864
rect 5632 30719 5684 30728
rect 5632 30685 5641 30719
rect 5641 30685 5675 30719
rect 5675 30685 5684 30719
rect 5632 30676 5684 30685
rect 8300 30608 8352 30660
rect 3802 30438 3854 30490
rect 3866 30438 3918 30490
rect 3930 30438 3982 30490
rect 3994 30438 4046 30490
rect 4058 30438 4110 30490
rect 3066 29894 3118 29946
rect 3130 29894 3182 29946
rect 3194 29894 3246 29946
rect 3258 29894 3310 29946
rect 3322 29894 3374 29946
rect 8300 29656 8352 29708
rect 5448 29631 5500 29640
rect 5448 29597 5457 29631
rect 5457 29597 5491 29631
rect 5491 29597 5500 29631
rect 5448 29588 5500 29597
rect 848 29452 900 29504
rect 5356 29495 5408 29504
rect 5356 29461 5365 29495
rect 5365 29461 5399 29495
rect 5399 29461 5408 29495
rect 5356 29452 5408 29461
rect 3802 29350 3854 29402
rect 3866 29350 3918 29402
rect 3930 29350 3982 29402
rect 3994 29350 4046 29402
rect 4058 29350 4110 29402
rect 3066 28806 3118 28858
rect 3130 28806 3182 28858
rect 3194 28806 3246 28858
rect 3258 28806 3310 28858
rect 3322 28806 3374 28858
rect 3802 28262 3854 28314
rect 3866 28262 3918 28314
rect 3930 28262 3982 28314
rect 3994 28262 4046 28314
rect 4058 28262 4110 28314
rect 5080 28203 5132 28212
rect 5080 28169 5089 28203
rect 5089 28169 5123 28203
rect 5123 28169 5132 28203
rect 5080 28160 5132 28169
rect 5264 28203 5316 28212
rect 5264 28169 5273 28203
rect 5273 28169 5307 28203
rect 5307 28169 5316 28203
rect 5264 28160 5316 28169
rect 8300 27956 8352 28008
rect 848 27820 900 27872
rect 3066 27718 3118 27770
rect 3130 27718 3182 27770
rect 3194 27718 3246 27770
rect 3258 27718 3310 27770
rect 3322 27718 3374 27770
rect 3802 27174 3854 27226
rect 3866 27174 3918 27226
rect 3930 27174 3982 27226
rect 3994 27174 4046 27226
rect 4058 27174 4110 27226
rect 8300 27072 8352 27124
rect 5264 27047 5316 27056
rect 5264 27013 5273 27047
rect 5273 27013 5307 27047
rect 5307 27013 5316 27047
rect 5264 27004 5316 27013
rect 1308 26936 1360 26988
rect 5540 26775 5592 26784
rect 5540 26741 5549 26775
rect 5549 26741 5583 26775
rect 5583 26741 5592 26775
rect 5540 26732 5592 26741
rect 3066 26630 3118 26682
rect 3130 26630 3182 26682
rect 3194 26630 3246 26682
rect 3258 26630 3310 26682
rect 3322 26630 3374 26682
rect 3802 26086 3854 26138
rect 3866 26086 3918 26138
rect 3930 26086 3982 26138
rect 3994 26086 4046 26138
rect 4058 26086 4110 26138
rect 3066 25542 3118 25594
rect 3130 25542 3182 25594
rect 3194 25542 3246 25594
rect 3258 25542 3310 25594
rect 3322 25542 3374 25594
rect 5816 25440 5868 25492
rect 8300 25372 8352 25424
rect 1216 25236 1268 25288
rect 6368 25100 6420 25152
rect 3802 24998 3854 25050
rect 3866 24998 3918 25050
rect 3930 24998 3982 25050
rect 3994 24998 4046 25050
rect 4058 24998 4110 25050
rect 3066 24454 3118 24506
rect 3130 24454 3182 24506
rect 3194 24454 3246 24506
rect 3258 24454 3310 24506
rect 3322 24454 3374 24506
rect 8300 24284 8352 24336
rect 1308 24148 1360 24200
rect 3802 23910 3854 23962
rect 3866 23910 3918 23962
rect 3930 23910 3982 23962
rect 3994 23910 4046 23962
rect 4058 23910 4110 23962
rect 3066 23366 3118 23418
rect 3130 23366 3182 23418
rect 3194 23366 3246 23418
rect 3258 23366 3310 23418
rect 3322 23366 3374 23418
rect 3802 22822 3854 22874
rect 3866 22822 3918 22874
rect 3930 22822 3982 22874
rect 3994 22822 4046 22874
rect 4058 22822 4110 22874
rect 1308 22584 1360 22636
rect 8300 22448 8352 22500
rect 3066 22278 3118 22330
rect 3130 22278 3182 22330
rect 3194 22278 3246 22330
rect 3258 22278 3310 22330
rect 3322 22278 3374 22330
rect 3802 21734 3854 21786
rect 3866 21734 3918 21786
rect 3930 21734 3982 21786
rect 3994 21734 4046 21786
rect 4058 21734 4110 21786
rect 8300 21632 8352 21684
rect 1308 21496 1360 21548
rect 3066 21190 3118 21242
rect 3130 21190 3182 21242
rect 3194 21190 3246 21242
rect 3258 21190 3310 21242
rect 3322 21190 3374 21242
rect 3802 20646 3854 20698
rect 3866 20646 3918 20698
rect 3930 20646 3982 20698
rect 3994 20646 4046 20698
rect 4058 20646 4110 20698
rect 3066 20102 3118 20154
rect 3130 20102 3182 20154
rect 3194 20102 3246 20154
rect 3258 20102 3310 20154
rect 3322 20102 3374 20154
rect 8300 20000 8352 20052
rect 1216 19796 1268 19848
rect 3802 19558 3854 19610
rect 3866 19558 3918 19610
rect 3930 19558 3982 19610
rect 3994 19558 4046 19610
rect 4058 19558 4110 19610
rect 3066 19014 3118 19066
rect 3130 19014 3182 19066
rect 3194 19014 3246 19066
rect 3258 19014 3310 19066
rect 3322 19014 3374 19066
rect 8300 18844 8352 18896
rect 1308 18708 1360 18760
rect 3802 18470 3854 18522
rect 3866 18470 3918 18522
rect 3930 18470 3982 18522
rect 3994 18470 4046 18522
rect 4058 18470 4110 18522
rect 3066 17926 3118 17978
rect 3130 17926 3182 17978
rect 3194 17926 3246 17978
rect 3258 17926 3310 17978
rect 3322 17926 3374 17978
rect 3802 17382 3854 17434
rect 3866 17382 3918 17434
rect 3930 17382 3982 17434
rect 3994 17382 4046 17434
rect 4058 17382 4110 17434
rect 1308 17144 1360 17196
rect 8300 17008 8352 17060
rect 3066 16838 3118 16890
rect 3130 16838 3182 16890
rect 3194 16838 3246 16890
rect 3258 16838 3310 16890
rect 3322 16838 3374 16890
rect 3802 16294 3854 16346
rect 3866 16294 3918 16346
rect 3930 16294 3982 16346
rect 3994 16294 4046 16346
rect 4058 16294 4110 16346
rect 8300 16192 8352 16244
rect 1308 16056 1360 16108
rect 3066 15750 3118 15802
rect 3130 15750 3182 15802
rect 3194 15750 3246 15802
rect 3258 15750 3310 15802
rect 3322 15750 3374 15802
rect 3802 15206 3854 15258
rect 3866 15206 3918 15258
rect 3930 15206 3982 15258
rect 3994 15206 4046 15258
rect 4058 15206 4110 15258
rect 3066 14662 3118 14714
rect 3130 14662 3182 14714
rect 3194 14662 3246 14714
rect 3258 14662 3310 14714
rect 3322 14662 3374 14714
rect 8300 14560 8352 14612
rect 1216 14356 1268 14408
rect 3802 14118 3854 14170
rect 3866 14118 3918 14170
rect 3930 14118 3982 14170
rect 3994 14118 4046 14170
rect 4058 14118 4110 14170
rect 3066 13574 3118 13626
rect 3130 13574 3182 13626
rect 3194 13574 3246 13626
rect 3258 13574 3310 13626
rect 3322 13574 3374 13626
rect 8300 13404 8352 13456
rect 1308 13268 1360 13320
rect 3802 13030 3854 13082
rect 3866 13030 3918 13082
rect 3930 13030 3982 13082
rect 3994 13030 4046 13082
rect 4058 13030 4110 13082
rect 3066 12486 3118 12538
rect 3130 12486 3182 12538
rect 3194 12486 3246 12538
rect 3258 12486 3310 12538
rect 3322 12486 3374 12538
rect 3802 11942 3854 11994
rect 3866 11942 3918 11994
rect 3930 11942 3982 11994
rect 3994 11942 4046 11994
rect 4058 11942 4110 11994
rect 1308 11704 1360 11756
rect 8300 11568 8352 11620
rect 3066 11398 3118 11450
rect 3130 11398 3182 11450
rect 3194 11398 3246 11450
rect 3258 11398 3310 11450
rect 3322 11398 3374 11450
rect 3802 10854 3854 10906
rect 3866 10854 3918 10906
rect 3930 10854 3982 10906
rect 3994 10854 4046 10906
rect 4058 10854 4110 10906
rect 3066 10310 3118 10362
rect 3130 10310 3182 10362
rect 3194 10310 3246 10362
rect 3258 10310 3310 10362
rect 3322 10310 3374 10362
rect 3802 9766 3854 9818
rect 3866 9766 3918 9818
rect 3930 9766 3982 9818
rect 3994 9766 4046 9818
rect 4058 9766 4110 9818
rect 46756 9596 46808 9648
rect 48688 9596 48740 9648
rect 86868 9460 86920 9512
rect 88156 9460 88208 9512
rect 3066 9222 3118 9274
rect 3130 9222 3182 9274
rect 3194 9222 3246 9274
rect 3258 9222 3310 9274
rect 3322 9222 3374 9274
rect 88064 8780 88116 8832
rect 89168 8780 89220 8832
rect 3802 8678 3854 8730
rect 3866 8678 3918 8730
rect 3930 8678 3982 8730
rect 3994 8678 4046 8730
rect 4058 8678 4110 8730
rect 47584 8576 47636 8628
rect 49332 8576 49384 8628
rect 5356 8236 5408 8288
rect 3066 8134 3118 8186
rect 3130 8134 3182 8186
rect 3194 8134 3246 8186
rect 3258 8134 3310 8186
rect 3322 8134 3374 8186
rect 8208 8168 8260 8220
rect 12716 8168 12768 8220
rect 48688 8168 48740 8220
rect 53840 8168 53892 8220
rect 84752 8236 84804 8288
rect 87236 8236 87288 8288
rect 86040 8168 86092 8220
rect 6828 8100 6880 8152
rect 8024 8100 8076 8152
rect 10508 8100 10560 8152
rect 11612 8032 11664 8084
rect 5448 7964 5500 8016
rect 47400 7964 47452 8016
rect 5540 7896 5592 7948
rect 47676 7896 47728 7948
rect 4988 7828 5040 7880
rect 47952 7828 48004 7880
rect 5632 7760 5684 7812
rect 47492 7760 47544 7812
rect 85304 7760 85356 7812
rect 6368 7692 6420 7744
rect 84752 7692 84804 7744
rect 3802 7590 3854 7642
rect 3866 7590 3918 7642
rect 3930 7590 3982 7642
rect 3994 7590 4046 7642
rect 4058 7590 4110 7642
rect 6184 7624 6236 7676
rect 85672 7624 85724 7676
rect 6276 7556 6328 7608
rect 85764 7556 85816 7608
rect 3066 7046 3118 7098
rect 3130 7046 3182 7098
rect 3194 7046 3246 7098
rect 3258 7046 3310 7098
rect 3322 7046 3374 7098
rect 3802 6502 3854 6554
rect 3866 6502 3918 6554
rect 3930 6502 3982 6554
rect 3994 6502 4046 6554
rect 4058 6502 4110 6554
rect 48228 6196 48280 6248
rect 50252 6196 50304 6248
rect 10876 6128 10928 6180
rect 50804 6128 50856 6180
rect 3066 5958 3118 6010
rect 3130 5958 3182 6010
rect 3194 5958 3246 6010
rect 3258 5958 3310 6010
rect 3322 5958 3374 6010
rect 72950 5958 73002 6010
rect 73014 5958 73066 6010
rect 73078 5958 73130 6010
rect 73142 5958 73194 6010
rect 73206 5958 73258 6010
rect 10876 5899 10928 5908
rect 10876 5865 10885 5899
rect 10885 5865 10919 5899
rect 10919 5865 10928 5899
rect 10876 5856 10928 5865
rect 12992 5899 13044 5908
rect 12992 5865 13001 5899
rect 13001 5865 13035 5899
rect 13035 5865 13044 5899
rect 12992 5856 13044 5865
rect 15108 5856 15160 5908
rect 49700 5899 49752 5908
rect 49700 5865 49709 5899
rect 49709 5865 49743 5899
rect 49743 5865 49752 5899
rect 49700 5856 49752 5865
rect 50252 5899 50304 5908
rect 50252 5865 50261 5899
rect 50261 5865 50295 5899
rect 50295 5865 50304 5899
rect 50252 5856 50304 5865
rect 50804 5899 50856 5908
rect 50804 5865 50813 5899
rect 50813 5865 50847 5899
rect 50847 5865 50856 5899
rect 50804 5856 50856 5865
rect 46940 5788 46992 5840
rect 47860 5788 47912 5840
rect 84752 5899 84804 5908
rect 84752 5865 84761 5899
rect 84761 5865 84795 5899
rect 84795 5865 84804 5899
rect 84752 5856 84804 5865
rect 85028 5856 85080 5908
rect 85120 5831 85172 5840
rect 85120 5797 85129 5831
rect 85129 5797 85163 5831
rect 85163 5797 85172 5831
rect 85120 5788 85172 5797
rect 85304 5899 85356 5908
rect 85304 5865 85313 5899
rect 85313 5865 85347 5899
rect 85347 5865 85356 5899
rect 85304 5856 85356 5865
rect 86316 5899 86368 5908
rect 86316 5865 86325 5899
rect 86325 5865 86359 5899
rect 86359 5865 86368 5899
rect 86316 5856 86368 5865
rect 86592 5899 86644 5908
rect 86592 5865 86601 5899
rect 86601 5865 86635 5899
rect 86635 5865 86644 5899
rect 86592 5856 86644 5865
rect 88064 5899 88116 5908
rect 88064 5865 88073 5899
rect 88073 5865 88107 5899
rect 88107 5865 88116 5899
rect 88064 5856 88116 5865
rect 88524 5856 88576 5908
rect 43444 5720 43496 5772
rect 47768 5720 47820 5772
rect 86868 5720 86920 5772
rect 89260 5788 89312 5840
rect 88984 5720 89036 5772
rect 9772 5695 9824 5704
rect 9772 5661 9781 5695
rect 9781 5661 9815 5695
rect 9815 5661 9824 5695
rect 9772 5652 9824 5661
rect 46940 5652 46992 5704
rect 11980 5627 12032 5636
rect 11980 5593 11989 5627
rect 11989 5593 12023 5627
rect 12023 5593 12032 5627
rect 11980 5584 12032 5593
rect 13360 5584 13412 5636
rect 48044 5652 48096 5704
rect 86316 5652 86368 5704
rect 86408 5695 86460 5704
rect 86408 5661 86417 5695
rect 86417 5661 86451 5695
rect 86451 5661 86460 5695
rect 86408 5652 86460 5661
rect 87052 5652 87104 5704
rect 87144 5695 87196 5704
rect 87144 5661 87153 5695
rect 87153 5661 87187 5695
rect 87187 5661 87196 5695
rect 87144 5652 87196 5661
rect 87512 5695 87564 5704
rect 87512 5661 87521 5695
rect 87521 5661 87555 5695
rect 87555 5661 87564 5695
rect 87512 5652 87564 5661
rect 87696 5652 87748 5704
rect 88248 5695 88300 5704
rect 88248 5661 88257 5695
rect 88257 5661 88291 5695
rect 88291 5661 88300 5695
rect 88248 5652 88300 5661
rect 51908 5627 51960 5636
rect 51908 5593 51917 5627
rect 51917 5593 51951 5627
rect 51951 5593 51960 5627
rect 51908 5584 51960 5593
rect 85580 5627 85632 5636
rect 85580 5593 85589 5627
rect 85589 5593 85623 5627
rect 85623 5593 85632 5627
rect 85580 5584 85632 5593
rect 86500 5584 86552 5636
rect 43444 5516 43496 5568
rect 53012 5559 53064 5568
rect 53012 5525 53021 5559
rect 53021 5525 53055 5559
rect 53055 5525 53064 5559
rect 53012 5516 53064 5525
rect 89076 5516 89128 5568
rect 3802 5414 3854 5466
rect 3866 5414 3918 5466
rect 3930 5414 3982 5466
rect 3994 5414 4046 5466
rect 4058 5414 4110 5466
rect 37610 5414 37662 5466
rect 37674 5414 37726 5466
rect 37738 5414 37790 5466
rect 37802 5414 37854 5466
rect 37866 5414 37918 5466
rect 73610 5414 73662 5466
rect 73674 5414 73726 5466
rect 73738 5414 73790 5466
rect 73802 5414 73854 5466
rect 73866 5414 73918 5466
rect 85672 5312 85724 5364
rect 86040 5355 86092 5364
rect 86040 5321 86049 5355
rect 86049 5321 86083 5355
rect 86083 5321 86092 5355
rect 86040 5312 86092 5321
rect 86500 5355 86552 5364
rect 86500 5321 86509 5355
rect 86509 5321 86543 5355
rect 86543 5321 86552 5355
rect 86500 5312 86552 5321
rect 86684 5355 86736 5364
rect 86684 5321 86693 5355
rect 86693 5321 86727 5355
rect 86727 5321 86736 5355
rect 86684 5312 86736 5321
rect 86776 5244 86828 5296
rect 87972 5244 88024 5296
rect 88432 5355 88484 5364
rect 88432 5321 88441 5355
rect 88441 5321 88475 5355
rect 88475 5321 88484 5355
rect 88432 5312 88484 5321
rect 88892 5244 88944 5296
rect 83924 5108 83976 5160
rect 87420 5176 87472 5228
rect 87880 5219 87932 5228
rect 87880 5185 87889 5219
rect 87889 5185 87923 5219
rect 87923 5185 87932 5219
rect 87880 5176 87932 5185
rect 88248 5219 88300 5228
rect 88248 5185 88257 5219
rect 88257 5185 88291 5219
rect 88291 5185 88300 5219
rect 88248 5176 88300 5185
rect 88340 5108 88392 5160
rect 53840 5040 53892 5092
rect 89352 5040 89404 5092
rect 88708 4972 88760 5024
rect 36950 4870 37002 4922
rect 37014 4870 37066 4922
rect 37078 4870 37130 4922
rect 37142 4870 37194 4922
rect 37206 4870 37258 4922
rect 72950 4870 73002 4922
rect 73014 4870 73066 4922
rect 73078 4870 73130 4922
rect 73142 4870 73194 4922
rect 73206 4870 73258 4922
rect 85764 4768 85816 4820
rect 87236 4811 87288 4820
rect 87236 4777 87245 4811
rect 87245 4777 87279 4811
rect 87279 4777 87288 4811
rect 87236 4768 87288 4777
rect 88156 4768 88208 4820
rect 89444 4768 89496 4820
rect 87696 4743 87748 4752
rect 87696 4709 87705 4743
rect 87705 4709 87739 4743
rect 87739 4709 87748 4743
rect 87696 4700 87748 4709
rect 88800 4700 88852 4752
rect 88340 4632 88392 4684
rect 87788 4564 87840 4616
rect 88616 4564 88668 4616
rect 47216 4496 47268 4548
rect 86960 4539 87012 4548
rect 86960 4505 86969 4539
rect 86969 4505 87003 4539
rect 87003 4505 87012 4539
rect 86960 4496 87012 4505
rect 46848 4428 46900 4480
rect 37610 4326 37662 4378
rect 37674 4326 37726 4378
rect 37738 4326 37790 4378
rect 37802 4326 37854 4378
rect 37866 4326 37918 4378
rect 73610 4326 73662 4378
rect 73674 4326 73726 4378
rect 73738 4326 73790 4378
rect 73802 4326 73854 4378
rect 73866 4326 73918 4378
rect 88156 4267 88208 4276
rect 88156 4233 88165 4267
rect 88165 4233 88199 4267
rect 88199 4233 88208 4267
rect 88156 4224 88208 4233
rect 36950 3782 37002 3834
rect 37014 3782 37066 3834
rect 37078 3782 37130 3834
rect 37142 3782 37194 3834
rect 37206 3782 37258 3834
rect 72950 3782 73002 3834
rect 73014 3782 73066 3834
rect 73078 3782 73130 3834
rect 73142 3782 73194 3834
rect 73206 3782 73258 3834
rect 37610 3238 37662 3290
rect 37674 3238 37726 3290
rect 37738 3238 37790 3290
rect 37802 3238 37854 3290
rect 37866 3238 37918 3290
rect 73610 3238 73662 3290
rect 73674 3238 73726 3290
rect 73738 3238 73790 3290
rect 73802 3238 73854 3290
rect 73866 3238 73918 3290
rect 36950 2694 37002 2746
rect 37014 2694 37066 2746
rect 37078 2694 37130 2746
rect 37142 2694 37194 2746
rect 37206 2694 37258 2746
rect 72950 2694 73002 2746
rect 73014 2694 73066 2746
rect 73078 2694 73130 2746
rect 73142 2694 73194 2746
rect 73206 2694 73258 2746
rect 8300 2592 8352 2644
rect 10876 2592 10928 2644
rect 13360 2635 13412 2644
rect 13360 2601 13369 2635
rect 13369 2601 13403 2635
rect 13403 2601 13412 2635
rect 13360 2592 13412 2601
rect 15108 2635 15160 2644
rect 8116 2524 8168 2576
rect 15108 2601 15117 2635
rect 15117 2601 15151 2635
rect 15151 2601 15160 2635
rect 15108 2592 15160 2601
rect 31024 2635 31076 2644
rect 31024 2601 31033 2635
rect 31033 2601 31067 2635
rect 31067 2601 31076 2635
rect 31024 2592 31076 2601
rect 31852 2635 31904 2644
rect 31852 2601 31861 2635
rect 31861 2601 31895 2635
rect 31895 2601 31904 2635
rect 31852 2592 31904 2601
rect 32956 2635 33008 2644
rect 32956 2601 32965 2635
rect 32965 2601 32999 2635
rect 32999 2601 33008 2635
rect 32956 2592 33008 2601
rect 34244 2635 34296 2644
rect 34244 2601 34253 2635
rect 34253 2601 34287 2635
rect 34287 2601 34296 2635
rect 34244 2592 34296 2601
rect 35072 2635 35124 2644
rect 35072 2601 35081 2635
rect 35081 2601 35115 2635
rect 35115 2601 35124 2635
rect 35072 2592 35124 2601
rect 36176 2635 36228 2644
rect 36176 2601 36185 2635
rect 36185 2601 36219 2635
rect 36219 2601 36228 2635
rect 36176 2592 36228 2601
rect 37464 2635 37516 2644
rect 37464 2601 37473 2635
rect 37473 2601 37507 2635
rect 37507 2601 37516 2635
rect 37464 2592 37516 2601
rect 42800 2635 42852 2644
rect 42800 2601 42809 2635
rect 42809 2601 42843 2635
rect 42843 2601 42852 2635
rect 42800 2592 42852 2601
rect 45192 2635 45244 2644
rect 45192 2601 45201 2635
rect 45201 2601 45235 2635
rect 45235 2601 45244 2635
rect 45192 2592 45244 2601
rect 70952 2635 71004 2644
rect 70952 2601 70961 2635
rect 70961 2601 70995 2635
rect 70995 2601 71004 2635
rect 70952 2592 71004 2601
rect 71780 2635 71832 2644
rect 71780 2601 71789 2635
rect 71789 2601 71823 2635
rect 71823 2601 71832 2635
rect 71780 2592 71832 2601
rect 72792 2592 72844 2644
rect 74172 2635 74224 2644
rect 74172 2601 74181 2635
rect 74181 2601 74215 2635
rect 74215 2601 74224 2635
rect 74172 2592 74224 2601
rect 75092 2592 75144 2644
rect 76288 2635 76340 2644
rect 76288 2601 76297 2635
rect 76297 2601 76331 2635
rect 76331 2601 76340 2635
rect 76288 2592 76340 2601
rect 77392 2635 77444 2644
rect 77392 2601 77401 2635
rect 77401 2601 77435 2635
rect 77435 2601 77444 2635
rect 77392 2592 77444 2601
rect 39856 2567 39908 2576
rect 39856 2533 39865 2567
rect 39865 2533 39899 2567
rect 39899 2533 39908 2567
rect 39856 2524 39908 2533
rect 40684 2567 40736 2576
rect 40684 2533 40693 2567
rect 40693 2533 40727 2567
rect 40727 2533 40736 2567
rect 40684 2524 40736 2533
rect 41972 2567 42024 2576
rect 41972 2533 41981 2567
rect 41981 2533 42015 2567
rect 42015 2533 42024 2567
rect 41972 2524 42024 2533
rect 43904 2567 43956 2576
rect 43904 2533 43913 2567
rect 43913 2533 43947 2567
rect 43947 2533 43956 2567
rect 43904 2524 43956 2533
rect 79600 2567 79652 2576
rect 79600 2533 79609 2567
rect 79609 2533 79643 2567
rect 79643 2533 79652 2567
rect 79600 2524 79652 2533
rect 80612 2567 80664 2576
rect 80612 2533 80621 2567
rect 80621 2533 80655 2567
rect 80655 2533 80664 2567
rect 80612 2524 80664 2533
rect 81900 2567 81952 2576
rect 81900 2533 81909 2567
rect 81909 2533 81943 2567
rect 81943 2533 81952 2567
rect 81900 2524 81952 2533
rect 82820 2524 82872 2576
rect 38384 2456 38436 2508
rect 78404 2456 78456 2508
rect 15568 2431 15620 2440
rect 15568 2397 15577 2431
rect 15577 2397 15611 2431
rect 15611 2397 15620 2431
rect 15568 2388 15620 2397
rect 16488 2431 16540 2440
rect 16488 2397 16497 2431
rect 16497 2397 16531 2431
rect 16531 2397 16540 2431
rect 16488 2388 16540 2397
rect 17500 2431 17552 2440
rect 17500 2397 17509 2431
rect 17509 2397 17543 2431
rect 17543 2397 17552 2431
rect 17500 2388 17552 2397
rect 18788 2431 18840 2440
rect 18788 2397 18797 2431
rect 18797 2397 18831 2431
rect 18831 2397 18840 2431
rect 18788 2388 18840 2397
rect 19708 2431 19760 2440
rect 19708 2397 19717 2431
rect 19717 2397 19751 2431
rect 19751 2397 19760 2431
rect 19708 2388 19760 2397
rect 20720 2431 20772 2440
rect 20720 2397 20729 2431
rect 20729 2397 20763 2431
rect 20763 2397 20772 2431
rect 20720 2388 20772 2397
rect 22008 2431 22060 2440
rect 22008 2397 22017 2431
rect 22017 2397 22051 2431
rect 22051 2397 22060 2431
rect 22008 2388 22060 2397
rect 23296 2431 23348 2440
rect 23296 2397 23305 2431
rect 23305 2397 23339 2431
rect 23339 2397 23348 2431
rect 23296 2388 23348 2397
rect 24216 2431 24268 2440
rect 24216 2397 24225 2431
rect 24225 2397 24259 2431
rect 24259 2397 24268 2431
rect 24216 2388 24268 2397
rect 25228 2431 25280 2440
rect 25228 2397 25237 2431
rect 25237 2397 25271 2431
rect 25271 2397 25280 2431
rect 25228 2388 25280 2397
rect 26516 2431 26568 2440
rect 26516 2397 26525 2431
rect 26525 2397 26559 2431
rect 26559 2397 26568 2431
rect 26516 2388 26568 2397
rect 27436 2431 27488 2440
rect 27436 2397 27445 2431
rect 27445 2397 27479 2431
rect 27479 2397 27488 2431
rect 27436 2388 27488 2397
rect 28448 2431 28500 2440
rect 28448 2397 28457 2431
rect 28457 2397 28491 2431
rect 28491 2397 28500 2431
rect 28448 2388 28500 2397
rect 29736 2431 29788 2440
rect 29736 2397 29745 2431
rect 29745 2397 29779 2431
rect 29779 2397 29788 2431
rect 29736 2388 29788 2397
rect 10968 2320 11020 2372
rect 7748 2295 7800 2304
rect 7748 2261 7757 2295
rect 7757 2261 7791 2295
rect 7791 2261 7800 2295
rect 7748 2252 7800 2261
rect 8392 2295 8444 2304
rect 8392 2261 8401 2295
rect 8401 2261 8435 2295
rect 8435 2261 8444 2295
rect 8392 2252 8444 2261
rect 12256 2295 12308 2304
rect 12256 2261 12265 2295
rect 12265 2261 12299 2295
rect 12299 2261 12308 2295
rect 12256 2252 12308 2261
rect 13544 2252 13596 2304
rect 39304 2320 39356 2372
rect 15476 2252 15528 2304
rect 16120 2252 16172 2304
rect 17408 2252 17460 2304
rect 18696 2252 18748 2304
rect 19340 2252 19392 2304
rect 20628 2252 20680 2304
rect 21916 2252 21968 2304
rect 23204 2252 23256 2304
rect 23848 2252 23900 2304
rect 25136 2252 25188 2304
rect 26424 2252 26476 2304
rect 27068 2252 27120 2304
rect 28356 2252 28408 2304
rect 29644 2252 29696 2304
rect 30932 2295 30984 2304
rect 30932 2261 30941 2295
rect 30941 2261 30975 2295
rect 30975 2261 30984 2295
rect 30932 2252 30984 2261
rect 31576 2295 31628 2304
rect 31576 2261 31585 2295
rect 31585 2261 31619 2295
rect 31619 2261 31628 2295
rect 31576 2252 31628 2261
rect 32864 2295 32916 2304
rect 32864 2261 32873 2295
rect 32873 2261 32907 2295
rect 32907 2261 32916 2295
rect 32864 2252 32916 2261
rect 34152 2295 34204 2304
rect 34152 2261 34161 2295
rect 34161 2261 34195 2295
rect 34195 2261 34204 2295
rect 34152 2252 34204 2261
rect 34796 2295 34848 2304
rect 34796 2261 34805 2295
rect 34805 2261 34839 2295
rect 34839 2261 34848 2295
rect 34796 2252 34848 2261
rect 36084 2295 36136 2304
rect 36084 2261 36093 2295
rect 36093 2261 36127 2295
rect 36127 2261 36136 2295
rect 36084 2252 36136 2261
rect 37372 2295 37424 2304
rect 37372 2261 37381 2295
rect 37381 2261 37415 2295
rect 37415 2261 37424 2295
rect 37372 2252 37424 2261
rect 38660 2295 38712 2304
rect 38660 2261 38669 2295
rect 38669 2261 38703 2295
rect 38703 2261 38712 2295
rect 38660 2252 38712 2261
rect 40592 2295 40644 2304
rect 40592 2261 40601 2295
rect 40601 2261 40635 2295
rect 40635 2261 40644 2295
rect 40592 2252 40644 2261
rect 41880 2295 41932 2304
rect 41880 2261 41889 2295
rect 41889 2261 41923 2295
rect 41923 2261 41932 2295
rect 41880 2252 41932 2261
rect 42524 2295 42576 2304
rect 42524 2261 42533 2295
rect 42533 2261 42567 2295
rect 42567 2261 42576 2295
rect 42524 2252 42576 2261
rect 43812 2295 43864 2304
rect 43812 2261 43821 2295
rect 43821 2261 43855 2295
rect 43855 2261 43864 2295
rect 55496 2431 55548 2440
rect 55496 2397 55505 2431
rect 55505 2397 55539 2431
rect 55539 2397 55548 2431
rect 55496 2388 55548 2397
rect 56416 2431 56468 2440
rect 56416 2397 56425 2431
rect 56425 2397 56459 2431
rect 56459 2397 56468 2431
rect 56416 2388 56468 2397
rect 57428 2431 57480 2440
rect 57428 2397 57437 2431
rect 57437 2397 57471 2431
rect 57471 2397 57480 2431
rect 57428 2388 57480 2397
rect 58716 2431 58768 2440
rect 58716 2397 58725 2431
rect 58725 2397 58759 2431
rect 58759 2397 58768 2431
rect 58716 2388 58768 2397
rect 59636 2388 59688 2440
rect 60740 2388 60792 2440
rect 61936 2431 61988 2440
rect 61936 2397 61945 2431
rect 61945 2397 61979 2431
rect 61979 2397 61988 2431
rect 61936 2388 61988 2397
rect 63224 2431 63276 2440
rect 63224 2397 63233 2431
rect 63233 2397 63267 2431
rect 63267 2397 63276 2431
rect 63224 2388 63276 2397
rect 64144 2431 64196 2440
rect 64144 2397 64153 2431
rect 64153 2397 64187 2431
rect 64187 2397 64196 2431
rect 64144 2388 64196 2397
rect 65156 2431 65208 2440
rect 65156 2397 65165 2431
rect 65165 2397 65199 2431
rect 65199 2397 65208 2431
rect 65156 2388 65208 2397
rect 66444 2431 66496 2440
rect 66444 2397 66453 2431
rect 66453 2397 66487 2431
rect 66487 2397 66496 2431
rect 66444 2388 66496 2397
rect 67364 2388 67416 2440
rect 68376 2431 68428 2440
rect 68376 2397 68385 2431
rect 68385 2397 68419 2431
rect 68419 2397 68428 2431
rect 68376 2388 68428 2397
rect 69664 2431 69716 2440
rect 69664 2397 69673 2431
rect 69673 2397 69707 2431
rect 69707 2397 69716 2431
rect 69664 2388 69716 2397
rect 79232 2320 79284 2372
rect 43812 2252 43864 2261
rect 45100 2295 45152 2304
rect 45100 2261 45109 2295
rect 45109 2261 45143 2295
rect 45143 2261 45152 2295
rect 45100 2252 45152 2261
rect 55404 2252 55456 2304
rect 56048 2252 56100 2304
rect 57336 2252 57388 2304
rect 58624 2252 58676 2304
rect 59912 2252 59964 2304
rect 60556 2252 60608 2304
rect 61844 2252 61896 2304
rect 63132 2252 63184 2304
rect 63776 2252 63828 2304
rect 65064 2252 65116 2304
rect 66352 2252 66404 2304
rect 67640 2252 67692 2304
rect 68284 2252 68336 2304
rect 69572 2252 69624 2304
rect 70860 2295 70912 2304
rect 70860 2261 70869 2295
rect 70869 2261 70903 2295
rect 70903 2261 70912 2295
rect 70860 2252 70912 2261
rect 71504 2295 71556 2304
rect 71504 2261 71513 2295
rect 71513 2261 71547 2295
rect 71547 2261 71556 2295
rect 71504 2252 71556 2261
rect 72792 2295 72844 2304
rect 72792 2261 72801 2295
rect 72801 2261 72835 2295
rect 72835 2261 72844 2295
rect 72792 2252 72844 2261
rect 74080 2295 74132 2304
rect 74080 2261 74089 2295
rect 74089 2261 74123 2295
rect 74123 2261 74132 2295
rect 74080 2252 74132 2261
rect 75368 2295 75420 2304
rect 75368 2261 75377 2295
rect 75377 2261 75411 2295
rect 75411 2261 75420 2295
rect 75368 2252 75420 2261
rect 76012 2295 76064 2304
rect 76012 2261 76021 2295
rect 76021 2261 76055 2295
rect 76055 2261 76064 2295
rect 76012 2252 76064 2261
rect 77300 2295 77352 2304
rect 77300 2261 77309 2295
rect 77309 2261 77343 2295
rect 77343 2261 77352 2295
rect 77300 2252 77352 2261
rect 78588 2295 78640 2304
rect 78588 2261 78597 2295
rect 78597 2261 78631 2295
rect 78631 2261 78640 2295
rect 78588 2252 78640 2261
rect 80520 2295 80572 2304
rect 80520 2261 80529 2295
rect 80529 2261 80563 2295
rect 80563 2261 80572 2295
rect 80520 2252 80572 2261
rect 81808 2295 81860 2304
rect 81808 2261 81817 2295
rect 81817 2261 81851 2295
rect 81851 2261 81860 2295
rect 81808 2252 81860 2261
rect 83096 2295 83148 2304
rect 83096 2261 83105 2295
rect 83105 2261 83139 2295
rect 83139 2261 83148 2295
rect 83096 2252 83148 2261
rect 37610 2150 37662 2202
rect 37674 2150 37726 2202
rect 37738 2150 37790 2202
rect 37802 2150 37854 2202
rect 37866 2150 37918 2202
rect 73610 2150 73662 2202
rect 73674 2150 73726 2202
rect 73738 2150 73790 2202
rect 73802 2150 73854 2202
rect 73866 2150 73918 2202
<< metal2 >>
rect 8390 97322 8446 98000
rect 14830 97322 14886 98000
rect 8390 97294 8708 97322
rect 8390 97200 8446 97294
rect 8680 95674 8708 97294
rect 14752 97294 14886 97322
rect 14752 95674 14780 97294
rect 14830 97200 14886 97294
rect 15474 97322 15530 98000
rect 16762 97322 16818 98000
rect 18050 97322 18106 98000
rect 15474 97294 15608 97322
rect 15474 97200 15530 97294
rect 8668 95668 8720 95674
rect 8668 95610 8720 95616
rect 14740 95668 14792 95674
rect 14740 95610 14792 95616
rect 15580 95538 15608 97294
rect 16684 97294 16818 97322
rect 16684 95674 16712 97294
rect 16762 97200 16818 97294
rect 17972 97294 18106 97322
rect 17972 95674 18000 97294
rect 18050 97200 18106 97294
rect 19338 97322 19394 98000
rect 19982 97322 20038 98000
rect 21270 97322 21326 98000
rect 22558 97322 22614 98000
rect 23202 97322 23258 98000
rect 24490 97322 24546 98000
rect 25778 97322 25834 98000
rect 27066 97322 27122 98000
rect 27710 97322 27766 98000
rect 19338 97294 19472 97322
rect 19338 97200 19394 97294
rect 19444 95674 19472 97294
rect 19982 97294 20392 97322
rect 19982 97200 20038 97294
rect 20364 95674 20392 97294
rect 21192 97294 21326 97322
rect 21192 95674 21220 97294
rect 21270 97200 21326 97294
rect 22480 97294 22614 97322
rect 22480 95674 22508 97294
rect 22558 97200 22614 97294
rect 23124 97294 23258 97322
rect 23124 95674 23152 97294
rect 23202 97200 23258 97294
rect 24412 97294 24546 97322
rect 24412 95674 24440 97294
rect 24490 97200 24546 97294
rect 25700 97294 25834 97322
rect 25700 95674 25728 97294
rect 25778 97200 25834 97294
rect 26988 97294 27122 97322
rect 26988 95674 27016 97294
rect 27066 97200 27122 97294
rect 27632 97294 27766 97322
rect 27632 95674 27660 97294
rect 27710 97200 27766 97294
rect 28998 97322 29054 98000
rect 30286 97322 30342 98000
rect 28998 97294 29132 97322
rect 28998 97200 29054 97294
rect 29104 95674 29132 97294
rect 30208 97294 30342 97322
rect 30208 95674 30236 97294
rect 30286 97200 30342 97294
rect 30930 97322 30986 98000
rect 32218 97322 32274 98000
rect 33506 97322 33562 98000
rect 34794 97322 34850 98000
rect 35438 97322 35494 98000
rect 36726 97322 36782 98000
rect 38014 97322 38070 98000
rect 38658 97322 38714 98000
rect 39946 97322 40002 98000
rect 30930 97294 31156 97322
rect 30930 97200 30986 97294
rect 31128 95674 31156 97294
rect 32218 97294 32536 97322
rect 32218 97200 32274 97294
rect 32508 95674 32536 97294
rect 33506 97294 33824 97322
rect 33506 97200 33562 97294
rect 33796 95674 33824 97294
rect 34794 97294 35112 97322
rect 34794 97200 34850 97294
rect 35084 95674 35112 97294
rect 35438 97294 35664 97322
rect 35438 97200 35494 97294
rect 35636 95674 35664 97294
rect 36726 97294 37044 97322
rect 36726 97200 36782 97294
rect 37016 95674 37044 97294
rect 38014 97294 38332 97322
rect 38014 97200 38070 97294
rect 37610 95772 37918 95781
rect 37610 95770 37616 95772
rect 37672 95770 37696 95772
rect 37752 95770 37776 95772
rect 37832 95770 37856 95772
rect 37912 95770 37918 95772
rect 37672 95718 37674 95770
rect 37854 95718 37856 95770
rect 37610 95716 37616 95718
rect 37672 95716 37696 95718
rect 37752 95716 37776 95718
rect 37832 95716 37856 95718
rect 37912 95716 37918 95718
rect 37610 95707 37918 95716
rect 38304 95674 38332 97294
rect 38658 97294 38884 97322
rect 38658 97200 38714 97294
rect 38856 95674 38884 97294
rect 39868 97294 40002 97322
rect 39868 95674 39896 97294
rect 39946 97200 40002 97294
rect 41234 97322 41290 98000
rect 42522 97322 42578 98000
rect 43166 97322 43222 98000
rect 43442 97336 43498 97345
rect 41234 97294 41368 97322
rect 41234 97200 41290 97294
rect 41340 95674 41368 97294
rect 42522 97294 42748 97322
rect 42522 97200 42578 97294
rect 42720 95674 42748 97294
rect 43166 97294 43392 97322
rect 43166 97200 43222 97294
rect 43364 95674 43392 97294
rect 43442 97271 43498 97280
rect 44454 97322 44510 98000
rect 49330 97336 49386 97345
rect 44454 97294 44772 97322
rect 16672 95668 16724 95674
rect 16672 95610 16724 95616
rect 17960 95668 18012 95674
rect 17960 95610 18012 95616
rect 19432 95668 19484 95674
rect 19432 95610 19484 95616
rect 20352 95668 20404 95674
rect 20352 95610 20404 95616
rect 21180 95668 21232 95674
rect 21180 95610 21232 95616
rect 22468 95668 22520 95674
rect 22468 95610 22520 95616
rect 23112 95668 23164 95674
rect 23112 95610 23164 95616
rect 24400 95668 24452 95674
rect 24400 95610 24452 95616
rect 25688 95668 25740 95674
rect 25688 95610 25740 95616
rect 26976 95668 27028 95674
rect 26976 95610 27028 95616
rect 27620 95668 27672 95674
rect 27620 95610 27672 95616
rect 29092 95668 29144 95674
rect 29092 95610 29144 95616
rect 30196 95668 30248 95674
rect 30196 95610 30248 95616
rect 31116 95668 31168 95674
rect 31116 95610 31168 95616
rect 32496 95668 32548 95674
rect 32496 95610 32548 95616
rect 33784 95668 33836 95674
rect 33784 95610 33836 95616
rect 35072 95668 35124 95674
rect 35072 95610 35124 95616
rect 35624 95668 35676 95674
rect 35624 95610 35676 95616
rect 37004 95668 37056 95674
rect 37004 95610 37056 95616
rect 38292 95668 38344 95674
rect 38292 95610 38344 95616
rect 38844 95668 38896 95674
rect 38844 95610 38896 95616
rect 39856 95668 39908 95674
rect 39856 95610 39908 95616
rect 41328 95668 41380 95674
rect 41328 95610 41380 95616
rect 42708 95668 42760 95674
rect 42708 95610 42760 95616
rect 43352 95668 43404 95674
rect 43352 95610 43404 95616
rect 8484 95532 8536 95538
rect 8484 95474 8536 95480
rect 15568 95532 15620 95538
rect 15568 95474 15620 95480
rect 30104 95532 30156 95538
rect 30104 95474 30156 95480
rect 31300 95532 31352 95538
rect 31300 95474 31352 95480
rect 32312 95532 32364 95538
rect 32312 95474 32364 95480
rect 33600 95532 33652 95538
rect 33600 95474 33652 95480
rect 34888 95532 34940 95538
rect 34888 95474 34940 95480
rect 35808 95532 35860 95538
rect 35808 95474 35860 95480
rect 36820 95532 36872 95538
rect 36820 95474 36872 95480
rect 38108 95532 38160 95538
rect 38108 95474 38160 95480
rect 39028 95532 39080 95538
rect 39028 95474 39080 95480
rect 40040 95532 40092 95538
rect 40040 95474 40092 95480
rect 41328 95532 41380 95538
rect 41328 95474 41380 95480
rect 42616 95532 42668 95538
rect 42616 95474 42668 95480
rect 8496 95305 8524 95474
rect 19064 95464 19116 95470
rect 19064 95406 19116 95412
rect 23572 95464 23624 95470
rect 23572 95406 23624 95412
rect 14648 95328 14700 95334
rect 8482 95296 8538 95305
rect 14648 95270 14700 95276
rect 15752 95328 15804 95334
rect 15752 95270 15804 95276
rect 17040 95328 17092 95334
rect 17040 95270 17092 95276
rect 18328 95328 18380 95334
rect 18328 95270 18380 95276
rect 8482 95231 8538 95240
rect 3066 91964 3374 91973
rect 3066 91962 3072 91964
rect 3128 91962 3152 91964
rect 3208 91962 3232 91964
rect 3288 91962 3312 91964
rect 3368 91962 3374 91964
rect 3128 91910 3130 91962
rect 3310 91910 3312 91962
rect 3066 91908 3072 91910
rect 3128 91908 3152 91910
rect 3208 91908 3232 91910
rect 3288 91908 3312 91910
rect 3368 91908 3374 91910
rect 3066 91899 3374 91908
rect 5632 91588 5684 91594
rect 5632 91530 5684 91536
rect 10324 91588 10376 91594
rect 10324 91530 10376 91536
rect 3802 91420 4110 91429
rect 3802 91418 3808 91420
rect 3864 91418 3888 91420
rect 3944 91418 3968 91420
rect 4024 91418 4048 91420
rect 4104 91418 4110 91420
rect 3864 91366 3866 91418
rect 4046 91366 4048 91418
rect 3802 91364 3808 91366
rect 3864 91364 3888 91366
rect 3944 91364 3968 91366
rect 4024 91364 4048 91366
rect 4104 91364 4110 91366
rect 3802 91355 4110 91364
rect 3066 90876 3374 90885
rect 3066 90874 3072 90876
rect 3128 90874 3152 90876
rect 3208 90874 3232 90876
rect 3288 90874 3312 90876
rect 3368 90874 3374 90876
rect 3128 90822 3130 90874
rect 3310 90822 3312 90874
rect 3066 90820 3072 90822
rect 3128 90820 3152 90822
rect 3208 90820 3232 90822
rect 3288 90820 3312 90822
rect 3368 90820 3374 90822
rect 3066 90811 3374 90820
rect 3802 90332 4110 90341
rect 3802 90330 3808 90332
rect 3864 90330 3888 90332
rect 3944 90330 3968 90332
rect 4024 90330 4048 90332
rect 4104 90330 4110 90332
rect 3864 90278 3866 90330
rect 4046 90278 4048 90330
rect 3802 90276 3808 90278
rect 3864 90276 3888 90278
rect 3944 90276 3968 90278
rect 4024 90276 4048 90278
rect 4104 90276 4110 90278
rect 3802 90267 4110 90276
rect 3066 89788 3374 89797
rect 3066 89786 3072 89788
rect 3128 89786 3152 89788
rect 3208 89786 3232 89788
rect 3288 89786 3312 89788
rect 3368 89786 3374 89788
rect 3128 89734 3130 89786
rect 3310 89734 3312 89786
rect 3066 89732 3072 89734
rect 3128 89732 3152 89734
rect 3208 89732 3232 89734
rect 3288 89732 3312 89734
rect 3368 89732 3374 89734
rect 3066 89723 3374 89732
rect 5172 89344 5224 89350
rect 5172 89286 5224 89292
rect 3802 89244 4110 89253
rect 3802 89242 3808 89244
rect 3864 89242 3888 89244
rect 3944 89242 3968 89244
rect 4024 89242 4048 89244
rect 4104 89242 4110 89244
rect 3864 89190 3866 89242
rect 4046 89190 4048 89242
rect 3802 89188 3808 89190
rect 3864 89188 3888 89190
rect 3944 89188 3968 89190
rect 4024 89188 4048 89190
rect 4104 89188 4110 89190
rect 3802 89179 4110 89188
rect 5080 89004 5132 89010
rect 5080 88946 5132 88952
rect 3066 88700 3374 88709
rect 3066 88698 3072 88700
rect 3128 88698 3152 88700
rect 3208 88698 3232 88700
rect 3288 88698 3312 88700
rect 3368 88698 3374 88700
rect 3128 88646 3130 88698
rect 3310 88646 3312 88698
rect 3066 88644 3072 88646
rect 3128 88644 3152 88646
rect 3208 88644 3232 88646
rect 3288 88644 3312 88646
rect 3368 88644 3374 88646
rect 3066 88635 3374 88644
rect 3802 88156 4110 88165
rect 3802 88154 3808 88156
rect 3864 88154 3888 88156
rect 3944 88154 3968 88156
rect 4024 88154 4048 88156
rect 4104 88154 4110 88156
rect 3864 88102 3866 88154
rect 4046 88102 4048 88154
rect 3802 88100 3808 88102
rect 3864 88100 3888 88102
rect 3944 88100 3968 88102
rect 4024 88100 4048 88102
rect 4104 88100 4110 88102
rect 3802 88091 4110 88100
rect 3066 87612 3374 87621
rect 3066 87610 3072 87612
rect 3128 87610 3152 87612
rect 3208 87610 3232 87612
rect 3288 87610 3312 87612
rect 3368 87610 3374 87612
rect 3128 87558 3130 87610
rect 3310 87558 3312 87610
rect 3066 87556 3072 87558
rect 3128 87556 3152 87558
rect 3208 87556 3232 87558
rect 3288 87556 3312 87558
rect 3368 87556 3374 87558
rect 3066 87547 3374 87556
rect 3802 87068 4110 87077
rect 3802 87066 3808 87068
rect 3864 87066 3888 87068
rect 3944 87066 3968 87068
rect 4024 87066 4048 87068
rect 4104 87066 4110 87068
rect 3864 87014 3866 87066
rect 4046 87014 4048 87066
rect 3802 87012 3808 87014
rect 3864 87012 3888 87014
rect 3944 87012 3968 87014
rect 4024 87012 4048 87014
rect 4104 87012 4110 87014
rect 3802 87003 4110 87012
rect 848 86624 900 86630
rect 846 86592 848 86601
rect 900 86592 902 86601
rect 846 86527 902 86536
rect 3066 86524 3374 86533
rect 3066 86522 3072 86524
rect 3128 86522 3152 86524
rect 3208 86522 3232 86524
rect 3288 86522 3312 86524
rect 3368 86522 3374 86524
rect 3128 86470 3130 86522
rect 3310 86470 3312 86522
rect 3066 86468 3072 86470
rect 3128 86468 3152 86470
rect 3208 86468 3232 86470
rect 3288 86468 3312 86470
rect 3368 86468 3374 86470
rect 3066 86459 3374 86468
rect 3802 85980 4110 85989
rect 3802 85978 3808 85980
rect 3864 85978 3888 85980
rect 3944 85978 3968 85980
rect 4024 85978 4048 85980
rect 4104 85978 4110 85980
rect 3864 85926 3866 85978
rect 4046 85926 4048 85978
rect 3802 85924 3808 85926
rect 3864 85924 3888 85926
rect 3944 85924 3968 85926
rect 4024 85924 4048 85926
rect 4104 85924 4110 85926
rect 3802 85915 4110 85924
rect 3066 85436 3374 85445
rect 3066 85434 3072 85436
rect 3128 85434 3152 85436
rect 3208 85434 3232 85436
rect 3288 85434 3312 85436
rect 3368 85434 3374 85436
rect 3128 85382 3130 85434
rect 3310 85382 3312 85434
rect 3066 85380 3072 85382
rect 3128 85380 3152 85382
rect 3208 85380 3232 85382
rect 3288 85380 3312 85382
rect 3368 85380 3374 85382
rect 3066 85371 3374 85380
rect 848 85264 900 85270
rect 846 85232 848 85241
rect 900 85232 902 85241
rect 846 85167 902 85176
rect 3802 84892 4110 84901
rect 3802 84890 3808 84892
rect 3864 84890 3888 84892
rect 3944 84890 3968 84892
rect 4024 84890 4048 84892
rect 4104 84890 4110 84892
rect 3864 84838 3866 84890
rect 4046 84838 4048 84890
rect 3802 84836 3808 84838
rect 3864 84836 3888 84838
rect 3944 84836 3968 84838
rect 4024 84836 4048 84838
rect 4104 84836 4110 84838
rect 3802 84827 4110 84836
rect 3066 84348 3374 84357
rect 3066 84346 3072 84348
rect 3128 84346 3152 84348
rect 3208 84346 3232 84348
rect 3288 84346 3312 84348
rect 3368 84346 3374 84348
rect 3128 84294 3130 84346
rect 3310 84294 3312 84346
rect 3066 84292 3072 84294
rect 3128 84292 3152 84294
rect 3208 84292 3232 84294
rect 3288 84292 3312 84294
rect 3368 84292 3374 84294
rect 3066 84283 3374 84292
rect 848 83904 900 83910
rect 846 83872 848 83881
rect 900 83872 902 83881
rect 846 83807 902 83816
rect 3802 83804 4110 83813
rect 3802 83802 3808 83804
rect 3864 83802 3888 83804
rect 3944 83802 3968 83804
rect 4024 83802 4048 83804
rect 4104 83802 4110 83804
rect 3864 83750 3866 83802
rect 4046 83750 4048 83802
rect 3802 83748 3808 83750
rect 3864 83748 3888 83750
rect 3944 83748 3968 83750
rect 4024 83748 4048 83750
rect 4104 83748 4110 83750
rect 3802 83739 4110 83748
rect 3066 83260 3374 83269
rect 3066 83258 3072 83260
rect 3128 83258 3152 83260
rect 3208 83258 3232 83260
rect 3288 83258 3312 83260
rect 3368 83258 3374 83260
rect 3128 83206 3130 83258
rect 3310 83206 3312 83258
rect 3066 83204 3072 83206
rect 3128 83204 3152 83206
rect 3208 83204 3232 83206
rect 3288 83204 3312 83206
rect 3368 83204 3374 83206
rect 3066 83195 3374 83204
rect 3802 82716 4110 82725
rect 3802 82714 3808 82716
rect 3864 82714 3888 82716
rect 3944 82714 3968 82716
rect 4024 82714 4048 82716
rect 4104 82714 4110 82716
rect 3864 82662 3866 82714
rect 4046 82662 4048 82714
rect 3802 82660 3808 82662
rect 3864 82660 3888 82662
rect 3944 82660 3968 82662
rect 4024 82660 4048 82662
rect 4104 82660 4110 82662
rect 3802 82651 4110 82660
rect 848 82272 900 82278
rect 846 82240 848 82249
rect 900 82240 902 82249
rect 846 82175 902 82184
rect 3066 82172 3374 82181
rect 3066 82170 3072 82172
rect 3128 82170 3152 82172
rect 3208 82170 3232 82172
rect 3288 82170 3312 82172
rect 3368 82170 3374 82172
rect 3128 82118 3130 82170
rect 3310 82118 3312 82170
rect 3066 82116 3072 82118
rect 3128 82116 3152 82118
rect 3208 82116 3232 82118
rect 3288 82116 3312 82118
rect 3368 82116 3374 82118
rect 3066 82107 3374 82116
rect 3802 81628 4110 81637
rect 3802 81626 3808 81628
rect 3864 81626 3888 81628
rect 3944 81626 3968 81628
rect 4024 81626 4048 81628
rect 4104 81626 4110 81628
rect 3864 81574 3866 81626
rect 4046 81574 4048 81626
rect 3802 81572 3808 81574
rect 3864 81572 3888 81574
rect 3944 81572 3968 81574
rect 4024 81572 4048 81574
rect 4104 81572 4110 81574
rect 3802 81563 4110 81572
rect 848 81184 900 81190
rect 846 81152 848 81161
rect 900 81152 902 81161
rect 846 81087 902 81096
rect 3066 81084 3374 81093
rect 3066 81082 3072 81084
rect 3128 81082 3152 81084
rect 3208 81082 3232 81084
rect 3288 81082 3312 81084
rect 3368 81082 3374 81084
rect 3128 81030 3130 81082
rect 3310 81030 3312 81082
rect 3066 81028 3072 81030
rect 3128 81028 3152 81030
rect 3208 81028 3232 81030
rect 3288 81028 3312 81030
rect 3368 81028 3374 81030
rect 3066 81019 3374 81028
rect 3802 80540 4110 80549
rect 3802 80538 3808 80540
rect 3864 80538 3888 80540
rect 3944 80538 3968 80540
rect 4024 80538 4048 80540
rect 4104 80538 4110 80540
rect 3864 80486 3866 80538
rect 4046 80486 4048 80538
rect 3802 80484 3808 80486
rect 3864 80484 3888 80486
rect 3944 80484 3968 80486
rect 4024 80484 4048 80486
rect 4104 80484 4110 80486
rect 3802 80475 4110 80484
rect 3066 79996 3374 80005
rect 3066 79994 3072 79996
rect 3128 79994 3152 79996
rect 3208 79994 3232 79996
rect 3288 79994 3312 79996
rect 3368 79994 3374 79996
rect 3128 79942 3130 79994
rect 3310 79942 3312 79994
rect 3066 79940 3072 79942
rect 3128 79940 3152 79942
rect 3208 79940 3232 79942
rect 3288 79940 3312 79942
rect 3368 79940 3374 79942
rect 3066 79931 3374 79940
rect 848 79552 900 79558
rect 846 79520 848 79529
rect 900 79520 902 79529
rect 846 79455 902 79464
rect 3802 79452 4110 79461
rect 3802 79450 3808 79452
rect 3864 79450 3888 79452
rect 3944 79450 3968 79452
rect 4024 79450 4048 79452
rect 4104 79450 4110 79452
rect 3864 79398 3866 79450
rect 4046 79398 4048 79450
rect 3802 79396 3808 79398
rect 3864 79396 3888 79398
rect 3944 79396 3968 79398
rect 4024 79396 4048 79398
rect 4104 79396 4110 79398
rect 3802 79387 4110 79396
rect 3066 78908 3374 78917
rect 3066 78906 3072 78908
rect 3128 78906 3152 78908
rect 3208 78906 3232 78908
rect 3288 78906 3312 78908
rect 3368 78906 3374 78908
rect 3128 78854 3130 78906
rect 3310 78854 3312 78906
rect 3066 78852 3072 78854
rect 3128 78852 3152 78854
rect 3208 78852 3232 78854
rect 3288 78852 3312 78854
rect 3368 78852 3374 78854
rect 3066 78843 3374 78852
rect 848 78464 900 78470
rect 846 78432 848 78441
rect 900 78432 902 78441
rect 846 78367 902 78376
rect 3802 78364 4110 78373
rect 3802 78362 3808 78364
rect 3864 78362 3888 78364
rect 3944 78362 3968 78364
rect 4024 78362 4048 78364
rect 4104 78362 4110 78364
rect 3864 78310 3866 78362
rect 4046 78310 4048 78362
rect 3802 78308 3808 78310
rect 3864 78308 3888 78310
rect 3944 78308 3968 78310
rect 4024 78308 4048 78310
rect 4104 78308 4110 78310
rect 3802 78299 4110 78308
rect 3066 77820 3374 77829
rect 3066 77818 3072 77820
rect 3128 77818 3152 77820
rect 3208 77818 3232 77820
rect 3288 77818 3312 77820
rect 3368 77818 3374 77820
rect 3128 77766 3130 77818
rect 3310 77766 3312 77818
rect 3066 77764 3072 77766
rect 3128 77764 3152 77766
rect 3208 77764 3232 77766
rect 3288 77764 3312 77766
rect 3368 77764 3374 77766
rect 3066 77755 3374 77764
rect 3802 77276 4110 77285
rect 3802 77274 3808 77276
rect 3864 77274 3888 77276
rect 3944 77274 3968 77276
rect 4024 77274 4048 77276
rect 4104 77274 4110 77276
rect 3864 77222 3866 77274
rect 4046 77222 4048 77274
rect 3802 77220 3808 77222
rect 3864 77220 3888 77222
rect 3944 77220 3968 77222
rect 4024 77220 4048 77222
rect 4104 77220 4110 77222
rect 3802 77211 4110 77220
rect 848 76832 900 76838
rect 846 76800 848 76809
rect 900 76800 902 76809
rect 846 76735 902 76744
rect 3066 76732 3374 76741
rect 3066 76730 3072 76732
rect 3128 76730 3152 76732
rect 3208 76730 3232 76732
rect 3288 76730 3312 76732
rect 3368 76730 3374 76732
rect 3128 76678 3130 76730
rect 3310 76678 3312 76730
rect 3066 76676 3072 76678
rect 3128 76676 3152 76678
rect 3208 76676 3232 76678
rect 3288 76676 3312 76678
rect 3368 76676 3374 76678
rect 3066 76667 3374 76676
rect 3802 76188 4110 76197
rect 3802 76186 3808 76188
rect 3864 76186 3888 76188
rect 3944 76186 3968 76188
rect 4024 76186 4048 76188
rect 4104 76186 4110 76188
rect 3864 76134 3866 76186
rect 4046 76134 4048 76186
rect 3802 76132 3808 76134
rect 3864 76132 3888 76134
rect 3944 76132 3968 76134
rect 4024 76132 4048 76134
rect 4104 76132 4110 76134
rect 3802 76123 4110 76132
rect 848 76084 900 76090
rect 848 76026 900 76032
rect 860 75721 888 76026
rect 846 75712 902 75721
rect 846 75647 902 75656
rect 3066 75644 3374 75653
rect 3066 75642 3072 75644
rect 3128 75642 3152 75644
rect 3208 75642 3232 75644
rect 3288 75642 3312 75644
rect 3368 75642 3374 75644
rect 3128 75590 3130 75642
rect 3310 75590 3312 75642
rect 3066 75588 3072 75590
rect 3128 75588 3152 75590
rect 3208 75588 3232 75590
rect 3288 75588 3312 75590
rect 3368 75588 3374 75590
rect 3066 75579 3374 75588
rect 3802 75100 4110 75109
rect 3802 75098 3808 75100
rect 3864 75098 3888 75100
rect 3944 75098 3968 75100
rect 4024 75098 4048 75100
rect 4104 75098 4110 75100
rect 3864 75046 3866 75098
rect 4046 75046 4048 75098
rect 3802 75044 3808 75046
rect 3864 75044 3888 75046
rect 3944 75044 3968 75046
rect 4024 75044 4048 75046
rect 4104 75044 4110 75046
rect 3802 75035 4110 75044
rect 3066 74556 3374 74565
rect 3066 74554 3072 74556
rect 3128 74554 3152 74556
rect 3208 74554 3232 74556
rect 3288 74554 3312 74556
rect 3368 74554 3374 74556
rect 3128 74502 3130 74554
rect 3310 74502 3312 74554
rect 3066 74500 3072 74502
rect 3128 74500 3152 74502
rect 3208 74500 3232 74502
rect 3288 74500 3312 74502
rect 3368 74500 3374 74502
rect 3066 74491 3374 74500
rect 848 74112 900 74118
rect 846 74080 848 74089
rect 900 74080 902 74089
rect 846 74015 902 74024
rect 3802 74012 4110 74021
rect 3802 74010 3808 74012
rect 3864 74010 3888 74012
rect 3944 74010 3968 74012
rect 4024 74010 4048 74012
rect 4104 74010 4110 74012
rect 3864 73958 3866 74010
rect 4046 73958 4048 74010
rect 3802 73956 3808 73958
rect 3864 73956 3888 73958
rect 3944 73956 3968 73958
rect 4024 73956 4048 73958
rect 4104 73956 4110 73958
rect 3802 73947 4110 73956
rect 3066 73468 3374 73477
rect 3066 73466 3072 73468
rect 3128 73466 3152 73468
rect 3208 73466 3232 73468
rect 3288 73466 3312 73468
rect 3368 73466 3374 73468
rect 3128 73414 3130 73466
rect 3310 73414 3312 73466
rect 3066 73412 3072 73414
rect 3128 73412 3152 73414
rect 3208 73412 3232 73414
rect 3288 73412 3312 73414
rect 3368 73412 3374 73414
rect 3066 73403 3374 73412
rect 848 73024 900 73030
rect 846 72992 848 73001
rect 900 72992 902 73001
rect 846 72927 902 72936
rect 3802 72924 4110 72933
rect 3802 72922 3808 72924
rect 3864 72922 3888 72924
rect 3944 72922 3968 72924
rect 4024 72922 4048 72924
rect 4104 72922 4110 72924
rect 3864 72870 3866 72922
rect 4046 72870 4048 72922
rect 3802 72868 3808 72870
rect 3864 72868 3888 72870
rect 3944 72868 3968 72870
rect 4024 72868 4048 72870
rect 4104 72868 4110 72870
rect 3802 72859 4110 72868
rect 3066 72380 3374 72389
rect 3066 72378 3072 72380
rect 3128 72378 3152 72380
rect 3208 72378 3232 72380
rect 3288 72378 3312 72380
rect 3368 72378 3374 72380
rect 3128 72326 3130 72378
rect 3310 72326 3312 72378
rect 3066 72324 3072 72326
rect 3128 72324 3152 72326
rect 3208 72324 3232 72326
rect 3288 72324 3312 72326
rect 3368 72324 3374 72326
rect 3066 72315 3374 72324
rect 3802 71836 4110 71845
rect 3802 71834 3808 71836
rect 3864 71834 3888 71836
rect 3944 71834 3968 71836
rect 4024 71834 4048 71836
rect 4104 71834 4110 71836
rect 3864 71782 3866 71834
rect 4046 71782 4048 71834
rect 3802 71780 3808 71782
rect 3864 71780 3888 71782
rect 3944 71780 3968 71782
rect 4024 71780 4048 71782
rect 4104 71780 4110 71782
rect 3802 71771 4110 71780
rect 4620 71460 4672 71466
rect 4620 71402 4672 71408
rect 848 71392 900 71398
rect 846 71360 848 71369
rect 900 71360 902 71369
rect 846 71295 902 71304
rect 3066 71292 3374 71301
rect 3066 71290 3072 71292
rect 3128 71290 3152 71292
rect 3208 71290 3232 71292
rect 3288 71290 3312 71292
rect 3368 71290 3374 71292
rect 3128 71238 3130 71290
rect 3310 71238 3312 71290
rect 3066 71236 3072 71238
rect 3128 71236 3152 71238
rect 3208 71236 3232 71238
rect 3288 71236 3312 71238
rect 3368 71236 3374 71238
rect 3066 71227 3374 71236
rect 3802 70748 4110 70757
rect 3802 70746 3808 70748
rect 3864 70746 3888 70748
rect 3944 70746 3968 70748
rect 4024 70746 4048 70748
rect 4104 70746 4110 70748
rect 3864 70694 3866 70746
rect 4046 70694 4048 70746
rect 3802 70692 3808 70694
rect 3864 70692 3888 70694
rect 3944 70692 3968 70694
rect 4024 70692 4048 70694
rect 4104 70692 4110 70694
rect 3802 70683 4110 70692
rect 848 70644 900 70650
rect 848 70586 900 70592
rect 860 70281 888 70586
rect 846 70272 902 70281
rect 846 70207 902 70216
rect 3066 70204 3374 70213
rect 3066 70202 3072 70204
rect 3128 70202 3152 70204
rect 3208 70202 3232 70204
rect 3288 70202 3312 70204
rect 3368 70202 3374 70204
rect 3128 70150 3130 70202
rect 3310 70150 3312 70202
rect 3066 70148 3072 70150
rect 3128 70148 3152 70150
rect 3208 70148 3232 70150
rect 3288 70148 3312 70150
rect 3368 70148 3374 70150
rect 3066 70139 3374 70148
rect 3802 69660 4110 69669
rect 3802 69658 3808 69660
rect 3864 69658 3888 69660
rect 3944 69658 3968 69660
rect 4024 69658 4048 69660
rect 4104 69658 4110 69660
rect 3864 69606 3866 69658
rect 4046 69606 4048 69658
rect 3802 69604 3808 69606
rect 3864 69604 3888 69606
rect 3944 69604 3968 69606
rect 4024 69604 4048 69606
rect 4104 69604 4110 69606
rect 3802 69595 4110 69604
rect 3066 69116 3374 69125
rect 3066 69114 3072 69116
rect 3128 69114 3152 69116
rect 3208 69114 3232 69116
rect 3288 69114 3312 69116
rect 3368 69114 3374 69116
rect 3128 69062 3130 69114
rect 3310 69062 3312 69114
rect 3066 69060 3072 69062
rect 3128 69060 3152 69062
rect 3208 69060 3232 69062
rect 3288 69060 3312 69062
rect 3368 69060 3374 69062
rect 3066 69051 3374 69060
rect 1216 68808 1268 68814
rect 1214 68776 1216 68785
rect 1268 68776 1270 68785
rect 1214 68711 1270 68720
rect 3802 68572 4110 68581
rect 3802 68570 3808 68572
rect 3864 68570 3888 68572
rect 3944 68570 3968 68572
rect 4024 68570 4048 68572
rect 4104 68570 4110 68572
rect 3864 68518 3866 68570
rect 4046 68518 4048 68570
rect 3802 68516 3808 68518
rect 3864 68516 3888 68518
rect 3944 68516 3968 68518
rect 4024 68516 4048 68518
rect 4104 68516 4110 68518
rect 3802 68507 4110 68516
rect 3066 68028 3374 68037
rect 3066 68026 3072 68028
rect 3128 68026 3152 68028
rect 3208 68026 3232 68028
rect 3288 68026 3312 68028
rect 3368 68026 3374 68028
rect 3128 67974 3130 68026
rect 3310 67974 3312 68026
rect 3066 67972 3072 67974
rect 3128 67972 3152 67974
rect 3208 67972 3232 67974
rect 3288 67972 3312 67974
rect 3368 67972 3374 67974
rect 3066 67963 3374 67972
rect 1308 67720 1360 67726
rect 1308 67662 1360 67668
rect 1320 67425 1348 67662
rect 3802 67484 4110 67493
rect 3802 67482 3808 67484
rect 3864 67482 3888 67484
rect 3944 67482 3968 67484
rect 4024 67482 4048 67484
rect 4104 67482 4110 67484
rect 3864 67430 3866 67482
rect 4046 67430 4048 67482
rect 3802 67428 3808 67430
rect 3864 67428 3888 67430
rect 3944 67428 3968 67430
rect 4024 67428 4048 67430
rect 4104 67428 4110 67430
rect 1306 67416 1362 67425
rect 3802 67419 4110 67428
rect 1306 67351 1362 67360
rect 3066 66940 3374 66949
rect 3066 66938 3072 66940
rect 3128 66938 3152 66940
rect 3208 66938 3232 66940
rect 3288 66938 3312 66940
rect 3368 66938 3374 66940
rect 3128 66886 3130 66938
rect 3310 66886 3312 66938
rect 3066 66884 3072 66886
rect 3128 66884 3152 66886
rect 3208 66884 3232 66886
rect 3288 66884 3312 66886
rect 3368 66884 3374 66886
rect 3066 66875 3374 66884
rect 3802 66396 4110 66405
rect 3802 66394 3808 66396
rect 3864 66394 3888 66396
rect 3944 66394 3968 66396
rect 4024 66394 4048 66396
rect 4104 66394 4110 66396
rect 3864 66342 3866 66394
rect 4046 66342 4048 66394
rect 3802 66340 3808 66342
rect 3864 66340 3888 66342
rect 3944 66340 3968 66342
rect 4024 66340 4048 66342
rect 4104 66340 4110 66342
rect 3802 66331 4110 66340
rect 1308 66156 1360 66162
rect 1308 66098 1360 66104
rect 1320 66065 1348 66098
rect 1306 66056 1362 66065
rect 1306 65991 1362 66000
rect 3066 65852 3374 65861
rect 3066 65850 3072 65852
rect 3128 65850 3152 65852
rect 3208 65850 3232 65852
rect 3288 65850 3312 65852
rect 3368 65850 3374 65852
rect 3128 65798 3130 65850
rect 3310 65798 3312 65850
rect 3066 65796 3072 65798
rect 3128 65796 3152 65798
rect 3208 65796 3232 65798
rect 3288 65796 3312 65798
rect 3368 65796 3374 65798
rect 3066 65787 3374 65796
rect 3802 65308 4110 65317
rect 3802 65306 3808 65308
rect 3864 65306 3888 65308
rect 3944 65306 3968 65308
rect 4024 65306 4048 65308
rect 4104 65306 4110 65308
rect 3864 65254 3866 65306
rect 4046 65254 4048 65306
rect 3802 65252 3808 65254
rect 3864 65252 3888 65254
rect 3944 65252 3968 65254
rect 4024 65252 4048 65254
rect 4104 65252 4110 65254
rect 3802 65243 4110 65252
rect 1308 65068 1360 65074
rect 1308 65010 1360 65016
rect 1320 64705 1348 65010
rect 3066 64764 3374 64773
rect 3066 64762 3072 64764
rect 3128 64762 3152 64764
rect 3208 64762 3232 64764
rect 3288 64762 3312 64764
rect 3368 64762 3374 64764
rect 3128 64710 3130 64762
rect 3310 64710 3312 64762
rect 3066 64708 3072 64710
rect 3128 64708 3152 64710
rect 3208 64708 3232 64710
rect 3288 64708 3312 64710
rect 3368 64708 3374 64710
rect 1306 64696 1362 64705
rect 3066 64699 3374 64708
rect 1306 64631 1362 64640
rect 3802 64220 4110 64229
rect 3802 64218 3808 64220
rect 3864 64218 3888 64220
rect 3944 64218 3968 64220
rect 4024 64218 4048 64220
rect 4104 64218 4110 64220
rect 3864 64166 3866 64218
rect 4046 64166 4048 64218
rect 3802 64164 3808 64166
rect 3864 64164 3888 64166
rect 3944 64164 3968 64166
rect 4024 64164 4048 64166
rect 4104 64164 4110 64166
rect 3802 64155 4110 64164
rect 3066 63676 3374 63685
rect 3066 63674 3072 63676
rect 3128 63674 3152 63676
rect 3208 63674 3232 63676
rect 3288 63674 3312 63676
rect 3368 63674 3374 63676
rect 3128 63622 3130 63674
rect 3310 63622 3312 63674
rect 3066 63620 3072 63622
rect 3128 63620 3152 63622
rect 3208 63620 3232 63622
rect 3288 63620 3312 63622
rect 3368 63620 3374 63622
rect 3066 63611 3374 63620
rect 1216 63368 1268 63374
rect 1214 63336 1216 63345
rect 1268 63336 1270 63345
rect 1214 63271 1270 63280
rect 4528 63232 4580 63238
rect 4528 63174 4580 63180
rect 3802 63132 4110 63141
rect 3802 63130 3808 63132
rect 3864 63130 3888 63132
rect 3944 63130 3968 63132
rect 4024 63130 4048 63132
rect 4104 63130 4110 63132
rect 3864 63078 3866 63130
rect 4046 63078 4048 63130
rect 3802 63076 3808 63078
rect 3864 63076 3888 63078
rect 3944 63076 3968 63078
rect 4024 63076 4048 63078
rect 4104 63076 4110 63078
rect 3802 63067 4110 63076
rect 3066 62588 3374 62597
rect 3066 62586 3072 62588
rect 3128 62586 3152 62588
rect 3208 62586 3232 62588
rect 3288 62586 3312 62588
rect 3368 62586 3374 62588
rect 3128 62534 3130 62586
rect 3310 62534 3312 62586
rect 3066 62532 3072 62534
rect 3128 62532 3152 62534
rect 3208 62532 3232 62534
rect 3288 62532 3312 62534
rect 3368 62532 3374 62534
rect 3066 62523 3374 62532
rect 1308 62280 1360 62286
rect 1308 62222 1360 62228
rect 1320 61985 1348 62222
rect 3802 62044 4110 62053
rect 3802 62042 3808 62044
rect 3864 62042 3888 62044
rect 3944 62042 3968 62044
rect 4024 62042 4048 62044
rect 4104 62042 4110 62044
rect 3864 61990 3866 62042
rect 4046 61990 4048 62042
rect 3802 61988 3808 61990
rect 3864 61988 3888 61990
rect 3944 61988 3968 61990
rect 4024 61988 4048 61990
rect 4104 61988 4110 61990
rect 1306 61976 1362 61985
rect 3802 61979 4110 61988
rect 1306 61911 1362 61920
rect 1308 61804 1360 61810
rect 1308 61746 1360 61752
rect 1320 61305 1348 61746
rect 3066 61500 3374 61509
rect 3066 61498 3072 61500
rect 3128 61498 3152 61500
rect 3208 61498 3232 61500
rect 3288 61498 3312 61500
rect 3368 61498 3374 61500
rect 3128 61446 3130 61498
rect 3310 61446 3312 61498
rect 3066 61444 3072 61446
rect 3128 61444 3152 61446
rect 3208 61444 3232 61446
rect 3288 61444 3312 61446
rect 3368 61444 3374 61446
rect 3066 61435 3374 61444
rect 1306 61296 1362 61305
rect 1306 61231 1362 61240
rect 3802 60956 4110 60965
rect 3802 60954 3808 60956
rect 3864 60954 3888 60956
rect 3944 60954 3968 60956
rect 4024 60954 4048 60956
rect 4104 60954 4110 60956
rect 3864 60902 3866 60954
rect 4046 60902 4048 60954
rect 3802 60900 3808 60902
rect 3864 60900 3888 60902
rect 3944 60900 3968 60902
rect 4024 60900 4048 60902
rect 4104 60900 4110 60902
rect 3802 60891 4110 60900
rect 848 60512 900 60518
rect 846 60480 848 60489
rect 900 60480 902 60489
rect 846 60415 902 60424
rect 3066 60412 3374 60421
rect 3066 60410 3072 60412
rect 3128 60410 3152 60412
rect 3208 60410 3232 60412
rect 3288 60410 3312 60412
rect 3368 60410 3374 60412
rect 3128 60358 3130 60410
rect 3310 60358 3312 60410
rect 3066 60356 3072 60358
rect 3128 60356 3152 60358
rect 3208 60356 3232 60358
rect 3288 60356 3312 60358
rect 3368 60356 3374 60358
rect 3066 60347 3374 60356
rect 1216 60104 1268 60110
rect 1216 60046 1268 60052
rect 1228 59945 1256 60046
rect 1214 59936 1270 59945
rect 1214 59871 1270 59880
rect 3802 59868 4110 59877
rect 3802 59866 3808 59868
rect 3864 59866 3888 59868
rect 3944 59866 3968 59868
rect 4024 59866 4048 59868
rect 4104 59866 4110 59868
rect 3864 59814 3866 59866
rect 4046 59814 4048 59866
rect 3802 59812 3808 59814
rect 3864 59812 3888 59814
rect 3944 59812 3968 59814
rect 4024 59812 4048 59814
rect 4104 59812 4110 59814
rect 3802 59803 4110 59812
rect 848 59424 900 59430
rect 848 59366 900 59372
rect 860 59129 888 59366
rect 3066 59324 3374 59333
rect 3066 59322 3072 59324
rect 3128 59322 3152 59324
rect 3208 59322 3232 59324
rect 3288 59322 3312 59324
rect 3368 59322 3374 59324
rect 3128 59270 3130 59322
rect 3310 59270 3312 59322
rect 3066 59268 3072 59270
rect 3128 59268 3152 59270
rect 3208 59268 3232 59270
rect 3288 59268 3312 59270
rect 3368 59268 3374 59270
rect 3066 59259 3374 59268
rect 846 59120 902 59129
rect 846 59055 902 59064
rect 1308 59016 1360 59022
rect 1308 58958 1360 58964
rect 1320 58585 1348 58958
rect 3802 58780 4110 58789
rect 3802 58778 3808 58780
rect 3864 58778 3888 58780
rect 3944 58778 3968 58780
rect 4024 58778 4048 58780
rect 4104 58778 4110 58780
rect 3864 58726 3866 58778
rect 4046 58726 4048 58778
rect 3802 58724 3808 58726
rect 3864 58724 3888 58726
rect 3944 58724 3968 58726
rect 4024 58724 4048 58726
rect 4104 58724 4110 58726
rect 3802 58715 4110 58724
rect 1306 58576 1362 58585
rect 1306 58511 1362 58520
rect 3066 58236 3374 58245
rect 3066 58234 3072 58236
rect 3128 58234 3152 58236
rect 3208 58234 3232 58236
rect 3288 58234 3312 58236
rect 3368 58234 3374 58236
rect 3128 58182 3130 58234
rect 3310 58182 3312 58234
rect 3066 58180 3072 58182
rect 3128 58180 3152 58182
rect 3208 58180 3232 58182
rect 3288 58180 3312 58182
rect 3368 58180 3374 58182
rect 3066 58171 3374 58180
rect 848 57996 900 58002
rect 848 57938 900 57944
rect 860 57769 888 57938
rect 846 57760 902 57769
rect 846 57695 902 57704
rect 3802 57692 4110 57701
rect 3802 57690 3808 57692
rect 3864 57690 3888 57692
rect 3944 57690 3968 57692
rect 4024 57690 4048 57692
rect 4104 57690 4110 57692
rect 3864 57638 3866 57690
rect 4046 57638 4048 57690
rect 3802 57636 3808 57638
rect 3864 57636 3888 57638
rect 3944 57636 3968 57638
rect 4024 57636 4048 57638
rect 4104 57636 4110 57638
rect 3802 57627 4110 57636
rect 1308 57452 1360 57458
rect 1308 57394 1360 57400
rect 1320 57225 1348 57394
rect 1306 57216 1362 57225
rect 1306 57151 1362 57160
rect 3066 57148 3374 57157
rect 3066 57146 3072 57148
rect 3128 57146 3152 57148
rect 3208 57146 3232 57148
rect 3288 57146 3312 57148
rect 3368 57146 3374 57148
rect 3128 57094 3130 57146
rect 3310 57094 3312 57146
rect 3066 57092 3072 57094
rect 3128 57092 3152 57094
rect 3208 57092 3232 57094
rect 3288 57092 3312 57094
rect 3368 57092 3374 57094
rect 3066 57083 3374 57092
rect 848 56840 900 56846
rect 848 56782 900 56788
rect 860 56409 888 56782
rect 3802 56604 4110 56613
rect 3802 56602 3808 56604
rect 3864 56602 3888 56604
rect 3944 56602 3968 56604
rect 4024 56602 4048 56604
rect 4104 56602 4110 56604
rect 3864 56550 3866 56602
rect 4046 56550 4048 56602
rect 3802 56548 3808 56550
rect 3864 56548 3888 56550
rect 3944 56548 3968 56550
rect 4024 56548 4048 56550
rect 4104 56548 4110 56550
rect 3802 56539 4110 56548
rect 846 56400 902 56409
rect 846 56335 902 56344
rect 1308 56364 1360 56370
rect 1308 56306 1360 56312
rect 1320 55865 1348 56306
rect 3066 56060 3374 56069
rect 3066 56058 3072 56060
rect 3128 56058 3152 56060
rect 3208 56058 3232 56060
rect 3288 56058 3312 56060
rect 3368 56058 3374 56060
rect 3128 56006 3130 56058
rect 3310 56006 3312 56058
rect 3066 56004 3072 56006
rect 3128 56004 3152 56006
rect 3208 56004 3232 56006
rect 3288 56004 3312 56006
rect 3368 56004 3374 56006
rect 3066 55995 3374 56004
rect 1306 55856 1362 55865
rect 1306 55791 1362 55800
rect 3802 55516 4110 55525
rect 3802 55514 3808 55516
rect 3864 55514 3888 55516
rect 3944 55514 3968 55516
rect 4024 55514 4048 55516
rect 4104 55514 4110 55516
rect 3864 55462 3866 55514
rect 4046 55462 4048 55514
rect 3802 55460 3808 55462
rect 3864 55460 3888 55462
rect 3944 55460 3968 55462
rect 4024 55460 4048 55462
rect 4104 55460 4110 55462
rect 3802 55451 4110 55460
rect 848 55072 900 55078
rect 846 55040 848 55049
rect 900 55040 902 55049
rect 846 54975 902 54984
rect 3066 54972 3374 54981
rect 3066 54970 3072 54972
rect 3128 54970 3152 54972
rect 3208 54970 3232 54972
rect 3288 54970 3312 54972
rect 3368 54970 3374 54972
rect 3128 54918 3130 54970
rect 3310 54918 3312 54970
rect 3066 54916 3072 54918
rect 3128 54916 3152 54918
rect 3208 54916 3232 54918
rect 3288 54916 3312 54918
rect 3368 54916 3374 54918
rect 3066 54907 3374 54916
rect 1216 54664 1268 54670
rect 1216 54606 1268 54612
rect 1228 54505 1256 54606
rect 1214 54496 1270 54505
rect 1214 54431 1270 54440
rect 3802 54428 4110 54437
rect 3802 54426 3808 54428
rect 3864 54426 3888 54428
rect 3944 54426 3968 54428
rect 4024 54426 4048 54428
rect 4104 54426 4110 54428
rect 3864 54374 3866 54426
rect 4046 54374 4048 54426
rect 3802 54372 3808 54374
rect 3864 54372 3888 54374
rect 3944 54372 3968 54374
rect 4024 54372 4048 54374
rect 4104 54372 4110 54374
rect 3802 54363 4110 54372
rect 848 53984 900 53990
rect 848 53926 900 53932
rect 860 53689 888 53926
rect 3066 53884 3374 53893
rect 3066 53882 3072 53884
rect 3128 53882 3152 53884
rect 3208 53882 3232 53884
rect 3288 53882 3312 53884
rect 3368 53882 3374 53884
rect 3128 53830 3130 53882
rect 3310 53830 3312 53882
rect 3066 53828 3072 53830
rect 3128 53828 3152 53830
rect 3208 53828 3232 53830
rect 3288 53828 3312 53830
rect 3368 53828 3374 53830
rect 3066 53819 3374 53828
rect 846 53680 902 53689
rect 846 53615 902 53624
rect 1308 53576 1360 53582
rect 1308 53518 1360 53524
rect 1320 53145 1348 53518
rect 3802 53340 4110 53349
rect 3802 53338 3808 53340
rect 3864 53338 3888 53340
rect 3944 53338 3968 53340
rect 4024 53338 4048 53340
rect 4104 53338 4110 53340
rect 3864 53286 3866 53338
rect 4046 53286 4048 53338
rect 3802 53284 3808 53286
rect 3864 53284 3888 53286
rect 3944 53284 3968 53286
rect 4024 53284 4048 53286
rect 4104 53284 4110 53286
rect 3802 53275 4110 53284
rect 1306 53136 1362 53145
rect 1306 53071 1362 53080
rect 3066 52796 3374 52805
rect 3066 52794 3072 52796
rect 3128 52794 3152 52796
rect 3208 52794 3232 52796
rect 3288 52794 3312 52796
rect 3368 52794 3374 52796
rect 3128 52742 3130 52794
rect 3310 52742 3312 52794
rect 3066 52740 3072 52742
rect 3128 52740 3152 52742
rect 3208 52740 3232 52742
rect 3288 52740 3312 52742
rect 3368 52740 3374 52742
rect 3066 52731 3374 52740
rect 848 52488 900 52494
rect 848 52430 900 52436
rect 860 52329 888 52430
rect 846 52320 902 52329
rect 846 52255 902 52264
rect 3802 52252 4110 52261
rect 3802 52250 3808 52252
rect 3864 52250 3888 52252
rect 3944 52250 3968 52252
rect 4024 52250 4048 52252
rect 4104 52250 4110 52252
rect 3864 52198 3866 52250
rect 4046 52198 4048 52250
rect 3802 52196 3808 52198
rect 3864 52196 3888 52198
rect 3944 52196 3968 52198
rect 4024 52196 4048 52198
rect 4104 52196 4110 52198
rect 3802 52187 4110 52196
rect 848 51944 900 51950
rect 846 51912 848 51921
rect 900 51912 902 51921
rect 846 51847 902 51856
rect 3066 51708 3374 51717
rect 3066 51706 3072 51708
rect 3128 51706 3152 51708
rect 3208 51706 3232 51708
rect 3288 51706 3312 51708
rect 3368 51706 3374 51708
rect 3128 51654 3130 51706
rect 3310 51654 3312 51706
rect 3066 51652 3072 51654
rect 3128 51652 3152 51654
rect 3208 51652 3232 51654
rect 3288 51652 3312 51654
rect 3368 51652 3374 51654
rect 3066 51643 3374 51652
rect 1032 51400 1084 51406
rect 1032 51342 1084 51348
rect 1582 51368 1638 51377
rect 1044 51105 1072 51342
rect 1582 51303 1638 51312
rect 1030 51096 1086 51105
rect 1030 51031 1086 51040
rect 1400 50720 1452 50726
rect 1400 50662 1452 50668
rect 1412 50561 1440 50662
rect 1398 50552 1454 50561
rect 1398 50487 1454 50496
rect 1400 49632 1452 49638
rect 1400 49574 1452 49580
rect 1412 49473 1440 49574
rect 1398 49464 1454 49473
rect 1398 49399 1454 49408
rect 1400 49360 1452 49366
rect 1398 49328 1400 49337
rect 1452 49328 1454 49337
rect 1398 49263 1454 49272
rect 1596 48890 1624 51303
rect 3802 51164 4110 51173
rect 3802 51162 3808 51164
rect 3864 51162 3888 51164
rect 3944 51162 3968 51164
rect 4024 51162 4048 51164
rect 4104 51162 4110 51164
rect 3864 51110 3866 51162
rect 4046 51110 4048 51162
rect 3802 51108 3808 51110
rect 3864 51108 3888 51110
rect 3944 51108 3968 51110
rect 4024 51108 4048 51110
rect 4104 51108 4110 51110
rect 3802 51099 4110 51108
rect 3066 50620 3374 50629
rect 3066 50618 3072 50620
rect 3128 50618 3152 50620
rect 3208 50618 3232 50620
rect 3288 50618 3312 50620
rect 3368 50618 3374 50620
rect 3128 50566 3130 50618
rect 3310 50566 3312 50618
rect 3066 50564 3072 50566
rect 3128 50564 3152 50566
rect 3208 50564 3232 50566
rect 3288 50564 3312 50566
rect 3368 50564 3374 50566
rect 3066 50555 3374 50564
rect 3802 50076 4110 50085
rect 3802 50074 3808 50076
rect 3864 50074 3888 50076
rect 3944 50074 3968 50076
rect 4024 50074 4048 50076
rect 4104 50074 4110 50076
rect 3864 50022 3866 50074
rect 4046 50022 4048 50074
rect 3802 50020 3808 50022
rect 3864 50020 3888 50022
rect 3944 50020 3968 50022
rect 4024 50020 4048 50022
rect 4104 50020 4110 50022
rect 3802 50011 4110 50020
rect 3066 49532 3374 49541
rect 3066 49530 3072 49532
rect 3128 49530 3152 49532
rect 3208 49530 3232 49532
rect 3288 49530 3312 49532
rect 3368 49530 3374 49532
rect 3128 49478 3130 49530
rect 3310 49478 3312 49530
rect 3066 49476 3072 49478
rect 3128 49476 3152 49478
rect 3208 49476 3232 49478
rect 3288 49476 3312 49478
rect 3368 49476 3374 49478
rect 3066 49467 3374 49476
rect 4540 49337 4568 63174
rect 4632 49910 4660 71402
rect 5092 70650 5120 88946
rect 5080 70644 5132 70650
rect 5080 70586 5132 70592
rect 4896 66156 4948 66162
rect 4896 66098 4948 66104
rect 4908 65958 4936 66098
rect 4896 65952 4948 65958
rect 4896 65894 4948 65900
rect 4908 60058 4936 65894
rect 5184 60722 5212 89286
rect 5356 89140 5408 89146
rect 5356 89082 5408 89088
rect 5264 88392 5316 88398
rect 5264 88334 5316 88340
rect 5276 62490 5304 88334
rect 5368 65210 5396 89082
rect 5448 89072 5500 89078
rect 5448 89014 5500 89020
rect 5460 67862 5488 89014
rect 5540 75948 5592 75954
rect 5540 75890 5592 75896
rect 5552 75721 5580 75890
rect 5538 75712 5594 75721
rect 5538 75647 5594 75656
rect 5540 70508 5592 70514
rect 5540 70450 5592 70456
rect 5552 70281 5580 70450
rect 5538 70272 5594 70281
rect 5538 70207 5594 70216
rect 5448 67856 5500 67862
rect 5448 67798 5500 67804
rect 5540 67856 5592 67862
rect 5540 67798 5592 67804
rect 5552 67697 5580 67798
rect 5538 67688 5594 67697
rect 5538 67623 5594 67632
rect 5356 65204 5408 65210
rect 5356 65146 5408 65152
rect 5538 64968 5594 64977
rect 5538 64903 5540 64912
rect 5592 64903 5594 64912
rect 5540 64874 5592 64880
rect 5264 62484 5316 62490
rect 5264 62426 5316 62432
rect 5276 62286 5304 62426
rect 5540 62416 5592 62422
rect 5540 62358 5592 62364
rect 5264 62280 5316 62286
rect 5264 62222 5316 62228
rect 5552 62121 5580 62358
rect 5538 62112 5594 62121
rect 5538 62047 5594 62056
rect 5172 60716 5224 60722
rect 5172 60658 5224 60664
rect 4816 60030 4936 60058
rect 4712 54324 4764 54330
rect 4712 54266 4764 54272
rect 4620 49904 4672 49910
rect 4620 49846 4672 49852
rect 4526 49328 4582 49337
rect 4526 49263 4582 49272
rect 4724 49201 4752 54266
rect 4816 50289 4844 60030
rect 5264 59628 5316 59634
rect 5264 59570 5316 59576
rect 5276 59430 5304 59570
rect 5264 59424 5316 59430
rect 5264 59366 5316 59372
rect 5080 56364 5132 56370
rect 5080 56306 5132 56312
rect 5092 56166 5120 56306
rect 5080 56160 5132 56166
rect 5080 56102 5132 56108
rect 4896 55412 4948 55418
rect 4896 55354 4948 55360
rect 4908 54330 4936 55354
rect 4896 54324 4948 54330
rect 4896 54266 4948 54272
rect 5092 54210 5120 56102
rect 4908 54182 5120 54210
rect 4802 50280 4858 50289
rect 4802 50215 4858 50224
rect 4908 49434 4936 54182
rect 5276 54074 5304 59366
rect 5448 57792 5500 57798
rect 5448 57734 5500 57740
rect 5000 54046 5304 54074
rect 5000 49609 5028 54046
rect 5080 53984 5132 53990
rect 5080 53926 5132 53932
rect 4986 49600 5042 49609
rect 4986 49535 5042 49544
rect 4896 49428 4948 49434
rect 4896 49370 4948 49376
rect 4710 49192 4766 49201
rect 4710 49127 4766 49136
rect 5092 49065 5120 53926
rect 5172 52488 5224 52494
rect 5172 52430 5224 52436
rect 5184 49094 5212 52430
rect 5264 51264 5316 51270
rect 5264 51206 5316 51212
rect 5276 49162 5304 51206
rect 5356 50924 5408 50930
rect 5356 50866 5408 50872
rect 5264 49156 5316 49162
rect 5264 49098 5316 49104
rect 5172 49088 5224 49094
rect 5078 49056 5134 49065
rect 5172 49030 5224 49036
rect 3802 48988 4110 48997
rect 5078 48991 5134 49000
rect 3802 48986 3808 48988
rect 3864 48986 3888 48988
rect 3944 48986 3968 48988
rect 4024 48986 4048 48988
rect 4104 48986 4110 48988
rect 3864 48934 3866 48986
rect 4046 48934 4048 48986
rect 3802 48932 3808 48934
rect 3864 48932 3888 48934
rect 3944 48932 3968 48934
rect 4024 48932 4048 48934
rect 4104 48932 4110 48934
rect 3802 48923 4110 48932
rect 5368 48890 5396 50866
rect 5460 50561 5488 57734
rect 5644 57594 5672 91530
rect 10336 88890 10364 91530
rect 11612 91520 11664 91526
rect 11612 91462 11664 91468
rect 12532 91520 12584 91526
rect 12532 91462 12584 91468
rect 13544 91520 13596 91526
rect 13544 91462 13596 91468
rect 11624 91254 11652 91462
rect 12544 91322 12572 91462
rect 12532 91316 12584 91322
rect 12532 91258 12584 91264
rect 11612 91248 11664 91254
rect 11612 91190 11664 91196
rect 11624 88890 11652 91190
rect 12544 89714 12572 91258
rect 10258 88862 10364 88890
rect 11362 88862 11652 88890
rect 12452 89686 12572 89714
rect 12452 88876 12480 89686
rect 13556 88890 13584 91462
rect 13556 88876 13768 88890
rect 14660 88876 14688 95270
rect 15764 88876 15792 95270
rect 17052 88890 17080 95270
rect 18340 88890 18368 95270
rect 13570 88862 13768 88876
rect 16882 88862 17080 88890
rect 17986 88862 18368 88890
rect 19076 88876 19104 95406
rect 22652 95396 22704 95402
rect 22652 95338 22704 95344
rect 20168 95328 20220 95334
rect 20168 95270 20220 95276
rect 21548 95328 21600 95334
rect 21548 95270 21600 95276
rect 20180 88876 20208 95270
rect 21560 88890 21588 95270
rect 22664 88890 22692 95338
rect 23584 88890 23612 95406
rect 25872 95396 25924 95402
rect 25872 95338 25924 95344
rect 27160 95396 27212 95402
rect 27160 95338 27212 95344
rect 24768 95328 24820 95334
rect 24768 95270 24820 95276
rect 24780 88890 24808 95270
rect 25884 88890 25912 95338
rect 27172 88890 27200 95338
rect 27988 95328 28040 95334
rect 27988 95270 28040 95276
rect 29092 95328 29144 95334
rect 29092 95270 29144 95276
rect 28000 88890 28028 95270
rect 29104 88890 29132 95270
rect 21298 88862 21588 88890
rect 22402 88862 22692 88890
rect 23506 88862 23612 88890
rect 24610 88862 24808 88890
rect 25714 88862 25912 88890
rect 26818 88862 27200 88890
rect 27922 88862 28028 88890
rect 29026 88862 29132 88890
rect 30116 88876 30144 95474
rect 30472 92064 30524 92070
rect 30472 92006 30524 92012
rect 30484 91526 30512 92006
rect 30472 91520 30524 91526
rect 30472 91462 30524 91468
rect 31312 88890 31340 95474
rect 31234 88862 31340 88890
rect 32324 88876 32352 95474
rect 32404 92132 32456 92138
rect 32404 92074 32456 92080
rect 32416 91662 32444 92074
rect 32404 91656 32456 91662
rect 32404 91598 32456 91604
rect 33612 88890 33640 95474
rect 34900 88890 34928 95474
rect 35820 88890 35848 95474
rect 36832 88890 36860 95474
rect 36950 95228 37258 95237
rect 36950 95226 36956 95228
rect 37012 95226 37036 95228
rect 37092 95226 37116 95228
rect 37172 95226 37196 95228
rect 37252 95226 37258 95228
rect 37012 95174 37014 95226
rect 37194 95174 37196 95226
rect 36950 95172 36956 95174
rect 37012 95172 37036 95174
rect 37092 95172 37116 95174
rect 37172 95172 37196 95174
rect 37252 95172 37258 95174
rect 36950 95163 37258 95172
rect 37610 94684 37918 94693
rect 37610 94682 37616 94684
rect 37672 94682 37696 94684
rect 37752 94682 37776 94684
rect 37832 94682 37856 94684
rect 37912 94682 37918 94684
rect 37672 94630 37674 94682
rect 37854 94630 37856 94682
rect 37610 94628 37616 94630
rect 37672 94628 37696 94630
rect 37752 94628 37776 94630
rect 37832 94628 37856 94630
rect 37912 94628 37918 94630
rect 37610 94619 37918 94628
rect 36950 94140 37258 94149
rect 36950 94138 36956 94140
rect 37012 94138 37036 94140
rect 37092 94138 37116 94140
rect 37172 94138 37196 94140
rect 37252 94138 37258 94140
rect 37012 94086 37014 94138
rect 37194 94086 37196 94138
rect 36950 94084 36956 94086
rect 37012 94084 37036 94086
rect 37092 94084 37116 94086
rect 37172 94084 37196 94086
rect 37252 94084 37258 94086
rect 36950 94075 37258 94084
rect 37610 93596 37918 93605
rect 37610 93594 37616 93596
rect 37672 93594 37696 93596
rect 37752 93594 37776 93596
rect 37832 93594 37856 93596
rect 37912 93594 37918 93596
rect 37672 93542 37674 93594
rect 37854 93542 37856 93594
rect 37610 93540 37616 93542
rect 37672 93540 37696 93542
rect 37752 93540 37776 93542
rect 37832 93540 37856 93542
rect 37912 93540 37918 93542
rect 37610 93531 37918 93540
rect 36950 93052 37258 93061
rect 36950 93050 36956 93052
rect 37012 93050 37036 93052
rect 37092 93050 37116 93052
rect 37172 93050 37196 93052
rect 37252 93050 37258 93052
rect 37012 92998 37014 93050
rect 37194 92998 37196 93050
rect 36950 92996 36956 92998
rect 37012 92996 37036 92998
rect 37092 92996 37116 92998
rect 37172 92996 37196 92998
rect 37252 92996 37258 92998
rect 36950 92987 37258 92996
rect 37610 92508 37918 92517
rect 37610 92506 37616 92508
rect 37672 92506 37696 92508
rect 37752 92506 37776 92508
rect 37832 92506 37856 92508
rect 37912 92506 37918 92508
rect 37672 92454 37674 92506
rect 37854 92454 37856 92506
rect 37610 92452 37616 92454
rect 37672 92452 37696 92454
rect 37752 92452 37776 92454
rect 37832 92452 37856 92454
rect 37912 92452 37918 92454
rect 37610 92443 37918 92452
rect 36950 91964 37258 91973
rect 36950 91962 36956 91964
rect 37012 91962 37036 91964
rect 37092 91962 37116 91964
rect 37172 91962 37196 91964
rect 37252 91962 37258 91964
rect 37012 91910 37014 91962
rect 37194 91910 37196 91962
rect 36950 91908 36956 91910
rect 37012 91908 37036 91910
rect 37092 91908 37116 91910
rect 37172 91908 37196 91910
rect 37252 91908 37258 91910
rect 36950 91899 37258 91908
rect 37610 91420 37918 91429
rect 37610 91418 37616 91420
rect 37672 91418 37696 91420
rect 37752 91418 37776 91420
rect 37832 91418 37856 91420
rect 37912 91418 37918 91420
rect 37672 91366 37674 91418
rect 37854 91366 37856 91418
rect 37610 91364 37616 91366
rect 37672 91364 37696 91366
rect 37752 91364 37776 91366
rect 37832 91364 37856 91366
rect 37912 91364 37918 91366
rect 37610 91355 37918 91364
rect 38120 88890 38148 95474
rect 39040 88890 39068 95474
rect 33442 88862 33640 88890
rect 34546 88862 34928 88890
rect 35650 88862 35848 88890
rect 36754 88862 36860 88890
rect 37858 88862 38148 88890
rect 38962 88862 39068 88890
rect 40052 88876 40080 95474
rect 41340 88890 41368 95474
rect 42628 88890 42656 95474
rect 43456 91594 43484 97271
rect 44454 97200 44510 97294
rect 44744 95674 44772 97294
rect 49606 97322 49662 98000
rect 50894 97322 50950 98000
rect 49386 97294 49662 97322
rect 49330 97271 49386 97280
rect 49606 97200 49662 97294
rect 50816 97294 50950 97322
rect 50816 95674 50844 97294
rect 50894 97200 50950 97294
rect 52182 97322 52238 98000
rect 54758 97322 54814 98000
rect 56046 97322 56102 98000
rect 56690 97322 56746 98000
rect 57978 97322 58034 98000
rect 59266 97322 59322 98000
rect 52182 97294 52316 97322
rect 52182 97200 52238 97294
rect 44732 95668 44784 95674
rect 44732 95610 44784 95616
rect 50804 95668 50856 95674
rect 50804 95610 50856 95616
rect 52288 95538 52316 97294
rect 54758 97294 54984 97322
rect 54758 97200 54814 97294
rect 54956 95606 54984 97294
rect 56046 97294 56456 97322
rect 56046 97200 56102 97294
rect 56428 95674 56456 97294
rect 56690 97294 57008 97322
rect 56690 97200 56746 97294
rect 56980 95674 57008 97294
rect 57978 97294 58112 97322
rect 57978 97200 58034 97294
rect 58084 95674 58112 97294
rect 59188 97294 59322 97322
rect 59188 95674 59216 97294
rect 59266 97200 59322 97294
rect 59910 97322 59966 98000
rect 61198 97322 61254 98000
rect 62486 97322 62542 98000
rect 63774 97322 63830 98000
rect 59910 97294 60044 97322
rect 59910 97200 59966 97294
rect 56416 95668 56468 95674
rect 56416 95610 56468 95616
rect 56968 95668 57020 95674
rect 56968 95610 57020 95616
rect 58072 95668 58124 95674
rect 58072 95610 58124 95616
rect 59176 95668 59228 95674
rect 59176 95610 59228 95616
rect 54944 95600 54996 95606
rect 54944 95542 54996 95548
rect 60016 95538 60044 97294
rect 61120 97294 61254 97322
rect 61120 95674 61148 97294
rect 61198 97200 61254 97294
rect 62408 97294 62542 97322
rect 62408 95674 62436 97294
rect 62486 97200 62542 97294
rect 63696 97294 63830 97322
rect 63696 95674 63724 97294
rect 63774 97200 63830 97294
rect 64418 97322 64474 98000
rect 65706 97322 65762 98000
rect 66994 97322 67050 98000
rect 64418 97294 64644 97322
rect 64418 97200 64474 97294
rect 64616 95674 64644 97294
rect 65628 97294 65762 97322
rect 65628 95674 65656 97294
rect 65706 97200 65762 97294
rect 66916 97294 67050 97322
rect 66916 95674 66944 97294
rect 66994 97200 67050 97294
rect 67638 97322 67694 98000
rect 68926 97322 68982 98000
rect 67638 97294 67772 97322
rect 67638 97200 67694 97294
rect 67744 95674 67772 97294
rect 68848 97294 68982 97322
rect 68848 95674 68876 97294
rect 68926 97200 68982 97294
rect 70214 97322 70270 98000
rect 71502 97322 71558 98000
rect 72146 97322 72202 98000
rect 73434 97322 73490 98000
rect 74722 97322 74778 98000
rect 75366 97322 75422 98000
rect 76654 97322 76710 98000
rect 77942 97322 77998 98000
rect 79230 97322 79286 98000
rect 79874 97322 79930 98000
rect 81162 97322 81218 98000
rect 82450 97322 82506 98000
rect 70214 97294 70348 97322
rect 70214 97200 70270 97294
rect 70320 95674 70348 97294
rect 71502 97294 71728 97322
rect 71502 97200 71558 97294
rect 71700 95674 71728 97294
rect 72146 97294 72464 97322
rect 72146 97200 72202 97294
rect 72436 95674 72464 97294
rect 73434 97294 73568 97322
rect 73434 97200 73490 97294
rect 73540 95674 73568 97294
rect 74722 97294 75040 97322
rect 74722 97200 74778 97294
rect 73610 95772 73918 95781
rect 73610 95770 73616 95772
rect 73672 95770 73696 95772
rect 73752 95770 73776 95772
rect 73832 95770 73856 95772
rect 73912 95770 73918 95772
rect 73672 95718 73674 95770
rect 73854 95718 73856 95770
rect 73610 95716 73616 95718
rect 73672 95716 73696 95718
rect 73752 95716 73776 95718
rect 73832 95716 73856 95718
rect 73912 95716 73918 95718
rect 73610 95707 73918 95716
rect 75012 95674 75040 97294
rect 75366 97294 75592 97322
rect 75366 97200 75422 97294
rect 75564 95674 75592 97294
rect 76654 97294 76972 97322
rect 76654 97200 76710 97294
rect 76944 95674 76972 97294
rect 77942 97294 78260 97322
rect 77942 97200 77998 97294
rect 78232 95674 78260 97294
rect 79230 97294 79548 97322
rect 79230 97200 79286 97294
rect 79520 95674 79548 97294
rect 79874 97294 80008 97322
rect 79874 97200 79930 97294
rect 79980 95674 80008 97294
rect 81162 97294 81388 97322
rect 81162 97200 81218 97294
rect 81360 95674 81388 97294
rect 82450 97294 82768 97322
rect 82450 97200 82506 97294
rect 82740 95674 82768 97294
rect 61108 95668 61160 95674
rect 61108 95610 61160 95616
rect 62396 95668 62448 95674
rect 62396 95610 62448 95616
rect 63684 95668 63736 95674
rect 63684 95610 63736 95616
rect 64604 95668 64656 95674
rect 64604 95610 64656 95616
rect 65616 95668 65668 95674
rect 65616 95610 65668 95616
rect 66904 95668 66956 95674
rect 66904 95610 66956 95616
rect 67732 95668 67784 95674
rect 67732 95610 67784 95616
rect 68836 95668 68888 95674
rect 68836 95610 68888 95616
rect 70308 95668 70360 95674
rect 70308 95610 70360 95616
rect 71688 95668 71740 95674
rect 71688 95610 71740 95616
rect 72424 95668 72476 95674
rect 72424 95610 72476 95616
rect 73528 95668 73580 95674
rect 73528 95610 73580 95616
rect 75000 95668 75052 95674
rect 75000 95610 75052 95616
rect 75552 95668 75604 95674
rect 75552 95610 75604 95616
rect 76932 95668 76984 95674
rect 76932 95610 76984 95616
rect 78220 95668 78272 95674
rect 78220 95610 78272 95616
rect 79508 95668 79560 95674
rect 79508 95610 79560 95616
rect 79968 95668 80020 95674
rect 79968 95610 80020 95616
rect 81348 95668 81400 95674
rect 81348 95610 81400 95616
rect 82728 95668 82780 95674
rect 82728 95610 82780 95616
rect 43536 95532 43588 95538
rect 43536 95474 43588 95480
rect 44548 95532 44600 95538
rect 44548 95474 44600 95480
rect 52276 95532 52328 95538
rect 52276 95474 52328 95480
rect 60004 95532 60056 95538
rect 60004 95474 60056 95480
rect 70308 95532 70360 95538
rect 70308 95474 70360 95480
rect 71228 95532 71280 95538
rect 71228 95474 71280 95480
rect 72240 95532 72292 95538
rect 72240 95474 72292 95480
rect 73528 95532 73580 95538
rect 73528 95474 73580 95480
rect 74816 95532 74868 95538
rect 74816 95474 74868 95480
rect 75736 95532 75788 95538
rect 75736 95474 75788 95480
rect 76748 95532 76800 95538
rect 76748 95474 76800 95480
rect 78036 95532 78088 95538
rect 78036 95474 78088 95480
rect 78956 95532 79008 95538
rect 78956 95474 79008 95480
rect 80060 95532 80112 95538
rect 80060 95474 80112 95480
rect 81256 95532 81308 95538
rect 81256 95474 81308 95480
rect 82544 95532 82596 95538
rect 82544 95474 82596 95480
rect 43444 91588 43496 91594
rect 43444 91530 43496 91536
rect 43548 88890 43576 95474
rect 44560 88890 44588 95474
rect 52288 95130 52316 95474
rect 52368 95464 52420 95470
rect 52368 95406 52420 95412
rect 53748 95464 53800 95470
rect 53748 95406 53800 95412
rect 59084 95464 59136 95470
rect 59084 95406 59136 95412
rect 63500 95464 63552 95470
rect 63500 95406 63552 95412
rect 52276 95124 52328 95130
rect 52276 95066 52328 95072
rect 47492 92268 47544 92274
rect 47492 92210 47544 92216
rect 47400 92200 47452 92206
rect 46846 92168 46902 92177
rect 47400 92142 47452 92148
rect 46846 92103 46902 92112
rect 46754 91624 46810 91633
rect 46754 91559 46810 91568
rect 41170 88862 41368 88890
rect 42274 88862 42656 88890
rect 43378 88862 43576 88890
rect 44482 88862 44588 88890
rect 6736 88528 6788 88534
rect 6736 88470 6788 88476
rect 5908 71596 5960 71602
rect 5908 71538 5960 71544
rect 5816 70508 5868 70514
rect 5816 70450 5868 70456
rect 5724 67924 5776 67930
rect 5724 67866 5776 67872
rect 5736 67561 5764 67866
rect 5722 67552 5778 67561
rect 5722 67487 5778 67496
rect 5828 67402 5856 70450
rect 5736 67374 5856 67402
rect 5632 57588 5684 57594
rect 5632 57530 5684 57536
rect 5540 57248 5592 57254
rect 5540 57190 5592 57196
rect 5552 56710 5580 57190
rect 5644 56846 5672 57530
rect 5632 56840 5684 56846
rect 5632 56782 5684 56788
rect 5540 56704 5592 56710
rect 5540 56646 5592 56652
rect 5446 50552 5502 50561
rect 5446 50487 5502 50496
rect 1584 48884 1636 48890
rect 1584 48826 1636 48832
rect 5356 48884 5408 48890
rect 5356 48826 5408 48832
rect 1308 48748 1360 48754
rect 1308 48690 1360 48696
rect 1320 48385 1348 48690
rect 5172 48612 5224 48618
rect 5172 48554 5224 48560
rect 3066 48444 3374 48453
rect 3066 48442 3072 48444
rect 3128 48442 3152 48444
rect 3208 48442 3232 48444
rect 3288 48442 3312 48444
rect 3368 48442 3374 48444
rect 3128 48390 3130 48442
rect 3310 48390 3312 48442
rect 3066 48388 3072 48390
rect 3128 48388 3152 48390
rect 3208 48388 3232 48390
rect 3288 48388 3312 48390
rect 3368 48388 3374 48390
rect 1306 48376 1362 48385
rect 3066 48379 3374 48388
rect 1306 48311 1362 48320
rect 4710 48376 4766 48385
rect 4710 48311 4766 48320
rect 1400 48136 1452 48142
rect 1400 48078 1452 48084
rect 1412 47977 1440 48078
rect 1398 47968 1454 47977
rect 1398 47903 1454 47912
rect 3802 47900 4110 47909
rect 3802 47898 3808 47900
rect 3864 47898 3888 47900
rect 3944 47898 3968 47900
rect 4024 47898 4048 47900
rect 4104 47898 4110 47900
rect 3864 47846 3866 47898
rect 4046 47846 4048 47898
rect 3802 47844 3808 47846
rect 3864 47844 3888 47846
rect 3944 47844 3968 47846
rect 4024 47844 4048 47846
rect 4104 47844 4110 47846
rect 3802 47835 4110 47844
rect 4618 47832 4674 47841
rect 4618 47767 4674 47776
rect 3066 47356 3374 47365
rect 3066 47354 3072 47356
rect 3128 47354 3152 47356
rect 3208 47354 3232 47356
rect 3288 47354 3312 47356
rect 3368 47354 3374 47356
rect 3128 47302 3130 47354
rect 3310 47302 3312 47354
rect 3066 47300 3072 47302
rect 3128 47300 3152 47302
rect 3208 47300 3232 47302
rect 3288 47300 3312 47302
rect 3368 47300 3374 47302
rect 3066 47291 3374 47300
rect 1400 47048 1452 47054
rect 1398 47016 1400 47025
rect 1452 47016 1454 47025
rect 1398 46951 1454 46960
rect 3802 46812 4110 46821
rect 3802 46810 3808 46812
rect 3864 46810 3888 46812
rect 3944 46810 3968 46812
rect 4024 46810 4048 46812
rect 4104 46810 4110 46812
rect 3864 46758 3866 46810
rect 4046 46758 4048 46810
rect 3802 46756 3808 46758
rect 3864 46756 3888 46758
rect 3944 46756 3968 46758
rect 4024 46756 4048 46758
rect 4104 46756 4110 46758
rect 3802 46747 4110 46756
rect 1400 46368 1452 46374
rect 1398 46336 1400 46345
rect 1452 46336 1454 46345
rect 1398 46271 1454 46280
rect 3066 46268 3374 46277
rect 3066 46266 3072 46268
rect 3128 46266 3152 46268
rect 3208 46266 3232 46268
rect 3288 46266 3312 46268
rect 3368 46266 3374 46268
rect 3128 46214 3130 46266
rect 3310 46214 3312 46266
rect 3066 46212 3072 46214
rect 3128 46212 3152 46214
rect 3208 46212 3232 46214
rect 3288 46212 3312 46214
rect 3368 46212 3374 46214
rect 3066 46203 3374 46212
rect 1492 45824 1544 45830
rect 1490 45792 1492 45801
rect 1544 45792 1546 45801
rect 1490 45727 1546 45736
rect 3802 45724 4110 45733
rect 3802 45722 3808 45724
rect 3864 45722 3888 45724
rect 3944 45722 3968 45724
rect 4024 45722 4048 45724
rect 4104 45722 4110 45724
rect 3864 45670 3866 45722
rect 4046 45670 4048 45722
rect 3802 45668 3808 45670
rect 3864 45668 3888 45670
rect 3944 45668 3968 45670
rect 4024 45668 4048 45670
rect 4104 45668 4110 45670
rect 3802 45659 4110 45668
rect 1400 45280 1452 45286
rect 1400 45222 1452 45228
rect 1412 45121 1440 45222
rect 3066 45180 3374 45189
rect 3066 45178 3072 45180
rect 3128 45178 3152 45180
rect 3208 45178 3232 45180
rect 3288 45178 3312 45180
rect 3368 45178 3374 45180
rect 3128 45126 3130 45178
rect 3310 45126 3312 45178
rect 3066 45124 3072 45126
rect 3128 45124 3152 45126
rect 3208 45124 3232 45126
rect 3288 45124 3312 45126
rect 3368 45124 3374 45126
rect 1398 45112 1454 45121
rect 3066 45115 3374 45124
rect 1398 45047 1454 45056
rect 3802 44636 4110 44645
rect 3802 44634 3808 44636
rect 3864 44634 3888 44636
rect 3944 44634 3968 44636
rect 4024 44634 4048 44636
rect 4104 44634 4110 44636
rect 3864 44582 3866 44634
rect 4046 44582 4048 44634
rect 3802 44580 3808 44582
rect 3864 44580 3888 44582
rect 3944 44580 3968 44582
rect 4024 44580 4048 44582
rect 4104 44580 4110 44582
rect 3802 44571 4110 44580
rect 1490 44296 1546 44305
rect 1490 44231 1492 44240
rect 1544 44231 1546 44240
rect 1492 44202 1544 44208
rect 3066 44092 3374 44101
rect 3066 44090 3072 44092
rect 3128 44090 3152 44092
rect 3208 44090 3232 44092
rect 3288 44090 3312 44092
rect 3368 44090 3374 44092
rect 3128 44038 3130 44090
rect 3310 44038 3312 44090
rect 3066 44036 3072 44038
rect 3128 44036 3152 44038
rect 3208 44036 3232 44038
rect 3288 44036 3312 44038
rect 3368 44036 3374 44038
rect 3066 44027 3374 44036
rect 1216 43716 1268 43722
rect 1216 43658 1268 43664
rect 1228 43625 1256 43658
rect 1214 43616 1270 43625
rect 1214 43551 1270 43560
rect 3802 43548 4110 43557
rect 3802 43546 3808 43548
rect 3864 43546 3888 43548
rect 3944 43546 3968 43548
rect 4024 43546 4048 43548
rect 4104 43546 4110 43548
rect 3864 43494 3866 43546
rect 4046 43494 4048 43546
rect 3802 43492 3808 43494
rect 3864 43492 3888 43494
rect 3944 43492 3968 43494
rect 4024 43492 4048 43494
rect 4104 43492 4110 43494
rect 3802 43483 4110 43492
rect 1492 43104 1544 43110
rect 1490 43072 1492 43081
rect 1544 43072 1546 43081
rect 1490 43007 1546 43016
rect 3066 43004 3374 43013
rect 3066 43002 3072 43004
rect 3128 43002 3152 43004
rect 3208 43002 3232 43004
rect 3288 43002 3312 43004
rect 3368 43002 3374 43004
rect 3128 42950 3130 43002
rect 3310 42950 3312 43002
rect 3066 42948 3072 42950
rect 3128 42948 3152 42950
rect 3208 42948 3232 42950
rect 3288 42948 3312 42950
rect 3368 42948 3374 42950
rect 3066 42939 3374 42948
rect 3802 42460 4110 42469
rect 3802 42458 3808 42460
rect 3864 42458 3888 42460
rect 3944 42458 3968 42460
rect 4024 42458 4048 42460
rect 4104 42458 4110 42460
rect 3864 42406 3866 42458
rect 4046 42406 4048 42458
rect 3802 42404 3808 42406
rect 3864 42404 3888 42406
rect 3944 42404 3968 42406
rect 4024 42404 4048 42406
rect 4104 42404 4110 42406
rect 3802 42395 4110 42404
rect 3066 41916 3374 41925
rect 3066 41914 3072 41916
rect 3128 41914 3152 41916
rect 3208 41914 3232 41916
rect 3288 41914 3312 41916
rect 3368 41914 3374 41916
rect 3128 41862 3130 41914
rect 3310 41862 3312 41914
rect 3066 41860 3072 41862
rect 3128 41860 3152 41862
rect 3208 41860 3232 41862
rect 3288 41860 3312 41862
rect 3368 41860 3374 41862
rect 3066 41851 3374 41860
rect 1490 41576 1546 41585
rect 1490 41511 1546 41520
rect 1504 41478 1532 41511
rect 1492 41472 1544 41478
rect 1492 41414 1544 41420
rect 3802 41372 4110 41381
rect 3802 41370 3808 41372
rect 3864 41370 3888 41372
rect 3944 41370 3968 41372
rect 4024 41370 4048 41372
rect 4104 41370 4110 41372
rect 3864 41318 3866 41370
rect 4046 41318 4048 41370
rect 3802 41316 3808 41318
rect 3864 41316 3888 41318
rect 3944 41316 3968 41318
rect 4024 41316 4048 41318
rect 4104 41316 4110 41318
rect 3802 41307 4110 41316
rect 3066 40828 3374 40837
rect 3066 40826 3072 40828
rect 3128 40826 3152 40828
rect 3208 40826 3232 40828
rect 3288 40826 3312 40828
rect 3368 40826 3374 40828
rect 3128 40774 3130 40826
rect 3310 40774 3312 40826
rect 3066 40772 3072 40774
rect 3128 40772 3152 40774
rect 3208 40772 3232 40774
rect 3288 40772 3312 40774
rect 3368 40772 3374 40774
rect 3066 40763 3374 40772
rect 848 40384 900 40390
rect 846 40352 848 40361
rect 900 40352 902 40361
rect 846 40287 902 40296
rect 3802 40284 4110 40293
rect 3802 40282 3808 40284
rect 3864 40282 3888 40284
rect 3944 40282 3968 40284
rect 4024 40282 4048 40284
rect 4104 40282 4110 40284
rect 3864 40230 3866 40282
rect 4046 40230 4048 40282
rect 3802 40228 3808 40230
rect 3864 40228 3888 40230
rect 3944 40228 3968 40230
rect 4024 40228 4048 40230
rect 4104 40228 4110 40230
rect 3802 40219 4110 40228
rect 3066 39740 3374 39749
rect 3066 39738 3072 39740
rect 3128 39738 3152 39740
rect 3208 39738 3232 39740
rect 3288 39738 3312 39740
rect 3368 39738 3374 39740
rect 3128 39686 3130 39738
rect 3310 39686 3312 39738
rect 3066 39684 3072 39686
rect 3128 39684 3152 39686
rect 3208 39684 3232 39686
rect 3288 39684 3312 39686
rect 3368 39684 3374 39686
rect 3066 39675 3374 39684
rect 3802 39196 4110 39205
rect 3802 39194 3808 39196
rect 3864 39194 3888 39196
rect 3944 39194 3968 39196
rect 4024 39194 4048 39196
rect 4104 39194 4110 39196
rect 3864 39142 3866 39194
rect 4046 39142 4048 39194
rect 3802 39140 3808 39142
rect 3864 39140 3888 39142
rect 3944 39140 3968 39142
rect 4024 39140 4048 39142
rect 4104 39140 4110 39142
rect 3802 39131 4110 39140
rect 848 38752 900 38758
rect 846 38720 848 38729
rect 900 38720 902 38729
rect 846 38655 902 38664
rect 3066 38652 3374 38661
rect 3066 38650 3072 38652
rect 3128 38650 3152 38652
rect 3208 38650 3232 38652
rect 3288 38650 3312 38652
rect 3368 38650 3374 38652
rect 3128 38598 3130 38650
rect 3310 38598 3312 38650
rect 3066 38596 3072 38598
rect 3128 38596 3152 38598
rect 3208 38596 3232 38598
rect 3288 38596 3312 38598
rect 3368 38596 3374 38598
rect 3066 38587 3374 38596
rect 3802 38108 4110 38117
rect 3802 38106 3808 38108
rect 3864 38106 3888 38108
rect 3944 38106 3968 38108
rect 4024 38106 4048 38108
rect 4104 38106 4110 38108
rect 3864 38054 3866 38106
rect 4046 38054 4048 38106
rect 3802 38052 3808 38054
rect 3864 38052 3888 38054
rect 3944 38052 3968 38054
rect 4024 38052 4048 38054
rect 4104 38052 4110 38054
rect 3802 38043 4110 38052
rect 848 37664 900 37670
rect 846 37632 848 37641
rect 900 37632 902 37641
rect 846 37567 902 37576
rect 3066 37564 3374 37573
rect 3066 37562 3072 37564
rect 3128 37562 3152 37564
rect 3208 37562 3232 37564
rect 3288 37562 3312 37564
rect 3368 37562 3374 37564
rect 3128 37510 3130 37562
rect 3310 37510 3312 37562
rect 3066 37508 3072 37510
rect 3128 37508 3152 37510
rect 3208 37508 3232 37510
rect 3288 37508 3312 37510
rect 3368 37508 3374 37510
rect 3066 37499 3374 37508
rect 3802 37020 4110 37029
rect 3802 37018 3808 37020
rect 3864 37018 3888 37020
rect 3944 37018 3968 37020
rect 4024 37018 4048 37020
rect 4104 37018 4110 37020
rect 3864 36966 3866 37018
rect 4046 36966 4048 37018
rect 3802 36964 3808 36966
rect 3864 36964 3888 36966
rect 3944 36964 3968 36966
rect 4024 36964 4048 36966
rect 4104 36964 4110 36966
rect 3802 36955 4110 36964
rect 3066 36476 3374 36485
rect 3066 36474 3072 36476
rect 3128 36474 3152 36476
rect 3208 36474 3232 36476
rect 3288 36474 3312 36476
rect 3368 36474 3374 36476
rect 3128 36422 3130 36474
rect 3310 36422 3312 36474
rect 3066 36420 3072 36422
rect 3128 36420 3152 36422
rect 3208 36420 3232 36422
rect 3288 36420 3312 36422
rect 3368 36420 3374 36422
rect 3066 36411 3374 36420
rect 4632 36378 4660 47767
rect 4620 36372 4672 36378
rect 4620 36314 4672 36320
rect 848 36304 900 36310
rect 846 36272 848 36281
rect 900 36272 902 36281
rect 846 36207 902 36216
rect 3802 35932 4110 35941
rect 3802 35930 3808 35932
rect 3864 35930 3888 35932
rect 3944 35930 3968 35932
rect 4024 35930 4048 35932
rect 4104 35930 4110 35932
rect 3864 35878 3866 35930
rect 4046 35878 4048 35930
rect 3802 35876 3808 35878
rect 3864 35876 3888 35878
rect 3944 35876 3968 35878
rect 4024 35876 4048 35878
rect 4104 35876 4110 35878
rect 3802 35867 4110 35876
rect 3066 35388 3374 35397
rect 3066 35386 3072 35388
rect 3128 35386 3152 35388
rect 3208 35386 3232 35388
rect 3288 35386 3312 35388
rect 3368 35386 3374 35388
rect 3128 35334 3130 35386
rect 3310 35334 3312 35386
rect 3066 35332 3072 35334
rect 3128 35332 3152 35334
rect 3208 35332 3232 35334
rect 3288 35332 3312 35334
rect 3368 35332 3374 35334
rect 3066 35323 3374 35332
rect 848 34944 900 34950
rect 846 34912 848 34921
rect 900 34912 902 34921
rect 846 34847 902 34856
rect 3802 34844 4110 34853
rect 3802 34842 3808 34844
rect 3864 34842 3888 34844
rect 3944 34842 3968 34844
rect 4024 34842 4048 34844
rect 4104 34842 4110 34844
rect 3864 34790 3866 34842
rect 4046 34790 4048 34842
rect 3802 34788 3808 34790
rect 3864 34788 3888 34790
rect 3944 34788 3968 34790
rect 4024 34788 4048 34790
rect 4104 34788 4110 34790
rect 3802 34779 4110 34788
rect 3066 34300 3374 34309
rect 3066 34298 3072 34300
rect 3128 34298 3152 34300
rect 3208 34298 3232 34300
rect 3288 34298 3312 34300
rect 3368 34298 3374 34300
rect 3128 34246 3130 34298
rect 3310 34246 3312 34298
rect 3066 34244 3072 34246
rect 3128 34244 3152 34246
rect 3208 34244 3232 34246
rect 3288 34244 3312 34246
rect 3368 34244 3374 34246
rect 3066 34235 3374 34244
rect 3802 33756 4110 33765
rect 3802 33754 3808 33756
rect 3864 33754 3888 33756
rect 3944 33754 3968 33756
rect 4024 33754 4048 33756
rect 4104 33754 4110 33756
rect 3864 33702 3866 33754
rect 4046 33702 4048 33754
rect 3802 33700 3808 33702
rect 3864 33700 3888 33702
rect 3944 33700 3968 33702
rect 4024 33700 4048 33702
rect 4104 33700 4110 33702
rect 3802 33691 4110 33700
rect 848 33312 900 33318
rect 846 33280 848 33289
rect 900 33280 902 33289
rect 846 33215 902 33224
rect 3066 33212 3374 33221
rect 3066 33210 3072 33212
rect 3128 33210 3152 33212
rect 3208 33210 3232 33212
rect 3288 33210 3312 33212
rect 3368 33210 3374 33212
rect 3128 33158 3130 33210
rect 3310 33158 3312 33210
rect 3066 33156 3072 33158
rect 3128 33156 3152 33158
rect 3208 33156 3232 33158
rect 3288 33156 3312 33158
rect 3368 33156 3374 33158
rect 3066 33147 3374 33156
rect 3802 32668 4110 32677
rect 3802 32666 3808 32668
rect 3864 32666 3888 32668
rect 3944 32666 3968 32668
rect 4024 32666 4048 32668
rect 4104 32666 4110 32668
rect 3864 32614 3866 32666
rect 4046 32614 4048 32666
rect 3802 32612 3808 32614
rect 3864 32612 3888 32614
rect 3944 32612 3968 32614
rect 4024 32612 4048 32614
rect 4104 32612 4110 32614
rect 3802 32603 4110 32612
rect 848 32224 900 32230
rect 846 32192 848 32201
rect 900 32192 902 32201
rect 846 32127 902 32136
rect 3066 32124 3374 32133
rect 3066 32122 3072 32124
rect 3128 32122 3152 32124
rect 3208 32122 3232 32124
rect 3288 32122 3312 32124
rect 3368 32122 3374 32124
rect 3128 32070 3130 32122
rect 3310 32070 3312 32122
rect 3066 32068 3072 32070
rect 3128 32068 3152 32070
rect 3208 32068 3232 32070
rect 3288 32068 3312 32070
rect 3368 32068 3374 32070
rect 3066 32059 3374 32068
rect 3802 31580 4110 31589
rect 3802 31578 3808 31580
rect 3864 31578 3888 31580
rect 3944 31578 3968 31580
rect 4024 31578 4048 31580
rect 4104 31578 4110 31580
rect 3864 31526 3866 31578
rect 4046 31526 4048 31578
rect 3802 31524 3808 31526
rect 3864 31524 3888 31526
rect 3944 31524 3968 31526
rect 4024 31524 4048 31526
rect 4104 31524 4110 31526
rect 3802 31515 4110 31524
rect 3066 31036 3374 31045
rect 3066 31034 3072 31036
rect 3128 31034 3152 31036
rect 3208 31034 3232 31036
rect 3288 31034 3312 31036
rect 3368 31034 3374 31036
rect 3128 30982 3130 31034
rect 3310 30982 3312 31034
rect 3066 30980 3072 30982
rect 3128 30980 3152 30982
rect 3208 30980 3232 30982
rect 3288 30980 3312 30982
rect 3368 30980 3374 30982
rect 3066 30971 3374 30980
rect 4724 30938 4752 48311
rect 4986 48104 5042 48113
rect 4986 48039 5042 48048
rect 4894 47968 4950 47977
rect 4894 47903 4950 47912
rect 4804 46504 4856 46510
rect 4804 46446 4856 46452
rect 4816 32570 4844 46446
rect 4908 40730 4936 47903
rect 4896 40724 4948 40730
rect 4896 40666 4948 40672
rect 4908 40458 4936 40666
rect 4896 40452 4948 40458
rect 4896 40394 4948 40400
rect 5000 39098 5028 48039
rect 5080 47660 5132 47666
rect 5080 47602 5132 47608
rect 5092 41818 5120 47602
rect 5080 41812 5132 41818
rect 5080 41754 5132 41760
rect 5092 41546 5120 41754
rect 5080 41540 5132 41546
rect 5080 41482 5132 41488
rect 5184 41414 5212 48554
rect 5448 47456 5500 47462
rect 5448 47398 5500 47404
rect 5354 47152 5410 47161
rect 5354 47087 5410 47096
rect 5262 46472 5318 46481
rect 5262 46407 5318 46416
rect 5092 41386 5212 41414
rect 4988 39092 5040 39098
rect 4988 39034 5040 39040
rect 4988 34944 5040 34950
rect 4988 34886 5040 34892
rect 4804 32564 4856 32570
rect 4804 32506 4856 32512
rect 4816 32434 4844 32506
rect 4804 32428 4856 32434
rect 4804 32370 4856 32376
rect 4712 30932 4764 30938
rect 4712 30874 4764 30880
rect 848 30864 900 30870
rect 846 30832 848 30841
rect 900 30832 902 30841
rect 846 30767 902 30776
rect 3802 30492 4110 30501
rect 3802 30490 3808 30492
rect 3864 30490 3888 30492
rect 3944 30490 3968 30492
rect 4024 30490 4048 30492
rect 4104 30490 4110 30492
rect 3864 30438 3866 30490
rect 4046 30438 4048 30490
rect 3802 30436 3808 30438
rect 3864 30436 3888 30438
rect 3944 30436 3968 30438
rect 4024 30436 4048 30438
rect 4104 30436 4110 30438
rect 3802 30427 4110 30436
rect 3066 29948 3374 29957
rect 3066 29946 3072 29948
rect 3128 29946 3152 29948
rect 3208 29946 3232 29948
rect 3288 29946 3312 29948
rect 3368 29946 3374 29948
rect 3128 29894 3130 29946
rect 3310 29894 3312 29946
rect 3066 29892 3072 29894
rect 3128 29892 3152 29894
rect 3208 29892 3232 29894
rect 3288 29892 3312 29894
rect 3368 29892 3374 29894
rect 3066 29883 3374 29892
rect 848 29504 900 29510
rect 846 29472 848 29481
rect 900 29472 902 29481
rect 846 29407 902 29416
rect 3802 29404 4110 29413
rect 3802 29402 3808 29404
rect 3864 29402 3888 29404
rect 3944 29402 3968 29404
rect 4024 29402 4048 29404
rect 4104 29402 4110 29404
rect 3864 29350 3866 29402
rect 4046 29350 4048 29402
rect 3802 29348 3808 29350
rect 3864 29348 3888 29350
rect 3944 29348 3968 29350
rect 4024 29348 4048 29350
rect 4104 29348 4110 29350
rect 3802 29339 4110 29348
rect 3066 28860 3374 28869
rect 3066 28858 3072 28860
rect 3128 28858 3152 28860
rect 3208 28858 3232 28860
rect 3288 28858 3312 28860
rect 3368 28858 3374 28860
rect 3128 28806 3130 28858
rect 3310 28806 3312 28858
rect 3066 28804 3072 28806
rect 3128 28804 3152 28806
rect 3208 28804 3232 28806
rect 3288 28804 3312 28806
rect 3368 28804 3374 28806
rect 3066 28795 3374 28804
rect 3802 28316 4110 28325
rect 3802 28314 3808 28316
rect 3864 28314 3888 28316
rect 3944 28314 3968 28316
rect 4024 28314 4048 28316
rect 4104 28314 4110 28316
rect 3864 28262 3866 28314
rect 4046 28262 4048 28314
rect 3802 28260 3808 28262
rect 3864 28260 3888 28262
rect 3944 28260 3968 28262
rect 4024 28260 4048 28262
rect 4104 28260 4110 28262
rect 3802 28251 4110 28260
rect 848 27872 900 27878
rect 846 27840 848 27849
rect 900 27840 902 27849
rect 846 27775 902 27784
rect 3066 27772 3374 27781
rect 3066 27770 3072 27772
rect 3128 27770 3152 27772
rect 3208 27770 3232 27772
rect 3288 27770 3312 27772
rect 3368 27770 3374 27772
rect 3128 27718 3130 27770
rect 3310 27718 3312 27770
rect 3066 27716 3072 27718
rect 3128 27716 3152 27718
rect 3208 27716 3232 27718
rect 3288 27716 3312 27718
rect 3368 27716 3374 27718
rect 3066 27707 3374 27716
rect 3802 27228 4110 27237
rect 3802 27226 3808 27228
rect 3864 27226 3888 27228
rect 3944 27226 3968 27228
rect 4024 27226 4048 27228
rect 4104 27226 4110 27228
rect 3864 27174 3866 27226
rect 4046 27174 4048 27226
rect 3802 27172 3808 27174
rect 3864 27172 3888 27174
rect 3944 27172 3968 27174
rect 4024 27172 4048 27174
rect 4104 27172 4110 27174
rect 3802 27163 4110 27172
rect 1308 26988 1360 26994
rect 1308 26930 1360 26936
rect 1320 26625 1348 26930
rect 3066 26684 3374 26693
rect 3066 26682 3072 26684
rect 3128 26682 3152 26684
rect 3208 26682 3232 26684
rect 3288 26682 3312 26684
rect 3368 26682 3374 26684
rect 3128 26630 3130 26682
rect 3310 26630 3312 26682
rect 3066 26628 3072 26630
rect 3128 26628 3152 26630
rect 3208 26628 3232 26630
rect 3288 26628 3312 26630
rect 3368 26628 3374 26630
rect 1306 26616 1362 26625
rect 3066 26619 3374 26628
rect 1306 26551 1362 26560
rect 3802 26140 4110 26149
rect 3802 26138 3808 26140
rect 3864 26138 3888 26140
rect 3944 26138 3968 26140
rect 4024 26138 4048 26140
rect 4104 26138 4110 26140
rect 3864 26086 3866 26138
rect 4046 26086 4048 26138
rect 3802 26084 3808 26086
rect 3864 26084 3888 26086
rect 3944 26084 3968 26086
rect 4024 26084 4048 26086
rect 4104 26084 4110 26086
rect 3802 26075 4110 26084
rect 3066 25596 3374 25605
rect 3066 25594 3072 25596
rect 3128 25594 3152 25596
rect 3208 25594 3232 25596
rect 3288 25594 3312 25596
rect 3368 25594 3374 25596
rect 3128 25542 3130 25594
rect 3310 25542 3312 25594
rect 3066 25540 3072 25542
rect 3128 25540 3152 25542
rect 3208 25540 3232 25542
rect 3288 25540 3312 25542
rect 3368 25540 3374 25542
rect 3066 25531 3374 25540
rect 1216 25288 1268 25294
rect 1214 25256 1216 25265
rect 1268 25256 1270 25265
rect 1214 25191 1270 25200
rect 3802 25052 4110 25061
rect 3802 25050 3808 25052
rect 3864 25050 3888 25052
rect 3944 25050 3968 25052
rect 4024 25050 4048 25052
rect 4104 25050 4110 25052
rect 3864 24998 3866 25050
rect 4046 24998 4048 25050
rect 3802 24996 3808 24998
rect 3864 24996 3888 24998
rect 3944 24996 3968 24998
rect 4024 24996 4048 24998
rect 4104 24996 4110 24998
rect 3802 24987 4110 24996
rect 3066 24508 3374 24517
rect 3066 24506 3072 24508
rect 3128 24506 3152 24508
rect 3208 24506 3232 24508
rect 3288 24506 3312 24508
rect 3368 24506 3374 24508
rect 3128 24454 3130 24506
rect 3310 24454 3312 24506
rect 3066 24452 3072 24454
rect 3128 24452 3152 24454
rect 3208 24452 3232 24454
rect 3288 24452 3312 24454
rect 3368 24452 3374 24454
rect 3066 24443 3374 24452
rect 1308 24200 1360 24206
rect 1308 24142 1360 24148
rect 1320 23905 1348 24142
rect 3802 23964 4110 23973
rect 3802 23962 3808 23964
rect 3864 23962 3888 23964
rect 3944 23962 3968 23964
rect 4024 23962 4048 23964
rect 4104 23962 4110 23964
rect 3864 23910 3866 23962
rect 4046 23910 4048 23962
rect 3802 23908 3808 23910
rect 3864 23908 3888 23910
rect 3944 23908 3968 23910
rect 4024 23908 4048 23910
rect 4104 23908 4110 23910
rect 1306 23896 1362 23905
rect 3802 23899 4110 23908
rect 1306 23831 1362 23840
rect 3066 23420 3374 23429
rect 3066 23418 3072 23420
rect 3128 23418 3152 23420
rect 3208 23418 3232 23420
rect 3288 23418 3312 23420
rect 3368 23418 3374 23420
rect 3128 23366 3130 23418
rect 3310 23366 3312 23418
rect 3066 23364 3072 23366
rect 3128 23364 3152 23366
rect 3208 23364 3232 23366
rect 3288 23364 3312 23366
rect 3368 23364 3374 23366
rect 3066 23355 3374 23364
rect 3802 22876 4110 22885
rect 3802 22874 3808 22876
rect 3864 22874 3888 22876
rect 3944 22874 3968 22876
rect 4024 22874 4048 22876
rect 4104 22874 4110 22876
rect 3864 22822 3866 22874
rect 4046 22822 4048 22874
rect 3802 22820 3808 22822
rect 3864 22820 3888 22822
rect 3944 22820 3968 22822
rect 4024 22820 4048 22822
rect 4104 22820 4110 22822
rect 3802 22811 4110 22820
rect 1308 22636 1360 22642
rect 1308 22578 1360 22584
rect 1320 22545 1348 22578
rect 1306 22536 1362 22545
rect 1306 22471 1362 22480
rect 3066 22332 3374 22341
rect 3066 22330 3072 22332
rect 3128 22330 3152 22332
rect 3208 22330 3232 22332
rect 3288 22330 3312 22332
rect 3368 22330 3374 22332
rect 3128 22278 3130 22330
rect 3310 22278 3312 22330
rect 3066 22276 3072 22278
rect 3128 22276 3152 22278
rect 3208 22276 3232 22278
rect 3288 22276 3312 22278
rect 3368 22276 3374 22278
rect 3066 22267 3374 22276
rect 3802 21788 4110 21797
rect 3802 21786 3808 21788
rect 3864 21786 3888 21788
rect 3944 21786 3968 21788
rect 4024 21786 4048 21788
rect 4104 21786 4110 21788
rect 3864 21734 3866 21786
rect 4046 21734 4048 21786
rect 3802 21732 3808 21734
rect 3864 21732 3888 21734
rect 3944 21732 3968 21734
rect 4024 21732 4048 21734
rect 4104 21732 4110 21734
rect 3802 21723 4110 21732
rect 1308 21548 1360 21554
rect 1308 21490 1360 21496
rect 1320 21185 1348 21490
rect 3066 21244 3374 21253
rect 3066 21242 3072 21244
rect 3128 21242 3152 21244
rect 3208 21242 3232 21244
rect 3288 21242 3312 21244
rect 3368 21242 3374 21244
rect 3128 21190 3130 21242
rect 3310 21190 3312 21242
rect 3066 21188 3072 21190
rect 3128 21188 3152 21190
rect 3208 21188 3232 21190
rect 3288 21188 3312 21190
rect 3368 21188 3374 21190
rect 1306 21176 1362 21185
rect 3066 21179 3374 21188
rect 1306 21111 1362 21120
rect 3802 20700 4110 20709
rect 3802 20698 3808 20700
rect 3864 20698 3888 20700
rect 3944 20698 3968 20700
rect 4024 20698 4048 20700
rect 4104 20698 4110 20700
rect 3864 20646 3866 20698
rect 4046 20646 4048 20698
rect 3802 20644 3808 20646
rect 3864 20644 3888 20646
rect 3944 20644 3968 20646
rect 4024 20644 4048 20646
rect 4104 20644 4110 20646
rect 3802 20635 4110 20644
rect 3066 20156 3374 20165
rect 3066 20154 3072 20156
rect 3128 20154 3152 20156
rect 3208 20154 3232 20156
rect 3288 20154 3312 20156
rect 3368 20154 3374 20156
rect 3128 20102 3130 20154
rect 3310 20102 3312 20154
rect 3066 20100 3072 20102
rect 3128 20100 3152 20102
rect 3208 20100 3232 20102
rect 3288 20100 3312 20102
rect 3368 20100 3374 20102
rect 3066 20091 3374 20100
rect 1216 19848 1268 19854
rect 1214 19816 1216 19825
rect 1268 19816 1270 19825
rect 1214 19751 1270 19760
rect 3802 19612 4110 19621
rect 3802 19610 3808 19612
rect 3864 19610 3888 19612
rect 3944 19610 3968 19612
rect 4024 19610 4048 19612
rect 4104 19610 4110 19612
rect 3864 19558 3866 19610
rect 4046 19558 4048 19610
rect 3802 19556 3808 19558
rect 3864 19556 3888 19558
rect 3944 19556 3968 19558
rect 4024 19556 4048 19558
rect 4104 19556 4110 19558
rect 3802 19547 4110 19556
rect 3066 19068 3374 19077
rect 3066 19066 3072 19068
rect 3128 19066 3152 19068
rect 3208 19066 3232 19068
rect 3288 19066 3312 19068
rect 3368 19066 3374 19068
rect 3128 19014 3130 19066
rect 3310 19014 3312 19066
rect 3066 19012 3072 19014
rect 3128 19012 3152 19014
rect 3208 19012 3232 19014
rect 3288 19012 3312 19014
rect 3368 19012 3374 19014
rect 3066 19003 3374 19012
rect 1308 18760 1360 18766
rect 1308 18702 1360 18708
rect 1320 18465 1348 18702
rect 3802 18524 4110 18533
rect 3802 18522 3808 18524
rect 3864 18522 3888 18524
rect 3944 18522 3968 18524
rect 4024 18522 4048 18524
rect 4104 18522 4110 18524
rect 3864 18470 3866 18522
rect 4046 18470 4048 18522
rect 3802 18468 3808 18470
rect 3864 18468 3888 18470
rect 3944 18468 3968 18470
rect 4024 18468 4048 18470
rect 4104 18468 4110 18470
rect 1306 18456 1362 18465
rect 3802 18459 4110 18468
rect 1306 18391 1362 18400
rect 3066 17980 3374 17989
rect 3066 17978 3072 17980
rect 3128 17978 3152 17980
rect 3208 17978 3232 17980
rect 3288 17978 3312 17980
rect 3368 17978 3374 17980
rect 3128 17926 3130 17978
rect 3310 17926 3312 17978
rect 3066 17924 3072 17926
rect 3128 17924 3152 17926
rect 3208 17924 3232 17926
rect 3288 17924 3312 17926
rect 3368 17924 3374 17926
rect 3066 17915 3374 17924
rect 3802 17436 4110 17445
rect 3802 17434 3808 17436
rect 3864 17434 3888 17436
rect 3944 17434 3968 17436
rect 4024 17434 4048 17436
rect 4104 17434 4110 17436
rect 3864 17382 3866 17434
rect 4046 17382 4048 17434
rect 3802 17380 3808 17382
rect 3864 17380 3888 17382
rect 3944 17380 3968 17382
rect 4024 17380 4048 17382
rect 4104 17380 4110 17382
rect 3802 17371 4110 17380
rect 1308 17196 1360 17202
rect 1308 17138 1360 17144
rect 1320 17105 1348 17138
rect 1306 17096 1362 17105
rect 1306 17031 1362 17040
rect 3066 16892 3374 16901
rect 3066 16890 3072 16892
rect 3128 16890 3152 16892
rect 3208 16890 3232 16892
rect 3288 16890 3312 16892
rect 3368 16890 3374 16892
rect 3128 16838 3130 16890
rect 3310 16838 3312 16890
rect 3066 16836 3072 16838
rect 3128 16836 3152 16838
rect 3208 16836 3232 16838
rect 3288 16836 3312 16838
rect 3368 16836 3374 16838
rect 3066 16827 3374 16836
rect 3802 16348 4110 16357
rect 3802 16346 3808 16348
rect 3864 16346 3888 16348
rect 3944 16346 3968 16348
rect 4024 16346 4048 16348
rect 4104 16346 4110 16348
rect 3864 16294 3866 16346
rect 4046 16294 4048 16346
rect 3802 16292 3808 16294
rect 3864 16292 3888 16294
rect 3944 16292 3968 16294
rect 4024 16292 4048 16294
rect 4104 16292 4110 16294
rect 3802 16283 4110 16292
rect 1308 16108 1360 16114
rect 1308 16050 1360 16056
rect 1320 15745 1348 16050
rect 3066 15804 3374 15813
rect 3066 15802 3072 15804
rect 3128 15802 3152 15804
rect 3208 15802 3232 15804
rect 3288 15802 3312 15804
rect 3368 15802 3374 15804
rect 3128 15750 3130 15802
rect 3310 15750 3312 15802
rect 3066 15748 3072 15750
rect 3128 15748 3152 15750
rect 3208 15748 3232 15750
rect 3288 15748 3312 15750
rect 3368 15748 3374 15750
rect 1306 15736 1362 15745
rect 3066 15739 3374 15748
rect 1306 15671 1362 15680
rect 3802 15260 4110 15269
rect 3802 15258 3808 15260
rect 3864 15258 3888 15260
rect 3944 15258 3968 15260
rect 4024 15258 4048 15260
rect 4104 15258 4110 15260
rect 3864 15206 3866 15258
rect 4046 15206 4048 15258
rect 3802 15204 3808 15206
rect 3864 15204 3888 15206
rect 3944 15204 3968 15206
rect 4024 15204 4048 15206
rect 4104 15204 4110 15206
rect 3802 15195 4110 15204
rect 3066 14716 3374 14725
rect 3066 14714 3072 14716
rect 3128 14714 3152 14716
rect 3208 14714 3232 14716
rect 3288 14714 3312 14716
rect 3368 14714 3374 14716
rect 3128 14662 3130 14714
rect 3310 14662 3312 14714
rect 3066 14660 3072 14662
rect 3128 14660 3152 14662
rect 3208 14660 3232 14662
rect 3288 14660 3312 14662
rect 3368 14660 3374 14662
rect 3066 14651 3374 14660
rect 1216 14408 1268 14414
rect 1214 14376 1216 14385
rect 1268 14376 1270 14385
rect 1214 14311 1270 14320
rect 3802 14172 4110 14181
rect 3802 14170 3808 14172
rect 3864 14170 3888 14172
rect 3944 14170 3968 14172
rect 4024 14170 4048 14172
rect 4104 14170 4110 14172
rect 3864 14118 3866 14170
rect 4046 14118 4048 14170
rect 3802 14116 3808 14118
rect 3864 14116 3888 14118
rect 3944 14116 3968 14118
rect 4024 14116 4048 14118
rect 4104 14116 4110 14118
rect 3802 14107 4110 14116
rect 3066 13628 3374 13637
rect 3066 13626 3072 13628
rect 3128 13626 3152 13628
rect 3208 13626 3232 13628
rect 3288 13626 3312 13628
rect 3368 13626 3374 13628
rect 3128 13574 3130 13626
rect 3310 13574 3312 13626
rect 3066 13572 3072 13574
rect 3128 13572 3152 13574
rect 3208 13572 3232 13574
rect 3288 13572 3312 13574
rect 3368 13572 3374 13574
rect 3066 13563 3374 13572
rect 1308 13320 1360 13326
rect 1308 13262 1360 13268
rect 1320 13025 1348 13262
rect 3802 13084 4110 13093
rect 3802 13082 3808 13084
rect 3864 13082 3888 13084
rect 3944 13082 3968 13084
rect 4024 13082 4048 13084
rect 4104 13082 4110 13084
rect 3864 13030 3866 13082
rect 4046 13030 4048 13082
rect 3802 13028 3808 13030
rect 3864 13028 3888 13030
rect 3944 13028 3968 13030
rect 4024 13028 4048 13030
rect 4104 13028 4110 13030
rect 1306 13016 1362 13025
rect 3802 13019 4110 13028
rect 1306 12951 1362 12960
rect 3066 12540 3374 12549
rect 3066 12538 3072 12540
rect 3128 12538 3152 12540
rect 3208 12538 3232 12540
rect 3288 12538 3312 12540
rect 3368 12538 3374 12540
rect 3128 12486 3130 12538
rect 3310 12486 3312 12538
rect 3066 12484 3072 12486
rect 3128 12484 3152 12486
rect 3208 12484 3232 12486
rect 3288 12484 3312 12486
rect 3368 12484 3374 12486
rect 3066 12475 3374 12484
rect 3802 11996 4110 12005
rect 3802 11994 3808 11996
rect 3864 11994 3888 11996
rect 3944 11994 3968 11996
rect 4024 11994 4048 11996
rect 4104 11994 4110 11996
rect 3864 11942 3866 11994
rect 4046 11942 4048 11994
rect 3802 11940 3808 11942
rect 3864 11940 3888 11942
rect 3944 11940 3968 11942
rect 4024 11940 4048 11942
rect 4104 11940 4110 11942
rect 3802 11931 4110 11940
rect 1308 11756 1360 11762
rect 1308 11698 1360 11704
rect 1320 11665 1348 11698
rect 1306 11656 1362 11665
rect 1306 11591 1362 11600
rect 3066 11452 3374 11461
rect 3066 11450 3072 11452
rect 3128 11450 3152 11452
rect 3208 11450 3232 11452
rect 3288 11450 3312 11452
rect 3368 11450 3374 11452
rect 3128 11398 3130 11450
rect 3310 11398 3312 11450
rect 3066 11396 3072 11398
rect 3128 11396 3152 11398
rect 3208 11396 3232 11398
rect 3288 11396 3312 11398
rect 3368 11396 3374 11398
rect 3066 11387 3374 11396
rect 3802 10908 4110 10917
rect 3802 10906 3808 10908
rect 3864 10906 3888 10908
rect 3944 10906 3968 10908
rect 4024 10906 4048 10908
rect 4104 10906 4110 10908
rect 3864 10854 3866 10906
rect 4046 10854 4048 10906
rect 3802 10852 3808 10854
rect 3864 10852 3888 10854
rect 3944 10852 3968 10854
rect 4024 10852 4048 10854
rect 4104 10852 4110 10854
rect 3802 10843 4110 10852
rect 3066 10364 3374 10373
rect 3066 10362 3072 10364
rect 3128 10362 3152 10364
rect 3208 10362 3232 10364
rect 3288 10362 3312 10364
rect 3368 10362 3374 10364
rect 3128 10310 3130 10362
rect 3310 10310 3312 10362
rect 3066 10308 3072 10310
rect 3128 10308 3152 10310
rect 3208 10308 3232 10310
rect 3288 10308 3312 10310
rect 3368 10308 3374 10310
rect 3066 10299 3374 10308
rect 3802 9820 4110 9829
rect 3802 9818 3808 9820
rect 3864 9818 3888 9820
rect 3944 9818 3968 9820
rect 4024 9818 4048 9820
rect 4104 9818 4110 9820
rect 3864 9766 3866 9818
rect 4046 9766 4048 9818
rect 3802 9764 3808 9766
rect 3864 9764 3888 9766
rect 3944 9764 3968 9766
rect 4024 9764 4048 9766
rect 4104 9764 4110 9766
rect 3802 9755 4110 9764
rect 3066 9276 3374 9285
rect 3066 9274 3072 9276
rect 3128 9274 3152 9276
rect 3208 9274 3232 9276
rect 3288 9274 3312 9276
rect 3368 9274 3374 9276
rect 3128 9222 3130 9274
rect 3310 9222 3312 9274
rect 3066 9220 3072 9222
rect 3128 9220 3152 9222
rect 3208 9220 3232 9222
rect 3288 9220 3312 9222
rect 3368 9220 3374 9222
rect 3066 9211 3374 9220
rect 3802 8732 4110 8741
rect 3802 8730 3808 8732
rect 3864 8730 3888 8732
rect 3944 8730 3968 8732
rect 4024 8730 4048 8732
rect 4104 8730 4110 8732
rect 3864 8678 3866 8730
rect 4046 8678 4048 8730
rect 3802 8676 3808 8678
rect 3864 8676 3888 8678
rect 3944 8676 3968 8678
rect 4024 8676 4048 8678
rect 4104 8676 4110 8678
rect 3802 8667 4110 8676
rect 3066 8188 3374 8197
rect 3066 8186 3072 8188
rect 3128 8186 3152 8188
rect 3208 8186 3232 8188
rect 3288 8186 3312 8188
rect 3368 8186 3374 8188
rect 3128 8134 3130 8186
rect 3310 8134 3312 8186
rect 3066 8132 3072 8134
rect 3128 8132 3152 8134
rect 3208 8132 3232 8134
rect 3288 8132 3312 8134
rect 3368 8132 3374 8134
rect 3066 8123 3374 8132
rect 5000 7886 5028 34886
rect 5092 28218 5120 41386
rect 5276 28218 5304 46407
rect 5368 40730 5396 47087
rect 5460 44402 5488 47398
rect 5552 47258 5580 56646
rect 5632 50856 5684 50862
rect 5632 50798 5684 50804
rect 5644 50522 5672 50798
rect 5632 50516 5684 50522
rect 5632 50458 5684 50464
rect 5736 48278 5764 67374
rect 5920 67266 5948 71538
rect 6184 68740 6236 68746
rect 6184 68682 6236 68688
rect 6092 68672 6144 68678
rect 6092 68614 6144 68620
rect 5828 67238 5948 67266
rect 5828 49706 5856 67238
rect 5908 65000 5960 65006
rect 5908 64942 5960 64948
rect 5920 64841 5948 64942
rect 5906 64832 5962 64841
rect 5906 64767 5962 64776
rect 5906 62248 5962 62257
rect 5906 62183 5962 62192
rect 5920 62150 5948 62183
rect 5908 62144 5960 62150
rect 5908 62086 5960 62092
rect 5908 59424 5960 59430
rect 5908 59366 5960 59372
rect 5816 49700 5868 49706
rect 5816 49642 5868 49648
rect 5920 48822 5948 59366
rect 6104 49774 6132 68614
rect 6196 51074 6224 68682
rect 6748 64874 6776 88470
rect 13740 88466 13768 88862
rect 13728 88460 13780 88466
rect 13728 88402 13780 88408
rect 8300 86828 8352 86834
rect 8300 86770 8352 86776
rect 8312 86737 8340 86770
rect 8298 86728 8354 86737
rect 8298 86663 8354 86672
rect 8298 85368 8354 85377
rect 8298 85303 8354 85312
rect 8312 85134 8340 85303
rect 8300 85128 8352 85134
rect 8300 85070 8352 85076
rect 8300 84040 8352 84046
rect 8298 84008 8300 84017
rect 8352 84008 8354 84017
rect 8298 83943 8354 83952
rect 8298 82648 8354 82657
rect 8298 82583 8354 82592
rect 8312 82482 8340 82583
rect 8300 82476 8352 82482
rect 8300 82418 8352 82424
rect 8300 81388 8352 81394
rect 8300 81330 8352 81336
rect 8312 81297 8340 81330
rect 8298 81288 8354 81297
rect 8298 81223 8354 81232
rect 8298 79928 8354 79937
rect 8298 79863 8354 79872
rect 8312 79694 8340 79863
rect 8300 79688 8352 79694
rect 8300 79630 8352 79636
rect 8300 78600 8352 78606
rect 8298 78568 8300 78577
rect 8352 78568 8354 78577
rect 8298 78503 8354 78512
rect 8298 77208 8354 77217
rect 8298 77143 8354 77152
rect 8312 77042 8340 77143
rect 8300 77036 8352 77042
rect 8300 76978 8352 76984
rect 8298 74488 8354 74497
rect 8298 74423 8354 74432
rect 8312 74254 8340 74423
rect 8300 74248 8352 74254
rect 8300 74190 8352 74196
rect 8300 73160 8352 73166
rect 8298 73128 8300 73137
rect 8352 73128 8354 73137
rect 8298 73063 8354 73072
rect 8298 71768 8354 71777
rect 8298 71703 8354 71712
rect 8312 71670 8340 71703
rect 8300 71664 8352 71670
rect 8300 71606 8352 71612
rect 8300 68944 8352 68950
rect 8300 68886 8352 68892
rect 8312 68649 8340 68886
rect 8298 68640 8354 68649
rect 8298 68575 8354 68584
rect 8300 66020 8352 66026
rect 8300 65962 8352 65968
rect 7564 65952 7616 65958
rect 8312 65929 8340 65962
rect 7564 65894 7616 65900
rect 8298 65920 8354 65929
rect 6656 64846 6776 64874
rect 6196 51046 6316 51074
rect 6092 49768 6144 49774
rect 6092 49710 6144 49716
rect 5908 48816 5960 48822
rect 5908 48758 5960 48764
rect 6184 48680 6236 48686
rect 6184 48622 6236 48628
rect 5724 48272 5776 48278
rect 5724 48214 5776 48220
rect 5632 47728 5684 47734
rect 5632 47670 5684 47676
rect 5540 47252 5592 47258
rect 5540 47194 5592 47200
rect 5448 44396 5500 44402
rect 5448 44338 5500 44344
rect 5356 40724 5408 40730
rect 5356 40666 5408 40672
rect 5644 33522 5672 47670
rect 6092 47320 6144 47326
rect 6092 47262 6144 47268
rect 6104 44282 6132 47262
rect 5736 44254 6132 44282
rect 5736 37874 5764 44254
rect 6196 41414 6224 48622
rect 6288 48210 6316 51046
rect 6552 50992 6604 50998
rect 6552 50934 6604 50940
rect 6460 49836 6512 49842
rect 6460 49778 6512 49784
rect 6276 48204 6328 48210
rect 6276 48146 6328 48152
rect 6366 47696 6422 47705
rect 6366 47631 6422 47640
rect 6276 47116 6328 47122
rect 6276 47058 6328 47064
rect 5828 41386 6224 41414
rect 5724 37868 5776 37874
rect 5724 37810 5776 37816
rect 5632 33516 5684 33522
rect 5632 33458 5684 33464
rect 5632 30728 5684 30734
rect 5632 30670 5684 30676
rect 5448 29640 5500 29646
rect 5448 29582 5500 29588
rect 5356 29504 5408 29510
rect 5356 29446 5408 29452
rect 5080 28212 5132 28218
rect 5080 28154 5132 28160
rect 5264 28212 5316 28218
rect 5264 28154 5316 28160
rect 5262 27160 5318 27169
rect 5262 27095 5318 27104
rect 5276 27062 5304 27095
rect 5264 27056 5316 27062
rect 5264 26998 5316 27004
rect 5368 8294 5396 29446
rect 5356 8288 5408 8294
rect 5356 8230 5408 8236
rect 5460 8022 5488 29582
rect 5540 26784 5592 26790
rect 5540 26726 5592 26732
rect 5448 8016 5500 8022
rect 5448 7958 5500 7964
rect 5552 7954 5580 26726
rect 5540 7948 5592 7954
rect 5540 7890 5592 7896
rect 4988 7880 5040 7886
rect 4988 7822 5040 7828
rect 5644 7818 5672 30670
rect 5828 25498 5856 41386
rect 6288 35086 6316 47058
rect 6380 38010 6408 47631
rect 6472 41750 6500 49778
rect 6564 48754 6592 50934
rect 6656 50794 6684 64846
rect 7196 57792 7248 57798
rect 7196 57734 7248 57740
rect 6736 56160 6788 56166
rect 6736 56102 6788 56108
rect 6748 50998 6776 56102
rect 6828 55412 6880 55418
rect 6828 55354 6880 55360
rect 6736 50992 6788 50998
rect 6736 50934 6788 50940
rect 6644 50788 6696 50794
rect 6644 50730 6696 50736
rect 6656 50658 6684 50730
rect 6736 50720 6788 50726
rect 6736 50662 6788 50668
rect 6644 50652 6696 50658
rect 6644 50594 6696 50600
rect 6644 50516 6696 50522
rect 6644 50458 6696 50464
rect 6552 48748 6604 48754
rect 6552 48690 6604 48696
rect 6552 47388 6604 47394
rect 6552 47330 6604 47336
rect 6564 44538 6592 47330
rect 6552 44532 6604 44538
rect 6552 44474 6604 44480
rect 6460 41744 6512 41750
rect 6460 41686 6512 41692
rect 6656 41414 6684 50458
rect 6748 48074 6776 50662
rect 6840 49638 6868 55354
rect 6828 49632 6880 49638
rect 6828 49574 6880 49580
rect 7208 49230 7236 57734
rect 7576 50998 7604 65894
rect 8298 65855 8354 65864
rect 8300 63504 8352 63510
rect 8300 63446 8352 63452
rect 7656 63232 7708 63238
rect 8312 63209 8340 63446
rect 7656 63174 7708 63180
rect 8298 63200 8354 63209
rect 7564 50992 7616 50998
rect 7564 50934 7616 50940
rect 7668 49366 7696 63174
rect 8298 63135 8354 63144
rect 8300 61668 8352 61674
rect 8300 61610 8352 61616
rect 8312 61305 8340 61610
rect 8298 61296 8354 61305
rect 8298 61231 8354 61240
rect 7840 60512 7892 60518
rect 7840 60454 7892 60460
rect 7656 49360 7708 49366
rect 7656 49302 7708 49308
rect 7852 49298 7880 60454
rect 8300 60036 8352 60042
rect 8300 59978 8352 59984
rect 8312 59945 8340 59978
rect 8298 59936 8354 59945
rect 8298 59871 8354 59880
rect 8300 59152 8352 59158
rect 8300 59094 8352 59100
rect 8312 58585 8340 59094
rect 8298 58576 8354 58585
rect 8298 58511 8354 58520
rect 8300 57316 8352 57322
rect 8300 57258 8352 57264
rect 8312 57225 8340 57258
rect 8298 57216 8354 57225
rect 8298 57151 8354 57160
rect 8300 56228 8352 56234
rect 8300 56170 8352 56176
rect 8312 55865 8340 56170
rect 8298 55856 8354 55865
rect 8298 55791 8354 55800
rect 8300 54596 8352 54602
rect 8300 54538 8352 54544
rect 8312 54505 8340 54538
rect 8298 54496 8354 54505
rect 8298 54431 8354 54440
rect 7932 53984 7984 53990
rect 7932 53926 7984 53932
rect 7944 50862 7972 53926
rect 8300 53712 8352 53718
rect 8300 53654 8352 53660
rect 8312 53145 8340 53654
rect 8298 53136 8354 53145
rect 8298 53071 8354 53080
rect 8208 52624 8260 52630
rect 8208 52566 8260 52572
rect 7932 50856 7984 50862
rect 7932 50798 7984 50804
rect 8220 50590 8248 52566
rect 9600 50658 9706 50674
rect 9588 50652 9706 50658
rect 9640 50646 9706 50652
rect 9588 50594 9640 50600
rect 8208 50584 8260 50590
rect 46768 50561 46796 91559
rect 46860 50658 46888 92103
rect 47308 89684 47360 89690
rect 47308 89626 47360 89632
rect 47320 88398 47348 89626
rect 47308 88392 47360 88398
rect 47306 88360 47308 88369
rect 47360 88360 47362 88369
rect 47306 88295 47362 88304
rect 46848 50652 46900 50658
rect 46848 50594 46900 50600
rect 46754 50552 46810 50561
rect 8208 50526 8260 50532
rect 11624 50522 12296 50538
rect 11612 50516 12296 50522
rect 11664 50510 12296 50516
rect 11612 50458 11664 50464
rect 8208 50312 8260 50318
rect 8208 50254 8260 50260
rect 8024 50176 8076 50182
rect 8024 50118 8076 50124
rect 8036 49978 8064 50118
rect 8024 49972 8076 49978
rect 8024 49914 8076 49920
rect 7840 49292 7892 49298
rect 7840 49234 7892 49240
rect 7196 49224 7248 49230
rect 7196 49166 7248 49172
rect 7012 48476 7064 48482
rect 7012 48418 7064 48424
rect 6736 48068 6788 48074
rect 6736 48010 6788 48016
rect 6920 47592 6972 47598
rect 6920 47534 6972 47540
rect 6828 46708 6880 46714
rect 6828 46650 6880 46656
rect 6840 43994 6868 46650
rect 6828 43988 6880 43994
rect 6828 43930 6880 43936
rect 6932 43314 6960 47534
rect 7024 43450 7052 48418
rect 7562 47288 7618 47297
rect 7562 47223 7618 47232
rect 7012 43444 7064 43450
rect 7012 43386 7064 43392
rect 6920 43308 6972 43314
rect 6920 43250 6972 43256
rect 6656 41386 6868 41414
rect 6368 38004 6420 38010
rect 6368 37946 6420 37952
rect 6276 35080 6328 35086
rect 6276 35022 6328 35028
rect 6184 33312 6236 33318
rect 6184 33254 6236 33260
rect 5816 25492 5868 25498
rect 5816 25434 5868 25440
rect 5632 7812 5684 7818
rect 5632 7754 5684 7760
rect 6196 7682 6224 33254
rect 6276 32224 6328 32230
rect 6276 32166 6328 32172
rect 6184 7676 6236 7682
rect 3802 7644 4110 7653
rect 3802 7642 3808 7644
rect 3864 7642 3888 7644
rect 3944 7642 3968 7644
rect 4024 7642 4048 7644
rect 4104 7642 4110 7644
rect 3864 7590 3866 7642
rect 4046 7590 4048 7642
rect 6184 7618 6236 7624
rect 6288 7614 6316 32166
rect 6368 25152 6420 25158
rect 6368 25094 6420 25100
rect 6380 7750 6408 25094
rect 6840 8158 6868 41386
rect 7576 36174 7604 47223
rect 7840 47184 7892 47190
rect 7840 47126 7892 47132
rect 7852 38962 7880 47126
rect 7840 38956 7892 38962
rect 7840 38898 7892 38904
rect 7564 36168 7616 36174
rect 7564 36110 7616 36116
rect 8036 8158 8064 49914
rect 8114 10024 8170 10033
rect 8114 9959 8170 9968
rect 6828 8152 6880 8158
rect 6828 8094 6880 8100
rect 8024 8152 8076 8158
rect 8024 8094 8076 8100
rect 6368 7744 6420 7750
rect 6368 7686 6420 7692
rect 3802 7588 3808 7590
rect 3864 7588 3888 7590
rect 3944 7588 3968 7590
rect 4024 7588 4048 7590
rect 4104 7588 4110 7590
rect 3802 7579 4110 7588
rect 6276 7608 6328 7614
rect 6276 7550 6328 7556
rect 3066 7100 3374 7109
rect 3066 7098 3072 7100
rect 3128 7098 3152 7100
rect 3208 7098 3232 7100
rect 3288 7098 3312 7100
rect 3368 7098 3374 7100
rect 3128 7046 3130 7098
rect 3310 7046 3312 7098
rect 3066 7044 3072 7046
rect 3128 7044 3152 7046
rect 3208 7044 3232 7046
rect 3288 7044 3312 7046
rect 3368 7044 3374 7046
rect 3066 7035 3374 7044
rect 3802 6556 4110 6565
rect 3802 6554 3808 6556
rect 3864 6554 3888 6556
rect 3944 6554 3968 6556
rect 4024 6554 4048 6556
rect 4104 6554 4110 6556
rect 3864 6502 3866 6554
rect 4046 6502 4048 6554
rect 3802 6500 3808 6502
rect 3864 6500 3888 6502
rect 3944 6500 3968 6502
rect 4024 6500 4048 6502
rect 4104 6500 4110 6502
rect 3802 6491 4110 6500
rect 3066 6012 3374 6021
rect 3066 6010 3072 6012
rect 3128 6010 3152 6012
rect 3208 6010 3232 6012
rect 3288 6010 3312 6012
rect 3368 6010 3374 6012
rect 3128 5958 3130 6010
rect 3310 5958 3312 6010
rect 3066 5956 3072 5958
rect 3128 5956 3152 5958
rect 3208 5956 3232 5958
rect 3288 5956 3312 5958
rect 3368 5956 3374 5958
rect 3066 5947 3374 5956
rect 3802 5468 4110 5477
rect 3802 5466 3808 5468
rect 3864 5466 3888 5468
rect 3944 5466 3968 5468
rect 4024 5466 4048 5468
rect 4104 5466 4110 5468
rect 3864 5414 3866 5466
rect 4046 5414 4048 5466
rect 3802 5412 3808 5414
rect 3864 5412 3888 5414
rect 3944 5412 3968 5414
rect 4024 5412 4048 5414
rect 4104 5412 4110 5414
rect 3802 5403 4110 5412
rect 8128 2582 8156 9959
rect 8220 8226 8248 50254
rect 12268 50250 12296 50510
rect 46754 50487 46810 50496
rect 46754 50416 46810 50425
rect 46754 50351 46810 50360
rect 13084 50312 13136 50318
rect 13018 50260 13084 50266
rect 13018 50254 13136 50260
rect 12256 50244 12308 50250
rect 13018 50238 13124 50254
rect 12256 50186 12308 50192
rect 10876 50176 10928 50182
rect 10520 50124 10876 50130
rect 10520 50118 10928 50124
rect 10520 50102 10916 50118
rect 10520 49978 10548 50102
rect 10508 49972 10560 49978
rect 10508 49914 10560 49920
rect 9680 49768 9732 49774
rect 8390 49736 8446 49745
rect 9680 49710 9732 49716
rect 8390 49671 8446 49680
rect 8404 46102 8432 49671
rect 9692 48142 9720 49710
rect 15212 48362 15240 50116
rect 15120 48334 15240 48362
rect 16040 50102 16330 50130
rect 17144 50102 17434 50130
rect 18248 50102 18538 50130
rect 19352 50102 19642 50130
rect 9680 48136 9732 48142
rect 9680 48078 9732 48084
rect 10508 47592 10560 47598
rect 10508 47534 10560 47540
rect 11244 47592 11296 47598
rect 11244 47534 11296 47540
rect 10520 47326 10548 47534
rect 11152 47456 11204 47462
rect 11152 47398 11204 47404
rect 10416 47320 10468 47326
rect 10416 47262 10468 47268
rect 10508 47320 10560 47326
rect 10508 47262 10560 47268
rect 10232 47252 10284 47258
rect 10232 47194 10284 47200
rect 9680 46980 9732 46986
rect 9680 46922 9732 46928
rect 9692 46442 9720 46922
rect 10244 46866 10272 47194
rect 10428 47190 10456 47262
rect 10416 47184 10468 47190
rect 10416 47126 10468 47132
rect 11164 47054 11192 47398
rect 11060 47048 11112 47054
rect 11060 46990 11112 46996
rect 11152 47048 11204 47054
rect 11256 47025 11284 47534
rect 11428 47524 11480 47530
rect 11428 47466 11480 47472
rect 11152 46990 11204 46996
rect 11242 47016 11298 47025
rect 11072 46866 11100 46990
rect 11440 46986 11468 47466
rect 11242 46951 11298 46960
rect 11428 46980 11480 46986
rect 11428 46922 11480 46928
rect 12532 46912 12584 46918
rect 10244 46852 10364 46866
rect 10258 46838 10364 46852
rect 11072 46838 11744 46866
rect 12466 46860 12532 46866
rect 15120 46866 15148 48334
rect 16040 46866 16068 50102
rect 17144 46866 17172 50102
rect 18248 46866 18276 50102
rect 19352 48314 19380 50102
rect 20732 48314 20760 50116
rect 19260 48286 19380 48314
rect 20640 48286 20760 48314
rect 21560 50102 21850 50130
rect 22664 50102 22954 50130
rect 23768 50102 24058 50130
rect 24872 50102 25162 50130
rect 19260 46866 19288 48286
rect 20640 46866 20668 48286
rect 21560 46866 21588 50102
rect 22664 46866 22692 50102
rect 23768 46866 23796 50102
rect 24872 48314 24900 50102
rect 26252 48314 26280 50116
rect 24780 48286 24900 48314
rect 26160 48286 26280 48314
rect 27080 50102 27370 50130
rect 28184 50102 28474 50130
rect 29288 50102 29578 50130
rect 30392 50102 30682 50130
rect 24780 46866 24808 48286
rect 26160 46866 26188 48286
rect 27080 46866 27108 50102
rect 28184 46866 28212 50102
rect 29288 46866 29316 50102
rect 30392 48314 30420 50102
rect 31772 48314 31800 50116
rect 30300 48286 30420 48314
rect 31680 48286 31800 48314
rect 32600 50102 32890 50130
rect 33704 50102 33994 50130
rect 34808 50102 35098 50130
rect 35912 50102 36202 50130
rect 30300 46866 30328 48286
rect 31680 46866 31708 48286
rect 32600 46866 32628 50102
rect 33704 46866 33732 50102
rect 34808 46866 34836 50102
rect 35912 48314 35940 50102
rect 37292 48314 37320 50116
rect 35820 48286 35940 48314
rect 37200 48286 37320 48314
rect 38120 50102 38410 50130
rect 39224 50102 39514 50130
rect 40328 50102 40618 50130
rect 41432 50102 41722 50130
rect 35820 46866 35848 48286
rect 37200 46866 37228 48286
rect 38120 46866 38148 50102
rect 39224 46866 39252 50102
rect 40328 46866 40356 50102
rect 40682 49328 40738 49337
rect 40682 49263 40738 49272
rect 40696 48929 40724 49263
rect 40682 48920 40738 48929
rect 40682 48855 40738 48864
rect 41432 48314 41460 50102
rect 42812 48314 42840 50116
rect 41340 48286 41460 48314
rect 42720 48286 42840 48314
rect 43640 50102 43930 50130
rect 44744 50102 45034 50130
rect 41340 46866 41368 48286
rect 42720 46866 42748 48286
rect 43640 46866 43668 50102
rect 44744 46866 44772 50102
rect 46768 48074 46796 50351
rect 46860 50289 46888 50594
rect 46846 50280 46902 50289
rect 47412 50250 47440 92142
rect 47504 50454 47532 92210
rect 52380 92138 52408 95406
rect 52460 92200 52512 92206
rect 52460 92142 52512 92148
rect 51080 92132 51132 92138
rect 51080 92074 51132 92080
rect 52368 92132 52420 92138
rect 52368 92074 52420 92080
rect 50252 92064 50304 92070
rect 50252 92006 50304 92012
rect 50264 91866 50292 92006
rect 50252 91860 50304 91866
rect 50252 91802 50304 91808
rect 47952 91724 48004 91730
rect 47952 91666 48004 91672
rect 47768 91588 47820 91594
rect 47768 91530 47820 91536
rect 47676 91520 47728 91526
rect 47676 91462 47728 91468
rect 47584 88460 47636 88466
rect 47584 88402 47636 88408
rect 47492 50448 47544 50454
rect 47492 50390 47544 50396
rect 46846 50215 46902 50224
rect 47400 50244 47452 50250
rect 47400 50186 47452 50192
rect 46848 49836 46900 49842
rect 46848 49778 46900 49784
rect 46860 48890 46888 49778
rect 47214 49736 47270 49745
rect 47214 49671 47270 49680
rect 46848 48884 46900 48890
rect 46848 48826 46900 48832
rect 46756 48068 46808 48074
rect 46756 48010 46808 48016
rect 46848 47592 46900 47598
rect 46846 47560 46848 47569
rect 46900 47560 46902 47569
rect 46846 47495 46902 47504
rect 46754 47424 46810 47433
rect 46754 47359 46810 47368
rect 12466 46854 12584 46860
rect 12466 46838 12572 46854
rect 14674 46838 15148 46866
rect 15778 46838 16068 46866
rect 16882 46838 17172 46866
rect 17986 46838 18276 46866
rect 19090 46838 19288 46866
rect 20194 46838 20668 46866
rect 21298 46838 21588 46866
rect 22402 46838 22692 46866
rect 23506 46838 23796 46866
rect 24610 46838 24808 46866
rect 25714 46838 26188 46866
rect 26818 46838 27108 46866
rect 27922 46838 28212 46866
rect 29026 46838 29316 46866
rect 30130 46838 30328 46866
rect 31234 46838 31708 46866
rect 32338 46838 32628 46866
rect 33442 46838 33732 46866
rect 34546 46838 34836 46866
rect 35650 46838 35848 46866
rect 36754 46838 37228 46866
rect 37858 46838 38148 46866
rect 38962 46838 39252 46866
rect 40066 46838 40356 46866
rect 41170 46838 41368 46866
rect 42274 46838 42748 46866
rect 43378 46838 43668 46866
rect 44482 46838 44772 46866
rect 10336 46510 10364 46838
rect 11716 46646 11744 46838
rect 11704 46640 11756 46646
rect 11704 46582 11756 46588
rect 10324 46504 10376 46510
rect 10324 46446 10376 46452
rect 12544 46442 12572 46838
rect 13280 46714 13570 46730
rect 13268 46708 13570 46714
rect 13320 46702 13570 46708
rect 13268 46650 13320 46656
rect 9680 46436 9732 46442
rect 9680 46378 9732 46384
rect 12532 46436 12584 46442
rect 12532 46378 12584 46384
rect 8392 46096 8444 46102
rect 8298 46064 8354 46073
rect 8392 46038 8444 46044
rect 8298 45999 8354 46008
rect 8312 45966 8340 45999
rect 8300 45960 8352 45966
rect 8300 45902 8352 45908
rect 8300 44328 8352 44334
rect 8298 44296 8300 44305
rect 8352 44296 8354 44305
rect 8298 44231 8354 44240
rect 8300 43376 8352 43382
rect 8298 43344 8300 43353
rect 8352 43344 8354 43353
rect 8298 43279 8354 43288
rect 8300 41608 8352 41614
rect 8298 41576 8300 41585
rect 8352 41576 8354 41585
rect 8298 41511 8354 41520
rect 8298 40624 8354 40633
rect 8298 40559 8354 40568
rect 8312 40526 8340 40559
rect 8300 40520 8352 40526
rect 8300 40462 8352 40468
rect 8300 38888 8352 38894
rect 8298 38856 8300 38865
rect 8352 38856 8354 38865
rect 8298 38791 8354 38800
rect 8300 37936 8352 37942
rect 8298 37904 8300 37913
rect 8352 37904 8354 37913
rect 8298 37839 8354 37848
rect 8298 36136 8354 36145
rect 8298 36071 8300 36080
rect 8352 36071 8354 36080
rect 8300 36042 8352 36048
rect 8298 35184 8354 35193
rect 8298 35119 8300 35128
rect 8352 35119 8354 35128
rect 8300 35090 8352 35096
rect 8300 33448 8352 33454
rect 8298 33416 8300 33425
rect 8352 33416 8354 33425
rect 8298 33351 8354 33360
rect 8300 32496 8352 32502
rect 8298 32464 8300 32473
rect 8352 32464 8354 32473
rect 8298 32399 8354 32408
rect 8298 30696 8354 30705
rect 8298 30631 8300 30640
rect 8352 30631 8354 30640
rect 8300 30602 8352 30608
rect 8298 29744 8354 29753
rect 8298 29679 8300 29688
rect 8352 29679 8354 29688
rect 8300 29650 8352 29656
rect 8300 28008 8352 28014
rect 8298 27976 8300 27985
rect 8352 27976 8354 27985
rect 8298 27911 8354 27920
rect 8300 27124 8352 27130
rect 8300 27066 8352 27072
rect 8312 27033 8340 27066
rect 8298 27024 8354 27033
rect 8298 26959 8354 26968
rect 8298 25664 8354 25673
rect 8298 25599 8354 25608
rect 8312 25430 8340 25599
rect 8300 25424 8352 25430
rect 8300 25366 8352 25372
rect 8300 24336 8352 24342
rect 8298 24304 8300 24313
rect 8352 24304 8354 24313
rect 8298 24239 8354 24248
rect 8298 22536 8354 22545
rect 8298 22471 8300 22480
rect 8352 22471 8354 22480
rect 8300 22442 8352 22448
rect 8300 21684 8352 21690
rect 8300 21626 8352 21632
rect 8312 21593 8340 21626
rect 8298 21584 8354 21593
rect 8298 21519 8354 21528
rect 8298 20224 8354 20233
rect 8298 20159 8354 20168
rect 8312 20058 8340 20159
rect 8300 20052 8352 20058
rect 8300 19994 8352 20000
rect 8300 18896 8352 18902
rect 8298 18864 8300 18873
rect 8352 18864 8354 18873
rect 8298 18799 8354 18808
rect 8298 17096 8354 17105
rect 8298 17031 8300 17040
rect 8352 17031 8354 17040
rect 8300 17002 8352 17008
rect 8300 16244 8352 16250
rect 8300 16186 8352 16192
rect 8312 16153 8340 16186
rect 8298 16144 8354 16153
rect 8298 16079 8354 16088
rect 8298 14784 8354 14793
rect 8298 14719 8354 14728
rect 8312 14618 8340 14719
rect 8300 14612 8352 14618
rect 8300 14554 8352 14560
rect 8300 13456 8352 13462
rect 8298 13424 8300 13433
rect 8352 13424 8354 13433
rect 8298 13359 8354 13368
rect 8298 11656 8354 11665
rect 8298 11591 8300 11600
rect 8352 11591 8354 11600
rect 8300 11562 8352 11568
rect 46768 9654 46796 47359
rect 46756 9648 46808 9654
rect 46756 9590 46808 9596
rect 8298 8664 8354 8673
rect 8298 8599 8354 8608
rect 8208 8220 8260 8226
rect 8208 8162 8260 8168
rect 8312 2650 8340 8599
rect 12728 8228 13018 8242
rect 12728 8226 13032 8228
rect 12716 8220 13032 8226
rect 12768 8214 13032 8220
rect 12716 8162 12768 8168
rect 10508 8152 10560 8158
rect 9706 8078 9812 8106
rect 10560 8100 10916 8106
rect 10508 8094 10916 8100
rect 10520 8078 10916 8094
rect 11624 8090 12020 8106
rect 9784 5710 9812 8078
rect 10888 6186 10916 8078
rect 11612 8084 12020 8090
rect 11664 8078 12020 8084
rect 11612 8026 11664 8032
rect 10876 6180 10928 6186
rect 10876 6122 10928 6128
rect 10888 5914 10916 6122
rect 10876 5908 10928 5914
rect 10876 5850 10928 5856
rect 9772 5704 9824 5710
rect 9772 5646 9824 5652
rect 10888 2650 10916 5850
rect 11992 5642 12020 8078
rect 13004 5914 13032 8214
rect 15226 8078 15608 8106
rect 16330 8078 16528 8106
rect 17434 8078 17540 8106
rect 18538 8078 18828 8106
rect 19642 8078 19748 8106
rect 12992 5908 13044 5914
rect 12992 5850 13044 5856
rect 15108 5908 15160 5914
rect 15108 5850 15160 5856
rect 11980 5636 12032 5642
rect 11980 5578 12032 5584
rect 13360 5636 13412 5642
rect 13360 5578 13412 5584
rect 13372 2650 13400 5578
rect 15120 2650 15148 5850
rect 8300 2644 8352 2650
rect 8300 2586 8352 2592
rect 10876 2644 10928 2650
rect 10876 2586 10928 2592
rect 13360 2644 13412 2650
rect 13360 2586 13412 2592
rect 15108 2644 15160 2650
rect 15108 2586 15160 2592
rect 8116 2576 8168 2582
rect 8116 2518 8168 2524
rect 15580 2446 15608 8078
rect 16500 2446 16528 8078
rect 17512 2446 17540 8078
rect 18800 2446 18828 8078
rect 19720 2446 19748 8078
rect 20732 2446 20760 8092
rect 21850 8078 22048 8106
rect 22954 8078 23336 8106
rect 24058 8078 24256 8106
rect 25162 8078 25268 8106
rect 26266 8078 26556 8106
rect 27370 8078 27476 8106
rect 22020 2446 22048 8078
rect 23308 2446 23336 8078
rect 24228 2446 24256 8078
rect 25240 2446 25268 8078
rect 26528 2446 26556 8078
rect 27448 2446 27476 8078
rect 28460 2446 28488 8092
rect 29578 8078 29776 8106
rect 30682 8078 31064 8106
rect 31786 8078 31892 8106
rect 32890 8078 32996 8106
rect 33994 8078 34284 8106
rect 29748 2446 29776 8078
rect 31036 2650 31064 8078
rect 31864 2650 31892 8078
rect 32968 2650 32996 8078
rect 34256 2650 34284 8078
rect 35084 2650 35112 8092
rect 36188 2650 36216 8092
rect 37306 8078 37504 8106
rect 36950 4924 37258 4933
rect 36950 4922 36956 4924
rect 37012 4922 37036 4924
rect 37092 4922 37116 4924
rect 37172 4922 37196 4924
rect 37252 4922 37258 4924
rect 37012 4870 37014 4922
rect 37194 4870 37196 4922
rect 36950 4868 36956 4870
rect 37012 4868 37036 4870
rect 37092 4868 37116 4870
rect 37172 4868 37196 4870
rect 37252 4868 37258 4870
rect 36950 4859 37258 4868
rect 36950 3836 37258 3845
rect 36950 3834 36956 3836
rect 37012 3834 37036 3836
rect 37092 3834 37116 3836
rect 37172 3834 37196 3836
rect 37252 3834 37258 3836
rect 37012 3782 37014 3834
rect 37194 3782 37196 3834
rect 36950 3780 36956 3782
rect 37012 3780 37036 3782
rect 37092 3780 37116 3782
rect 37172 3780 37196 3782
rect 37252 3780 37258 3782
rect 36950 3771 37258 3780
rect 36950 2748 37258 2757
rect 36950 2746 36956 2748
rect 37012 2746 37036 2748
rect 37092 2746 37116 2748
rect 37172 2746 37196 2748
rect 37252 2746 37258 2748
rect 37012 2694 37014 2746
rect 37194 2694 37196 2746
rect 36950 2692 36956 2694
rect 37012 2692 37036 2694
rect 37092 2692 37116 2694
rect 37172 2692 37196 2694
rect 37252 2692 37258 2694
rect 36950 2683 37258 2692
rect 37476 2650 37504 8078
rect 37610 5468 37918 5477
rect 37610 5466 37616 5468
rect 37672 5466 37696 5468
rect 37752 5466 37776 5468
rect 37832 5466 37856 5468
rect 37912 5466 37918 5468
rect 37672 5414 37674 5466
rect 37854 5414 37856 5466
rect 37610 5412 37616 5414
rect 37672 5412 37696 5414
rect 37752 5412 37776 5414
rect 37832 5412 37856 5414
rect 37912 5412 37918 5414
rect 37610 5403 37918 5412
rect 37610 4380 37918 4389
rect 37610 4378 37616 4380
rect 37672 4378 37696 4380
rect 37752 4378 37776 4380
rect 37832 4378 37856 4380
rect 37912 4378 37918 4380
rect 37672 4326 37674 4378
rect 37854 4326 37856 4378
rect 37610 4324 37616 4326
rect 37672 4324 37696 4326
rect 37752 4324 37776 4326
rect 37832 4324 37856 4326
rect 37912 4324 37918 4326
rect 37610 4315 37918 4324
rect 37610 3292 37918 3301
rect 37610 3290 37616 3292
rect 37672 3290 37696 3292
rect 37752 3290 37776 3292
rect 37832 3290 37856 3292
rect 37912 3290 37918 3292
rect 37672 3238 37674 3290
rect 37854 3238 37856 3290
rect 37610 3236 37616 3238
rect 37672 3236 37696 3238
rect 37752 3236 37776 3238
rect 37832 3236 37856 3238
rect 37912 3236 37918 3238
rect 37610 3227 37918 3236
rect 31024 2644 31076 2650
rect 31024 2586 31076 2592
rect 31852 2644 31904 2650
rect 31852 2586 31904 2592
rect 32956 2644 33008 2650
rect 32956 2586 33008 2592
rect 34244 2644 34296 2650
rect 34244 2586 34296 2592
rect 35072 2644 35124 2650
rect 35072 2586 35124 2592
rect 36176 2644 36228 2650
rect 36176 2586 36228 2592
rect 37464 2644 37516 2650
rect 37464 2586 37516 2592
rect 38396 2514 38424 8092
rect 39514 8078 39896 8106
rect 40618 8078 40724 8106
rect 41722 8078 42012 8106
rect 39868 2582 39896 8078
rect 40696 2582 40724 8078
rect 41984 2582 42012 8078
rect 42812 2650 42840 8092
rect 43444 5772 43496 5778
rect 43444 5714 43496 5720
rect 43456 5574 43484 5714
rect 43444 5568 43496 5574
rect 43444 5510 43496 5516
rect 42800 2644 42852 2650
rect 42800 2586 42852 2592
rect 43916 2582 43944 8092
rect 45034 8078 45232 8106
rect 45204 2650 45232 8078
rect 46860 4486 46888 47495
rect 46940 5840 46992 5846
rect 46940 5782 46992 5788
rect 46952 5710 46980 5782
rect 46940 5704 46992 5710
rect 46940 5646 46992 5652
rect 47228 4554 47256 49671
rect 47492 47592 47544 47598
rect 47492 47534 47544 47540
rect 47398 46608 47454 46617
rect 47398 46543 47454 46552
rect 47412 8022 47440 46543
rect 47400 8016 47452 8022
rect 47400 7958 47452 7964
rect 47504 7818 47532 47534
rect 47596 8634 47624 88402
rect 47688 49842 47716 91462
rect 47780 50182 47808 91530
rect 47860 91180 47912 91186
rect 47860 91122 47912 91128
rect 47768 50176 47820 50182
rect 47768 50118 47820 50124
rect 47676 49836 47728 49842
rect 47676 49778 47728 49784
rect 47768 49496 47820 49502
rect 47768 49438 47820 49444
rect 47780 46714 47808 49438
rect 47872 49065 47900 91122
rect 47964 49094 47992 91666
rect 48136 91112 48188 91118
rect 48136 91054 48188 91060
rect 48044 90976 48096 90982
rect 48044 90918 48096 90924
rect 47952 49088 48004 49094
rect 47858 49056 47914 49065
rect 47952 49030 48004 49036
rect 47858 48991 47914 49000
rect 47952 48544 48004 48550
rect 47952 48486 48004 48492
rect 47768 46708 47820 46714
rect 47768 46650 47820 46656
rect 47676 46640 47728 46646
rect 47676 46582 47728 46588
rect 47584 8628 47636 8634
rect 47584 8570 47636 8576
rect 47688 7954 47716 46582
rect 47676 7948 47728 7954
rect 47676 7890 47728 7896
rect 47492 7812 47544 7818
rect 47492 7754 47544 7760
rect 47780 5778 47808 46650
rect 47860 46572 47912 46578
rect 47860 46514 47912 46520
rect 47872 5846 47900 46514
rect 47964 7886 47992 48486
rect 48056 46850 48084 90918
rect 48148 49162 48176 91054
rect 48228 91044 48280 91050
rect 48228 90986 48280 90992
rect 48240 49502 48268 90986
rect 50264 88876 50292 91802
rect 51092 91526 51120 92074
rect 52472 91594 52500 92142
rect 52644 92064 52696 92070
rect 52696 92012 52776 92018
rect 52644 92006 52776 92012
rect 52656 91990 52776 92006
rect 52748 91662 52776 91990
rect 53760 91662 53788 95406
rect 54668 95328 54720 95334
rect 54668 95270 54720 95276
rect 55956 95328 56008 95334
rect 55956 95270 56008 95276
rect 56876 95328 56928 95334
rect 56876 95270 56928 95276
rect 58256 95328 58308 95334
rect 58256 95270 58308 95276
rect 52736 91656 52788 91662
rect 52736 91598 52788 91604
rect 53748 91656 53800 91662
rect 53748 91598 53800 91604
rect 52460 91588 52512 91594
rect 52460 91530 52512 91536
rect 51080 91520 51132 91526
rect 51080 91462 51132 91468
rect 51092 91254 51120 91462
rect 51080 91248 51132 91254
rect 51080 91190 51132 91196
rect 51092 88890 51120 91190
rect 52472 91050 52500 91530
rect 52748 91322 52776 91598
rect 53840 91588 53892 91594
rect 53840 91530 53892 91536
rect 53748 91520 53800 91526
rect 53748 91462 53800 91468
rect 52736 91316 52788 91322
rect 52736 91258 52788 91264
rect 52460 91044 52512 91050
rect 52460 90986 52512 90992
rect 52748 88890 52776 91258
rect 51092 88862 51382 88890
rect 52486 88862 52776 88890
rect 53196 88528 53248 88534
rect 53760 88482 53788 91462
rect 53852 90982 53880 91530
rect 53840 90976 53892 90982
rect 53840 90918 53892 90924
rect 54680 88876 54708 95270
rect 55968 88890 55996 95270
rect 55798 88862 55996 88890
rect 56888 88876 56916 95270
rect 58268 88890 58296 95270
rect 58006 88862 58296 88890
rect 59096 88876 59124 95406
rect 62580 95396 62632 95402
rect 62580 95338 62632 95344
rect 60188 95328 60240 95334
rect 60188 95270 60240 95276
rect 61476 95328 61528 95334
rect 61476 95270 61528 95276
rect 60200 88876 60228 95270
rect 61488 88890 61516 95270
rect 62592 88890 62620 95338
rect 61318 88862 61516 88890
rect 62422 88862 62620 88890
rect 63512 88876 63540 95406
rect 65800 95396 65852 95402
rect 65800 95338 65852 95344
rect 67088 95396 67140 95402
rect 67088 95338 67140 95344
rect 64604 95328 64656 95334
rect 64604 95270 64656 95276
rect 64616 88876 64644 95270
rect 65812 88890 65840 95338
rect 67100 88890 67128 95338
rect 67916 95328 67968 95334
rect 67916 95270 67968 95276
rect 69020 95328 69072 95334
rect 69020 95270 69072 95276
rect 65734 88862 65840 88890
rect 66838 88862 67128 88890
rect 67928 88876 67956 95270
rect 69032 88876 69060 95270
rect 70320 88890 70348 95474
rect 70150 88862 70348 88890
rect 71240 88876 71268 95474
rect 72252 93854 72280 95474
rect 72950 95228 73258 95237
rect 72950 95226 72956 95228
rect 73012 95226 73036 95228
rect 73092 95226 73116 95228
rect 73172 95226 73196 95228
rect 73252 95226 73258 95228
rect 73012 95174 73014 95226
rect 73194 95174 73196 95226
rect 72950 95172 72956 95174
rect 73012 95172 73036 95174
rect 73092 95172 73116 95174
rect 73172 95172 73196 95174
rect 73252 95172 73258 95174
rect 72950 95163 73258 95172
rect 72950 94140 73258 94149
rect 72950 94138 72956 94140
rect 73012 94138 73036 94140
rect 73092 94138 73116 94140
rect 73172 94138 73196 94140
rect 73252 94138 73258 94140
rect 73012 94086 73014 94138
rect 73194 94086 73196 94138
rect 72950 94084 72956 94086
rect 73012 94084 73036 94086
rect 73092 94084 73116 94086
rect 73172 94084 73196 94086
rect 73252 94084 73258 94086
rect 72950 94075 73258 94084
rect 72252 93826 72372 93854
rect 72344 88876 72372 93826
rect 72950 93052 73258 93061
rect 72950 93050 72956 93052
rect 73012 93050 73036 93052
rect 73092 93050 73116 93052
rect 73172 93050 73196 93052
rect 73252 93050 73258 93052
rect 73012 92998 73014 93050
rect 73194 92998 73196 93050
rect 72950 92996 72956 92998
rect 73012 92996 73036 92998
rect 73092 92996 73116 92998
rect 73172 92996 73196 92998
rect 73252 92996 73258 92998
rect 72950 92987 73258 92996
rect 72950 91964 73258 91973
rect 72950 91962 72956 91964
rect 73012 91962 73036 91964
rect 73092 91962 73116 91964
rect 73172 91962 73196 91964
rect 73252 91962 73258 91964
rect 73012 91910 73014 91962
rect 73194 91910 73196 91962
rect 72950 91908 72956 91910
rect 73012 91908 73036 91910
rect 73092 91908 73116 91910
rect 73172 91908 73196 91910
rect 73252 91908 73258 91910
rect 72950 91899 73258 91908
rect 73540 88890 73568 95474
rect 73610 94684 73918 94693
rect 73610 94682 73616 94684
rect 73672 94682 73696 94684
rect 73752 94682 73776 94684
rect 73832 94682 73856 94684
rect 73912 94682 73918 94684
rect 73672 94630 73674 94682
rect 73854 94630 73856 94682
rect 73610 94628 73616 94630
rect 73672 94628 73696 94630
rect 73752 94628 73776 94630
rect 73832 94628 73856 94630
rect 73912 94628 73918 94630
rect 73610 94619 73918 94628
rect 73610 93596 73918 93605
rect 73610 93594 73616 93596
rect 73672 93594 73696 93596
rect 73752 93594 73776 93596
rect 73832 93594 73856 93596
rect 73912 93594 73918 93596
rect 73672 93542 73674 93594
rect 73854 93542 73856 93594
rect 73610 93540 73616 93542
rect 73672 93540 73696 93542
rect 73752 93540 73776 93542
rect 73832 93540 73856 93542
rect 73912 93540 73918 93542
rect 73610 93531 73918 93540
rect 73610 92508 73918 92517
rect 73610 92506 73616 92508
rect 73672 92506 73696 92508
rect 73752 92506 73776 92508
rect 73832 92506 73856 92508
rect 73912 92506 73918 92508
rect 73672 92454 73674 92506
rect 73854 92454 73856 92506
rect 73610 92452 73616 92454
rect 73672 92452 73696 92454
rect 73752 92452 73776 92454
rect 73832 92452 73856 92454
rect 73912 92452 73918 92454
rect 73610 92443 73918 92452
rect 73610 91420 73918 91429
rect 73610 91418 73616 91420
rect 73672 91418 73696 91420
rect 73752 91418 73776 91420
rect 73832 91418 73856 91420
rect 73912 91418 73918 91420
rect 73672 91366 73674 91418
rect 73854 91366 73856 91418
rect 73610 91364 73616 91366
rect 73672 91364 73696 91366
rect 73752 91364 73776 91366
rect 73832 91364 73856 91366
rect 73912 91364 73918 91366
rect 73610 91355 73918 91364
rect 74828 88890 74856 95474
rect 75748 88890 75776 95474
rect 73462 88862 73568 88890
rect 74566 88862 74856 88890
rect 75670 88862 75776 88890
rect 76760 88876 76788 95474
rect 78048 88890 78076 95474
rect 77878 88862 78076 88890
rect 78968 88876 78996 95474
rect 80072 88876 80100 95474
rect 81268 88890 81296 95474
rect 82556 88890 82584 95474
rect 88156 94240 88208 94246
rect 88156 94182 88208 94188
rect 88064 93696 88116 93702
rect 88064 93638 88116 93644
rect 87788 93220 87840 93226
rect 87788 93162 87840 93168
rect 87236 93152 87288 93158
rect 87236 93094 87288 93100
rect 87696 93152 87748 93158
rect 87696 93094 87748 93100
rect 83372 92948 83424 92954
rect 83372 92890 83424 92896
rect 81190 88862 81296 88890
rect 82294 88862 82584 88890
rect 83384 88876 83412 92890
rect 86408 92880 86460 92886
rect 86408 92822 86460 92828
rect 86774 92848 86830 92857
rect 86224 92200 86276 92206
rect 86222 92168 86224 92177
rect 86316 92200 86368 92206
rect 86276 92168 86278 92177
rect 86316 92142 86368 92148
rect 86222 92103 86278 92112
rect 85672 92064 85724 92070
rect 85672 92006 85724 92012
rect 85948 92064 86000 92070
rect 85948 92006 86000 92012
rect 86040 92064 86092 92070
rect 86040 92006 86092 92012
rect 84476 91656 84528 91662
rect 84476 91598 84528 91604
rect 85210 91624 85266 91633
rect 84488 88876 84516 91598
rect 85210 91559 85212 91568
rect 85264 91559 85266 91568
rect 85212 91530 85264 91536
rect 85028 91520 85080 91526
rect 85028 91462 85080 91468
rect 85396 91520 85448 91526
rect 85396 91462 85448 91468
rect 85040 89690 85068 91462
rect 85408 91186 85436 91462
rect 85396 91180 85448 91186
rect 85396 91122 85448 91128
rect 85028 89684 85080 89690
rect 85028 89626 85080 89632
rect 85684 89350 85712 92006
rect 85856 91656 85908 91662
rect 85856 91598 85908 91604
rect 85764 91520 85816 91526
rect 85764 91462 85816 91468
rect 85776 91118 85804 91462
rect 85764 91112 85816 91118
rect 85764 91054 85816 91060
rect 85868 89842 85896 91598
rect 85960 91225 85988 92006
rect 86052 91730 86080 92006
rect 86328 91866 86356 92142
rect 86316 91860 86368 91866
rect 86316 91802 86368 91808
rect 86040 91724 86092 91730
rect 86040 91666 86092 91672
rect 86316 91520 86368 91526
rect 86316 91462 86368 91468
rect 85946 91216 86002 91225
rect 85946 91151 86002 91160
rect 86038 89856 86094 89865
rect 85868 89814 86038 89842
rect 86038 89791 86094 89800
rect 85672 89344 85724 89350
rect 85672 89286 85724 89292
rect 53248 88476 53788 88482
rect 53196 88470 53788 88476
rect 53208 88454 53788 88470
rect 85684 88466 85712 89286
rect 86052 89078 86080 89791
rect 86040 89072 86092 89078
rect 86040 89014 86092 89020
rect 86328 89010 86356 91462
rect 86420 91361 86448 92822
rect 86774 92783 86776 92792
rect 86828 92783 86830 92792
rect 86776 92754 86828 92760
rect 87142 92712 87198 92721
rect 87142 92647 87144 92656
rect 87196 92647 87198 92656
rect 87144 92618 87196 92624
rect 86592 92608 86644 92614
rect 86590 92576 86592 92585
rect 87052 92608 87104 92614
rect 86644 92576 86646 92585
rect 86590 92511 86646 92520
rect 87050 92576 87052 92585
rect 87104 92576 87106 92585
rect 87050 92511 87106 92520
rect 87248 92274 87276 93094
rect 87328 92744 87380 92750
rect 87328 92686 87380 92692
rect 87236 92268 87288 92274
rect 87236 92210 87288 92216
rect 86500 92064 86552 92070
rect 86500 92006 86552 92012
rect 86684 92064 86736 92070
rect 86684 92006 86736 92012
rect 86776 92064 86828 92070
rect 86776 92006 86828 92012
rect 87052 92064 87104 92070
rect 87052 92006 87104 92012
rect 86406 91352 86462 91361
rect 86406 91287 86462 91296
rect 86512 89146 86540 92006
rect 86696 91633 86724 92006
rect 86682 91624 86738 91633
rect 86682 91559 86738 91568
rect 86684 91520 86736 91526
rect 86684 91462 86736 91468
rect 86500 89140 86552 89146
rect 86500 89082 86552 89088
rect 86316 89004 86368 89010
rect 86316 88946 86368 88952
rect 86328 88534 86356 88946
rect 86316 88528 86368 88534
rect 86512 88505 86540 89082
rect 86316 88470 86368 88476
rect 86498 88496 86554 88505
rect 85672 88460 85724 88466
rect 86498 88431 86554 88440
rect 85672 88402 85724 88408
rect 86696 81433 86724 91462
rect 86788 87281 86816 92006
rect 86868 88460 86920 88466
rect 86868 88402 86920 88408
rect 86774 87272 86830 87281
rect 86774 87207 86830 87216
rect 86880 85921 86908 88402
rect 86958 87000 87014 87009
rect 86958 86935 87014 86944
rect 86866 85912 86922 85921
rect 86866 85847 86922 85856
rect 86682 81424 86738 81433
rect 86682 81359 86738 81368
rect 86682 71360 86738 71369
rect 86682 71295 86738 71304
rect 85580 50652 85632 50658
rect 85580 50594 85632 50600
rect 85592 50561 85620 50594
rect 85578 50552 85634 50561
rect 85578 50487 85634 50496
rect 52644 50448 52696 50454
rect 52696 50396 53038 50402
rect 52644 50390 53038 50396
rect 52656 50374 53038 50390
rect 51552 50250 51934 50266
rect 51540 50244 51934 50250
rect 51592 50238 51934 50244
rect 51540 50186 51592 50192
rect 50436 50176 50488 50182
rect 50488 50124 50830 50130
rect 50436 50118 50830 50124
rect 49712 49842 49740 50116
rect 50448 50102 50830 50118
rect 49700 49836 49752 49842
rect 49700 49778 49752 49784
rect 48228 49496 48280 49502
rect 48228 49438 48280 49444
rect 48226 49328 48282 49337
rect 48226 49263 48282 49272
rect 48136 49156 48188 49162
rect 48136 49098 48188 49104
rect 48240 49094 48268 49263
rect 48228 49088 48280 49094
rect 48228 49030 48280 49036
rect 51172 47728 51224 47734
rect 51172 47670 51224 47676
rect 48136 47524 48188 47530
rect 48136 47466 48188 47472
rect 48044 46844 48096 46850
rect 48044 46786 48096 46792
rect 48056 46442 48084 46786
rect 48044 46436 48096 46442
rect 48044 46378 48096 46384
rect 47952 7880 48004 7886
rect 47952 7822 48004 7828
rect 47860 5840 47912 5846
rect 47860 5782 47912 5788
rect 47768 5772 47820 5778
rect 47768 5714 47820 5720
rect 48056 5710 48084 46378
rect 48148 46374 48176 47466
rect 51080 46708 51132 46714
rect 51080 46650 51132 46656
rect 51092 46617 51120 46650
rect 51078 46608 51134 46617
rect 51078 46543 51134 46552
rect 51184 46510 51212 47670
rect 55232 46866 55260 50116
rect 56060 50102 56350 50130
rect 57164 50102 57454 50130
rect 58268 50102 58558 50130
rect 59372 50102 59662 50130
rect 56060 46866 56088 50102
rect 57164 46866 57192 50102
rect 58268 46866 58296 50102
rect 59372 46866 59400 50102
rect 60752 46866 60780 50116
rect 61580 50102 61870 50130
rect 62684 50102 62974 50130
rect 63788 50102 64078 50130
rect 64892 50102 65182 50130
rect 61580 46866 61608 50102
rect 62684 46866 62712 50102
rect 63788 46866 63816 50102
rect 64892 46866 64920 50102
rect 66272 46866 66300 50116
rect 67100 50102 67390 50130
rect 68204 50102 68494 50130
rect 69308 50102 69598 50130
rect 70412 50102 70702 50130
rect 67100 46866 67128 50102
rect 68204 46866 68232 50102
rect 69308 46866 69336 50102
rect 70412 46866 70440 50102
rect 71792 46866 71820 50116
rect 72620 50102 72910 50130
rect 73724 50102 74014 50130
rect 74828 50102 75118 50130
rect 75932 50102 76222 50130
rect 72620 46866 72648 50102
rect 73724 46866 73752 50102
rect 74828 46866 74856 50102
rect 75932 46866 75960 50102
rect 77312 46866 77340 50116
rect 78140 50102 78430 50130
rect 79244 50102 79534 50130
rect 80348 50102 80638 50130
rect 81452 50102 81742 50130
rect 78140 46866 78168 50102
rect 79244 46866 79272 50102
rect 80348 46866 80376 50102
rect 81452 46866 81480 50102
rect 82832 46866 82860 50116
rect 83660 50102 83950 50130
rect 84764 50102 85054 50130
rect 83660 46866 83688 50102
rect 84764 46866 84792 50102
rect 86696 49910 86724 71295
rect 86774 68368 86830 68377
rect 86774 68303 86830 68312
rect 86684 49904 86736 49910
rect 86684 49846 86736 49852
rect 85578 49736 85634 49745
rect 85578 49671 85634 49680
rect 52486 46850 52592 46866
rect 52486 46844 52604 46850
rect 52486 46838 52552 46844
rect 54694 46838 55260 46866
rect 55798 46838 56088 46866
rect 56902 46838 57192 46866
rect 58006 46838 58296 46866
rect 59110 46838 59400 46866
rect 60214 46838 60780 46866
rect 61318 46838 61608 46866
rect 62422 46838 62712 46866
rect 63526 46838 63816 46866
rect 64630 46838 64920 46866
rect 65734 46838 66300 46866
rect 66838 46838 67128 46866
rect 67942 46838 68232 46866
rect 69046 46838 69336 46866
rect 70150 46838 70440 46866
rect 71254 46838 71820 46866
rect 72358 46838 72648 46866
rect 73462 46838 73752 46866
rect 74566 46838 74856 46866
rect 75670 46838 75960 46866
rect 76774 46838 77340 46866
rect 77878 46838 78168 46866
rect 78982 46838 79272 46866
rect 80086 46838 80376 46866
rect 81190 46838 81480 46866
rect 82294 46838 82860 46866
rect 83398 46838 83688 46866
rect 84502 46838 84792 46866
rect 52552 46786 52604 46792
rect 51448 46776 51500 46782
rect 51382 46724 51448 46730
rect 51382 46718 51500 46724
rect 51382 46702 51488 46718
rect 53208 46578 53590 46594
rect 53196 46572 53590 46578
rect 53248 46566 53590 46572
rect 53196 46514 53248 46520
rect 51172 46504 51224 46510
rect 49896 46442 50278 46458
rect 85592 46481 85620 49671
rect 86684 48476 86736 48482
rect 86684 48418 86736 48424
rect 51172 46446 51224 46452
rect 85578 46472 85634 46481
rect 48228 46436 48280 46442
rect 48228 46378 48280 46384
rect 49884 46436 50278 46442
rect 49936 46430 50278 46436
rect 85578 46407 85634 46416
rect 49884 46378 49936 46384
rect 48136 46368 48188 46374
rect 48136 46310 48188 46316
rect 48240 6254 48268 46378
rect 86696 43353 86724 48418
rect 86788 48210 86816 68303
rect 86972 57225 87000 86935
rect 87064 78577 87092 92006
rect 87248 91866 87276 92210
rect 87236 91860 87288 91866
rect 87236 91802 87288 91808
rect 87340 91594 87368 92686
rect 87604 92676 87656 92682
rect 87604 92618 87656 92624
rect 87512 92608 87564 92614
rect 87512 92550 87564 92556
rect 87524 92138 87552 92550
rect 87512 92132 87564 92138
rect 87512 92074 87564 92080
rect 87420 92064 87472 92070
rect 87420 92006 87472 92012
rect 87144 91588 87196 91594
rect 87144 91530 87196 91536
rect 87328 91588 87380 91594
rect 87328 91530 87380 91536
rect 87156 87961 87184 91530
rect 87142 87952 87198 87961
rect 87142 87887 87198 87896
rect 87340 87825 87368 91530
rect 87326 87816 87382 87825
rect 87326 87751 87382 87760
rect 87142 87136 87198 87145
rect 87142 87071 87198 87080
rect 87050 78568 87106 78577
rect 87050 78503 87106 78512
rect 87156 71641 87184 87071
rect 87432 75721 87460 92006
rect 87616 91730 87644 92618
rect 87708 92410 87736 93094
rect 87696 92404 87748 92410
rect 87696 92346 87748 92352
rect 87800 92274 87828 93162
rect 87880 93152 87932 93158
rect 87880 93094 87932 93100
rect 87788 92268 87840 92274
rect 87788 92210 87840 92216
rect 87800 92177 87828 92210
rect 87786 92168 87842 92177
rect 87696 92132 87748 92138
rect 87786 92103 87842 92112
rect 87696 92074 87748 92080
rect 87604 91724 87656 91730
rect 87604 91666 87656 91672
rect 87512 91588 87564 91594
rect 87512 91530 87564 91536
rect 87524 85241 87552 91530
rect 87602 87272 87658 87281
rect 87602 87207 87658 87216
rect 87510 85232 87566 85241
rect 87510 85167 87566 85176
rect 87616 80054 87644 87207
rect 87708 86601 87736 92074
rect 87892 91594 87920 93094
rect 87972 92744 88024 92750
rect 87970 92712 87972 92721
rect 88024 92712 88026 92721
rect 88076 92682 88104 93638
rect 87970 92647 88026 92656
rect 88064 92676 88116 92682
rect 88064 92618 88116 92624
rect 88168 92614 88196 94182
rect 88616 93968 88668 93974
rect 88616 93910 88668 93916
rect 88340 93900 88392 93906
rect 88340 93842 88392 93848
rect 88524 93900 88576 93906
rect 88524 93842 88576 93848
rect 88628 93854 88656 93910
rect 88156 92608 88208 92614
rect 88156 92550 88208 92556
rect 88352 92206 88380 93842
rect 88536 93378 88564 93842
rect 88628 93826 88748 93854
rect 88536 93350 88656 93378
rect 88524 93220 88576 93226
rect 88524 93162 88576 93168
rect 88432 92608 88484 92614
rect 88432 92550 88484 92556
rect 88340 92200 88392 92206
rect 88340 92142 88392 92148
rect 88064 92132 88116 92138
rect 88064 92074 88116 92080
rect 87880 91588 87932 91594
rect 87880 91530 87932 91536
rect 87972 91520 88024 91526
rect 87972 91462 88024 91468
rect 87694 86592 87750 86601
rect 87694 86527 87750 86536
rect 87984 82521 88012 91462
rect 88076 83881 88104 92074
rect 88340 91792 88392 91798
rect 88340 91734 88392 91740
rect 88248 91588 88300 91594
rect 88248 91530 88300 91536
rect 88062 83872 88118 83881
rect 88062 83807 88118 83816
rect 87970 82512 88026 82521
rect 87970 82447 88026 82456
rect 87524 80026 87644 80054
rect 87418 75712 87474 75721
rect 87418 75647 87474 75656
rect 87524 74361 87552 80026
rect 88260 79801 88288 91530
rect 88352 88505 88380 91734
rect 88444 89185 88472 92550
rect 88536 91662 88564 93162
rect 88524 91656 88576 91662
rect 88524 91598 88576 91604
rect 88628 91594 88656 93350
rect 88720 92342 88748 93826
rect 88800 93152 88852 93158
rect 88800 93094 88852 93100
rect 88708 92336 88760 92342
rect 88708 92278 88760 92284
rect 88708 92200 88760 92206
rect 88708 92142 88760 92148
rect 88616 91588 88668 91594
rect 88616 91530 88668 91536
rect 88524 91520 88576 91526
rect 88524 91462 88576 91468
rect 88430 89176 88486 89185
rect 88430 89111 88486 89120
rect 88338 88496 88394 88505
rect 88338 88431 88394 88440
rect 88338 87408 88394 87417
rect 88338 87343 88394 87352
rect 88246 79792 88302 79801
rect 88246 79727 88302 79736
rect 87510 74352 87566 74361
rect 87510 74287 87566 74296
rect 87142 71632 87198 71641
rect 87142 71567 87198 71576
rect 88352 68921 88380 87343
rect 88536 85105 88564 91462
rect 88616 88528 88668 88534
rect 88616 88470 88668 88476
rect 88522 85096 88578 85105
rect 88522 85031 88578 85040
rect 88432 81796 88484 81802
rect 88432 81738 88484 81744
rect 88444 73001 88472 81738
rect 88628 80054 88656 88470
rect 88720 86465 88748 92142
rect 88812 92070 88840 93094
rect 89352 92676 89404 92682
rect 89352 92618 89404 92624
rect 89260 92404 89312 92410
rect 89260 92346 89312 92352
rect 88800 92064 88852 92070
rect 88800 92006 88852 92012
rect 88706 86456 88762 86465
rect 88706 86391 88762 86400
rect 88812 81802 88840 92006
rect 89168 91860 89220 91866
rect 89168 91802 89220 91808
rect 89076 91724 89128 91730
rect 89076 91666 89128 91672
rect 88984 91656 89036 91662
rect 88984 91598 89036 91604
rect 88996 82385 89024 91598
rect 88982 82376 89038 82385
rect 88982 82311 89038 82320
rect 88800 81796 88852 81802
rect 88800 81738 88852 81744
rect 89088 81025 89116 91666
rect 89074 81016 89130 81025
rect 89074 80951 89130 80960
rect 88536 80026 88656 80054
rect 88430 72992 88486 73001
rect 88430 72927 88486 72936
rect 88536 70281 88564 80026
rect 89180 78305 89208 91802
rect 89166 78296 89222 78305
rect 89166 78231 89222 78240
rect 89168 77104 89220 77110
rect 89168 77046 89220 77052
rect 89180 76945 89208 77046
rect 89166 76936 89222 76945
rect 89166 76871 89222 76880
rect 89166 75576 89222 75585
rect 89272 75562 89300 92346
rect 89364 77110 89392 92618
rect 89536 92268 89588 92274
rect 89536 92210 89588 92216
rect 89444 91588 89496 91594
rect 89444 91530 89496 91536
rect 89456 79937 89484 91530
rect 89548 83473 89576 92210
rect 89534 83464 89590 83473
rect 89534 83399 89590 83408
rect 89442 79928 89498 79937
rect 89442 79863 89498 79872
rect 89352 77104 89404 77110
rect 89352 77046 89404 77052
rect 89222 75534 89300 75562
rect 89166 75511 89222 75520
rect 89074 71496 89130 71505
rect 89074 71431 89130 71440
rect 89088 70394 89116 71431
rect 89088 70366 89208 70394
rect 88522 70272 88578 70281
rect 88522 70207 88578 70216
rect 88338 68912 88394 68921
rect 88338 68847 88394 68856
rect 88982 68776 89038 68785
rect 88982 68711 89038 68720
rect 87602 64696 87658 64705
rect 87602 64631 87658 64640
rect 87050 61568 87106 61577
rect 87050 61503 87106 61512
rect 86958 57216 87014 57225
rect 86958 57151 87014 57160
rect 87064 55214 87092 61503
rect 87142 58032 87198 58041
rect 87142 57967 87198 57976
rect 86972 55186 87092 55214
rect 86972 50289 87000 55186
rect 87156 51218 87184 57967
rect 87418 56672 87474 56681
rect 87418 56607 87474 56616
rect 87326 53952 87382 53961
rect 87326 53887 87382 53896
rect 87234 52592 87290 52601
rect 87234 52527 87290 52536
rect 87064 51190 87184 51218
rect 87064 50697 87092 51190
rect 87142 51096 87198 51105
rect 87142 51031 87144 51040
rect 87196 51031 87198 51040
rect 87144 51002 87196 51008
rect 87142 50960 87198 50969
rect 87142 50895 87198 50904
rect 87050 50688 87106 50697
rect 87050 50623 87106 50632
rect 86958 50280 87014 50289
rect 86958 50215 87014 50224
rect 86868 49768 86920 49774
rect 86868 49710 86920 49716
rect 86776 48204 86828 48210
rect 86776 48146 86828 48152
rect 86682 43344 86738 43353
rect 86682 43279 86738 43288
rect 86880 41993 86908 49710
rect 87156 49162 87184 50895
rect 87248 49337 87276 52527
rect 87234 49328 87290 49337
rect 87234 49263 87290 49272
rect 87144 49156 87196 49162
rect 87144 49098 87196 49104
rect 87340 49065 87368 53887
rect 87432 49434 87460 56607
rect 87616 50833 87644 64631
rect 88890 63336 88946 63345
rect 88890 63271 88946 63280
rect 87694 61976 87750 61985
rect 87694 61911 87750 61920
rect 87602 50824 87658 50833
rect 87602 50759 87658 50768
rect 87708 49473 87736 61911
rect 88798 60616 88854 60625
rect 88798 60551 88854 60560
rect 87786 59256 87842 59265
rect 87786 59191 87842 59200
rect 87694 49464 87750 49473
rect 87420 49428 87472 49434
rect 87694 49399 87750 49408
rect 87420 49370 87472 49376
rect 87326 49056 87382 49065
rect 87326 48991 87382 49000
rect 87800 48822 87828 59191
rect 88614 57896 88670 57905
rect 88614 57831 88670 57840
rect 88522 55176 88578 55185
rect 88522 55111 88578 55120
rect 88338 53816 88394 53825
rect 88338 53751 88394 53760
rect 88352 50862 88380 53751
rect 88430 52456 88486 52465
rect 88430 52391 88486 52400
rect 88340 50856 88392 50862
rect 88340 50798 88392 50804
rect 88444 50590 88472 52391
rect 88432 50584 88484 50590
rect 88432 50526 88484 50532
rect 88536 49638 88564 55111
rect 88524 49632 88576 49638
rect 88524 49574 88576 49580
rect 88628 49230 88656 57831
rect 88706 56536 88762 56545
rect 88706 56471 88762 56480
rect 88616 49224 88668 49230
rect 88616 49166 88668 49172
rect 87788 48816 87840 48822
rect 87788 48758 87840 48764
rect 88720 48754 88748 56471
rect 88812 49298 88840 60551
rect 88904 49366 88932 63271
rect 88892 49360 88944 49366
rect 88892 49302 88944 49308
rect 88800 49292 88852 49298
rect 88800 49234 88852 49240
rect 88708 48748 88760 48754
rect 88708 48690 88760 48696
rect 87328 48544 87380 48550
rect 87328 48486 87380 48492
rect 87050 47696 87106 47705
rect 87050 47631 87106 47640
rect 86960 47388 87012 47394
rect 86960 47330 87012 47336
rect 86972 44305 87000 47330
rect 86958 44296 87014 44305
rect 86958 44231 87014 44240
rect 86866 41984 86922 41993
rect 86866 41919 86922 41928
rect 86682 27976 86738 27985
rect 86682 27911 86738 27920
rect 86590 13696 86646 13705
rect 86590 13631 86646 13640
rect 48688 9648 48740 9654
rect 48688 9590 48740 9596
rect 48700 8226 48728 9590
rect 86406 8664 86462 8673
rect 49332 8628 49384 8634
rect 86604 8650 86632 13631
rect 86406 8599 86462 8608
rect 86512 8622 86632 8650
rect 49332 8570 49384 8576
rect 48688 8220 48740 8226
rect 48688 8162 48740 8168
rect 49344 8106 49372 8570
rect 86038 8392 86094 8401
rect 86038 8327 86094 8336
rect 84752 8288 84804 8294
rect 84752 8230 84804 8236
rect 85670 8256 85726 8265
rect 53840 8220 53892 8226
rect 53840 8162 53892 8168
rect 49344 8092 49726 8106
rect 49344 8078 49740 8092
rect 48228 6248 48280 6254
rect 48228 6190 48280 6196
rect 49712 5914 49740 8078
rect 50252 6248 50304 6254
rect 50252 6190 50304 6196
rect 50264 5914 50292 6190
rect 50816 6186 50844 8092
rect 50804 6180 50856 6186
rect 50804 6122 50856 6128
rect 50816 5914 50844 6122
rect 49700 5908 49752 5914
rect 49700 5850 49752 5856
rect 50252 5908 50304 5914
rect 50252 5850 50304 5856
rect 50804 5908 50856 5914
rect 50804 5850 50856 5856
rect 48044 5704 48096 5710
rect 48044 5646 48096 5652
rect 51920 5642 51948 8092
rect 51908 5636 51960 5642
rect 51908 5578 51960 5584
rect 53024 5574 53052 8092
rect 53012 5568 53064 5574
rect 53012 5510 53064 5516
rect 53852 5098 53880 8162
rect 55246 8078 55536 8106
rect 56350 8078 56456 8106
rect 53840 5092 53892 5098
rect 53840 5034 53892 5040
rect 47216 4548 47268 4554
rect 47216 4490 47268 4496
rect 46848 4480 46900 4486
rect 46848 4422 46900 4428
rect 45192 2644 45244 2650
rect 45192 2586 45244 2592
rect 39856 2576 39908 2582
rect 39856 2518 39908 2524
rect 40684 2576 40736 2582
rect 40684 2518 40736 2524
rect 41972 2576 42024 2582
rect 41972 2518 42024 2524
rect 43904 2576 43956 2582
rect 43904 2518 43956 2524
rect 38384 2508 38436 2514
rect 38384 2450 38436 2456
rect 55508 2446 55536 8078
rect 56428 2446 56456 8078
rect 57440 2446 57468 8092
rect 58558 8078 58756 8106
rect 58728 2446 58756 8078
rect 59648 2446 59676 8092
rect 60752 2446 60780 8092
rect 61870 8078 61976 8106
rect 62974 8078 63264 8106
rect 64078 8078 64184 8106
rect 61948 2446 61976 8078
rect 63236 2446 63264 8078
rect 64156 2446 64184 8078
rect 65168 2446 65196 8092
rect 66286 8078 66484 8106
rect 66456 2446 66484 8078
rect 67376 2446 67404 8092
rect 68480 6914 68508 8092
rect 69598 8078 69704 8106
rect 70702 8078 70992 8106
rect 68388 6886 68508 6914
rect 68388 2446 68416 6886
rect 69676 2446 69704 8078
rect 70964 2650 70992 8078
rect 71792 2650 71820 8092
rect 72896 6914 72924 8092
rect 74014 8078 74212 8106
rect 72804 6886 72924 6914
rect 72804 2650 72832 6886
rect 72950 6012 73258 6021
rect 72950 6010 72956 6012
rect 73012 6010 73036 6012
rect 73092 6010 73116 6012
rect 73172 6010 73196 6012
rect 73252 6010 73258 6012
rect 73012 5958 73014 6010
rect 73194 5958 73196 6010
rect 72950 5956 72956 5958
rect 73012 5956 73036 5958
rect 73092 5956 73116 5958
rect 73172 5956 73196 5958
rect 73252 5956 73258 5958
rect 72950 5947 73258 5956
rect 73610 5468 73918 5477
rect 73610 5466 73616 5468
rect 73672 5466 73696 5468
rect 73752 5466 73776 5468
rect 73832 5466 73856 5468
rect 73912 5466 73918 5468
rect 73672 5414 73674 5466
rect 73854 5414 73856 5466
rect 73610 5412 73616 5414
rect 73672 5412 73696 5414
rect 73752 5412 73776 5414
rect 73832 5412 73856 5414
rect 73912 5412 73918 5414
rect 73610 5403 73918 5412
rect 72950 4924 73258 4933
rect 72950 4922 72956 4924
rect 73012 4922 73036 4924
rect 73092 4922 73116 4924
rect 73172 4922 73196 4924
rect 73252 4922 73258 4924
rect 73012 4870 73014 4922
rect 73194 4870 73196 4922
rect 72950 4868 72956 4870
rect 73012 4868 73036 4870
rect 73092 4868 73116 4870
rect 73172 4868 73196 4870
rect 73252 4868 73258 4870
rect 72950 4859 73258 4868
rect 73610 4380 73918 4389
rect 73610 4378 73616 4380
rect 73672 4378 73696 4380
rect 73752 4378 73776 4380
rect 73832 4378 73856 4380
rect 73912 4378 73918 4380
rect 73672 4326 73674 4378
rect 73854 4326 73856 4378
rect 73610 4324 73616 4326
rect 73672 4324 73696 4326
rect 73752 4324 73776 4326
rect 73832 4324 73856 4326
rect 73912 4324 73918 4326
rect 73610 4315 73918 4324
rect 72950 3836 73258 3845
rect 72950 3834 72956 3836
rect 73012 3834 73036 3836
rect 73092 3834 73116 3836
rect 73172 3834 73196 3836
rect 73252 3834 73258 3836
rect 73012 3782 73014 3834
rect 73194 3782 73196 3834
rect 72950 3780 72956 3782
rect 73012 3780 73036 3782
rect 73092 3780 73116 3782
rect 73172 3780 73196 3782
rect 73252 3780 73258 3782
rect 72950 3771 73258 3780
rect 73610 3292 73918 3301
rect 73610 3290 73616 3292
rect 73672 3290 73696 3292
rect 73752 3290 73776 3292
rect 73832 3290 73856 3292
rect 73912 3290 73918 3292
rect 73672 3238 73674 3290
rect 73854 3238 73856 3290
rect 73610 3236 73616 3238
rect 73672 3236 73696 3238
rect 73752 3236 73776 3238
rect 73832 3236 73856 3238
rect 73912 3236 73918 3238
rect 73610 3227 73918 3236
rect 72950 2748 73258 2757
rect 72950 2746 72956 2748
rect 73012 2746 73036 2748
rect 73092 2746 73116 2748
rect 73172 2746 73196 2748
rect 73252 2746 73258 2748
rect 73012 2694 73014 2746
rect 73194 2694 73196 2746
rect 72950 2692 72956 2694
rect 73012 2692 73036 2694
rect 73092 2692 73116 2694
rect 73172 2692 73196 2694
rect 73252 2692 73258 2694
rect 72950 2683 73258 2692
rect 74184 2650 74212 8078
rect 75104 2650 75132 8092
rect 76222 8078 76328 8106
rect 77326 8078 77432 8106
rect 76300 2650 76328 8078
rect 77404 2650 77432 8078
rect 70952 2644 71004 2650
rect 70952 2586 71004 2592
rect 71780 2644 71832 2650
rect 71780 2586 71832 2592
rect 72792 2644 72844 2650
rect 72792 2586 72844 2592
rect 74172 2644 74224 2650
rect 74172 2586 74224 2592
rect 75092 2644 75144 2650
rect 75092 2586 75144 2592
rect 76288 2644 76340 2650
rect 76288 2586 76340 2592
rect 77392 2644 77444 2650
rect 77392 2586 77444 2592
rect 78416 2514 78444 8092
rect 79534 8078 79640 8106
rect 79612 2582 79640 8078
rect 80624 2582 80652 8092
rect 81742 8078 81940 8106
rect 81912 2582 81940 8078
rect 82832 2582 82860 8092
rect 83936 5166 83964 8092
rect 84764 7750 84792 8230
rect 86052 8226 86080 8327
rect 85670 8191 85726 8200
rect 86040 8220 86092 8226
rect 84752 7744 84804 7750
rect 84752 7686 84804 7692
rect 84764 5914 84792 7686
rect 85040 5914 85068 8092
rect 85304 7812 85356 7818
rect 85304 7754 85356 7760
rect 85316 5914 85344 7754
rect 85684 7682 85712 8191
rect 86040 8162 86092 8168
rect 85762 7984 85818 7993
rect 85762 7919 85818 7928
rect 85672 7676 85724 7682
rect 85672 7618 85724 7624
rect 84752 5908 84804 5914
rect 84752 5850 84804 5856
rect 85028 5908 85080 5914
rect 85028 5850 85080 5856
rect 85304 5908 85356 5914
rect 85304 5850 85356 5856
rect 85120 5840 85172 5846
rect 85118 5808 85120 5817
rect 85172 5808 85174 5817
rect 85118 5743 85174 5752
rect 85578 5672 85634 5681
rect 85578 5607 85580 5616
rect 85632 5607 85634 5616
rect 85580 5578 85632 5584
rect 85684 5370 85712 7618
rect 85776 7614 85804 7919
rect 85764 7608 85816 7614
rect 85764 7550 85816 7556
rect 85672 5364 85724 5370
rect 85672 5306 85724 5312
rect 83924 5160 83976 5166
rect 83924 5102 83976 5108
rect 85776 4826 85804 7550
rect 86052 5370 86080 8162
rect 86314 8120 86370 8129
rect 86314 8055 86370 8064
rect 86328 5914 86356 8055
rect 86316 5908 86368 5914
rect 86316 5850 86368 5856
rect 86328 5710 86356 5850
rect 86420 5710 86448 8599
rect 86316 5704 86368 5710
rect 86316 5646 86368 5652
rect 86408 5704 86460 5710
rect 86408 5646 86460 5652
rect 86512 5642 86540 8622
rect 86590 8528 86646 8537
rect 86590 8463 86646 8472
rect 86604 5914 86632 8463
rect 86592 5908 86644 5914
rect 86592 5850 86644 5856
rect 86500 5636 86552 5642
rect 86500 5578 86552 5584
rect 86498 5400 86554 5409
rect 86040 5364 86092 5370
rect 86696 5370 86724 27911
rect 86972 9602 87000 44231
rect 87064 39681 87092 47631
rect 87234 47424 87290 47433
rect 87234 47359 87290 47368
rect 87142 46608 87198 46617
rect 87142 46543 87198 46552
rect 87050 39672 87106 39681
rect 87050 39607 87106 39616
rect 87156 28257 87184 46543
rect 87248 37777 87276 47359
rect 87234 37768 87290 37777
rect 87234 37703 87290 37712
rect 87340 35057 87368 48486
rect 88996 48142 89024 68711
rect 89074 66056 89130 66065
rect 89074 65991 89130 66000
rect 89088 50998 89116 65991
rect 89076 50992 89128 50998
rect 89076 50934 89128 50940
rect 89180 49706 89208 70366
rect 89258 69864 89314 69873
rect 89258 69799 89314 69808
rect 89168 49700 89220 49706
rect 89168 49642 89220 49648
rect 89076 48612 89128 48618
rect 89076 48554 89128 48560
rect 88984 48136 89036 48142
rect 88984 48078 89036 48084
rect 88062 47968 88118 47977
rect 88062 47903 88118 47912
rect 87510 47832 87566 47841
rect 87510 47767 87566 47776
rect 87418 43208 87474 43217
rect 87418 43143 87474 43152
rect 87326 35048 87382 35057
rect 87326 34983 87382 34992
rect 87142 28248 87198 28257
rect 87142 28183 87198 28192
rect 87234 25528 87290 25537
rect 87234 25463 87290 25472
rect 87142 17368 87198 17377
rect 87142 17303 87198 17312
rect 87050 15464 87106 15473
rect 87050 15399 87106 15408
rect 86788 9574 87000 9602
rect 86498 5335 86500 5344
rect 86040 5306 86092 5312
rect 86552 5335 86554 5344
rect 86684 5364 86736 5370
rect 86500 5306 86552 5312
rect 86684 5306 86736 5312
rect 86788 5302 86816 9574
rect 86868 9512 86920 9518
rect 86868 9454 86920 9460
rect 86880 5778 86908 9454
rect 86868 5772 86920 5778
rect 86868 5714 86920 5720
rect 87064 5710 87092 15399
rect 87156 5710 87184 17303
rect 87248 8294 87276 25463
rect 87432 22094 87460 43143
rect 87524 36417 87552 47767
rect 87696 47184 87748 47190
rect 87696 47126 87748 47132
rect 87604 46572 87656 46578
rect 87604 46514 87656 46520
rect 87510 36408 87566 36417
rect 87510 36343 87566 36352
rect 87616 26625 87644 46514
rect 87708 37505 87736 47126
rect 87878 40760 87934 40769
rect 87878 40695 87934 40704
rect 87694 37496 87750 37505
rect 87694 37431 87750 37440
rect 87892 26897 87920 40695
rect 88076 40225 88104 47903
rect 88708 47660 88760 47666
rect 88708 47602 88760 47608
rect 88340 47456 88392 47462
rect 88340 47398 88392 47404
rect 88352 45665 88380 47398
rect 88524 47320 88576 47326
rect 88524 47262 88576 47268
rect 88432 47048 88484 47054
rect 88432 46990 88484 46996
rect 88338 45656 88394 45665
rect 88338 45591 88394 45600
rect 88444 45554 88472 46990
rect 88352 45526 88472 45554
rect 88352 44305 88380 45526
rect 88338 44296 88394 44305
rect 88338 44231 88394 44240
rect 88536 42945 88564 47262
rect 88616 47252 88668 47258
rect 88616 47194 88668 47200
rect 88522 42936 88578 42945
rect 88522 42871 88578 42880
rect 88338 41848 88394 41857
rect 88338 41783 88394 41792
rect 88062 40216 88118 40225
rect 88062 40151 88118 40160
rect 87970 29608 88026 29617
rect 87970 29543 88026 29552
rect 87878 26888 87934 26897
rect 87878 26823 87934 26832
rect 87602 26616 87658 26625
rect 87602 26551 87658 26560
rect 87340 22066 87460 22094
rect 87340 12617 87368 22066
rect 87510 20088 87566 20097
rect 87510 20023 87566 20032
rect 87418 13288 87474 13297
rect 87418 13223 87474 13232
rect 87326 12608 87382 12617
rect 87326 12543 87382 12552
rect 87236 8288 87288 8294
rect 87236 8230 87288 8236
rect 87052 5704 87104 5710
rect 87052 5646 87104 5652
rect 87144 5704 87196 5710
rect 87144 5646 87196 5652
rect 86776 5296 86828 5302
rect 86776 5238 86828 5244
rect 87432 5234 87460 13223
rect 87524 5710 87552 20023
rect 87878 18728 87934 18737
rect 87878 18663 87934 18672
rect 87786 11928 87842 11937
rect 87786 11863 87842 11872
rect 87512 5704 87564 5710
rect 87512 5646 87564 5652
rect 87696 5704 87748 5710
rect 87696 5646 87748 5652
rect 87420 5228 87472 5234
rect 87420 5170 87472 5176
rect 87234 4856 87290 4865
rect 85764 4820 85816 4826
rect 87234 4791 87236 4800
rect 85764 4762 85816 4768
rect 87288 4791 87290 4800
rect 87236 4762 87288 4768
rect 87708 4758 87736 5646
rect 87696 4752 87748 4758
rect 87696 4694 87748 4700
rect 87800 4622 87828 11863
rect 87892 5234 87920 18663
rect 87984 11121 88012 29543
rect 88352 12434 88380 41783
rect 88628 38865 88656 47194
rect 88720 41585 88748 47602
rect 88890 47288 88946 47297
rect 88890 47223 88946 47232
rect 88800 47116 88852 47122
rect 88800 47058 88852 47064
rect 88706 41576 88762 41585
rect 88706 41511 88762 41520
rect 88812 41138 88840 47058
rect 88800 41132 88852 41138
rect 88800 41074 88852 41080
rect 88904 41018 88932 47223
rect 88984 46504 89036 46510
rect 88984 46446 89036 46452
rect 88720 40990 88932 41018
rect 88614 38856 88670 38865
rect 88614 38791 88670 38800
rect 88720 36145 88748 40990
rect 88800 40860 88852 40866
rect 88800 40802 88852 40808
rect 88706 36136 88762 36145
rect 88706 36071 88762 36080
rect 88812 34785 88840 40802
rect 88892 40724 88944 40730
rect 88892 40666 88944 40672
rect 88798 34776 88854 34785
rect 88798 34711 88854 34720
rect 88904 32065 88932 40666
rect 88996 33425 89024 46446
rect 88982 33416 89038 33425
rect 88982 33351 89038 33360
rect 88890 32056 88946 32065
rect 88890 31991 88946 32000
rect 89088 27985 89116 48554
rect 89272 48278 89300 69799
rect 89350 67144 89406 67153
rect 89350 67079 89406 67088
rect 89364 50153 89392 67079
rect 89350 50144 89406 50153
rect 89350 50079 89406 50088
rect 89352 48680 89404 48686
rect 89352 48622 89404 48628
rect 89260 48272 89312 48278
rect 89260 48214 89312 48220
rect 89168 47524 89220 47530
rect 89168 47466 89220 47472
rect 89180 40730 89208 47466
rect 89260 46640 89312 46646
rect 89260 46582 89312 46588
rect 89168 40724 89220 40730
rect 89168 40666 89220 40672
rect 89168 40588 89220 40594
rect 89168 40530 89220 40536
rect 89180 30705 89208 40530
rect 89166 30696 89222 30705
rect 89166 30631 89222 30640
rect 89166 29336 89222 29345
rect 89272 29322 89300 46582
rect 89222 29294 89300 29322
rect 89166 29271 89222 29280
rect 89074 27976 89130 27985
rect 89074 27911 89130 27920
rect 89364 26234 89392 48622
rect 89444 47592 89496 47598
rect 89444 47534 89496 47540
rect 89456 40594 89484 47534
rect 89444 40588 89496 40594
rect 89444 40530 89496 40536
rect 89180 26206 89392 26234
rect 89180 25265 89208 26206
rect 89166 25256 89222 25265
rect 89166 25191 89222 25200
rect 89074 22536 89130 22545
rect 89074 22471 89130 22480
rect 89088 22094 89116 22471
rect 89088 22066 89208 22094
rect 88430 21176 88486 21185
rect 88430 21111 88486 21120
rect 88168 12406 88380 12434
rect 87970 11112 88026 11121
rect 87970 11047 88026 11056
rect 87970 10568 88026 10577
rect 87970 10503 88026 10512
rect 87984 5302 88012 10503
rect 88168 9518 88196 12406
rect 88246 9616 88302 9625
rect 88246 9551 88302 9560
rect 88156 9512 88208 9518
rect 88156 9454 88208 9460
rect 88064 8832 88116 8838
rect 88064 8774 88116 8780
rect 88076 5914 88104 8774
rect 88064 5908 88116 5914
rect 88064 5850 88116 5856
rect 88260 5710 88288 9551
rect 88338 8936 88394 8945
rect 88338 8871 88394 8880
rect 88248 5704 88300 5710
rect 88168 5652 88248 5658
rect 88168 5646 88300 5652
rect 88168 5630 88288 5646
rect 87972 5296 88024 5302
rect 87972 5238 88024 5244
rect 87880 5228 87932 5234
rect 87880 5170 87932 5176
rect 88168 4826 88196 5630
rect 88246 5536 88302 5545
rect 88246 5471 88302 5480
rect 88260 5234 88288 5471
rect 88248 5228 88300 5234
rect 88248 5170 88300 5176
rect 88352 5166 88380 8871
rect 88444 5370 88472 21111
rect 89074 17096 89130 17105
rect 89074 17031 89130 17040
rect 88982 15736 89038 15745
rect 88982 15671 89038 15680
rect 88614 14648 88670 14657
rect 88614 14583 88670 14592
rect 88522 5944 88578 5953
rect 88522 5879 88524 5888
rect 88576 5879 88578 5888
rect 88524 5850 88576 5856
rect 88432 5364 88484 5370
rect 88432 5306 88484 5312
rect 88340 5160 88392 5166
rect 88340 5102 88392 5108
rect 88156 4820 88208 4826
rect 88156 4762 88208 4768
rect 87788 4616 87840 4622
rect 86958 4584 87014 4593
rect 87788 4558 87840 4564
rect 86958 4519 86960 4528
rect 87012 4519 87014 4528
rect 86960 4490 87012 4496
rect 88168 4282 88196 4762
rect 88352 4690 88380 5102
rect 88340 4684 88392 4690
rect 88340 4626 88392 4632
rect 88628 4622 88656 14583
rect 88890 13016 88946 13025
rect 88890 12951 88946 12960
rect 88798 11656 88854 11665
rect 88798 11591 88854 11600
rect 88706 10296 88762 10305
rect 88706 10231 88762 10240
rect 88720 5030 88748 10231
rect 88708 5024 88760 5030
rect 88708 4966 88760 4972
rect 88812 4758 88840 11591
rect 88904 5302 88932 12951
rect 88996 5778 89024 15671
rect 88984 5772 89036 5778
rect 88984 5714 89036 5720
rect 89088 5574 89116 17031
rect 89180 8838 89208 22066
rect 89258 19544 89314 19553
rect 89258 19479 89314 19488
rect 89168 8832 89220 8838
rect 89168 8774 89220 8780
rect 89272 5846 89300 19479
rect 89350 18184 89406 18193
rect 89350 18119 89406 18128
rect 89260 5840 89312 5846
rect 89260 5782 89312 5788
rect 89076 5568 89128 5574
rect 89076 5510 89128 5516
rect 88892 5296 88944 5302
rect 88892 5238 88944 5244
rect 89364 5098 89392 18119
rect 89442 14104 89498 14113
rect 89442 14039 89498 14048
rect 89352 5092 89404 5098
rect 89352 5034 89404 5040
rect 89456 4826 89484 14039
rect 89444 4820 89496 4826
rect 89444 4762 89496 4768
rect 88800 4752 88852 4758
rect 88800 4694 88852 4700
rect 88616 4616 88668 4622
rect 88616 4558 88668 4564
rect 88156 4276 88208 4282
rect 88156 4218 88208 4224
rect 79600 2576 79652 2582
rect 79600 2518 79652 2524
rect 80612 2576 80664 2582
rect 80612 2518 80664 2524
rect 81900 2576 81952 2582
rect 81900 2518 81952 2524
rect 82820 2576 82872 2582
rect 82820 2518 82872 2524
rect 78404 2508 78456 2514
rect 78404 2450 78456 2456
rect 15568 2440 15620 2446
rect 15568 2382 15620 2388
rect 16488 2440 16540 2446
rect 16488 2382 16540 2388
rect 17500 2440 17552 2446
rect 17500 2382 17552 2388
rect 18788 2440 18840 2446
rect 18788 2382 18840 2388
rect 19708 2440 19760 2446
rect 19708 2382 19760 2388
rect 20720 2440 20772 2446
rect 20720 2382 20772 2388
rect 22008 2440 22060 2446
rect 22008 2382 22060 2388
rect 23296 2440 23348 2446
rect 23296 2382 23348 2388
rect 24216 2440 24268 2446
rect 24216 2382 24268 2388
rect 25228 2440 25280 2446
rect 25228 2382 25280 2388
rect 26516 2440 26568 2446
rect 26516 2382 26568 2388
rect 27436 2440 27488 2446
rect 27436 2382 27488 2388
rect 28448 2440 28500 2446
rect 28448 2382 28500 2388
rect 29736 2440 29788 2446
rect 29736 2382 29788 2388
rect 55496 2440 55548 2446
rect 55496 2382 55548 2388
rect 56416 2440 56468 2446
rect 56416 2382 56468 2388
rect 57428 2440 57480 2446
rect 57428 2382 57480 2388
rect 58716 2440 58768 2446
rect 58716 2382 58768 2388
rect 59636 2440 59688 2446
rect 59636 2382 59688 2388
rect 60740 2440 60792 2446
rect 60740 2382 60792 2388
rect 61936 2440 61988 2446
rect 61936 2382 61988 2388
rect 63224 2440 63276 2446
rect 63224 2382 63276 2388
rect 64144 2440 64196 2446
rect 64144 2382 64196 2388
rect 65156 2440 65208 2446
rect 65156 2382 65208 2388
rect 66444 2440 66496 2446
rect 66444 2382 66496 2388
rect 67364 2440 67416 2446
rect 67364 2382 67416 2388
rect 68376 2440 68428 2446
rect 68376 2382 68428 2388
rect 69664 2440 69716 2446
rect 69664 2382 69716 2388
rect 10968 2372 11020 2378
rect 10968 2314 11020 2320
rect 39304 2372 39356 2378
rect 39304 2314 39356 2320
rect 79232 2372 79284 2378
rect 79232 2314 79284 2320
rect 7748 2304 7800 2310
rect 7748 2246 7800 2252
rect 8392 2304 8444 2310
rect 8392 2246 8444 2252
rect 7760 800 7788 2246
rect 8404 800 8432 2246
rect 10980 800 11008 2314
rect 12256 2304 12308 2310
rect 12256 2246 12308 2252
rect 13544 2304 13596 2310
rect 13544 2246 13596 2252
rect 15476 2304 15528 2310
rect 15476 2246 15528 2252
rect 16120 2304 16172 2310
rect 16120 2246 16172 2252
rect 17408 2304 17460 2310
rect 17408 2246 17460 2252
rect 18696 2304 18748 2310
rect 18696 2246 18748 2252
rect 19340 2304 19392 2310
rect 19340 2246 19392 2252
rect 20628 2304 20680 2310
rect 20628 2246 20680 2252
rect 21916 2304 21968 2310
rect 21916 2246 21968 2252
rect 23204 2304 23256 2310
rect 23204 2246 23256 2252
rect 23848 2304 23900 2310
rect 23848 2246 23900 2252
rect 25136 2304 25188 2310
rect 25136 2246 25188 2252
rect 26424 2304 26476 2310
rect 26424 2246 26476 2252
rect 27068 2304 27120 2310
rect 27068 2246 27120 2252
rect 28356 2304 28408 2310
rect 28356 2246 28408 2252
rect 29644 2304 29696 2310
rect 29644 2246 29696 2252
rect 30932 2304 30984 2310
rect 30932 2246 30984 2252
rect 31576 2304 31628 2310
rect 31576 2246 31628 2252
rect 32864 2304 32916 2310
rect 32864 2246 32916 2252
rect 34152 2304 34204 2310
rect 34152 2246 34204 2252
rect 34796 2304 34848 2310
rect 34796 2246 34848 2252
rect 36084 2304 36136 2310
rect 36084 2246 36136 2252
rect 37372 2304 37424 2310
rect 37372 2246 37424 2252
rect 38660 2304 38712 2310
rect 38660 2246 38712 2252
rect 12268 800 12296 2246
rect 13556 800 13584 2246
rect 15488 800 15516 2246
rect 16132 800 16160 2246
rect 17420 800 17448 2246
rect 18708 800 18736 2246
rect 19352 800 19380 2246
rect 20640 800 20668 2246
rect 21928 800 21956 2246
rect 23216 800 23244 2246
rect 23860 800 23888 2246
rect 25148 800 25176 2246
rect 26436 800 26464 2246
rect 27080 800 27108 2246
rect 28368 800 28396 2246
rect 29656 800 29684 2246
rect 30944 800 30972 2246
rect 31588 800 31616 2246
rect 32876 800 32904 2246
rect 34164 800 34192 2246
rect 34808 800 34836 2246
rect 36096 800 36124 2246
rect 37384 800 37412 2246
rect 37610 2204 37918 2213
rect 37610 2202 37616 2204
rect 37672 2202 37696 2204
rect 37752 2202 37776 2204
rect 37832 2202 37856 2204
rect 37912 2202 37918 2204
rect 37672 2150 37674 2202
rect 37854 2150 37856 2202
rect 37610 2148 37616 2150
rect 37672 2148 37696 2150
rect 37752 2148 37776 2150
rect 37832 2148 37856 2150
rect 37912 2148 37918 2150
rect 37610 2139 37918 2148
rect 38672 800 38700 2246
rect 39316 800 39344 2314
rect 40592 2304 40644 2310
rect 40592 2246 40644 2252
rect 41880 2304 41932 2310
rect 41880 2246 41932 2252
rect 42524 2304 42576 2310
rect 42524 2246 42576 2252
rect 43812 2304 43864 2310
rect 43812 2246 43864 2252
rect 45100 2304 45152 2310
rect 45100 2246 45152 2252
rect 55404 2304 55456 2310
rect 55404 2246 55456 2252
rect 56048 2304 56100 2310
rect 56048 2246 56100 2252
rect 57336 2304 57388 2310
rect 57336 2246 57388 2252
rect 58624 2304 58676 2310
rect 58624 2246 58676 2252
rect 59912 2304 59964 2310
rect 59912 2246 59964 2252
rect 60556 2304 60608 2310
rect 60556 2246 60608 2252
rect 61844 2304 61896 2310
rect 61844 2246 61896 2252
rect 63132 2304 63184 2310
rect 63132 2246 63184 2252
rect 63776 2304 63828 2310
rect 63776 2246 63828 2252
rect 65064 2304 65116 2310
rect 65064 2246 65116 2252
rect 66352 2304 66404 2310
rect 66352 2246 66404 2252
rect 67640 2304 67692 2310
rect 67640 2246 67692 2252
rect 68284 2304 68336 2310
rect 68284 2246 68336 2252
rect 69572 2304 69624 2310
rect 69572 2246 69624 2252
rect 70860 2304 70912 2310
rect 70860 2246 70912 2252
rect 71504 2304 71556 2310
rect 71504 2246 71556 2252
rect 72792 2304 72844 2310
rect 72792 2246 72844 2252
rect 74080 2304 74132 2310
rect 74080 2246 74132 2252
rect 75368 2304 75420 2310
rect 75368 2246 75420 2252
rect 76012 2304 76064 2310
rect 76012 2246 76064 2252
rect 77300 2304 77352 2310
rect 77300 2246 77352 2252
rect 78588 2304 78640 2310
rect 78588 2246 78640 2252
rect 40604 800 40632 2246
rect 41892 800 41920 2246
rect 42536 800 42564 2246
rect 43824 800 43852 2246
rect 45112 800 45140 2246
rect 55416 800 55444 2246
rect 56060 800 56088 2246
rect 57348 800 57376 2246
rect 58636 800 58664 2246
rect 59924 800 59952 2246
rect 60568 800 60596 2246
rect 61856 800 61884 2246
rect 63144 800 63172 2246
rect 63788 800 63816 2246
rect 65076 800 65104 2246
rect 66364 800 66392 2246
rect 67652 800 67680 2246
rect 68296 800 68324 2246
rect 69584 800 69612 2246
rect 70872 800 70900 2246
rect 71516 800 71544 2246
rect 72804 800 72832 2246
rect 73610 2204 73918 2213
rect 73610 2202 73616 2204
rect 73672 2202 73696 2204
rect 73752 2202 73776 2204
rect 73832 2202 73856 2204
rect 73912 2202 73918 2204
rect 73672 2150 73674 2202
rect 73854 2150 73856 2202
rect 73610 2148 73616 2150
rect 73672 2148 73696 2150
rect 73752 2148 73776 2150
rect 73832 2148 73856 2150
rect 73912 2148 73918 2150
rect 73610 2139 73918 2148
rect 74092 800 74120 2246
rect 75380 800 75408 2246
rect 76024 800 76052 2246
rect 77312 800 77340 2246
rect 78600 800 78628 2246
rect 79244 800 79272 2314
rect 80520 2304 80572 2310
rect 80520 2246 80572 2252
rect 81808 2304 81860 2310
rect 81808 2246 81860 2252
rect 83096 2304 83148 2310
rect 83096 2246 83148 2252
rect 80532 800 80560 2246
rect 81820 800 81848 2246
rect 83108 800 83136 2246
rect 18 0 74 800
rect 662 0 718 800
rect 1306 0 1362 800
rect 1950 0 2006 800
rect 2594 0 2650 800
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 10966 0 11022 800
rect 11610 0 11666 800
rect 12254 0 12310 800
rect 13542 0 13598 800
rect 15474 0 15530 800
rect 16118 0 16174 800
rect 17406 0 17462 800
rect 18694 0 18750 800
rect 19338 0 19394 800
rect 20626 0 20682 800
rect 21914 0 21970 800
rect 23202 0 23258 800
rect 23846 0 23902 800
rect 25134 0 25190 800
rect 26422 0 26478 800
rect 27066 0 27122 800
rect 28354 0 28410 800
rect 29642 0 29698 800
rect 30930 0 30986 800
rect 31574 0 31630 800
rect 32862 0 32918 800
rect 34150 0 34206 800
rect 34794 0 34850 800
rect 36082 0 36138 800
rect 37370 0 37426 800
rect 38658 0 38714 800
rect 39302 0 39358 800
rect 40590 0 40646 800
rect 41878 0 41934 800
rect 42522 0 42578 800
rect 43810 0 43866 800
rect 45098 0 45154 800
rect 55402 0 55458 800
rect 56046 0 56102 800
rect 57334 0 57390 800
rect 58622 0 58678 800
rect 59910 0 59966 800
rect 60554 0 60610 800
rect 61842 0 61898 800
rect 63130 0 63186 800
rect 63774 0 63830 800
rect 65062 0 65118 800
rect 66350 0 66406 800
rect 67638 0 67694 800
rect 68282 0 68338 800
rect 69570 0 69626 800
rect 70858 0 70914 800
rect 71502 0 71558 800
rect 72790 0 72846 800
rect 74078 0 74134 800
rect 75366 0 75422 800
rect 76010 0 76066 800
rect 77298 0 77354 800
rect 78586 0 78642 800
rect 79230 0 79286 800
rect 80518 0 80574 800
rect 81806 0 81862 800
rect 83094 0 83150 800
<< via2 >>
rect 37616 95770 37672 95772
rect 37696 95770 37752 95772
rect 37776 95770 37832 95772
rect 37856 95770 37912 95772
rect 37616 95718 37662 95770
rect 37662 95718 37672 95770
rect 37696 95718 37726 95770
rect 37726 95718 37738 95770
rect 37738 95718 37752 95770
rect 37776 95718 37790 95770
rect 37790 95718 37802 95770
rect 37802 95718 37832 95770
rect 37856 95718 37866 95770
rect 37866 95718 37912 95770
rect 37616 95716 37672 95718
rect 37696 95716 37752 95718
rect 37776 95716 37832 95718
rect 37856 95716 37912 95718
rect 43442 97280 43498 97336
rect 8482 95240 8538 95296
rect 3072 91962 3128 91964
rect 3152 91962 3208 91964
rect 3232 91962 3288 91964
rect 3312 91962 3368 91964
rect 3072 91910 3118 91962
rect 3118 91910 3128 91962
rect 3152 91910 3182 91962
rect 3182 91910 3194 91962
rect 3194 91910 3208 91962
rect 3232 91910 3246 91962
rect 3246 91910 3258 91962
rect 3258 91910 3288 91962
rect 3312 91910 3322 91962
rect 3322 91910 3368 91962
rect 3072 91908 3128 91910
rect 3152 91908 3208 91910
rect 3232 91908 3288 91910
rect 3312 91908 3368 91910
rect 3808 91418 3864 91420
rect 3888 91418 3944 91420
rect 3968 91418 4024 91420
rect 4048 91418 4104 91420
rect 3808 91366 3854 91418
rect 3854 91366 3864 91418
rect 3888 91366 3918 91418
rect 3918 91366 3930 91418
rect 3930 91366 3944 91418
rect 3968 91366 3982 91418
rect 3982 91366 3994 91418
rect 3994 91366 4024 91418
rect 4048 91366 4058 91418
rect 4058 91366 4104 91418
rect 3808 91364 3864 91366
rect 3888 91364 3944 91366
rect 3968 91364 4024 91366
rect 4048 91364 4104 91366
rect 3072 90874 3128 90876
rect 3152 90874 3208 90876
rect 3232 90874 3288 90876
rect 3312 90874 3368 90876
rect 3072 90822 3118 90874
rect 3118 90822 3128 90874
rect 3152 90822 3182 90874
rect 3182 90822 3194 90874
rect 3194 90822 3208 90874
rect 3232 90822 3246 90874
rect 3246 90822 3258 90874
rect 3258 90822 3288 90874
rect 3312 90822 3322 90874
rect 3322 90822 3368 90874
rect 3072 90820 3128 90822
rect 3152 90820 3208 90822
rect 3232 90820 3288 90822
rect 3312 90820 3368 90822
rect 3808 90330 3864 90332
rect 3888 90330 3944 90332
rect 3968 90330 4024 90332
rect 4048 90330 4104 90332
rect 3808 90278 3854 90330
rect 3854 90278 3864 90330
rect 3888 90278 3918 90330
rect 3918 90278 3930 90330
rect 3930 90278 3944 90330
rect 3968 90278 3982 90330
rect 3982 90278 3994 90330
rect 3994 90278 4024 90330
rect 4048 90278 4058 90330
rect 4058 90278 4104 90330
rect 3808 90276 3864 90278
rect 3888 90276 3944 90278
rect 3968 90276 4024 90278
rect 4048 90276 4104 90278
rect 3072 89786 3128 89788
rect 3152 89786 3208 89788
rect 3232 89786 3288 89788
rect 3312 89786 3368 89788
rect 3072 89734 3118 89786
rect 3118 89734 3128 89786
rect 3152 89734 3182 89786
rect 3182 89734 3194 89786
rect 3194 89734 3208 89786
rect 3232 89734 3246 89786
rect 3246 89734 3258 89786
rect 3258 89734 3288 89786
rect 3312 89734 3322 89786
rect 3322 89734 3368 89786
rect 3072 89732 3128 89734
rect 3152 89732 3208 89734
rect 3232 89732 3288 89734
rect 3312 89732 3368 89734
rect 3808 89242 3864 89244
rect 3888 89242 3944 89244
rect 3968 89242 4024 89244
rect 4048 89242 4104 89244
rect 3808 89190 3854 89242
rect 3854 89190 3864 89242
rect 3888 89190 3918 89242
rect 3918 89190 3930 89242
rect 3930 89190 3944 89242
rect 3968 89190 3982 89242
rect 3982 89190 3994 89242
rect 3994 89190 4024 89242
rect 4048 89190 4058 89242
rect 4058 89190 4104 89242
rect 3808 89188 3864 89190
rect 3888 89188 3944 89190
rect 3968 89188 4024 89190
rect 4048 89188 4104 89190
rect 3072 88698 3128 88700
rect 3152 88698 3208 88700
rect 3232 88698 3288 88700
rect 3312 88698 3368 88700
rect 3072 88646 3118 88698
rect 3118 88646 3128 88698
rect 3152 88646 3182 88698
rect 3182 88646 3194 88698
rect 3194 88646 3208 88698
rect 3232 88646 3246 88698
rect 3246 88646 3258 88698
rect 3258 88646 3288 88698
rect 3312 88646 3322 88698
rect 3322 88646 3368 88698
rect 3072 88644 3128 88646
rect 3152 88644 3208 88646
rect 3232 88644 3288 88646
rect 3312 88644 3368 88646
rect 3808 88154 3864 88156
rect 3888 88154 3944 88156
rect 3968 88154 4024 88156
rect 4048 88154 4104 88156
rect 3808 88102 3854 88154
rect 3854 88102 3864 88154
rect 3888 88102 3918 88154
rect 3918 88102 3930 88154
rect 3930 88102 3944 88154
rect 3968 88102 3982 88154
rect 3982 88102 3994 88154
rect 3994 88102 4024 88154
rect 4048 88102 4058 88154
rect 4058 88102 4104 88154
rect 3808 88100 3864 88102
rect 3888 88100 3944 88102
rect 3968 88100 4024 88102
rect 4048 88100 4104 88102
rect 3072 87610 3128 87612
rect 3152 87610 3208 87612
rect 3232 87610 3288 87612
rect 3312 87610 3368 87612
rect 3072 87558 3118 87610
rect 3118 87558 3128 87610
rect 3152 87558 3182 87610
rect 3182 87558 3194 87610
rect 3194 87558 3208 87610
rect 3232 87558 3246 87610
rect 3246 87558 3258 87610
rect 3258 87558 3288 87610
rect 3312 87558 3322 87610
rect 3322 87558 3368 87610
rect 3072 87556 3128 87558
rect 3152 87556 3208 87558
rect 3232 87556 3288 87558
rect 3312 87556 3368 87558
rect 3808 87066 3864 87068
rect 3888 87066 3944 87068
rect 3968 87066 4024 87068
rect 4048 87066 4104 87068
rect 3808 87014 3854 87066
rect 3854 87014 3864 87066
rect 3888 87014 3918 87066
rect 3918 87014 3930 87066
rect 3930 87014 3944 87066
rect 3968 87014 3982 87066
rect 3982 87014 3994 87066
rect 3994 87014 4024 87066
rect 4048 87014 4058 87066
rect 4058 87014 4104 87066
rect 3808 87012 3864 87014
rect 3888 87012 3944 87014
rect 3968 87012 4024 87014
rect 4048 87012 4104 87014
rect 846 86572 848 86592
rect 848 86572 900 86592
rect 900 86572 902 86592
rect 846 86536 902 86572
rect 3072 86522 3128 86524
rect 3152 86522 3208 86524
rect 3232 86522 3288 86524
rect 3312 86522 3368 86524
rect 3072 86470 3118 86522
rect 3118 86470 3128 86522
rect 3152 86470 3182 86522
rect 3182 86470 3194 86522
rect 3194 86470 3208 86522
rect 3232 86470 3246 86522
rect 3246 86470 3258 86522
rect 3258 86470 3288 86522
rect 3312 86470 3322 86522
rect 3322 86470 3368 86522
rect 3072 86468 3128 86470
rect 3152 86468 3208 86470
rect 3232 86468 3288 86470
rect 3312 86468 3368 86470
rect 3808 85978 3864 85980
rect 3888 85978 3944 85980
rect 3968 85978 4024 85980
rect 4048 85978 4104 85980
rect 3808 85926 3854 85978
rect 3854 85926 3864 85978
rect 3888 85926 3918 85978
rect 3918 85926 3930 85978
rect 3930 85926 3944 85978
rect 3968 85926 3982 85978
rect 3982 85926 3994 85978
rect 3994 85926 4024 85978
rect 4048 85926 4058 85978
rect 4058 85926 4104 85978
rect 3808 85924 3864 85926
rect 3888 85924 3944 85926
rect 3968 85924 4024 85926
rect 4048 85924 4104 85926
rect 3072 85434 3128 85436
rect 3152 85434 3208 85436
rect 3232 85434 3288 85436
rect 3312 85434 3368 85436
rect 3072 85382 3118 85434
rect 3118 85382 3128 85434
rect 3152 85382 3182 85434
rect 3182 85382 3194 85434
rect 3194 85382 3208 85434
rect 3232 85382 3246 85434
rect 3246 85382 3258 85434
rect 3258 85382 3288 85434
rect 3312 85382 3322 85434
rect 3322 85382 3368 85434
rect 3072 85380 3128 85382
rect 3152 85380 3208 85382
rect 3232 85380 3288 85382
rect 3312 85380 3368 85382
rect 846 85212 848 85232
rect 848 85212 900 85232
rect 900 85212 902 85232
rect 846 85176 902 85212
rect 3808 84890 3864 84892
rect 3888 84890 3944 84892
rect 3968 84890 4024 84892
rect 4048 84890 4104 84892
rect 3808 84838 3854 84890
rect 3854 84838 3864 84890
rect 3888 84838 3918 84890
rect 3918 84838 3930 84890
rect 3930 84838 3944 84890
rect 3968 84838 3982 84890
rect 3982 84838 3994 84890
rect 3994 84838 4024 84890
rect 4048 84838 4058 84890
rect 4058 84838 4104 84890
rect 3808 84836 3864 84838
rect 3888 84836 3944 84838
rect 3968 84836 4024 84838
rect 4048 84836 4104 84838
rect 3072 84346 3128 84348
rect 3152 84346 3208 84348
rect 3232 84346 3288 84348
rect 3312 84346 3368 84348
rect 3072 84294 3118 84346
rect 3118 84294 3128 84346
rect 3152 84294 3182 84346
rect 3182 84294 3194 84346
rect 3194 84294 3208 84346
rect 3232 84294 3246 84346
rect 3246 84294 3258 84346
rect 3258 84294 3288 84346
rect 3312 84294 3322 84346
rect 3322 84294 3368 84346
rect 3072 84292 3128 84294
rect 3152 84292 3208 84294
rect 3232 84292 3288 84294
rect 3312 84292 3368 84294
rect 846 83852 848 83872
rect 848 83852 900 83872
rect 900 83852 902 83872
rect 846 83816 902 83852
rect 3808 83802 3864 83804
rect 3888 83802 3944 83804
rect 3968 83802 4024 83804
rect 4048 83802 4104 83804
rect 3808 83750 3854 83802
rect 3854 83750 3864 83802
rect 3888 83750 3918 83802
rect 3918 83750 3930 83802
rect 3930 83750 3944 83802
rect 3968 83750 3982 83802
rect 3982 83750 3994 83802
rect 3994 83750 4024 83802
rect 4048 83750 4058 83802
rect 4058 83750 4104 83802
rect 3808 83748 3864 83750
rect 3888 83748 3944 83750
rect 3968 83748 4024 83750
rect 4048 83748 4104 83750
rect 3072 83258 3128 83260
rect 3152 83258 3208 83260
rect 3232 83258 3288 83260
rect 3312 83258 3368 83260
rect 3072 83206 3118 83258
rect 3118 83206 3128 83258
rect 3152 83206 3182 83258
rect 3182 83206 3194 83258
rect 3194 83206 3208 83258
rect 3232 83206 3246 83258
rect 3246 83206 3258 83258
rect 3258 83206 3288 83258
rect 3312 83206 3322 83258
rect 3322 83206 3368 83258
rect 3072 83204 3128 83206
rect 3152 83204 3208 83206
rect 3232 83204 3288 83206
rect 3312 83204 3368 83206
rect 3808 82714 3864 82716
rect 3888 82714 3944 82716
rect 3968 82714 4024 82716
rect 4048 82714 4104 82716
rect 3808 82662 3854 82714
rect 3854 82662 3864 82714
rect 3888 82662 3918 82714
rect 3918 82662 3930 82714
rect 3930 82662 3944 82714
rect 3968 82662 3982 82714
rect 3982 82662 3994 82714
rect 3994 82662 4024 82714
rect 4048 82662 4058 82714
rect 4058 82662 4104 82714
rect 3808 82660 3864 82662
rect 3888 82660 3944 82662
rect 3968 82660 4024 82662
rect 4048 82660 4104 82662
rect 846 82220 848 82240
rect 848 82220 900 82240
rect 900 82220 902 82240
rect 846 82184 902 82220
rect 3072 82170 3128 82172
rect 3152 82170 3208 82172
rect 3232 82170 3288 82172
rect 3312 82170 3368 82172
rect 3072 82118 3118 82170
rect 3118 82118 3128 82170
rect 3152 82118 3182 82170
rect 3182 82118 3194 82170
rect 3194 82118 3208 82170
rect 3232 82118 3246 82170
rect 3246 82118 3258 82170
rect 3258 82118 3288 82170
rect 3312 82118 3322 82170
rect 3322 82118 3368 82170
rect 3072 82116 3128 82118
rect 3152 82116 3208 82118
rect 3232 82116 3288 82118
rect 3312 82116 3368 82118
rect 3808 81626 3864 81628
rect 3888 81626 3944 81628
rect 3968 81626 4024 81628
rect 4048 81626 4104 81628
rect 3808 81574 3854 81626
rect 3854 81574 3864 81626
rect 3888 81574 3918 81626
rect 3918 81574 3930 81626
rect 3930 81574 3944 81626
rect 3968 81574 3982 81626
rect 3982 81574 3994 81626
rect 3994 81574 4024 81626
rect 4048 81574 4058 81626
rect 4058 81574 4104 81626
rect 3808 81572 3864 81574
rect 3888 81572 3944 81574
rect 3968 81572 4024 81574
rect 4048 81572 4104 81574
rect 846 81132 848 81152
rect 848 81132 900 81152
rect 900 81132 902 81152
rect 846 81096 902 81132
rect 3072 81082 3128 81084
rect 3152 81082 3208 81084
rect 3232 81082 3288 81084
rect 3312 81082 3368 81084
rect 3072 81030 3118 81082
rect 3118 81030 3128 81082
rect 3152 81030 3182 81082
rect 3182 81030 3194 81082
rect 3194 81030 3208 81082
rect 3232 81030 3246 81082
rect 3246 81030 3258 81082
rect 3258 81030 3288 81082
rect 3312 81030 3322 81082
rect 3322 81030 3368 81082
rect 3072 81028 3128 81030
rect 3152 81028 3208 81030
rect 3232 81028 3288 81030
rect 3312 81028 3368 81030
rect 3808 80538 3864 80540
rect 3888 80538 3944 80540
rect 3968 80538 4024 80540
rect 4048 80538 4104 80540
rect 3808 80486 3854 80538
rect 3854 80486 3864 80538
rect 3888 80486 3918 80538
rect 3918 80486 3930 80538
rect 3930 80486 3944 80538
rect 3968 80486 3982 80538
rect 3982 80486 3994 80538
rect 3994 80486 4024 80538
rect 4048 80486 4058 80538
rect 4058 80486 4104 80538
rect 3808 80484 3864 80486
rect 3888 80484 3944 80486
rect 3968 80484 4024 80486
rect 4048 80484 4104 80486
rect 3072 79994 3128 79996
rect 3152 79994 3208 79996
rect 3232 79994 3288 79996
rect 3312 79994 3368 79996
rect 3072 79942 3118 79994
rect 3118 79942 3128 79994
rect 3152 79942 3182 79994
rect 3182 79942 3194 79994
rect 3194 79942 3208 79994
rect 3232 79942 3246 79994
rect 3246 79942 3258 79994
rect 3258 79942 3288 79994
rect 3312 79942 3322 79994
rect 3322 79942 3368 79994
rect 3072 79940 3128 79942
rect 3152 79940 3208 79942
rect 3232 79940 3288 79942
rect 3312 79940 3368 79942
rect 846 79500 848 79520
rect 848 79500 900 79520
rect 900 79500 902 79520
rect 846 79464 902 79500
rect 3808 79450 3864 79452
rect 3888 79450 3944 79452
rect 3968 79450 4024 79452
rect 4048 79450 4104 79452
rect 3808 79398 3854 79450
rect 3854 79398 3864 79450
rect 3888 79398 3918 79450
rect 3918 79398 3930 79450
rect 3930 79398 3944 79450
rect 3968 79398 3982 79450
rect 3982 79398 3994 79450
rect 3994 79398 4024 79450
rect 4048 79398 4058 79450
rect 4058 79398 4104 79450
rect 3808 79396 3864 79398
rect 3888 79396 3944 79398
rect 3968 79396 4024 79398
rect 4048 79396 4104 79398
rect 3072 78906 3128 78908
rect 3152 78906 3208 78908
rect 3232 78906 3288 78908
rect 3312 78906 3368 78908
rect 3072 78854 3118 78906
rect 3118 78854 3128 78906
rect 3152 78854 3182 78906
rect 3182 78854 3194 78906
rect 3194 78854 3208 78906
rect 3232 78854 3246 78906
rect 3246 78854 3258 78906
rect 3258 78854 3288 78906
rect 3312 78854 3322 78906
rect 3322 78854 3368 78906
rect 3072 78852 3128 78854
rect 3152 78852 3208 78854
rect 3232 78852 3288 78854
rect 3312 78852 3368 78854
rect 846 78412 848 78432
rect 848 78412 900 78432
rect 900 78412 902 78432
rect 846 78376 902 78412
rect 3808 78362 3864 78364
rect 3888 78362 3944 78364
rect 3968 78362 4024 78364
rect 4048 78362 4104 78364
rect 3808 78310 3854 78362
rect 3854 78310 3864 78362
rect 3888 78310 3918 78362
rect 3918 78310 3930 78362
rect 3930 78310 3944 78362
rect 3968 78310 3982 78362
rect 3982 78310 3994 78362
rect 3994 78310 4024 78362
rect 4048 78310 4058 78362
rect 4058 78310 4104 78362
rect 3808 78308 3864 78310
rect 3888 78308 3944 78310
rect 3968 78308 4024 78310
rect 4048 78308 4104 78310
rect 3072 77818 3128 77820
rect 3152 77818 3208 77820
rect 3232 77818 3288 77820
rect 3312 77818 3368 77820
rect 3072 77766 3118 77818
rect 3118 77766 3128 77818
rect 3152 77766 3182 77818
rect 3182 77766 3194 77818
rect 3194 77766 3208 77818
rect 3232 77766 3246 77818
rect 3246 77766 3258 77818
rect 3258 77766 3288 77818
rect 3312 77766 3322 77818
rect 3322 77766 3368 77818
rect 3072 77764 3128 77766
rect 3152 77764 3208 77766
rect 3232 77764 3288 77766
rect 3312 77764 3368 77766
rect 3808 77274 3864 77276
rect 3888 77274 3944 77276
rect 3968 77274 4024 77276
rect 4048 77274 4104 77276
rect 3808 77222 3854 77274
rect 3854 77222 3864 77274
rect 3888 77222 3918 77274
rect 3918 77222 3930 77274
rect 3930 77222 3944 77274
rect 3968 77222 3982 77274
rect 3982 77222 3994 77274
rect 3994 77222 4024 77274
rect 4048 77222 4058 77274
rect 4058 77222 4104 77274
rect 3808 77220 3864 77222
rect 3888 77220 3944 77222
rect 3968 77220 4024 77222
rect 4048 77220 4104 77222
rect 846 76780 848 76800
rect 848 76780 900 76800
rect 900 76780 902 76800
rect 846 76744 902 76780
rect 3072 76730 3128 76732
rect 3152 76730 3208 76732
rect 3232 76730 3288 76732
rect 3312 76730 3368 76732
rect 3072 76678 3118 76730
rect 3118 76678 3128 76730
rect 3152 76678 3182 76730
rect 3182 76678 3194 76730
rect 3194 76678 3208 76730
rect 3232 76678 3246 76730
rect 3246 76678 3258 76730
rect 3258 76678 3288 76730
rect 3312 76678 3322 76730
rect 3322 76678 3368 76730
rect 3072 76676 3128 76678
rect 3152 76676 3208 76678
rect 3232 76676 3288 76678
rect 3312 76676 3368 76678
rect 3808 76186 3864 76188
rect 3888 76186 3944 76188
rect 3968 76186 4024 76188
rect 4048 76186 4104 76188
rect 3808 76134 3854 76186
rect 3854 76134 3864 76186
rect 3888 76134 3918 76186
rect 3918 76134 3930 76186
rect 3930 76134 3944 76186
rect 3968 76134 3982 76186
rect 3982 76134 3994 76186
rect 3994 76134 4024 76186
rect 4048 76134 4058 76186
rect 4058 76134 4104 76186
rect 3808 76132 3864 76134
rect 3888 76132 3944 76134
rect 3968 76132 4024 76134
rect 4048 76132 4104 76134
rect 846 75656 902 75712
rect 3072 75642 3128 75644
rect 3152 75642 3208 75644
rect 3232 75642 3288 75644
rect 3312 75642 3368 75644
rect 3072 75590 3118 75642
rect 3118 75590 3128 75642
rect 3152 75590 3182 75642
rect 3182 75590 3194 75642
rect 3194 75590 3208 75642
rect 3232 75590 3246 75642
rect 3246 75590 3258 75642
rect 3258 75590 3288 75642
rect 3312 75590 3322 75642
rect 3322 75590 3368 75642
rect 3072 75588 3128 75590
rect 3152 75588 3208 75590
rect 3232 75588 3288 75590
rect 3312 75588 3368 75590
rect 3808 75098 3864 75100
rect 3888 75098 3944 75100
rect 3968 75098 4024 75100
rect 4048 75098 4104 75100
rect 3808 75046 3854 75098
rect 3854 75046 3864 75098
rect 3888 75046 3918 75098
rect 3918 75046 3930 75098
rect 3930 75046 3944 75098
rect 3968 75046 3982 75098
rect 3982 75046 3994 75098
rect 3994 75046 4024 75098
rect 4048 75046 4058 75098
rect 4058 75046 4104 75098
rect 3808 75044 3864 75046
rect 3888 75044 3944 75046
rect 3968 75044 4024 75046
rect 4048 75044 4104 75046
rect 3072 74554 3128 74556
rect 3152 74554 3208 74556
rect 3232 74554 3288 74556
rect 3312 74554 3368 74556
rect 3072 74502 3118 74554
rect 3118 74502 3128 74554
rect 3152 74502 3182 74554
rect 3182 74502 3194 74554
rect 3194 74502 3208 74554
rect 3232 74502 3246 74554
rect 3246 74502 3258 74554
rect 3258 74502 3288 74554
rect 3312 74502 3322 74554
rect 3322 74502 3368 74554
rect 3072 74500 3128 74502
rect 3152 74500 3208 74502
rect 3232 74500 3288 74502
rect 3312 74500 3368 74502
rect 846 74060 848 74080
rect 848 74060 900 74080
rect 900 74060 902 74080
rect 846 74024 902 74060
rect 3808 74010 3864 74012
rect 3888 74010 3944 74012
rect 3968 74010 4024 74012
rect 4048 74010 4104 74012
rect 3808 73958 3854 74010
rect 3854 73958 3864 74010
rect 3888 73958 3918 74010
rect 3918 73958 3930 74010
rect 3930 73958 3944 74010
rect 3968 73958 3982 74010
rect 3982 73958 3994 74010
rect 3994 73958 4024 74010
rect 4048 73958 4058 74010
rect 4058 73958 4104 74010
rect 3808 73956 3864 73958
rect 3888 73956 3944 73958
rect 3968 73956 4024 73958
rect 4048 73956 4104 73958
rect 3072 73466 3128 73468
rect 3152 73466 3208 73468
rect 3232 73466 3288 73468
rect 3312 73466 3368 73468
rect 3072 73414 3118 73466
rect 3118 73414 3128 73466
rect 3152 73414 3182 73466
rect 3182 73414 3194 73466
rect 3194 73414 3208 73466
rect 3232 73414 3246 73466
rect 3246 73414 3258 73466
rect 3258 73414 3288 73466
rect 3312 73414 3322 73466
rect 3322 73414 3368 73466
rect 3072 73412 3128 73414
rect 3152 73412 3208 73414
rect 3232 73412 3288 73414
rect 3312 73412 3368 73414
rect 846 72972 848 72992
rect 848 72972 900 72992
rect 900 72972 902 72992
rect 846 72936 902 72972
rect 3808 72922 3864 72924
rect 3888 72922 3944 72924
rect 3968 72922 4024 72924
rect 4048 72922 4104 72924
rect 3808 72870 3854 72922
rect 3854 72870 3864 72922
rect 3888 72870 3918 72922
rect 3918 72870 3930 72922
rect 3930 72870 3944 72922
rect 3968 72870 3982 72922
rect 3982 72870 3994 72922
rect 3994 72870 4024 72922
rect 4048 72870 4058 72922
rect 4058 72870 4104 72922
rect 3808 72868 3864 72870
rect 3888 72868 3944 72870
rect 3968 72868 4024 72870
rect 4048 72868 4104 72870
rect 3072 72378 3128 72380
rect 3152 72378 3208 72380
rect 3232 72378 3288 72380
rect 3312 72378 3368 72380
rect 3072 72326 3118 72378
rect 3118 72326 3128 72378
rect 3152 72326 3182 72378
rect 3182 72326 3194 72378
rect 3194 72326 3208 72378
rect 3232 72326 3246 72378
rect 3246 72326 3258 72378
rect 3258 72326 3288 72378
rect 3312 72326 3322 72378
rect 3322 72326 3368 72378
rect 3072 72324 3128 72326
rect 3152 72324 3208 72326
rect 3232 72324 3288 72326
rect 3312 72324 3368 72326
rect 3808 71834 3864 71836
rect 3888 71834 3944 71836
rect 3968 71834 4024 71836
rect 4048 71834 4104 71836
rect 3808 71782 3854 71834
rect 3854 71782 3864 71834
rect 3888 71782 3918 71834
rect 3918 71782 3930 71834
rect 3930 71782 3944 71834
rect 3968 71782 3982 71834
rect 3982 71782 3994 71834
rect 3994 71782 4024 71834
rect 4048 71782 4058 71834
rect 4058 71782 4104 71834
rect 3808 71780 3864 71782
rect 3888 71780 3944 71782
rect 3968 71780 4024 71782
rect 4048 71780 4104 71782
rect 846 71340 848 71360
rect 848 71340 900 71360
rect 900 71340 902 71360
rect 846 71304 902 71340
rect 3072 71290 3128 71292
rect 3152 71290 3208 71292
rect 3232 71290 3288 71292
rect 3312 71290 3368 71292
rect 3072 71238 3118 71290
rect 3118 71238 3128 71290
rect 3152 71238 3182 71290
rect 3182 71238 3194 71290
rect 3194 71238 3208 71290
rect 3232 71238 3246 71290
rect 3246 71238 3258 71290
rect 3258 71238 3288 71290
rect 3312 71238 3322 71290
rect 3322 71238 3368 71290
rect 3072 71236 3128 71238
rect 3152 71236 3208 71238
rect 3232 71236 3288 71238
rect 3312 71236 3368 71238
rect 3808 70746 3864 70748
rect 3888 70746 3944 70748
rect 3968 70746 4024 70748
rect 4048 70746 4104 70748
rect 3808 70694 3854 70746
rect 3854 70694 3864 70746
rect 3888 70694 3918 70746
rect 3918 70694 3930 70746
rect 3930 70694 3944 70746
rect 3968 70694 3982 70746
rect 3982 70694 3994 70746
rect 3994 70694 4024 70746
rect 4048 70694 4058 70746
rect 4058 70694 4104 70746
rect 3808 70692 3864 70694
rect 3888 70692 3944 70694
rect 3968 70692 4024 70694
rect 4048 70692 4104 70694
rect 846 70216 902 70272
rect 3072 70202 3128 70204
rect 3152 70202 3208 70204
rect 3232 70202 3288 70204
rect 3312 70202 3368 70204
rect 3072 70150 3118 70202
rect 3118 70150 3128 70202
rect 3152 70150 3182 70202
rect 3182 70150 3194 70202
rect 3194 70150 3208 70202
rect 3232 70150 3246 70202
rect 3246 70150 3258 70202
rect 3258 70150 3288 70202
rect 3312 70150 3322 70202
rect 3322 70150 3368 70202
rect 3072 70148 3128 70150
rect 3152 70148 3208 70150
rect 3232 70148 3288 70150
rect 3312 70148 3368 70150
rect 3808 69658 3864 69660
rect 3888 69658 3944 69660
rect 3968 69658 4024 69660
rect 4048 69658 4104 69660
rect 3808 69606 3854 69658
rect 3854 69606 3864 69658
rect 3888 69606 3918 69658
rect 3918 69606 3930 69658
rect 3930 69606 3944 69658
rect 3968 69606 3982 69658
rect 3982 69606 3994 69658
rect 3994 69606 4024 69658
rect 4048 69606 4058 69658
rect 4058 69606 4104 69658
rect 3808 69604 3864 69606
rect 3888 69604 3944 69606
rect 3968 69604 4024 69606
rect 4048 69604 4104 69606
rect 3072 69114 3128 69116
rect 3152 69114 3208 69116
rect 3232 69114 3288 69116
rect 3312 69114 3368 69116
rect 3072 69062 3118 69114
rect 3118 69062 3128 69114
rect 3152 69062 3182 69114
rect 3182 69062 3194 69114
rect 3194 69062 3208 69114
rect 3232 69062 3246 69114
rect 3246 69062 3258 69114
rect 3258 69062 3288 69114
rect 3312 69062 3322 69114
rect 3322 69062 3368 69114
rect 3072 69060 3128 69062
rect 3152 69060 3208 69062
rect 3232 69060 3288 69062
rect 3312 69060 3368 69062
rect 1214 68756 1216 68776
rect 1216 68756 1268 68776
rect 1268 68756 1270 68776
rect 1214 68720 1270 68756
rect 3808 68570 3864 68572
rect 3888 68570 3944 68572
rect 3968 68570 4024 68572
rect 4048 68570 4104 68572
rect 3808 68518 3854 68570
rect 3854 68518 3864 68570
rect 3888 68518 3918 68570
rect 3918 68518 3930 68570
rect 3930 68518 3944 68570
rect 3968 68518 3982 68570
rect 3982 68518 3994 68570
rect 3994 68518 4024 68570
rect 4048 68518 4058 68570
rect 4058 68518 4104 68570
rect 3808 68516 3864 68518
rect 3888 68516 3944 68518
rect 3968 68516 4024 68518
rect 4048 68516 4104 68518
rect 3072 68026 3128 68028
rect 3152 68026 3208 68028
rect 3232 68026 3288 68028
rect 3312 68026 3368 68028
rect 3072 67974 3118 68026
rect 3118 67974 3128 68026
rect 3152 67974 3182 68026
rect 3182 67974 3194 68026
rect 3194 67974 3208 68026
rect 3232 67974 3246 68026
rect 3246 67974 3258 68026
rect 3258 67974 3288 68026
rect 3312 67974 3322 68026
rect 3322 67974 3368 68026
rect 3072 67972 3128 67974
rect 3152 67972 3208 67974
rect 3232 67972 3288 67974
rect 3312 67972 3368 67974
rect 3808 67482 3864 67484
rect 3888 67482 3944 67484
rect 3968 67482 4024 67484
rect 4048 67482 4104 67484
rect 3808 67430 3854 67482
rect 3854 67430 3864 67482
rect 3888 67430 3918 67482
rect 3918 67430 3930 67482
rect 3930 67430 3944 67482
rect 3968 67430 3982 67482
rect 3982 67430 3994 67482
rect 3994 67430 4024 67482
rect 4048 67430 4058 67482
rect 4058 67430 4104 67482
rect 3808 67428 3864 67430
rect 3888 67428 3944 67430
rect 3968 67428 4024 67430
rect 4048 67428 4104 67430
rect 1306 67360 1362 67416
rect 3072 66938 3128 66940
rect 3152 66938 3208 66940
rect 3232 66938 3288 66940
rect 3312 66938 3368 66940
rect 3072 66886 3118 66938
rect 3118 66886 3128 66938
rect 3152 66886 3182 66938
rect 3182 66886 3194 66938
rect 3194 66886 3208 66938
rect 3232 66886 3246 66938
rect 3246 66886 3258 66938
rect 3258 66886 3288 66938
rect 3312 66886 3322 66938
rect 3322 66886 3368 66938
rect 3072 66884 3128 66886
rect 3152 66884 3208 66886
rect 3232 66884 3288 66886
rect 3312 66884 3368 66886
rect 3808 66394 3864 66396
rect 3888 66394 3944 66396
rect 3968 66394 4024 66396
rect 4048 66394 4104 66396
rect 3808 66342 3854 66394
rect 3854 66342 3864 66394
rect 3888 66342 3918 66394
rect 3918 66342 3930 66394
rect 3930 66342 3944 66394
rect 3968 66342 3982 66394
rect 3982 66342 3994 66394
rect 3994 66342 4024 66394
rect 4048 66342 4058 66394
rect 4058 66342 4104 66394
rect 3808 66340 3864 66342
rect 3888 66340 3944 66342
rect 3968 66340 4024 66342
rect 4048 66340 4104 66342
rect 1306 66000 1362 66056
rect 3072 65850 3128 65852
rect 3152 65850 3208 65852
rect 3232 65850 3288 65852
rect 3312 65850 3368 65852
rect 3072 65798 3118 65850
rect 3118 65798 3128 65850
rect 3152 65798 3182 65850
rect 3182 65798 3194 65850
rect 3194 65798 3208 65850
rect 3232 65798 3246 65850
rect 3246 65798 3258 65850
rect 3258 65798 3288 65850
rect 3312 65798 3322 65850
rect 3322 65798 3368 65850
rect 3072 65796 3128 65798
rect 3152 65796 3208 65798
rect 3232 65796 3288 65798
rect 3312 65796 3368 65798
rect 3808 65306 3864 65308
rect 3888 65306 3944 65308
rect 3968 65306 4024 65308
rect 4048 65306 4104 65308
rect 3808 65254 3854 65306
rect 3854 65254 3864 65306
rect 3888 65254 3918 65306
rect 3918 65254 3930 65306
rect 3930 65254 3944 65306
rect 3968 65254 3982 65306
rect 3982 65254 3994 65306
rect 3994 65254 4024 65306
rect 4048 65254 4058 65306
rect 4058 65254 4104 65306
rect 3808 65252 3864 65254
rect 3888 65252 3944 65254
rect 3968 65252 4024 65254
rect 4048 65252 4104 65254
rect 3072 64762 3128 64764
rect 3152 64762 3208 64764
rect 3232 64762 3288 64764
rect 3312 64762 3368 64764
rect 3072 64710 3118 64762
rect 3118 64710 3128 64762
rect 3152 64710 3182 64762
rect 3182 64710 3194 64762
rect 3194 64710 3208 64762
rect 3232 64710 3246 64762
rect 3246 64710 3258 64762
rect 3258 64710 3288 64762
rect 3312 64710 3322 64762
rect 3322 64710 3368 64762
rect 3072 64708 3128 64710
rect 3152 64708 3208 64710
rect 3232 64708 3288 64710
rect 3312 64708 3368 64710
rect 1306 64640 1362 64696
rect 3808 64218 3864 64220
rect 3888 64218 3944 64220
rect 3968 64218 4024 64220
rect 4048 64218 4104 64220
rect 3808 64166 3854 64218
rect 3854 64166 3864 64218
rect 3888 64166 3918 64218
rect 3918 64166 3930 64218
rect 3930 64166 3944 64218
rect 3968 64166 3982 64218
rect 3982 64166 3994 64218
rect 3994 64166 4024 64218
rect 4048 64166 4058 64218
rect 4058 64166 4104 64218
rect 3808 64164 3864 64166
rect 3888 64164 3944 64166
rect 3968 64164 4024 64166
rect 4048 64164 4104 64166
rect 3072 63674 3128 63676
rect 3152 63674 3208 63676
rect 3232 63674 3288 63676
rect 3312 63674 3368 63676
rect 3072 63622 3118 63674
rect 3118 63622 3128 63674
rect 3152 63622 3182 63674
rect 3182 63622 3194 63674
rect 3194 63622 3208 63674
rect 3232 63622 3246 63674
rect 3246 63622 3258 63674
rect 3258 63622 3288 63674
rect 3312 63622 3322 63674
rect 3322 63622 3368 63674
rect 3072 63620 3128 63622
rect 3152 63620 3208 63622
rect 3232 63620 3288 63622
rect 3312 63620 3368 63622
rect 1214 63316 1216 63336
rect 1216 63316 1268 63336
rect 1268 63316 1270 63336
rect 1214 63280 1270 63316
rect 3808 63130 3864 63132
rect 3888 63130 3944 63132
rect 3968 63130 4024 63132
rect 4048 63130 4104 63132
rect 3808 63078 3854 63130
rect 3854 63078 3864 63130
rect 3888 63078 3918 63130
rect 3918 63078 3930 63130
rect 3930 63078 3944 63130
rect 3968 63078 3982 63130
rect 3982 63078 3994 63130
rect 3994 63078 4024 63130
rect 4048 63078 4058 63130
rect 4058 63078 4104 63130
rect 3808 63076 3864 63078
rect 3888 63076 3944 63078
rect 3968 63076 4024 63078
rect 4048 63076 4104 63078
rect 3072 62586 3128 62588
rect 3152 62586 3208 62588
rect 3232 62586 3288 62588
rect 3312 62586 3368 62588
rect 3072 62534 3118 62586
rect 3118 62534 3128 62586
rect 3152 62534 3182 62586
rect 3182 62534 3194 62586
rect 3194 62534 3208 62586
rect 3232 62534 3246 62586
rect 3246 62534 3258 62586
rect 3258 62534 3288 62586
rect 3312 62534 3322 62586
rect 3322 62534 3368 62586
rect 3072 62532 3128 62534
rect 3152 62532 3208 62534
rect 3232 62532 3288 62534
rect 3312 62532 3368 62534
rect 3808 62042 3864 62044
rect 3888 62042 3944 62044
rect 3968 62042 4024 62044
rect 4048 62042 4104 62044
rect 3808 61990 3854 62042
rect 3854 61990 3864 62042
rect 3888 61990 3918 62042
rect 3918 61990 3930 62042
rect 3930 61990 3944 62042
rect 3968 61990 3982 62042
rect 3982 61990 3994 62042
rect 3994 61990 4024 62042
rect 4048 61990 4058 62042
rect 4058 61990 4104 62042
rect 3808 61988 3864 61990
rect 3888 61988 3944 61990
rect 3968 61988 4024 61990
rect 4048 61988 4104 61990
rect 1306 61920 1362 61976
rect 3072 61498 3128 61500
rect 3152 61498 3208 61500
rect 3232 61498 3288 61500
rect 3312 61498 3368 61500
rect 3072 61446 3118 61498
rect 3118 61446 3128 61498
rect 3152 61446 3182 61498
rect 3182 61446 3194 61498
rect 3194 61446 3208 61498
rect 3232 61446 3246 61498
rect 3246 61446 3258 61498
rect 3258 61446 3288 61498
rect 3312 61446 3322 61498
rect 3322 61446 3368 61498
rect 3072 61444 3128 61446
rect 3152 61444 3208 61446
rect 3232 61444 3288 61446
rect 3312 61444 3368 61446
rect 1306 61240 1362 61296
rect 3808 60954 3864 60956
rect 3888 60954 3944 60956
rect 3968 60954 4024 60956
rect 4048 60954 4104 60956
rect 3808 60902 3854 60954
rect 3854 60902 3864 60954
rect 3888 60902 3918 60954
rect 3918 60902 3930 60954
rect 3930 60902 3944 60954
rect 3968 60902 3982 60954
rect 3982 60902 3994 60954
rect 3994 60902 4024 60954
rect 4048 60902 4058 60954
rect 4058 60902 4104 60954
rect 3808 60900 3864 60902
rect 3888 60900 3944 60902
rect 3968 60900 4024 60902
rect 4048 60900 4104 60902
rect 846 60460 848 60480
rect 848 60460 900 60480
rect 900 60460 902 60480
rect 846 60424 902 60460
rect 3072 60410 3128 60412
rect 3152 60410 3208 60412
rect 3232 60410 3288 60412
rect 3312 60410 3368 60412
rect 3072 60358 3118 60410
rect 3118 60358 3128 60410
rect 3152 60358 3182 60410
rect 3182 60358 3194 60410
rect 3194 60358 3208 60410
rect 3232 60358 3246 60410
rect 3246 60358 3258 60410
rect 3258 60358 3288 60410
rect 3312 60358 3322 60410
rect 3322 60358 3368 60410
rect 3072 60356 3128 60358
rect 3152 60356 3208 60358
rect 3232 60356 3288 60358
rect 3312 60356 3368 60358
rect 1214 59880 1270 59936
rect 3808 59866 3864 59868
rect 3888 59866 3944 59868
rect 3968 59866 4024 59868
rect 4048 59866 4104 59868
rect 3808 59814 3854 59866
rect 3854 59814 3864 59866
rect 3888 59814 3918 59866
rect 3918 59814 3930 59866
rect 3930 59814 3944 59866
rect 3968 59814 3982 59866
rect 3982 59814 3994 59866
rect 3994 59814 4024 59866
rect 4048 59814 4058 59866
rect 4058 59814 4104 59866
rect 3808 59812 3864 59814
rect 3888 59812 3944 59814
rect 3968 59812 4024 59814
rect 4048 59812 4104 59814
rect 3072 59322 3128 59324
rect 3152 59322 3208 59324
rect 3232 59322 3288 59324
rect 3312 59322 3368 59324
rect 3072 59270 3118 59322
rect 3118 59270 3128 59322
rect 3152 59270 3182 59322
rect 3182 59270 3194 59322
rect 3194 59270 3208 59322
rect 3232 59270 3246 59322
rect 3246 59270 3258 59322
rect 3258 59270 3288 59322
rect 3312 59270 3322 59322
rect 3322 59270 3368 59322
rect 3072 59268 3128 59270
rect 3152 59268 3208 59270
rect 3232 59268 3288 59270
rect 3312 59268 3368 59270
rect 846 59064 902 59120
rect 3808 58778 3864 58780
rect 3888 58778 3944 58780
rect 3968 58778 4024 58780
rect 4048 58778 4104 58780
rect 3808 58726 3854 58778
rect 3854 58726 3864 58778
rect 3888 58726 3918 58778
rect 3918 58726 3930 58778
rect 3930 58726 3944 58778
rect 3968 58726 3982 58778
rect 3982 58726 3994 58778
rect 3994 58726 4024 58778
rect 4048 58726 4058 58778
rect 4058 58726 4104 58778
rect 3808 58724 3864 58726
rect 3888 58724 3944 58726
rect 3968 58724 4024 58726
rect 4048 58724 4104 58726
rect 1306 58520 1362 58576
rect 3072 58234 3128 58236
rect 3152 58234 3208 58236
rect 3232 58234 3288 58236
rect 3312 58234 3368 58236
rect 3072 58182 3118 58234
rect 3118 58182 3128 58234
rect 3152 58182 3182 58234
rect 3182 58182 3194 58234
rect 3194 58182 3208 58234
rect 3232 58182 3246 58234
rect 3246 58182 3258 58234
rect 3258 58182 3288 58234
rect 3312 58182 3322 58234
rect 3322 58182 3368 58234
rect 3072 58180 3128 58182
rect 3152 58180 3208 58182
rect 3232 58180 3288 58182
rect 3312 58180 3368 58182
rect 846 57704 902 57760
rect 3808 57690 3864 57692
rect 3888 57690 3944 57692
rect 3968 57690 4024 57692
rect 4048 57690 4104 57692
rect 3808 57638 3854 57690
rect 3854 57638 3864 57690
rect 3888 57638 3918 57690
rect 3918 57638 3930 57690
rect 3930 57638 3944 57690
rect 3968 57638 3982 57690
rect 3982 57638 3994 57690
rect 3994 57638 4024 57690
rect 4048 57638 4058 57690
rect 4058 57638 4104 57690
rect 3808 57636 3864 57638
rect 3888 57636 3944 57638
rect 3968 57636 4024 57638
rect 4048 57636 4104 57638
rect 1306 57160 1362 57216
rect 3072 57146 3128 57148
rect 3152 57146 3208 57148
rect 3232 57146 3288 57148
rect 3312 57146 3368 57148
rect 3072 57094 3118 57146
rect 3118 57094 3128 57146
rect 3152 57094 3182 57146
rect 3182 57094 3194 57146
rect 3194 57094 3208 57146
rect 3232 57094 3246 57146
rect 3246 57094 3258 57146
rect 3258 57094 3288 57146
rect 3312 57094 3322 57146
rect 3322 57094 3368 57146
rect 3072 57092 3128 57094
rect 3152 57092 3208 57094
rect 3232 57092 3288 57094
rect 3312 57092 3368 57094
rect 3808 56602 3864 56604
rect 3888 56602 3944 56604
rect 3968 56602 4024 56604
rect 4048 56602 4104 56604
rect 3808 56550 3854 56602
rect 3854 56550 3864 56602
rect 3888 56550 3918 56602
rect 3918 56550 3930 56602
rect 3930 56550 3944 56602
rect 3968 56550 3982 56602
rect 3982 56550 3994 56602
rect 3994 56550 4024 56602
rect 4048 56550 4058 56602
rect 4058 56550 4104 56602
rect 3808 56548 3864 56550
rect 3888 56548 3944 56550
rect 3968 56548 4024 56550
rect 4048 56548 4104 56550
rect 846 56344 902 56400
rect 3072 56058 3128 56060
rect 3152 56058 3208 56060
rect 3232 56058 3288 56060
rect 3312 56058 3368 56060
rect 3072 56006 3118 56058
rect 3118 56006 3128 56058
rect 3152 56006 3182 56058
rect 3182 56006 3194 56058
rect 3194 56006 3208 56058
rect 3232 56006 3246 56058
rect 3246 56006 3258 56058
rect 3258 56006 3288 56058
rect 3312 56006 3322 56058
rect 3322 56006 3368 56058
rect 3072 56004 3128 56006
rect 3152 56004 3208 56006
rect 3232 56004 3288 56006
rect 3312 56004 3368 56006
rect 1306 55800 1362 55856
rect 3808 55514 3864 55516
rect 3888 55514 3944 55516
rect 3968 55514 4024 55516
rect 4048 55514 4104 55516
rect 3808 55462 3854 55514
rect 3854 55462 3864 55514
rect 3888 55462 3918 55514
rect 3918 55462 3930 55514
rect 3930 55462 3944 55514
rect 3968 55462 3982 55514
rect 3982 55462 3994 55514
rect 3994 55462 4024 55514
rect 4048 55462 4058 55514
rect 4058 55462 4104 55514
rect 3808 55460 3864 55462
rect 3888 55460 3944 55462
rect 3968 55460 4024 55462
rect 4048 55460 4104 55462
rect 846 55020 848 55040
rect 848 55020 900 55040
rect 900 55020 902 55040
rect 846 54984 902 55020
rect 3072 54970 3128 54972
rect 3152 54970 3208 54972
rect 3232 54970 3288 54972
rect 3312 54970 3368 54972
rect 3072 54918 3118 54970
rect 3118 54918 3128 54970
rect 3152 54918 3182 54970
rect 3182 54918 3194 54970
rect 3194 54918 3208 54970
rect 3232 54918 3246 54970
rect 3246 54918 3258 54970
rect 3258 54918 3288 54970
rect 3312 54918 3322 54970
rect 3322 54918 3368 54970
rect 3072 54916 3128 54918
rect 3152 54916 3208 54918
rect 3232 54916 3288 54918
rect 3312 54916 3368 54918
rect 1214 54440 1270 54496
rect 3808 54426 3864 54428
rect 3888 54426 3944 54428
rect 3968 54426 4024 54428
rect 4048 54426 4104 54428
rect 3808 54374 3854 54426
rect 3854 54374 3864 54426
rect 3888 54374 3918 54426
rect 3918 54374 3930 54426
rect 3930 54374 3944 54426
rect 3968 54374 3982 54426
rect 3982 54374 3994 54426
rect 3994 54374 4024 54426
rect 4048 54374 4058 54426
rect 4058 54374 4104 54426
rect 3808 54372 3864 54374
rect 3888 54372 3944 54374
rect 3968 54372 4024 54374
rect 4048 54372 4104 54374
rect 3072 53882 3128 53884
rect 3152 53882 3208 53884
rect 3232 53882 3288 53884
rect 3312 53882 3368 53884
rect 3072 53830 3118 53882
rect 3118 53830 3128 53882
rect 3152 53830 3182 53882
rect 3182 53830 3194 53882
rect 3194 53830 3208 53882
rect 3232 53830 3246 53882
rect 3246 53830 3258 53882
rect 3258 53830 3288 53882
rect 3312 53830 3322 53882
rect 3322 53830 3368 53882
rect 3072 53828 3128 53830
rect 3152 53828 3208 53830
rect 3232 53828 3288 53830
rect 3312 53828 3368 53830
rect 846 53624 902 53680
rect 3808 53338 3864 53340
rect 3888 53338 3944 53340
rect 3968 53338 4024 53340
rect 4048 53338 4104 53340
rect 3808 53286 3854 53338
rect 3854 53286 3864 53338
rect 3888 53286 3918 53338
rect 3918 53286 3930 53338
rect 3930 53286 3944 53338
rect 3968 53286 3982 53338
rect 3982 53286 3994 53338
rect 3994 53286 4024 53338
rect 4048 53286 4058 53338
rect 4058 53286 4104 53338
rect 3808 53284 3864 53286
rect 3888 53284 3944 53286
rect 3968 53284 4024 53286
rect 4048 53284 4104 53286
rect 1306 53080 1362 53136
rect 3072 52794 3128 52796
rect 3152 52794 3208 52796
rect 3232 52794 3288 52796
rect 3312 52794 3368 52796
rect 3072 52742 3118 52794
rect 3118 52742 3128 52794
rect 3152 52742 3182 52794
rect 3182 52742 3194 52794
rect 3194 52742 3208 52794
rect 3232 52742 3246 52794
rect 3246 52742 3258 52794
rect 3258 52742 3288 52794
rect 3312 52742 3322 52794
rect 3322 52742 3368 52794
rect 3072 52740 3128 52742
rect 3152 52740 3208 52742
rect 3232 52740 3288 52742
rect 3312 52740 3368 52742
rect 846 52264 902 52320
rect 3808 52250 3864 52252
rect 3888 52250 3944 52252
rect 3968 52250 4024 52252
rect 4048 52250 4104 52252
rect 3808 52198 3854 52250
rect 3854 52198 3864 52250
rect 3888 52198 3918 52250
rect 3918 52198 3930 52250
rect 3930 52198 3944 52250
rect 3968 52198 3982 52250
rect 3982 52198 3994 52250
rect 3994 52198 4024 52250
rect 4048 52198 4058 52250
rect 4058 52198 4104 52250
rect 3808 52196 3864 52198
rect 3888 52196 3944 52198
rect 3968 52196 4024 52198
rect 4048 52196 4104 52198
rect 846 51892 848 51912
rect 848 51892 900 51912
rect 900 51892 902 51912
rect 846 51856 902 51892
rect 3072 51706 3128 51708
rect 3152 51706 3208 51708
rect 3232 51706 3288 51708
rect 3312 51706 3368 51708
rect 3072 51654 3118 51706
rect 3118 51654 3128 51706
rect 3152 51654 3182 51706
rect 3182 51654 3194 51706
rect 3194 51654 3208 51706
rect 3232 51654 3246 51706
rect 3246 51654 3258 51706
rect 3258 51654 3288 51706
rect 3312 51654 3322 51706
rect 3322 51654 3368 51706
rect 3072 51652 3128 51654
rect 3152 51652 3208 51654
rect 3232 51652 3288 51654
rect 3312 51652 3368 51654
rect 1582 51312 1638 51368
rect 1030 51040 1086 51096
rect 1398 50496 1454 50552
rect 1398 49408 1454 49464
rect 1398 49308 1400 49328
rect 1400 49308 1452 49328
rect 1452 49308 1454 49328
rect 1398 49272 1454 49308
rect 3808 51162 3864 51164
rect 3888 51162 3944 51164
rect 3968 51162 4024 51164
rect 4048 51162 4104 51164
rect 3808 51110 3854 51162
rect 3854 51110 3864 51162
rect 3888 51110 3918 51162
rect 3918 51110 3930 51162
rect 3930 51110 3944 51162
rect 3968 51110 3982 51162
rect 3982 51110 3994 51162
rect 3994 51110 4024 51162
rect 4048 51110 4058 51162
rect 4058 51110 4104 51162
rect 3808 51108 3864 51110
rect 3888 51108 3944 51110
rect 3968 51108 4024 51110
rect 4048 51108 4104 51110
rect 3072 50618 3128 50620
rect 3152 50618 3208 50620
rect 3232 50618 3288 50620
rect 3312 50618 3368 50620
rect 3072 50566 3118 50618
rect 3118 50566 3128 50618
rect 3152 50566 3182 50618
rect 3182 50566 3194 50618
rect 3194 50566 3208 50618
rect 3232 50566 3246 50618
rect 3246 50566 3258 50618
rect 3258 50566 3288 50618
rect 3312 50566 3322 50618
rect 3322 50566 3368 50618
rect 3072 50564 3128 50566
rect 3152 50564 3208 50566
rect 3232 50564 3288 50566
rect 3312 50564 3368 50566
rect 3808 50074 3864 50076
rect 3888 50074 3944 50076
rect 3968 50074 4024 50076
rect 4048 50074 4104 50076
rect 3808 50022 3854 50074
rect 3854 50022 3864 50074
rect 3888 50022 3918 50074
rect 3918 50022 3930 50074
rect 3930 50022 3944 50074
rect 3968 50022 3982 50074
rect 3982 50022 3994 50074
rect 3994 50022 4024 50074
rect 4048 50022 4058 50074
rect 4058 50022 4104 50074
rect 3808 50020 3864 50022
rect 3888 50020 3944 50022
rect 3968 50020 4024 50022
rect 4048 50020 4104 50022
rect 3072 49530 3128 49532
rect 3152 49530 3208 49532
rect 3232 49530 3288 49532
rect 3312 49530 3368 49532
rect 3072 49478 3118 49530
rect 3118 49478 3128 49530
rect 3152 49478 3182 49530
rect 3182 49478 3194 49530
rect 3194 49478 3208 49530
rect 3232 49478 3246 49530
rect 3246 49478 3258 49530
rect 3258 49478 3288 49530
rect 3312 49478 3322 49530
rect 3322 49478 3368 49530
rect 3072 49476 3128 49478
rect 3152 49476 3208 49478
rect 3232 49476 3288 49478
rect 3312 49476 3368 49478
rect 5538 75656 5594 75712
rect 5538 70216 5594 70272
rect 5538 67632 5594 67688
rect 5538 64932 5594 64968
rect 5538 64912 5540 64932
rect 5540 64912 5592 64932
rect 5592 64912 5594 64932
rect 5538 62056 5594 62112
rect 4526 49272 4582 49328
rect 4802 50224 4858 50280
rect 4986 49544 5042 49600
rect 4710 49136 4766 49192
rect 5078 49000 5134 49056
rect 3808 48986 3864 48988
rect 3888 48986 3944 48988
rect 3968 48986 4024 48988
rect 4048 48986 4104 48988
rect 3808 48934 3854 48986
rect 3854 48934 3864 48986
rect 3888 48934 3918 48986
rect 3918 48934 3930 48986
rect 3930 48934 3944 48986
rect 3968 48934 3982 48986
rect 3982 48934 3994 48986
rect 3994 48934 4024 48986
rect 4048 48934 4058 48986
rect 4058 48934 4104 48986
rect 3808 48932 3864 48934
rect 3888 48932 3944 48934
rect 3968 48932 4024 48934
rect 4048 48932 4104 48934
rect 36956 95226 37012 95228
rect 37036 95226 37092 95228
rect 37116 95226 37172 95228
rect 37196 95226 37252 95228
rect 36956 95174 37002 95226
rect 37002 95174 37012 95226
rect 37036 95174 37066 95226
rect 37066 95174 37078 95226
rect 37078 95174 37092 95226
rect 37116 95174 37130 95226
rect 37130 95174 37142 95226
rect 37142 95174 37172 95226
rect 37196 95174 37206 95226
rect 37206 95174 37252 95226
rect 36956 95172 37012 95174
rect 37036 95172 37092 95174
rect 37116 95172 37172 95174
rect 37196 95172 37252 95174
rect 37616 94682 37672 94684
rect 37696 94682 37752 94684
rect 37776 94682 37832 94684
rect 37856 94682 37912 94684
rect 37616 94630 37662 94682
rect 37662 94630 37672 94682
rect 37696 94630 37726 94682
rect 37726 94630 37738 94682
rect 37738 94630 37752 94682
rect 37776 94630 37790 94682
rect 37790 94630 37802 94682
rect 37802 94630 37832 94682
rect 37856 94630 37866 94682
rect 37866 94630 37912 94682
rect 37616 94628 37672 94630
rect 37696 94628 37752 94630
rect 37776 94628 37832 94630
rect 37856 94628 37912 94630
rect 36956 94138 37012 94140
rect 37036 94138 37092 94140
rect 37116 94138 37172 94140
rect 37196 94138 37252 94140
rect 36956 94086 37002 94138
rect 37002 94086 37012 94138
rect 37036 94086 37066 94138
rect 37066 94086 37078 94138
rect 37078 94086 37092 94138
rect 37116 94086 37130 94138
rect 37130 94086 37142 94138
rect 37142 94086 37172 94138
rect 37196 94086 37206 94138
rect 37206 94086 37252 94138
rect 36956 94084 37012 94086
rect 37036 94084 37092 94086
rect 37116 94084 37172 94086
rect 37196 94084 37252 94086
rect 37616 93594 37672 93596
rect 37696 93594 37752 93596
rect 37776 93594 37832 93596
rect 37856 93594 37912 93596
rect 37616 93542 37662 93594
rect 37662 93542 37672 93594
rect 37696 93542 37726 93594
rect 37726 93542 37738 93594
rect 37738 93542 37752 93594
rect 37776 93542 37790 93594
rect 37790 93542 37802 93594
rect 37802 93542 37832 93594
rect 37856 93542 37866 93594
rect 37866 93542 37912 93594
rect 37616 93540 37672 93542
rect 37696 93540 37752 93542
rect 37776 93540 37832 93542
rect 37856 93540 37912 93542
rect 36956 93050 37012 93052
rect 37036 93050 37092 93052
rect 37116 93050 37172 93052
rect 37196 93050 37252 93052
rect 36956 92998 37002 93050
rect 37002 92998 37012 93050
rect 37036 92998 37066 93050
rect 37066 92998 37078 93050
rect 37078 92998 37092 93050
rect 37116 92998 37130 93050
rect 37130 92998 37142 93050
rect 37142 92998 37172 93050
rect 37196 92998 37206 93050
rect 37206 92998 37252 93050
rect 36956 92996 37012 92998
rect 37036 92996 37092 92998
rect 37116 92996 37172 92998
rect 37196 92996 37252 92998
rect 37616 92506 37672 92508
rect 37696 92506 37752 92508
rect 37776 92506 37832 92508
rect 37856 92506 37912 92508
rect 37616 92454 37662 92506
rect 37662 92454 37672 92506
rect 37696 92454 37726 92506
rect 37726 92454 37738 92506
rect 37738 92454 37752 92506
rect 37776 92454 37790 92506
rect 37790 92454 37802 92506
rect 37802 92454 37832 92506
rect 37856 92454 37866 92506
rect 37866 92454 37912 92506
rect 37616 92452 37672 92454
rect 37696 92452 37752 92454
rect 37776 92452 37832 92454
rect 37856 92452 37912 92454
rect 36956 91962 37012 91964
rect 37036 91962 37092 91964
rect 37116 91962 37172 91964
rect 37196 91962 37252 91964
rect 36956 91910 37002 91962
rect 37002 91910 37012 91962
rect 37036 91910 37066 91962
rect 37066 91910 37078 91962
rect 37078 91910 37092 91962
rect 37116 91910 37130 91962
rect 37130 91910 37142 91962
rect 37142 91910 37172 91962
rect 37196 91910 37206 91962
rect 37206 91910 37252 91962
rect 36956 91908 37012 91910
rect 37036 91908 37092 91910
rect 37116 91908 37172 91910
rect 37196 91908 37252 91910
rect 37616 91418 37672 91420
rect 37696 91418 37752 91420
rect 37776 91418 37832 91420
rect 37856 91418 37912 91420
rect 37616 91366 37662 91418
rect 37662 91366 37672 91418
rect 37696 91366 37726 91418
rect 37726 91366 37738 91418
rect 37738 91366 37752 91418
rect 37776 91366 37790 91418
rect 37790 91366 37802 91418
rect 37802 91366 37832 91418
rect 37856 91366 37866 91418
rect 37866 91366 37912 91418
rect 37616 91364 37672 91366
rect 37696 91364 37752 91366
rect 37776 91364 37832 91366
rect 37856 91364 37912 91366
rect 49330 97280 49386 97336
rect 73616 95770 73672 95772
rect 73696 95770 73752 95772
rect 73776 95770 73832 95772
rect 73856 95770 73912 95772
rect 73616 95718 73662 95770
rect 73662 95718 73672 95770
rect 73696 95718 73726 95770
rect 73726 95718 73738 95770
rect 73738 95718 73752 95770
rect 73776 95718 73790 95770
rect 73790 95718 73802 95770
rect 73802 95718 73832 95770
rect 73856 95718 73866 95770
rect 73866 95718 73912 95770
rect 73616 95716 73672 95718
rect 73696 95716 73752 95718
rect 73776 95716 73832 95718
rect 73856 95716 73912 95718
rect 46846 92112 46902 92168
rect 46754 91568 46810 91624
rect 5722 67496 5778 67552
rect 5446 50496 5502 50552
rect 3072 48442 3128 48444
rect 3152 48442 3208 48444
rect 3232 48442 3288 48444
rect 3312 48442 3368 48444
rect 3072 48390 3118 48442
rect 3118 48390 3128 48442
rect 3152 48390 3182 48442
rect 3182 48390 3194 48442
rect 3194 48390 3208 48442
rect 3232 48390 3246 48442
rect 3246 48390 3258 48442
rect 3258 48390 3288 48442
rect 3312 48390 3322 48442
rect 3322 48390 3368 48442
rect 3072 48388 3128 48390
rect 3152 48388 3208 48390
rect 3232 48388 3288 48390
rect 3312 48388 3368 48390
rect 1306 48320 1362 48376
rect 4710 48320 4766 48376
rect 1398 47912 1454 47968
rect 3808 47898 3864 47900
rect 3888 47898 3944 47900
rect 3968 47898 4024 47900
rect 4048 47898 4104 47900
rect 3808 47846 3854 47898
rect 3854 47846 3864 47898
rect 3888 47846 3918 47898
rect 3918 47846 3930 47898
rect 3930 47846 3944 47898
rect 3968 47846 3982 47898
rect 3982 47846 3994 47898
rect 3994 47846 4024 47898
rect 4048 47846 4058 47898
rect 4058 47846 4104 47898
rect 3808 47844 3864 47846
rect 3888 47844 3944 47846
rect 3968 47844 4024 47846
rect 4048 47844 4104 47846
rect 4618 47776 4674 47832
rect 3072 47354 3128 47356
rect 3152 47354 3208 47356
rect 3232 47354 3288 47356
rect 3312 47354 3368 47356
rect 3072 47302 3118 47354
rect 3118 47302 3128 47354
rect 3152 47302 3182 47354
rect 3182 47302 3194 47354
rect 3194 47302 3208 47354
rect 3232 47302 3246 47354
rect 3246 47302 3258 47354
rect 3258 47302 3288 47354
rect 3312 47302 3322 47354
rect 3322 47302 3368 47354
rect 3072 47300 3128 47302
rect 3152 47300 3208 47302
rect 3232 47300 3288 47302
rect 3312 47300 3368 47302
rect 1398 46996 1400 47016
rect 1400 46996 1452 47016
rect 1452 46996 1454 47016
rect 1398 46960 1454 46996
rect 3808 46810 3864 46812
rect 3888 46810 3944 46812
rect 3968 46810 4024 46812
rect 4048 46810 4104 46812
rect 3808 46758 3854 46810
rect 3854 46758 3864 46810
rect 3888 46758 3918 46810
rect 3918 46758 3930 46810
rect 3930 46758 3944 46810
rect 3968 46758 3982 46810
rect 3982 46758 3994 46810
rect 3994 46758 4024 46810
rect 4048 46758 4058 46810
rect 4058 46758 4104 46810
rect 3808 46756 3864 46758
rect 3888 46756 3944 46758
rect 3968 46756 4024 46758
rect 4048 46756 4104 46758
rect 1398 46316 1400 46336
rect 1400 46316 1452 46336
rect 1452 46316 1454 46336
rect 1398 46280 1454 46316
rect 3072 46266 3128 46268
rect 3152 46266 3208 46268
rect 3232 46266 3288 46268
rect 3312 46266 3368 46268
rect 3072 46214 3118 46266
rect 3118 46214 3128 46266
rect 3152 46214 3182 46266
rect 3182 46214 3194 46266
rect 3194 46214 3208 46266
rect 3232 46214 3246 46266
rect 3246 46214 3258 46266
rect 3258 46214 3288 46266
rect 3312 46214 3322 46266
rect 3322 46214 3368 46266
rect 3072 46212 3128 46214
rect 3152 46212 3208 46214
rect 3232 46212 3288 46214
rect 3312 46212 3368 46214
rect 1490 45772 1492 45792
rect 1492 45772 1544 45792
rect 1544 45772 1546 45792
rect 1490 45736 1546 45772
rect 3808 45722 3864 45724
rect 3888 45722 3944 45724
rect 3968 45722 4024 45724
rect 4048 45722 4104 45724
rect 3808 45670 3854 45722
rect 3854 45670 3864 45722
rect 3888 45670 3918 45722
rect 3918 45670 3930 45722
rect 3930 45670 3944 45722
rect 3968 45670 3982 45722
rect 3982 45670 3994 45722
rect 3994 45670 4024 45722
rect 4048 45670 4058 45722
rect 4058 45670 4104 45722
rect 3808 45668 3864 45670
rect 3888 45668 3944 45670
rect 3968 45668 4024 45670
rect 4048 45668 4104 45670
rect 3072 45178 3128 45180
rect 3152 45178 3208 45180
rect 3232 45178 3288 45180
rect 3312 45178 3368 45180
rect 3072 45126 3118 45178
rect 3118 45126 3128 45178
rect 3152 45126 3182 45178
rect 3182 45126 3194 45178
rect 3194 45126 3208 45178
rect 3232 45126 3246 45178
rect 3246 45126 3258 45178
rect 3258 45126 3288 45178
rect 3312 45126 3322 45178
rect 3322 45126 3368 45178
rect 3072 45124 3128 45126
rect 3152 45124 3208 45126
rect 3232 45124 3288 45126
rect 3312 45124 3368 45126
rect 1398 45056 1454 45112
rect 3808 44634 3864 44636
rect 3888 44634 3944 44636
rect 3968 44634 4024 44636
rect 4048 44634 4104 44636
rect 3808 44582 3854 44634
rect 3854 44582 3864 44634
rect 3888 44582 3918 44634
rect 3918 44582 3930 44634
rect 3930 44582 3944 44634
rect 3968 44582 3982 44634
rect 3982 44582 3994 44634
rect 3994 44582 4024 44634
rect 4048 44582 4058 44634
rect 4058 44582 4104 44634
rect 3808 44580 3864 44582
rect 3888 44580 3944 44582
rect 3968 44580 4024 44582
rect 4048 44580 4104 44582
rect 1490 44260 1546 44296
rect 1490 44240 1492 44260
rect 1492 44240 1544 44260
rect 1544 44240 1546 44260
rect 3072 44090 3128 44092
rect 3152 44090 3208 44092
rect 3232 44090 3288 44092
rect 3312 44090 3368 44092
rect 3072 44038 3118 44090
rect 3118 44038 3128 44090
rect 3152 44038 3182 44090
rect 3182 44038 3194 44090
rect 3194 44038 3208 44090
rect 3232 44038 3246 44090
rect 3246 44038 3258 44090
rect 3258 44038 3288 44090
rect 3312 44038 3322 44090
rect 3322 44038 3368 44090
rect 3072 44036 3128 44038
rect 3152 44036 3208 44038
rect 3232 44036 3288 44038
rect 3312 44036 3368 44038
rect 1214 43560 1270 43616
rect 3808 43546 3864 43548
rect 3888 43546 3944 43548
rect 3968 43546 4024 43548
rect 4048 43546 4104 43548
rect 3808 43494 3854 43546
rect 3854 43494 3864 43546
rect 3888 43494 3918 43546
rect 3918 43494 3930 43546
rect 3930 43494 3944 43546
rect 3968 43494 3982 43546
rect 3982 43494 3994 43546
rect 3994 43494 4024 43546
rect 4048 43494 4058 43546
rect 4058 43494 4104 43546
rect 3808 43492 3864 43494
rect 3888 43492 3944 43494
rect 3968 43492 4024 43494
rect 4048 43492 4104 43494
rect 1490 43052 1492 43072
rect 1492 43052 1544 43072
rect 1544 43052 1546 43072
rect 1490 43016 1546 43052
rect 3072 43002 3128 43004
rect 3152 43002 3208 43004
rect 3232 43002 3288 43004
rect 3312 43002 3368 43004
rect 3072 42950 3118 43002
rect 3118 42950 3128 43002
rect 3152 42950 3182 43002
rect 3182 42950 3194 43002
rect 3194 42950 3208 43002
rect 3232 42950 3246 43002
rect 3246 42950 3258 43002
rect 3258 42950 3288 43002
rect 3312 42950 3322 43002
rect 3322 42950 3368 43002
rect 3072 42948 3128 42950
rect 3152 42948 3208 42950
rect 3232 42948 3288 42950
rect 3312 42948 3368 42950
rect 3808 42458 3864 42460
rect 3888 42458 3944 42460
rect 3968 42458 4024 42460
rect 4048 42458 4104 42460
rect 3808 42406 3854 42458
rect 3854 42406 3864 42458
rect 3888 42406 3918 42458
rect 3918 42406 3930 42458
rect 3930 42406 3944 42458
rect 3968 42406 3982 42458
rect 3982 42406 3994 42458
rect 3994 42406 4024 42458
rect 4048 42406 4058 42458
rect 4058 42406 4104 42458
rect 3808 42404 3864 42406
rect 3888 42404 3944 42406
rect 3968 42404 4024 42406
rect 4048 42404 4104 42406
rect 3072 41914 3128 41916
rect 3152 41914 3208 41916
rect 3232 41914 3288 41916
rect 3312 41914 3368 41916
rect 3072 41862 3118 41914
rect 3118 41862 3128 41914
rect 3152 41862 3182 41914
rect 3182 41862 3194 41914
rect 3194 41862 3208 41914
rect 3232 41862 3246 41914
rect 3246 41862 3258 41914
rect 3258 41862 3288 41914
rect 3312 41862 3322 41914
rect 3322 41862 3368 41914
rect 3072 41860 3128 41862
rect 3152 41860 3208 41862
rect 3232 41860 3288 41862
rect 3312 41860 3368 41862
rect 1490 41520 1546 41576
rect 3808 41370 3864 41372
rect 3888 41370 3944 41372
rect 3968 41370 4024 41372
rect 4048 41370 4104 41372
rect 3808 41318 3854 41370
rect 3854 41318 3864 41370
rect 3888 41318 3918 41370
rect 3918 41318 3930 41370
rect 3930 41318 3944 41370
rect 3968 41318 3982 41370
rect 3982 41318 3994 41370
rect 3994 41318 4024 41370
rect 4048 41318 4058 41370
rect 4058 41318 4104 41370
rect 3808 41316 3864 41318
rect 3888 41316 3944 41318
rect 3968 41316 4024 41318
rect 4048 41316 4104 41318
rect 3072 40826 3128 40828
rect 3152 40826 3208 40828
rect 3232 40826 3288 40828
rect 3312 40826 3368 40828
rect 3072 40774 3118 40826
rect 3118 40774 3128 40826
rect 3152 40774 3182 40826
rect 3182 40774 3194 40826
rect 3194 40774 3208 40826
rect 3232 40774 3246 40826
rect 3246 40774 3258 40826
rect 3258 40774 3288 40826
rect 3312 40774 3322 40826
rect 3322 40774 3368 40826
rect 3072 40772 3128 40774
rect 3152 40772 3208 40774
rect 3232 40772 3288 40774
rect 3312 40772 3368 40774
rect 846 40332 848 40352
rect 848 40332 900 40352
rect 900 40332 902 40352
rect 846 40296 902 40332
rect 3808 40282 3864 40284
rect 3888 40282 3944 40284
rect 3968 40282 4024 40284
rect 4048 40282 4104 40284
rect 3808 40230 3854 40282
rect 3854 40230 3864 40282
rect 3888 40230 3918 40282
rect 3918 40230 3930 40282
rect 3930 40230 3944 40282
rect 3968 40230 3982 40282
rect 3982 40230 3994 40282
rect 3994 40230 4024 40282
rect 4048 40230 4058 40282
rect 4058 40230 4104 40282
rect 3808 40228 3864 40230
rect 3888 40228 3944 40230
rect 3968 40228 4024 40230
rect 4048 40228 4104 40230
rect 3072 39738 3128 39740
rect 3152 39738 3208 39740
rect 3232 39738 3288 39740
rect 3312 39738 3368 39740
rect 3072 39686 3118 39738
rect 3118 39686 3128 39738
rect 3152 39686 3182 39738
rect 3182 39686 3194 39738
rect 3194 39686 3208 39738
rect 3232 39686 3246 39738
rect 3246 39686 3258 39738
rect 3258 39686 3288 39738
rect 3312 39686 3322 39738
rect 3322 39686 3368 39738
rect 3072 39684 3128 39686
rect 3152 39684 3208 39686
rect 3232 39684 3288 39686
rect 3312 39684 3368 39686
rect 3808 39194 3864 39196
rect 3888 39194 3944 39196
rect 3968 39194 4024 39196
rect 4048 39194 4104 39196
rect 3808 39142 3854 39194
rect 3854 39142 3864 39194
rect 3888 39142 3918 39194
rect 3918 39142 3930 39194
rect 3930 39142 3944 39194
rect 3968 39142 3982 39194
rect 3982 39142 3994 39194
rect 3994 39142 4024 39194
rect 4048 39142 4058 39194
rect 4058 39142 4104 39194
rect 3808 39140 3864 39142
rect 3888 39140 3944 39142
rect 3968 39140 4024 39142
rect 4048 39140 4104 39142
rect 846 38700 848 38720
rect 848 38700 900 38720
rect 900 38700 902 38720
rect 846 38664 902 38700
rect 3072 38650 3128 38652
rect 3152 38650 3208 38652
rect 3232 38650 3288 38652
rect 3312 38650 3368 38652
rect 3072 38598 3118 38650
rect 3118 38598 3128 38650
rect 3152 38598 3182 38650
rect 3182 38598 3194 38650
rect 3194 38598 3208 38650
rect 3232 38598 3246 38650
rect 3246 38598 3258 38650
rect 3258 38598 3288 38650
rect 3312 38598 3322 38650
rect 3322 38598 3368 38650
rect 3072 38596 3128 38598
rect 3152 38596 3208 38598
rect 3232 38596 3288 38598
rect 3312 38596 3368 38598
rect 3808 38106 3864 38108
rect 3888 38106 3944 38108
rect 3968 38106 4024 38108
rect 4048 38106 4104 38108
rect 3808 38054 3854 38106
rect 3854 38054 3864 38106
rect 3888 38054 3918 38106
rect 3918 38054 3930 38106
rect 3930 38054 3944 38106
rect 3968 38054 3982 38106
rect 3982 38054 3994 38106
rect 3994 38054 4024 38106
rect 4048 38054 4058 38106
rect 4058 38054 4104 38106
rect 3808 38052 3864 38054
rect 3888 38052 3944 38054
rect 3968 38052 4024 38054
rect 4048 38052 4104 38054
rect 846 37612 848 37632
rect 848 37612 900 37632
rect 900 37612 902 37632
rect 846 37576 902 37612
rect 3072 37562 3128 37564
rect 3152 37562 3208 37564
rect 3232 37562 3288 37564
rect 3312 37562 3368 37564
rect 3072 37510 3118 37562
rect 3118 37510 3128 37562
rect 3152 37510 3182 37562
rect 3182 37510 3194 37562
rect 3194 37510 3208 37562
rect 3232 37510 3246 37562
rect 3246 37510 3258 37562
rect 3258 37510 3288 37562
rect 3312 37510 3322 37562
rect 3322 37510 3368 37562
rect 3072 37508 3128 37510
rect 3152 37508 3208 37510
rect 3232 37508 3288 37510
rect 3312 37508 3368 37510
rect 3808 37018 3864 37020
rect 3888 37018 3944 37020
rect 3968 37018 4024 37020
rect 4048 37018 4104 37020
rect 3808 36966 3854 37018
rect 3854 36966 3864 37018
rect 3888 36966 3918 37018
rect 3918 36966 3930 37018
rect 3930 36966 3944 37018
rect 3968 36966 3982 37018
rect 3982 36966 3994 37018
rect 3994 36966 4024 37018
rect 4048 36966 4058 37018
rect 4058 36966 4104 37018
rect 3808 36964 3864 36966
rect 3888 36964 3944 36966
rect 3968 36964 4024 36966
rect 4048 36964 4104 36966
rect 3072 36474 3128 36476
rect 3152 36474 3208 36476
rect 3232 36474 3288 36476
rect 3312 36474 3368 36476
rect 3072 36422 3118 36474
rect 3118 36422 3128 36474
rect 3152 36422 3182 36474
rect 3182 36422 3194 36474
rect 3194 36422 3208 36474
rect 3232 36422 3246 36474
rect 3246 36422 3258 36474
rect 3258 36422 3288 36474
rect 3312 36422 3322 36474
rect 3322 36422 3368 36474
rect 3072 36420 3128 36422
rect 3152 36420 3208 36422
rect 3232 36420 3288 36422
rect 3312 36420 3368 36422
rect 846 36252 848 36272
rect 848 36252 900 36272
rect 900 36252 902 36272
rect 846 36216 902 36252
rect 3808 35930 3864 35932
rect 3888 35930 3944 35932
rect 3968 35930 4024 35932
rect 4048 35930 4104 35932
rect 3808 35878 3854 35930
rect 3854 35878 3864 35930
rect 3888 35878 3918 35930
rect 3918 35878 3930 35930
rect 3930 35878 3944 35930
rect 3968 35878 3982 35930
rect 3982 35878 3994 35930
rect 3994 35878 4024 35930
rect 4048 35878 4058 35930
rect 4058 35878 4104 35930
rect 3808 35876 3864 35878
rect 3888 35876 3944 35878
rect 3968 35876 4024 35878
rect 4048 35876 4104 35878
rect 3072 35386 3128 35388
rect 3152 35386 3208 35388
rect 3232 35386 3288 35388
rect 3312 35386 3368 35388
rect 3072 35334 3118 35386
rect 3118 35334 3128 35386
rect 3152 35334 3182 35386
rect 3182 35334 3194 35386
rect 3194 35334 3208 35386
rect 3232 35334 3246 35386
rect 3246 35334 3258 35386
rect 3258 35334 3288 35386
rect 3312 35334 3322 35386
rect 3322 35334 3368 35386
rect 3072 35332 3128 35334
rect 3152 35332 3208 35334
rect 3232 35332 3288 35334
rect 3312 35332 3368 35334
rect 846 34892 848 34912
rect 848 34892 900 34912
rect 900 34892 902 34912
rect 846 34856 902 34892
rect 3808 34842 3864 34844
rect 3888 34842 3944 34844
rect 3968 34842 4024 34844
rect 4048 34842 4104 34844
rect 3808 34790 3854 34842
rect 3854 34790 3864 34842
rect 3888 34790 3918 34842
rect 3918 34790 3930 34842
rect 3930 34790 3944 34842
rect 3968 34790 3982 34842
rect 3982 34790 3994 34842
rect 3994 34790 4024 34842
rect 4048 34790 4058 34842
rect 4058 34790 4104 34842
rect 3808 34788 3864 34790
rect 3888 34788 3944 34790
rect 3968 34788 4024 34790
rect 4048 34788 4104 34790
rect 3072 34298 3128 34300
rect 3152 34298 3208 34300
rect 3232 34298 3288 34300
rect 3312 34298 3368 34300
rect 3072 34246 3118 34298
rect 3118 34246 3128 34298
rect 3152 34246 3182 34298
rect 3182 34246 3194 34298
rect 3194 34246 3208 34298
rect 3232 34246 3246 34298
rect 3246 34246 3258 34298
rect 3258 34246 3288 34298
rect 3312 34246 3322 34298
rect 3322 34246 3368 34298
rect 3072 34244 3128 34246
rect 3152 34244 3208 34246
rect 3232 34244 3288 34246
rect 3312 34244 3368 34246
rect 3808 33754 3864 33756
rect 3888 33754 3944 33756
rect 3968 33754 4024 33756
rect 4048 33754 4104 33756
rect 3808 33702 3854 33754
rect 3854 33702 3864 33754
rect 3888 33702 3918 33754
rect 3918 33702 3930 33754
rect 3930 33702 3944 33754
rect 3968 33702 3982 33754
rect 3982 33702 3994 33754
rect 3994 33702 4024 33754
rect 4048 33702 4058 33754
rect 4058 33702 4104 33754
rect 3808 33700 3864 33702
rect 3888 33700 3944 33702
rect 3968 33700 4024 33702
rect 4048 33700 4104 33702
rect 846 33260 848 33280
rect 848 33260 900 33280
rect 900 33260 902 33280
rect 846 33224 902 33260
rect 3072 33210 3128 33212
rect 3152 33210 3208 33212
rect 3232 33210 3288 33212
rect 3312 33210 3368 33212
rect 3072 33158 3118 33210
rect 3118 33158 3128 33210
rect 3152 33158 3182 33210
rect 3182 33158 3194 33210
rect 3194 33158 3208 33210
rect 3232 33158 3246 33210
rect 3246 33158 3258 33210
rect 3258 33158 3288 33210
rect 3312 33158 3322 33210
rect 3322 33158 3368 33210
rect 3072 33156 3128 33158
rect 3152 33156 3208 33158
rect 3232 33156 3288 33158
rect 3312 33156 3368 33158
rect 3808 32666 3864 32668
rect 3888 32666 3944 32668
rect 3968 32666 4024 32668
rect 4048 32666 4104 32668
rect 3808 32614 3854 32666
rect 3854 32614 3864 32666
rect 3888 32614 3918 32666
rect 3918 32614 3930 32666
rect 3930 32614 3944 32666
rect 3968 32614 3982 32666
rect 3982 32614 3994 32666
rect 3994 32614 4024 32666
rect 4048 32614 4058 32666
rect 4058 32614 4104 32666
rect 3808 32612 3864 32614
rect 3888 32612 3944 32614
rect 3968 32612 4024 32614
rect 4048 32612 4104 32614
rect 846 32172 848 32192
rect 848 32172 900 32192
rect 900 32172 902 32192
rect 846 32136 902 32172
rect 3072 32122 3128 32124
rect 3152 32122 3208 32124
rect 3232 32122 3288 32124
rect 3312 32122 3368 32124
rect 3072 32070 3118 32122
rect 3118 32070 3128 32122
rect 3152 32070 3182 32122
rect 3182 32070 3194 32122
rect 3194 32070 3208 32122
rect 3232 32070 3246 32122
rect 3246 32070 3258 32122
rect 3258 32070 3288 32122
rect 3312 32070 3322 32122
rect 3322 32070 3368 32122
rect 3072 32068 3128 32070
rect 3152 32068 3208 32070
rect 3232 32068 3288 32070
rect 3312 32068 3368 32070
rect 3808 31578 3864 31580
rect 3888 31578 3944 31580
rect 3968 31578 4024 31580
rect 4048 31578 4104 31580
rect 3808 31526 3854 31578
rect 3854 31526 3864 31578
rect 3888 31526 3918 31578
rect 3918 31526 3930 31578
rect 3930 31526 3944 31578
rect 3968 31526 3982 31578
rect 3982 31526 3994 31578
rect 3994 31526 4024 31578
rect 4048 31526 4058 31578
rect 4058 31526 4104 31578
rect 3808 31524 3864 31526
rect 3888 31524 3944 31526
rect 3968 31524 4024 31526
rect 4048 31524 4104 31526
rect 3072 31034 3128 31036
rect 3152 31034 3208 31036
rect 3232 31034 3288 31036
rect 3312 31034 3368 31036
rect 3072 30982 3118 31034
rect 3118 30982 3128 31034
rect 3152 30982 3182 31034
rect 3182 30982 3194 31034
rect 3194 30982 3208 31034
rect 3232 30982 3246 31034
rect 3246 30982 3258 31034
rect 3258 30982 3288 31034
rect 3312 30982 3322 31034
rect 3322 30982 3368 31034
rect 3072 30980 3128 30982
rect 3152 30980 3208 30982
rect 3232 30980 3288 30982
rect 3312 30980 3368 30982
rect 4986 48048 5042 48104
rect 4894 47912 4950 47968
rect 5354 47096 5410 47152
rect 5262 46416 5318 46472
rect 846 30812 848 30832
rect 848 30812 900 30832
rect 900 30812 902 30832
rect 846 30776 902 30812
rect 3808 30490 3864 30492
rect 3888 30490 3944 30492
rect 3968 30490 4024 30492
rect 4048 30490 4104 30492
rect 3808 30438 3854 30490
rect 3854 30438 3864 30490
rect 3888 30438 3918 30490
rect 3918 30438 3930 30490
rect 3930 30438 3944 30490
rect 3968 30438 3982 30490
rect 3982 30438 3994 30490
rect 3994 30438 4024 30490
rect 4048 30438 4058 30490
rect 4058 30438 4104 30490
rect 3808 30436 3864 30438
rect 3888 30436 3944 30438
rect 3968 30436 4024 30438
rect 4048 30436 4104 30438
rect 3072 29946 3128 29948
rect 3152 29946 3208 29948
rect 3232 29946 3288 29948
rect 3312 29946 3368 29948
rect 3072 29894 3118 29946
rect 3118 29894 3128 29946
rect 3152 29894 3182 29946
rect 3182 29894 3194 29946
rect 3194 29894 3208 29946
rect 3232 29894 3246 29946
rect 3246 29894 3258 29946
rect 3258 29894 3288 29946
rect 3312 29894 3322 29946
rect 3322 29894 3368 29946
rect 3072 29892 3128 29894
rect 3152 29892 3208 29894
rect 3232 29892 3288 29894
rect 3312 29892 3368 29894
rect 846 29452 848 29472
rect 848 29452 900 29472
rect 900 29452 902 29472
rect 846 29416 902 29452
rect 3808 29402 3864 29404
rect 3888 29402 3944 29404
rect 3968 29402 4024 29404
rect 4048 29402 4104 29404
rect 3808 29350 3854 29402
rect 3854 29350 3864 29402
rect 3888 29350 3918 29402
rect 3918 29350 3930 29402
rect 3930 29350 3944 29402
rect 3968 29350 3982 29402
rect 3982 29350 3994 29402
rect 3994 29350 4024 29402
rect 4048 29350 4058 29402
rect 4058 29350 4104 29402
rect 3808 29348 3864 29350
rect 3888 29348 3944 29350
rect 3968 29348 4024 29350
rect 4048 29348 4104 29350
rect 3072 28858 3128 28860
rect 3152 28858 3208 28860
rect 3232 28858 3288 28860
rect 3312 28858 3368 28860
rect 3072 28806 3118 28858
rect 3118 28806 3128 28858
rect 3152 28806 3182 28858
rect 3182 28806 3194 28858
rect 3194 28806 3208 28858
rect 3232 28806 3246 28858
rect 3246 28806 3258 28858
rect 3258 28806 3288 28858
rect 3312 28806 3322 28858
rect 3322 28806 3368 28858
rect 3072 28804 3128 28806
rect 3152 28804 3208 28806
rect 3232 28804 3288 28806
rect 3312 28804 3368 28806
rect 3808 28314 3864 28316
rect 3888 28314 3944 28316
rect 3968 28314 4024 28316
rect 4048 28314 4104 28316
rect 3808 28262 3854 28314
rect 3854 28262 3864 28314
rect 3888 28262 3918 28314
rect 3918 28262 3930 28314
rect 3930 28262 3944 28314
rect 3968 28262 3982 28314
rect 3982 28262 3994 28314
rect 3994 28262 4024 28314
rect 4048 28262 4058 28314
rect 4058 28262 4104 28314
rect 3808 28260 3864 28262
rect 3888 28260 3944 28262
rect 3968 28260 4024 28262
rect 4048 28260 4104 28262
rect 846 27820 848 27840
rect 848 27820 900 27840
rect 900 27820 902 27840
rect 846 27784 902 27820
rect 3072 27770 3128 27772
rect 3152 27770 3208 27772
rect 3232 27770 3288 27772
rect 3312 27770 3368 27772
rect 3072 27718 3118 27770
rect 3118 27718 3128 27770
rect 3152 27718 3182 27770
rect 3182 27718 3194 27770
rect 3194 27718 3208 27770
rect 3232 27718 3246 27770
rect 3246 27718 3258 27770
rect 3258 27718 3288 27770
rect 3312 27718 3322 27770
rect 3322 27718 3368 27770
rect 3072 27716 3128 27718
rect 3152 27716 3208 27718
rect 3232 27716 3288 27718
rect 3312 27716 3368 27718
rect 3808 27226 3864 27228
rect 3888 27226 3944 27228
rect 3968 27226 4024 27228
rect 4048 27226 4104 27228
rect 3808 27174 3854 27226
rect 3854 27174 3864 27226
rect 3888 27174 3918 27226
rect 3918 27174 3930 27226
rect 3930 27174 3944 27226
rect 3968 27174 3982 27226
rect 3982 27174 3994 27226
rect 3994 27174 4024 27226
rect 4048 27174 4058 27226
rect 4058 27174 4104 27226
rect 3808 27172 3864 27174
rect 3888 27172 3944 27174
rect 3968 27172 4024 27174
rect 4048 27172 4104 27174
rect 3072 26682 3128 26684
rect 3152 26682 3208 26684
rect 3232 26682 3288 26684
rect 3312 26682 3368 26684
rect 3072 26630 3118 26682
rect 3118 26630 3128 26682
rect 3152 26630 3182 26682
rect 3182 26630 3194 26682
rect 3194 26630 3208 26682
rect 3232 26630 3246 26682
rect 3246 26630 3258 26682
rect 3258 26630 3288 26682
rect 3312 26630 3322 26682
rect 3322 26630 3368 26682
rect 3072 26628 3128 26630
rect 3152 26628 3208 26630
rect 3232 26628 3288 26630
rect 3312 26628 3368 26630
rect 1306 26560 1362 26616
rect 3808 26138 3864 26140
rect 3888 26138 3944 26140
rect 3968 26138 4024 26140
rect 4048 26138 4104 26140
rect 3808 26086 3854 26138
rect 3854 26086 3864 26138
rect 3888 26086 3918 26138
rect 3918 26086 3930 26138
rect 3930 26086 3944 26138
rect 3968 26086 3982 26138
rect 3982 26086 3994 26138
rect 3994 26086 4024 26138
rect 4048 26086 4058 26138
rect 4058 26086 4104 26138
rect 3808 26084 3864 26086
rect 3888 26084 3944 26086
rect 3968 26084 4024 26086
rect 4048 26084 4104 26086
rect 3072 25594 3128 25596
rect 3152 25594 3208 25596
rect 3232 25594 3288 25596
rect 3312 25594 3368 25596
rect 3072 25542 3118 25594
rect 3118 25542 3128 25594
rect 3152 25542 3182 25594
rect 3182 25542 3194 25594
rect 3194 25542 3208 25594
rect 3232 25542 3246 25594
rect 3246 25542 3258 25594
rect 3258 25542 3288 25594
rect 3312 25542 3322 25594
rect 3322 25542 3368 25594
rect 3072 25540 3128 25542
rect 3152 25540 3208 25542
rect 3232 25540 3288 25542
rect 3312 25540 3368 25542
rect 1214 25236 1216 25256
rect 1216 25236 1268 25256
rect 1268 25236 1270 25256
rect 1214 25200 1270 25236
rect 3808 25050 3864 25052
rect 3888 25050 3944 25052
rect 3968 25050 4024 25052
rect 4048 25050 4104 25052
rect 3808 24998 3854 25050
rect 3854 24998 3864 25050
rect 3888 24998 3918 25050
rect 3918 24998 3930 25050
rect 3930 24998 3944 25050
rect 3968 24998 3982 25050
rect 3982 24998 3994 25050
rect 3994 24998 4024 25050
rect 4048 24998 4058 25050
rect 4058 24998 4104 25050
rect 3808 24996 3864 24998
rect 3888 24996 3944 24998
rect 3968 24996 4024 24998
rect 4048 24996 4104 24998
rect 3072 24506 3128 24508
rect 3152 24506 3208 24508
rect 3232 24506 3288 24508
rect 3312 24506 3368 24508
rect 3072 24454 3118 24506
rect 3118 24454 3128 24506
rect 3152 24454 3182 24506
rect 3182 24454 3194 24506
rect 3194 24454 3208 24506
rect 3232 24454 3246 24506
rect 3246 24454 3258 24506
rect 3258 24454 3288 24506
rect 3312 24454 3322 24506
rect 3322 24454 3368 24506
rect 3072 24452 3128 24454
rect 3152 24452 3208 24454
rect 3232 24452 3288 24454
rect 3312 24452 3368 24454
rect 3808 23962 3864 23964
rect 3888 23962 3944 23964
rect 3968 23962 4024 23964
rect 4048 23962 4104 23964
rect 3808 23910 3854 23962
rect 3854 23910 3864 23962
rect 3888 23910 3918 23962
rect 3918 23910 3930 23962
rect 3930 23910 3944 23962
rect 3968 23910 3982 23962
rect 3982 23910 3994 23962
rect 3994 23910 4024 23962
rect 4048 23910 4058 23962
rect 4058 23910 4104 23962
rect 3808 23908 3864 23910
rect 3888 23908 3944 23910
rect 3968 23908 4024 23910
rect 4048 23908 4104 23910
rect 1306 23840 1362 23896
rect 3072 23418 3128 23420
rect 3152 23418 3208 23420
rect 3232 23418 3288 23420
rect 3312 23418 3368 23420
rect 3072 23366 3118 23418
rect 3118 23366 3128 23418
rect 3152 23366 3182 23418
rect 3182 23366 3194 23418
rect 3194 23366 3208 23418
rect 3232 23366 3246 23418
rect 3246 23366 3258 23418
rect 3258 23366 3288 23418
rect 3312 23366 3322 23418
rect 3322 23366 3368 23418
rect 3072 23364 3128 23366
rect 3152 23364 3208 23366
rect 3232 23364 3288 23366
rect 3312 23364 3368 23366
rect 3808 22874 3864 22876
rect 3888 22874 3944 22876
rect 3968 22874 4024 22876
rect 4048 22874 4104 22876
rect 3808 22822 3854 22874
rect 3854 22822 3864 22874
rect 3888 22822 3918 22874
rect 3918 22822 3930 22874
rect 3930 22822 3944 22874
rect 3968 22822 3982 22874
rect 3982 22822 3994 22874
rect 3994 22822 4024 22874
rect 4048 22822 4058 22874
rect 4058 22822 4104 22874
rect 3808 22820 3864 22822
rect 3888 22820 3944 22822
rect 3968 22820 4024 22822
rect 4048 22820 4104 22822
rect 1306 22480 1362 22536
rect 3072 22330 3128 22332
rect 3152 22330 3208 22332
rect 3232 22330 3288 22332
rect 3312 22330 3368 22332
rect 3072 22278 3118 22330
rect 3118 22278 3128 22330
rect 3152 22278 3182 22330
rect 3182 22278 3194 22330
rect 3194 22278 3208 22330
rect 3232 22278 3246 22330
rect 3246 22278 3258 22330
rect 3258 22278 3288 22330
rect 3312 22278 3322 22330
rect 3322 22278 3368 22330
rect 3072 22276 3128 22278
rect 3152 22276 3208 22278
rect 3232 22276 3288 22278
rect 3312 22276 3368 22278
rect 3808 21786 3864 21788
rect 3888 21786 3944 21788
rect 3968 21786 4024 21788
rect 4048 21786 4104 21788
rect 3808 21734 3854 21786
rect 3854 21734 3864 21786
rect 3888 21734 3918 21786
rect 3918 21734 3930 21786
rect 3930 21734 3944 21786
rect 3968 21734 3982 21786
rect 3982 21734 3994 21786
rect 3994 21734 4024 21786
rect 4048 21734 4058 21786
rect 4058 21734 4104 21786
rect 3808 21732 3864 21734
rect 3888 21732 3944 21734
rect 3968 21732 4024 21734
rect 4048 21732 4104 21734
rect 3072 21242 3128 21244
rect 3152 21242 3208 21244
rect 3232 21242 3288 21244
rect 3312 21242 3368 21244
rect 3072 21190 3118 21242
rect 3118 21190 3128 21242
rect 3152 21190 3182 21242
rect 3182 21190 3194 21242
rect 3194 21190 3208 21242
rect 3232 21190 3246 21242
rect 3246 21190 3258 21242
rect 3258 21190 3288 21242
rect 3312 21190 3322 21242
rect 3322 21190 3368 21242
rect 3072 21188 3128 21190
rect 3152 21188 3208 21190
rect 3232 21188 3288 21190
rect 3312 21188 3368 21190
rect 1306 21120 1362 21176
rect 3808 20698 3864 20700
rect 3888 20698 3944 20700
rect 3968 20698 4024 20700
rect 4048 20698 4104 20700
rect 3808 20646 3854 20698
rect 3854 20646 3864 20698
rect 3888 20646 3918 20698
rect 3918 20646 3930 20698
rect 3930 20646 3944 20698
rect 3968 20646 3982 20698
rect 3982 20646 3994 20698
rect 3994 20646 4024 20698
rect 4048 20646 4058 20698
rect 4058 20646 4104 20698
rect 3808 20644 3864 20646
rect 3888 20644 3944 20646
rect 3968 20644 4024 20646
rect 4048 20644 4104 20646
rect 3072 20154 3128 20156
rect 3152 20154 3208 20156
rect 3232 20154 3288 20156
rect 3312 20154 3368 20156
rect 3072 20102 3118 20154
rect 3118 20102 3128 20154
rect 3152 20102 3182 20154
rect 3182 20102 3194 20154
rect 3194 20102 3208 20154
rect 3232 20102 3246 20154
rect 3246 20102 3258 20154
rect 3258 20102 3288 20154
rect 3312 20102 3322 20154
rect 3322 20102 3368 20154
rect 3072 20100 3128 20102
rect 3152 20100 3208 20102
rect 3232 20100 3288 20102
rect 3312 20100 3368 20102
rect 1214 19796 1216 19816
rect 1216 19796 1268 19816
rect 1268 19796 1270 19816
rect 1214 19760 1270 19796
rect 3808 19610 3864 19612
rect 3888 19610 3944 19612
rect 3968 19610 4024 19612
rect 4048 19610 4104 19612
rect 3808 19558 3854 19610
rect 3854 19558 3864 19610
rect 3888 19558 3918 19610
rect 3918 19558 3930 19610
rect 3930 19558 3944 19610
rect 3968 19558 3982 19610
rect 3982 19558 3994 19610
rect 3994 19558 4024 19610
rect 4048 19558 4058 19610
rect 4058 19558 4104 19610
rect 3808 19556 3864 19558
rect 3888 19556 3944 19558
rect 3968 19556 4024 19558
rect 4048 19556 4104 19558
rect 3072 19066 3128 19068
rect 3152 19066 3208 19068
rect 3232 19066 3288 19068
rect 3312 19066 3368 19068
rect 3072 19014 3118 19066
rect 3118 19014 3128 19066
rect 3152 19014 3182 19066
rect 3182 19014 3194 19066
rect 3194 19014 3208 19066
rect 3232 19014 3246 19066
rect 3246 19014 3258 19066
rect 3258 19014 3288 19066
rect 3312 19014 3322 19066
rect 3322 19014 3368 19066
rect 3072 19012 3128 19014
rect 3152 19012 3208 19014
rect 3232 19012 3288 19014
rect 3312 19012 3368 19014
rect 3808 18522 3864 18524
rect 3888 18522 3944 18524
rect 3968 18522 4024 18524
rect 4048 18522 4104 18524
rect 3808 18470 3854 18522
rect 3854 18470 3864 18522
rect 3888 18470 3918 18522
rect 3918 18470 3930 18522
rect 3930 18470 3944 18522
rect 3968 18470 3982 18522
rect 3982 18470 3994 18522
rect 3994 18470 4024 18522
rect 4048 18470 4058 18522
rect 4058 18470 4104 18522
rect 3808 18468 3864 18470
rect 3888 18468 3944 18470
rect 3968 18468 4024 18470
rect 4048 18468 4104 18470
rect 1306 18400 1362 18456
rect 3072 17978 3128 17980
rect 3152 17978 3208 17980
rect 3232 17978 3288 17980
rect 3312 17978 3368 17980
rect 3072 17926 3118 17978
rect 3118 17926 3128 17978
rect 3152 17926 3182 17978
rect 3182 17926 3194 17978
rect 3194 17926 3208 17978
rect 3232 17926 3246 17978
rect 3246 17926 3258 17978
rect 3258 17926 3288 17978
rect 3312 17926 3322 17978
rect 3322 17926 3368 17978
rect 3072 17924 3128 17926
rect 3152 17924 3208 17926
rect 3232 17924 3288 17926
rect 3312 17924 3368 17926
rect 3808 17434 3864 17436
rect 3888 17434 3944 17436
rect 3968 17434 4024 17436
rect 4048 17434 4104 17436
rect 3808 17382 3854 17434
rect 3854 17382 3864 17434
rect 3888 17382 3918 17434
rect 3918 17382 3930 17434
rect 3930 17382 3944 17434
rect 3968 17382 3982 17434
rect 3982 17382 3994 17434
rect 3994 17382 4024 17434
rect 4048 17382 4058 17434
rect 4058 17382 4104 17434
rect 3808 17380 3864 17382
rect 3888 17380 3944 17382
rect 3968 17380 4024 17382
rect 4048 17380 4104 17382
rect 1306 17040 1362 17096
rect 3072 16890 3128 16892
rect 3152 16890 3208 16892
rect 3232 16890 3288 16892
rect 3312 16890 3368 16892
rect 3072 16838 3118 16890
rect 3118 16838 3128 16890
rect 3152 16838 3182 16890
rect 3182 16838 3194 16890
rect 3194 16838 3208 16890
rect 3232 16838 3246 16890
rect 3246 16838 3258 16890
rect 3258 16838 3288 16890
rect 3312 16838 3322 16890
rect 3322 16838 3368 16890
rect 3072 16836 3128 16838
rect 3152 16836 3208 16838
rect 3232 16836 3288 16838
rect 3312 16836 3368 16838
rect 3808 16346 3864 16348
rect 3888 16346 3944 16348
rect 3968 16346 4024 16348
rect 4048 16346 4104 16348
rect 3808 16294 3854 16346
rect 3854 16294 3864 16346
rect 3888 16294 3918 16346
rect 3918 16294 3930 16346
rect 3930 16294 3944 16346
rect 3968 16294 3982 16346
rect 3982 16294 3994 16346
rect 3994 16294 4024 16346
rect 4048 16294 4058 16346
rect 4058 16294 4104 16346
rect 3808 16292 3864 16294
rect 3888 16292 3944 16294
rect 3968 16292 4024 16294
rect 4048 16292 4104 16294
rect 3072 15802 3128 15804
rect 3152 15802 3208 15804
rect 3232 15802 3288 15804
rect 3312 15802 3368 15804
rect 3072 15750 3118 15802
rect 3118 15750 3128 15802
rect 3152 15750 3182 15802
rect 3182 15750 3194 15802
rect 3194 15750 3208 15802
rect 3232 15750 3246 15802
rect 3246 15750 3258 15802
rect 3258 15750 3288 15802
rect 3312 15750 3322 15802
rect 3322 15750 3368 15802
rect 3072 15748 3128 15750
rect 3152 15748 3208 15750
rect 3232 15748 3288 15750
rect 3312 15748 3368 15750
rect 1306 15680 1362 15736
rect 3808 15258 3864 15260
rect 3888 15258 3944 15260
rect 3968 15258 4024 15260
rect 4048 15258 4104 15260
rect 3808 15206 3854 15258
rect 3854 15206 3864 15258
rect 3888 15206 3918 15258
rect 3918 15206 3930 15258
rect 3930 15206 3944 15258
rect 3968 15206 3982 15258
rect 3982 15206 3994 15258
rect 3994 15206 4024 15258
rect 4048 15206 4058 15258
rect 4058 15206 4104 15258
rect 3808 15204 3864 15206
rect 3888 15204 3944 15206
rect 3968 15204 4024 15206
rect 4048 15204 4104 15206
rect 3072 14714 3128 14716
rect 3152 14714 3208 14716
rect 3232 14714 3288 14716
rect 3312 14714 3368 14716
rect 3072 14662 3118 14714
rect 3118 14662 3128 14714
rect 3152 14662 3182 14714
rect 3182 14662 3194 14714
rect 3194 14662 3208 14714
rect 3232 14662 3246 14714
rect 3246 14662 3258 14714
rect 3258 14662 3288 14714
rect 3312 14662 3322 14714
rect 3322 14662 3368 14714
rect 3072 14660 3128 14662
rect 3152 14660 3208 14662
rect 3232 14660 3288 14662
rect 3312 14660 3368 14662
rect 1214 14356 1216 14376
rect 1216 14356 1268 14376
rect 1268 14356 1270 14376
rect 1214 14320 1270 14356
rect 3808 14170 3864 14172
rect 3888 14170 3944 14172
rect 3968 14170 4024 14172
rect 4048 14170 4104 14172
rect 3808 14118 3854 14170
rect 3854 14118 3864 14170
rect 3888 14118 3918 14170
rect 3918 14118 3930 14170
rect 3930 14118 3944 14170
rect 3968 14118 3982 14170
rect 3982 14118 3994 14170
rect 3994 14118 4024 14170
rect 4048 14118 4058 14170
rect 4058 14118 4104 14170
rect 3808 14116 3864 14118
rect 3888 14116 3944 14118
rect 3968 14116 4024 14118
rect 4048 14116 4104 14118
rect 3072 13626 3128 13628
rect 3152 13626 3208 13628
rect 3232 13626 3288 13628
rect 3312 13626 3368 13628
rect 3072 13574 3118 13626
rect 3118 13574 3128 13626
rect 3152 13574 3182 13626
rect 3182 13574 3194 13626
rect 3194 13574 3208 13626
rect 3232 13574 3246 13626
rect 3246 13574 3258 13626
rect 3258 13574 3288 13626
rect 3312 13574 3322 13626
rect 3322 13574 3368 13626
rect 3072 13572 3128 13574
rect 3152 13572 3208 13574
rect 3232 13572 3288 13574
rect 3312 13572 3368 13574
rect 3808 13082 3864 13084
rect 3888 13082 3944 13084
rect 3968 13082 4024 13084
rect 4048 13082 4104 13084
rect 3808 13030 3854 13082
rect 3854 13030 3864 13082
rect 3888 13030 3918 13082
rect 3918 13030 3930 13082
rect 3930 13030 3944 13082
rect 3968 13030 3982 13082
rect 3982 13030 3994 13082
rect 3994 13030 4024 13082
rect 4048 13030 4058 13082
rect 4058 13030 4104 13082
rect 3808 13028 3864 13030
rect 3888 13028 3944 13030
rect 3968 13028 4024 13030
rect 4048 13028 4104 13030
rect 1306 12960 1362 13016
rect 3072 12538 3128 12540
rect 3152 12538 3208 12540
rect 3232 12538 3288 12540
rect 3312 12538 3368 12540
rect 3072 12486 3118 12538
rect 3118 12486 3128 12538
rect 3152 12486 3182 12538
rect 3182 12486 3194 12538
rect 3194 12486 3208 12538
rect 3232 12486 3246 12538
rect 3246 12486 3258 12538
rect 3258 12486 3288 12538
rect 3312 12486 3322 12538
rect 3322 12486 3368 12538
rect 3072 12484 3128 12486
rect 3152 12484 3208 12486
rect 3232 12484 3288 12486
rect 3312 12484 3368 12486
rect 3808 11994 3864 11996
rect 3888 11994 3944 11996
rect 3968 11994 4024 11996
rect 4048 11994 4104 11996
rect 3808 11942 3854 11994
rect 3854 11942 3864 11994
rect 3888 11942 3918 11994
rect 3918 11942 3930 11994
rect 3930 11942 3944 11994
rect 3968 11942 3982 11994
rect 3982 11942 3994 11994
rect 3994 11942 4024 11994
rect 4048 11942 4058 11994
rect 4058 11942 4104 11994
rect 3808 11940 3864 11942
rect 3888 11940 3944 11942
rect 3968 11940 4024 11942
rect 4048 11940 4104 11942
rect 1306 11600 1362 11656
rect 3072 11450 3128 11452
rect 3152 11450 3208 11452
rect 3232 11450 3288 11452
rect 3312 11450 3368 11452
rect 3072 11398 3118 11450
rect 3118 11398 3128 11450
rect 3152 11398 3182 11450
rect 3182 11398 3194 11450
rect 3194 11398 3208 11450
rect 3232 11398 3246 11450
rect 3246 11398 3258 11450
rect 3258 11398 3288 11450
rect 3312 11398 3322 11450
rect 3322 11398 3368 11450
rect 3072 11396 3128 11398
rect 3152 11396 3208 11398
rect 3232 11396 3288 11398
rect 3312 11396 3368 11398
rect 3808 10906 3864 10908
rect 3888 10906 3944 10908
rect 3968 10906 4024 10908
rect 4048 10906 4104 10908
rect 3808 10854 3854 10906
rect 3854 10854 3864 10906
rect 3888 10854 3918 10906
rect 3918 10854 3930 10906
rect 3930 10854 3944 10906
rect 3968 10854 3982 10906
rect 3982 10854 3994 10906
rect 3994 10854 4024 10906
rect 4048 10854 4058 10906
rect 4058 10854 4104 10906
rect 3808 10852 3864 10854
rect 3888 10852 3944 10854
rect 3968 10852 4024 10854
rect 4048 10852 4104 10854
rect 3072 10362 3128 10364
rect 3152 10362 3208 10364
rect 3232 10362 3288 10364
rect 3312 10362 3368 10364
rect 3072 10310 3118 10362
rect 3118 10310 3128 10362
rect 3152 10310 3182 10362
rect 3182 10310 3194 10362
rect 3194 10310 3208 10362
rect 3232 10310 3246 10362
rect 3246 10310 3258 10362
rect 3258 10310 3288 10362
rect 3312 10310 3322 10362
rect 3322 10310 3368 10362
rect 3072 10308 3128 10310
rect 3152 10308 3208 10310
rect 3232 10308 3288 10310
rect 3312 10308 3368 10310
rect 3808 9818 3864 9820
rect 3888 9818 3944 9820
rect 3968 9818 4024 9820
rect 4048 9818 4104 9820
rect 3808 9766 3854 9818
rect 3854 9766 3864 9818
rect 3888 9766 3918 9818
rect 3918 9766 3930 9818
rect 3930 9766 3944 9818
rect 3968 9766 3982 9818
rect 3982 9766 3994 9818
rect 3994 9766 4024 9818
rect 4048 9766 4058 9818
rect 4058 9766 4104 9818
rect 3808 9764 3864 9766
rect 3888 9764 3944 9766
rect 3968 9764 4024 9766
rect 4048 9764 4104 9766
rect 3072 9274 3128 9276
rect 3152 9274 3208 9276
rect 3232 9274 3288 9276
rect 3312 9274 3368 9276
rect 3072 9222 3118 9274
rect 3118 9222 3128 9274
rect 3152 9222 3182 9274
rect 3182 9222 3194 9274
rect 3194 9222 3208 9274
rect 3232 9222 3246 9274
rect 3246 9222 3258 9274
rect 3258 9222 3288 9274
rect 3312 9222 3322 9274
rect 3322 9222 3368 9274
rect 3072 9220 3128 9222
rect 3152 9220 3208 9222
rect 3232 9220 3288 9222
rect 3312 9220 3368 9222
rect 3808 8730 3864 8732
rect 3888 8730 3944 8732
rect 3968 8730 4024 8732
rect 4048 8730 4104 8732
rect 3808 8678 3854 8730
rect 3854 8678 3864 8730
rect 3888 8678 3918 8730
rect 3918 8678 3930 8730
rect 3930 8678 3944 8730
rect 3968 8678 3982 8730
rect 3982 8678 3994 8730
rect 3994 8678 4024 8730
rect 4048 8678 4058 8730
rect 4058 8678 4104 8730
rect 3808 8676 3864 8678
rect 3888 8676 3944 8678
rect 3968 8676 4024 8678
rect 4048 8676 4104 8678
rect 3072 8186 3128 8188
rect 3152 8186 3208 8188
rect 3232 8186 3288 8188
rect 3312 8186 3368 8188
rect 3072 8134 3118 8186
rect 3118 8134 3128 8186
rect 3152 8134 3182 8186
rect 3182 8134 3194 8186
rect 3194 8134 3208 8186
rect 3232 8134 3246 8186
rect 3246 8134 3258 8186
rect 3258 8134 3288 8186
rect 3312 8134 3322 8186
rect 3322 8134 3368 8186
rect 3072 8132 3128 8134
rect 3152 8132 3208 8134
rect 3232 8132 3288 8134
rect 3312 8132 3368 8134
rect 5906 64776 5962 64832
rect 5906 62192 5962 62248
rect 8298 86672 8354 86728
rect 8298 85312 8354 85368
rect 8298 83988 8300 84008
rect 8300 83988 8352 84008
rect 8352 83988 8354 84008
rect 8298 83952 8354 83988
rect 8298 82592 8354 82648
rect 8298 81232 8354 81288
rect 8298 79872 8354 79928
rect 8298 78548 8300 78568
rect 8300 78548 8352 78568
rect 8352 78548 8354 78568
rect 8298 78512 8354 78548
rect 8298 77152 8354 77208
rect 8298 74432 8354 74488
rect 8298 73108 8300 73128
rect 8300 73108 8352 73128
rect 8352 73108 8354 73128
rect 8298 73072 8354 73108
rect 8298 71712 8354 71768
rect 8298 68584 8354 68640
rect 6366 47640 6422 47696
rect 5262 27104 5318 27160
rect 8298 65864 8354 65920
rect 8298 63144 8354 63200
rect 8298 61240 8354 61296
rect 8298 59880 8354 59936
rect 8298 58520 8354 58576
rect 8298 57160 8354 57216
rect 8298 55800 8354 55856
rect 8298 54440 8354 54496
rect 8298 53080 8354 53136
rect 47306 88340 47308 88360
rect 47308 88340 47360 88360
rect 47360 88340 47362 88360
rect 47306 88304 47362 88340
rect 7562 47232 7618 47288
rect 3808 7642 3864 7644
rect 3888 7642 3944 7644
rect 3968 7642 4024 7644
rect 4048 7642 4104 7644
rect 3808 7590 3854 7642
rect 3854 7590 3864 7642
rect 3888 7590 3918 7642
rect 3918 7590 3930 7642
rect 3930 7590 3944 7642
rect 3968 7590 3982 7642
rect 3982 7590 3994 7642
rect 3994 7590 4024 7642
rect 4048 7590 4058 7642
rect 4058 7590 4104 7642
rect 8114 9968 8170 10024
rect 3808 7588 3864 7590
rect 3888 7588 3944 7590
rect 3968 7588 4024 7590
rect 4048 7588 4104 7590
rect 3072 7098 3128 7100
rect 3152 7098 3208 7100
rect 3232 7098 3288 7100
rect 3312 7098 3368 7100
rect 3072 7046 3118 7098
rect 3118 7046 3128 7098
rect 3152 7046 3182 7098
rect 3182 7046 3194 7098
rect 3194 7046 3208 7098
rect 3232 7046 3246 7098
rect 3246 7046 3258 7098
rect 3258 7046 3288 7098
rect 3312 7046 3322 7098
rect 3322 7046 3368 7098
rect 3072 7044 3128 7046
rect 3152 7044 3208 7046
rect 3232 7044 3288 7046
rect 3312 7044 3368 7046
rect 3808 6554 3864 6556
rect 3888 6554 3944 6556
rect 3968 6554 4024 6556
rect 4048 6554 4104 6556
rect 3808 6502 3854 6554
rect 3854 6502 3864 6554
rect 3888 6502 3918 6554
rect 3918 6502 3930 6554
rect 3930 6502 3944 6554
rect 3968 6502 3982 6554
rect 3982 6502 3994 6554
rect 3994 6502 4024 6554
rect 4048 6502 4058 6554
rect 4058 6502 4104 6554
rect 3808 6500 3864 6502
rect 3888 6500 3944 6502
rect 3968 6500 4024 6502
rect 4048 6500 4104 6502
rect 3072 6010 3128 6012
rect 3152 6010 3208 6012
rect 3232 6010 3288 6012
rect 3312 6010 3368 6012
rect 3072 5958 3118 6010
rect 3118 5958 3128 6010
rect 3152 5958 3182 6010
rect 3182 5958 3194 6010
rect 3194 5958 3208 6010
rect 3232 5958 3246 6010
rect 3246 5958 3258 6010
rect 3258 5958 3288 6010
rect 3312 5958 3322 6010
rect 3322 5958 3368 6010
rect 3072 5956 3128 5958
rect 3152 5956 3208 5958
rect 3232 5956 3288 5958
rect 3312 5956 3368 5958
rect 3808 5466 3864 5468
rect 3888 5466 3944 5468
rect 3968 5466 4024 5468
rect 4048 5466 4104 5468
rect 3808 5414 3854 5466
rect 3854 5414 3864 5466
rect 3888 5414 3918 5466
rect 3918 5414 3930 5466
rect 3930 5414 3944 5466
rect 3968 5414 3982 5466
rect 3982 5414 3994 5466
rect 3994 5414 4024 5466
rect 4048 5414 4058 5466
rect 4058 5414 4104 5466
rect 3808 5412 3864 5414
rect 3888 5412 3944 5414
rect 3968 5412 4024 5414
rect 4048 5412 4104 5414
rect 46754 50496 46810 50552
rect 46754 50360 46810 50416
rect 8390 49680 8446 49736
rect 11242 46960 11298 47016
rect 40682 49272 40738 49328
rect 40682 48864 40738 48920
rect 46846 50224 46902 50280
rect 47214 49680 47270 49736
rect 46846 47540 46848 47560
rect 46848 47540 46900 47560
rect 46900 47540 46902 47560
rect 46846 47504 46902 47540
rect 46754 47368 46810 47424
rect 8298 46008 8354 46064
rect 8298 44276 8300 44296
rect 8300 44276 8352 44296
rect 8352 44276 8354 44296
rect 8298 44240 8354 44276
rect 8298 43324 8300 43344
rect 8300 43324 8352 43344
rect 8352 43324 8354 43344
rect 8298 43288 8354 43324
rect 8298 41556 8300 41576
rect 8300 41556 8352 41576
rect 8352 41556 8354 41576
rect 8298 41520 8354 41556
rect 8298 40568 8354 40624
rect 8298 38836 8300 38856
rect 8300 38836 8352 38856
rect 8352 38836 8354 38856
rect 8298 38800 8354 38836
rect 8298 37884 8300 37904
rect 8300 37884 8352 37904
rect 8352 37884 8354 37904
rect 8298 37848 8354 37884
rect 8298 36100 8354 36136
rect 8298 36080 8300 36100
rect 8300 36080 8352 36100
rect 8352 36080 8354 36100
rect 8298 35148 8354 35184
rect 8298 35128 8300 35148
rect 8300 35128 8352 35148
rect 8352 35128 8354 35148
rect 8298 33396 8300 33416
rect 8300 33396 8352 33416
rect 8352 33396 8354 33416
rect 8298 33360 8354 33396
rect 8298 32444 8300 32464
rect 8300 32444 8352 32464
rect 8352 32444 8354 32464
rect 8298 32408 8354 32444
rect 8298 30660 8354 30696
rect 8298 30640 8300 30660
rect 8300 30640 8352 30660
rect 8352 30640 8354 30660
rect 8298 29708 8354 29744
rect 8298 29688 8300 29708
rect 8300 29688 8352 29708
rect 8352 29688 8354 29708
rect 8298 27956 8300 27976
rect 8300 27956 8352 27976
rect 8352 27956 8354 27976
rect 8298 27920 8354 27956
rect 8298 26968 8354 27024
rect 8298 25608 8354 25664
rect 8298 24284 8300 24304
rect 8300 24284 8352 24304
rect 8352 24284 8354 24304
rect 8298 24248 8354 24284
rect 8298 22500 8354 22536
rect 8298 22480 8300 22500
rect 8300 22480 8352 22500
rect 8352 22480 8354 22500
rect 8298 21528 8354 21584
rect 8298 20168 8354 20224
rect 8298 18844 8300 18864
rect 8300 18844 8352 18864
rect 8352 18844 8354 18864
rect 8298 18808 8354 18844
rect 8298 17060 8354 17096
rect 8298 17040 8300 17060
rect 8300 17040 8352 17060
rect 8352 17040 8354 17060
rect 8298 16088 8354 16144
rect 8298 14728 8354 14784
rect 8298 13404 8300 13424
rect 8300 13404 8352 13424
rect 8352 13404 8354 13424
rect 8298 13368 8354 13404
rect 8298 11620 8354 11656
rect 8298 11600 8300 11620
rect 8300 11600 8352 11620
rect 8352 11600 8354 11620
rect 8298 8608 8354 8664
rect 36956 4922 37012 4924
rect 37036 4922 37092 4924
rect 37116 4922 37172 4924
rect 37196 4922 37252 4924
rect 36956 4870 37002 4922
rect 37002 4870 37012 4922
rect 37036 4870 37066 4922
rect 37066 4870 37078 4922
rect 37078 4870 37092 4922
rect 37116 4870 37130 4922
rect 37130 4870 37142 4922
rect 37142 4870 37172 4922
rect 37196 4870 37206 4922
rect 37206 4870 37252 4922
rect 36956 4868 37012 4870
rect 37036 4868 37092 4870
rect 37116 4868 37172 4870
rect 37196 4868 37252 4870
rect 36956 3834 37012 3836
rect 37036 3834 37092 3836
rect 37116 3834 37172 3836
rect 37196 3834 37252 3836
rect 36956 3782 37002 3834
rect 37002 3782 37012 3834
rect 37036 3782 37066 3834
rect 37066 3782 37078 3834
rect 37078 3782 37092 3834
rect 37116 3782 37130 3834
rect 37130 3782 37142 3834
rect 37142 3782 37172 3834
rect 37196 3782 37206 3834
rect 37206 3782 37252 3834
rect 36956 3780 37012 3782
rect 37036 3780 37092 3782
rect 37116 3780 37172 3782
rect 37196 3780 37252 3782
rect 36956 2746 37012 2748
rect 37036 2746 37092 2748
rect 37116 2746 37172 2748
rect 37196 2746 37252 2748
rect 36956 2694 37002 2746
rect 37002 2694 37012 2746
rect 37036 2694 37066 2746
rect 37066 2694 37078 2746
rect 37078 2694 37092 2746
rect 37116 2694 37130 2746
rect 37130 2694 37142 2746
rect 37142 2694 37172 2746
rect 37196 2694 37206 2746
rect 37206 2694 37252 2746
rect 36956 2692 37012 2694
rect 37036 2692 37092 2694
rect 37116 2692 37172 2694
rect 37196 2692 37252 2694
rect 37616 5466 37672 5468
rect 37696 5466 37752 5468
rect 37776 5466 37832 5468
rect 37856 5466 37912 5468
rect 37616 5414 37662 5466
rect 37662 5414 37672 5466
rect 37696 5414 37726 5466
rect 37726 5414 37738 5466
rect 37738 5414 37752 5466
rect 37776 5414 37790 5466
rect 37790 5414 37802 5466
rect 37802 5414 37832 5466
rect 37856 5414 37866 5466
rect 37866 5414 37912 5466
rect 37616 5412 37672 5414
rect 37696 5412 37752 5414
rect 37776 5412 37832 5414
rect 37856 5412 37912 5414
rect 37616 4378 37672 4380
rect 37696 4378 37752 4380
rect 37776 4378 37832 4380
rect 37856 4378 37912 4380
rect 37616 4326 37662 4378
rect 37662 4326 37672 4378
rect 37696 4326 37726 4378
rect 37726 4326 37738 4378
rect 37738 4326 37752 4378
rect 37776 4326 37790 4378
rect 37790 4326 37802 4378
rect 37802 4326 37832 4378
rect 37856 4326 37866 4378
rect 37866 4326 37912 4378
rect 37616 4324 37672 4326
rect 37696 4324 37752 4326
rect 37776 4324 37832 4326
rect 37856 4324 37912 4326
rect 37616 3290 37672 3292
rect 37696 3290 37752 3292
rect 37776 3290 37832 3292
rect 37856 3290 37912 3292
rect 37616 3238 37662 3290
rect 37662 3238 37672 3290
rect 37696 3238 37726 3290
rect 37726 3238 37738 3290
rect 37738 3238 37752 3290
rect 37776 3238 37790 3290
rect 37790 3238 37802 3290
rect 37802 3238 37832 3290
rect 37856 3238 37866 3290
rect 37866 3238 37912 3290
rect 37616 3236 37672 3238
rect 37696 3236 37752 3238
rect 37776 3236 37832 3238
rect 37856 3236 37912 3238
rect 47398 46552 47454 46608
rect 47858 49000 47914 49056
rect 72956 95226 73012 95228
rect 73036 95226 73092 95228
rect 73116 95226 73172 95228
rect 73196 95226 73252 95228
rect 72956 95174 73002 95226
rect 73002 95174 73012 95226
rect 73036 95174 73066 95226
rect 73066 95174 73078 95226
rect 73078 95174 73092 95226
rect 73116 95174 73130 95226
rect 73130 95174 73142 95226
rect 73142 95174 73172 95226
rect 73196 95174 73206 95226
rect 73206 95174 73252 95226
rect 72956 95172 73012 95174
rect 73036 95172 73092 95174
rect 73116 95172 73172 95174
rect 73196 95172 73252 95174
rect 72956 94138 73012 94140
rect 73036 94138 73092 94140
rect 73116 94138 73172 94140
rect 73196 94138 73252 94140
rect 72956 94086 73002 94138
rect 73002 94086 73012 94138
rect 73036 94086 73066 94138
rect 73066 94086 73078 94138
rect 73078 94086 73092 94138
rect 73116 94086 73130 94138
rect 73130 94086 73142 94138
rect 73142 94086 73172 94138
rect 73196 94086 73206 94138
rect 73206 94086 73252 94138
rect 72956 94084 73012 94086
rect 73036 94084 73092 94086
rect 73116 94084 73172 94086
rect 73196 94084 73252 94086
rect 72956 93050 73012 93052
rect 73036 93050 73092 93052
rect 73116 93050 73172 93052
rect 73196 93050 73252 93052
rect 72956 92998 73002 93050
rect 73002 92998 73012 93050
rect 73036 92998 73066 93050
rect 73066 92998 73078 93050
rect 73078 92998 73092 93050
rect 73116 92998 73130 93050
rect 73130 92998 73142 93050
rect 73142 92998 73172 93050
rect 73196 92998 73206 93050
rect 73206 92998 73252 93050
rect 72956 92996 73012 92998
rect 73036 92996 73092 92998
rect 73116 92996 73172 92998
rect 73196 92996 73252 92998
rect 72956 91962 73012 91964
rect 73036 91962 73092 91964
rect 73116 91962 73172 91964
rect 73196 91962 73252 91964
rect 72956 91910 73002 91962
rect 73002 91910 73012 91962
rect 73036 91910 73066 91962
rect 73066 91910 73078 91962
rect 73078 91910 73092 91962
rect 73116 91910 73130 91962
rect 73130 91910 73142 91962
rect 73142 91910 73172 91962
rect 73196 91910 73206 91962
rect 73206 91910 73252 91962
rect 72956 91908 73012 91910
rect 73036 91908 73092 91910
rect 73116 91908 73172 91910
rect 73196 91908 73252 91910
rect 73616 94682 73672 94684
rect 73696 94682 73752 94684
rect 73776 94682 73832 94684
rect 73856 94682 73912 94684
rect 73616 94630 73662 94682
rect 73662 94630 73672 94682
rect 73696 94630 73726 94682
rect 73726 94630 73738 94682
rect 73738 94630 73752 94682
rect 73776 94630 73790 94682
rect 73790 94630 73802 94682
rect 73802 94630 73832 94682
rect 73856 94630 73866 94682
rect 73866 94630 73912 94682
rect 73616 94628 73672 94630
rect 73696 94628 73752 94630
rect 73776 94628 73832 94630
rect 73856 94628 73912 94630
rect 73616 93594 73672 93596
rect 73696 93594 73752 93596
rect 73776 93594 73832 93596
rect 73856 93594 73912 93596
rect 73616 93542 73662 93594
rect 73662 93542 73672 93594
rect 73696 93542 73726 93594
rect 73726 93542 73738 93594
rect 73738 93542 73752 93594
rect 73776 93542 73790 93594
rect 73790 93542 73802 93594
rect 73802 93542 73832 93594
rect 73856 93542 73866 93594
rect 73866 93542 73912 93594
rect 73616 93540 73672 93542
rect 73696 93540 73752 93542
rect 73776 93540 73832 93542
rect 73856 93540 73912 93542
rect 73616 92506 73672 92508
rect 73696 92506 73752 92508
rect 73776 92506 73832 92508
rect 73856 92506 73912 92508
rect 73616 92454 73662 92506
rect 73662 92454 73672 92506
rect 73696 92454 73726 92506
rect 73726 92454 73738 92506
rect 73738 92454 73752 92506
rect 73776 92454 73790 92506
rect 73790 92454 73802 92506
rect 73802 92454 73832 92506
rect 73856 92454 73866 92506
rect 73866 92454 73912 92506
rect 73616 92452 73672 92454
rect 73696 92452 73752 92454
rect 73776 92452 73832 92454
rect 73856 92452 73912 92454
rect 73616 91418 73672 91420
rect 73696 91418 73752 91420
rect 73776 91418 73832 91420
rect 73856 91418 73912 91420
rect 73616 91366 73662 91418
rect 73662 91366 73672 91418
rect 73696 91366 73726 91418
rect 73726 91366 73738 91418
rect 73738 91366 73752 91418
rect 73776 91366 73790 91418
rect 73790 91366 73802 91418
rect 73802 91366 73832 91418
rect 73856 91366 73866 91418
rect 73866 91366 73912 91418
rect 73616 91364 73672 91366
rect 73696 91364 73752 91366
rect 73776 91364 73832 91366
rect 73856 91364 73912 91366
rect 86222 92148 86224 92168
rect 86224 92148 86276 92168
rect 86276 92148 86278 92168
rect 86222 92112 86278 92148
rect 85210 91588 85266 91624
rect 85210 91568 85212 91588
rect 85212 91568 85264 91588
rect 85264 91568 85266 91588
rect 85946 91160 86002 91216
rect 86038 89800 86094 89856
rect 86774 92812 86830 92848
rect 86774 92792 86776 92812
rect 86776 92792 86828 92812
rect 86828 92792 86830 92812
rect 87142 92676 87198 92712
rect 87142 92656 87144 92676
rect 87144 92656 87196 92676
rect 87196 92656 87198 92676
rect 86590 92556 86592 92576
rect 86592 92556 86644 92576
rect 86644 92556 86646 92576
rect 86590 92520 86646 92556
rect 87050 92556 87052 92576
rect 87052 92556 87104 92576
rect 87104 92556 87106 92576
rect 87050 92520 87106 92556
rect 86406 91296 86462 91352
rect 86682 91568 86738 91624
rect 86498 88440 86554 88496
rect 86774 87216 86830 87272
rect 86958 86944 87014 87000
rect 86866 85856 86922 85912
rect 86682 81368 86738 81424
rect 86682 71304 86738 71360
rect 85578 50496 85634 50552
rect 48226 49272 48282 49328
rect 51078 46552 51134 46608
rect 86774 68312 86830 68368
rect 85578 49680 85634 49736
rect 85578 46416 85634 46472
rect 87142 87896 87198 87952
rect 87326 87760 87382 87816
rect 87142 87080 87198 87136
rect 87050 78512 87106 78568
rect 87786 92112 87842 92168
rect 87602 87216 87658 87272
rect 87510 85176 87566 85232
rect 87970 92692 87972 92712
rect 87972 92692 88024 92712
rect 88024 92692 88026 92712
rect 87970 92656 88026 92692
rect 87694 86536 87750 86592
rect 88062 83816 88118 83872
rect 87970 82456 88026 82512
rect 87418 75656 87474 75712
rect 88430 89120 88486 89176
rect 88338 88440 88394 88496
rect 88338 87352 88394 87408
rect 88246 79736 88302 79792
rect 87510 74296 87566 74352
rect 87142 71576 87198 71632
rect 88522 85040 88578 85096
rect 88706 86400 88762 86456
rect 88982 82320 89038 82376
rect 89074 80960 89130 81016
rect 88430 72936 88486 72992
rect 89166 78240 89222 78296
rect 89166 76880 89222 76936
rect 89166 75520 89222 75576
rect 89534 83408 89590 83464
rect 89442 79872 89498 79928
rect 89074 71440 89130 71496
rect 88522 70216 88578 70272
rect 88338 68856 88394 68912
rect 88982 68720 89038 68776
rect 87602 64640 87658 64696
rect 87050 61512 87106 61568
rect 86958 57160 87014 57216
rect 87142 57976 87198 58032
rect 87418 56616 87474 56672
rect 87326 53896 87382 53952
rect 87234 52536 87290 52592
rect 87142 51060 87198 51096
rect 87142 51040 87144 51060
rect 87144 51040 87196 51060
rect 87196 51040 87198 51060
rect 87142 50904 87198 50960
rect 87050 50632 87106 50688
rect 86958 50224 87014 50280
rect 86682 43288 86738 43344
rect 87234 49272 87290 49328
rect 88890 63280 88946 63336
rect 87694 61920 87750 61976
rect 87602 50768 87658 50824
rect 88798 60560 88854 60616
rect 87786 59200 87842 59256
rect 87694 49408 87750 49464
rect 87326 49000 87382 49056
rect 88614 57840 88670 57896
rect 88522 55120 88578 55176
rect 88338 53760 88394 53816
rect 88430 52400 88486 52456
rect 88706 56480 88762 56536
rect 87050 47640 87106 47696
rect 86958 44240 87014 44296
rect 86866 41928 86922 41984
rect 86682 27920 86738 27976
rect 86590 13640 86646 13696
rect 86406 8608 86462 8664
rect 86038 8336 86094 8392
rect 72956 6010 73012 6012
rect 73036 6010 73092 6012
rect 73116 6010 73172 6012
rect 73196 6010 73252 6012
rect 72956 5958 73002 6010
rect 73002 5958 73012 6010
rect 73036 5958 73066 6010
rect 73066 5958 73078 6010
rect 73078 5958 73092 6010
rect 73116 5958 73130 6010
rect 73130 5958 73142 6010
rect 73142 5958 73172 6010
rect 73196 5958 73206 6010
rect 73206 5958 73252 6010
rect 72956 5956 73012 5958
rect 73036 5956 73092 5958
rect 73116 5956 73172 5958
rect 73196 5956 73252 5958
rect 73616 5466 73672 5468
rect 73696 5466 73752 5468
rect 73776 5466 73832 5468
rect 73856 5466 73912 5468
rect 73616 5414 73662 5466
rect 73662 5414 73672 5466
rect 73696 5414 73726 5466
rect 73726 5414 73738 5466
rect 73738 5414 73752 5466
rect 73776 5414 73790 5466
rect 73790 5414 73802 5466
rect 73802 5414 73832 5466
rect 73856 5414 73866 5466
rect 73866 5414 73912 5466
rect 73616 5412 73672 5414
rect 73696 5412 73752 5414
rect 73776 5412 73832 5414
rect 73856 5412 73912 5414
rect 72956 4922 73012 4924
rect 73036 4922 73092 4924
rect 73116 4922 73172 4924
rect 73196 4922 73252 4924
rect 72956 4870 73002 4922
rect 73002 4870 73012 4922
rect 73036 4870 73066 4922
rect 73066 4870 73078 4922
rect 73078 4870 73092 4922
rect 73116 4870 73130 4922
rect 73130 4870 73142 4922
rect 73142 4870 73172 4922
rect 73196 4870 73206 4922
rect 73206 4870 73252 4922
rect 72956 4868 73012 4870
rect 73036 4868 73092 4870
rect 73116 4868 73172 4870
rect 73196 4868 73252 4870
rect 73616 4378 73672 4380
rect 73696 4378 73752 4380
rect 73776 4378 73832 4380
rect 73856 4378 73912 4380
rect 73616 4326 73662 4378
rect 73662 4326 73672 4378
rect 73696 4326 73726 4378
rect 73726 4326 73738 4378
rect 73738 4326 73752 4378
rect 73776 4326 73790 4378
rect 73790 4326 73802 4378
rect 73802 4326 73832 4378
rect 73856 4326 73866 4378
rect 73866 4326 73912 4378
rect 73616 4324 73672 4326
rect 73696 4324 73752 4326
rect 73776 4324 73832 4326
rect 73856 4324 73912 4326
rect 72956 3834 73012 3836
rect 73036 3834 73092 3836
rect 73116 3834 73172 3836
rect 73196 3834 73252 3836
rect 72956 3782 73002 3834
rect 73002 3782 73012 3834
rect 73036 3782 73066 3834
rect 73066 3782 73078 3834
rect 73078 3782 73092 3834
rect 73116 3782 73130 3834
rect 73130 3782 73142 3834
rect 73142 3782 73172 3834
rect 73196 3782 73206 3834
rect 73206 3782 73252 3834
rect 72956 3780 73012 3782
rect 73036 3780 73092 3782
rect 73116 3780 73172 3782
rect 73196 3780 73252 3782
rect 73616 3290 73672 3292
rect 73696 3290 73752 3292
rect 73776 3290 73832 3292
rect 73856 3290 73912 3292
rect 73616 3238 73662 3290
rect 73662 3238 73672 3290
rect 73696 3238 73726 3290
rect 73726 3238 73738 3290
rect 73738 3238 73752 3290
rect 73776 3238 73790 3290
rect 73790 3238 73802 3290
rect 73802 3238 73832 3290
rect 73856 3238 73866 3290
rect 73866 3238 73912 3290
rect 73616 3236 73672 3238
rect 73696 3236 73752 3238
rect 73776 3236 73832 3238
rect 73856 3236 73912 3238
rect 72956 2746 73012 2748
rect 73036 2746 73092 2748
rect 73116 2746 73172 2748
rect 73196 2746 73252 2748
rect 72956 2694 73002 2746
rect 73002 2694 73012 2746
rect 73036 2694 73066 2746
rect 73066 2694 73078 2746
rect 73078 2694 73092 2746
rect 73116 2694 73130 2746
rect 73130 2694 73142 2746
rect 73142 2694 73172 2746
rect 73196 2694 73206 2746
rect 73206 2694 73252 2746
rect 72956 2692 73012 2694
rect 73036 2692 73092 2694
rect 73116 2692 73172 2694
rect 73196 2692 73252 2694
rect 85670 8200 85726 8256
rect 85762 7928 85818 7984
rect 85118 5788 85120 5808
rect 85120 5788 85172 5808
rect 85172 5788 85174 5808
rect 85118 5752 85174 5788
rect 85578 5636 85634 5672
rect 85578 5616 85580 5636
rect 85580 5616 85632 5636
rect 85632 5616 85634 5636
rect 86314 8064 86370 8120
rect 86590 8472 86646 8528
rect 86498 5364 86554 5400
rect 87234 47368 87290 47424
rect 87142 46552 87198 46608
rect 87050 39616 87106 39672
rect 87234 37712 87290 37768
rect 89074 66000 89130 66056
rect 89258 69808 89314 69864
rect 88062 47912 88118 47968
rect 87510 47776 87566 47832
rect 87418 43152 87474 43208
rect 87326 34992 87382 35048
rect 87142 28192 87198 28248
rect 87234 25472 87290 25528
rect 87142 17312 87198 17368
rect 87050 15408 87106 15464
rect 86498 5344 86500 5364
rect 86500 5344 86552 5364
rect 86552 5344 86554 5364
rect 87510 36352 87566 36408
rect 87878 40704 87934 40760
rect 87694 37440 87750 37496
rect 88338 45600 88394 45656
rect 88338 44240 88394 44296
rect 88522 42880 88578 42936
rect 88338 41792 88394 41848
rect 88062 40160 88118 40216
rect 87970 29552 88026 29608
rect 87878 26832 87934 26888
rect 87602 26560 87658 26616
rect 87510 20032 87566 20088
rect 87418 13232 87474 13288
rect 87326 12552 87382 12608
rect 87878 18672 87934 18728
rect 87786 11872 87842 11928
rect 87234 4820 87290 4856
rect 87234 4800 87236 4820
rect 87236 4800 87288 4820
rect 87288 4800 87290 4820
rect 88890 47232 88946 47288
rect 88706 41520 88762 41576
rect 88614 38800 88670 38856
rect 88706 36080 88762 36136
rect 88798 34720 88854 34776
rect 88982 33360 89038 33416
rect 88890 32000 88946 32056
rect 89350 67088 89406 67144
rect 89350 50088 89406 50144
rect 89166 30640 89222 30696
rect 89166 29280 89222 29336
rect 89074 27920 89130 27976
rect 89166 25200 89222 25256
rect 89074 22480 89130 22536
rect 88430 21120 88486 21176
rect 87970 11056 88026 11112
rect 87970 10512 88026 10568
rect 88246 9560 88302 9616
rect 88338 8880 88394 8936
rect 88246 5480 88302 5536
rect 89074 17040 89130 17096
rect 88982 15680 89038 15736
rect 88614 14592 88670 14648
rect 88522 5908 88578 5944
rect 88522 5888 88524 5908
rect 88524 5888 88576 5908
rect 88576 5888 88578 5908
rect 86958 4548 87014 4584
rect 86958 4528 86960 4548
rect 86960 4528 87012 4548
rect 87012 4528 87014 4548
rect 88890 12960 88946 13016
rect 88798 11600 88854 11656
rect 88706 10240 88762 10296
rect 89258 19488 89314 19544
rect 89350 18128 89406 18184
rect 89442 14048 89498 14104
rect 37616 2202 37672 2204
rect 37696 2202 37752 2204
rect 37776 2202 37832 2204
rect 37856 2202 37912 2204
rect 37616 2150 37662 2202
rect 37662 2150 37672 2202
rect 37696 2150 37726 2202
rect 37726 2150 37738 2202
rect 37738 2150 37752 2202
rect 37776 2150 37790 2202
rect 37790 2150 37802 2202
rect 37802 2150 37832 2202
rect 37856 2150 37866 2202
rect 37866 2150 37912 2202
rect 37616 2148 37672 2150
rect 37696 2148 37752 2150
rect 37776 2148 37832 2150
rect 37856 2148 37912 2150
rect 73616 2202 73672 2204
rect 73696 2202 73752 2204
rect 73776 2202 73832 2204
rect 73856 2202 73912 2204
rect 73616 2150 73662 2202
rect 73662 2150 73672 2202
rect 73696 2150 73726 2202
rect 73726 2150 73738 2202
rect 73738 2150 73752 2202
rect 73776 2150 73790 2202
rect 73790 2150 73802 2202
rect 73802 2150 73832 2202
rect 73856 2150 73866 2202
rect 73866 2150 73912 2202
rect 73616 2148 73672 2150
rect 73696 2148 73752 2150
rect 73776 2148 73832 2150
rect 73856 2148 73912 2150
<< metal3 >>
rect 43437 97338 43503 97341
rect 49325 97338 49391 97341
rect 43437 97336 49391 97338
rect 43437 97280 43442 97336
rect 43498 97280 49330 97336
rect 49386 97280 49391 97336
rect 43437 97278 49391 97280
rect 43437 97275 43503 97278
rect 49325 97275 49391 97278
rect 37606 95776 37922 95777
rect 37606 95712 37612 95776
rect 37676 95712 37692 95776
rect 37756 95712 37772 95776
rect 37836 95712 37852 95776
rect 37916 95712 37922 95776
rect 37606 95711 37922 95712
rect 73606 95776 73922 95777
rect 73606 95712 73612 95776
rect 73676 95712 73692 95776
rect 73756 95712 73772 95776
rect 73836 95712 73852 95776
rect 73916 95712 73922 95776
rect 73606 95711 73922 95712
rect 8477 95300 8543 95301
rect 8477 95296 8524 95300
rect 8588 95298 8594 95300
rect 8477 95240 8482 95296
rect 8477 95236 8524 95240
rect 8588 95238 8634 95298
rect 8588 95236 8594 95238
rect 8477 95235 8543 95236
rect 36946 95232 37262 95233
rect 36946 95168 36952 95232
rect 37016 95168 37032 95232
rect 37096 95168 37112 95232
rect 37176 95168 37192 95232
rect 37256 95168 37262 95232
rect 36946 95167 37262 95168
rect 72946 95232 73262 95233
rect 72946 95168 72952 95232
rect 73016 95168 73032 95232
rect 73096 95168 73112 95232
rect 73176 95168 73192 95232
rect 73256 95168 73262 95232
rect 72946 95167 73262 95168
rect 37606 94688 37922 94689
rect 37606 94624 37612 94688
rect 37676 94624 37692 94688
rect 37756 94624 37772 94688
rect 37836 94624 37852 94688
rect 37916 94624 37922 94688
rect 37606 94623 37922 94624
rect 73606 94688 73922 94689
rect 73606 94624 73612 94688
rect 73676 94624 73692 94688
rect 73756 94624 73772 94688
rect 73836 94624 73852 94688
rect 73916 94624 73922 94688
rect 73606 94623 73922 94624
rect 36946 94144 37262 94145
rect 36946 94080 36952 94144
rect 37016 94080 37032 94144
rect 37096 94080 37112 94144
rect 37176 94080 37192 94144
rect 37256 94080 37262 94144
rect 36946 94079 37262 94080
rect 72946 94144 73262 94145
rect 72946 94080 72952 94144
rect 73016 94080 73032 94144
rect 73096 94080 73112 94144
rect 73176 94080 73192 94144
rect 73256 94080 73262 94144
rect 72946 94079 73262 94080
rect 37606 93600 37922 93601
rect 37606 93536 37612 93600
rect 37676 93536 37692 93600
rect 37756 93536 37772 93600
rect 37836 93536 37852 93600
rect 37916 93536 37922 93600
rect 37606 93535 37922 93536
rect 73606 93600 73922 93601
rect 73606 93536 73612 93600
rect 73676 93536 73692 93600
rect 73756 93536 73772 93600
rect 73836 93536 73852 93600
rect 73916 93536 73922 93600
rect 73606 93535 73922 93536
rect 36946 93056 37262 93057
rect 36946 92992 36952 93056
rect 37016 92992 37032 93056
rect 37096 92992 37112 93056
rect 37176 92992 37192 93056
rect 37256 92992 37262 93056
rect 36946 92991 37262 92992
rect 72946 93056 73262 93057
rect 72946 92992 72952 93056
rect 73016 92992 73032 93056
rect 73096 92992 73112 93056
rect 73176 92992 73192 93056
rect 73256 92992 73262 93056
rect 72946 92991 73262 92992
rect 48078 92788 48084 92852
rect 48148 92850 48154 92852
rect 86769 92850 86835 92853
rect 48148 92848 86835 92850
rect 48148 92792 86774 92848
rect 86830 92792 86835 92848
rect 48148 92790 86835 92792
rect 48148 92788 48154 92790
rect 86769 92787 86835 92790
rect 47526 92652 47532 92716
rect 47596 92714 47602 92716
rect 87137 92714 87203 92717
rect 47596 92712 87203 92714
rect 47596 92656 87142 92712
rect 87198 92656 87203 92712
rect 47596 92654 87203 92656
rect 47596 92652 47602 92654
rect 87137 92651 87203 92654
rect 87965 92714 88031 92717
rect 89110 92714 89116 92716
rect 87965 92712 89116 92714
rect 87965 92656 87970 92712
rect 88026 92656 89116 92712
rect 87965 92654 89116 92656
rect 87965 92651 88031 92654
rect 89110 92652 89116 92654
rect 89180 92652 89186 92716
rect 86585 92580 86651 92581
rect 86534 92578 86540 92580
rect 86494 92518 86540 92578
rect 86604 92576 86651 92580
rect 86646 92520 86651 92576
rect 86534 92516 86540 92518
rect 86604 92516 86651 92520
rect 86585 92515 86651 92516
rect 87045 92580 87111 92581
rect 87045 92576 87092 92580
rect 87156 92578 87162 92580
rect 87045 92520 87050 92576
rect 87045 92516 87092 92520
rect 87156 92518 87202 92578
rect 87156 92516 87162 92518
rect 87045 92515 87111 92516
rect 37606 92512 37922 92513
rect 37606 92448 37612 92512
rect 37676 92448 37692 92512
rect 37756 92448 37772 92512
rect 37836 92448 37852 92512
rect 37916 92448 37922 92512
rect 37606 92447 37922 92448
rect 73606 92512 73922 92513
rect 73606 92448 73612 92512
rect 73676 92448 73692 92512
rect 73756 92448 73772 92512
rect 73836 92448 73852 92512
rect 73916 92448 73922 92512
rect 73606 92447 73922 92448
rect 46841 92170 46907 92173
rect 86217 92170 86283 92173
rect 46841 92168 86283 92170
rect 46841 92112 46846 92168
rect 46902 92112 86222 92168
rect 86278 92112 86283 92168
rect 46841 92110 86283 92112
rect 46841 92107 46907 92110
rect 86217 92107 86283 92110
rect 87781 92170 87847 92173
rect 89294 92170 89300 92172
rect 87781 92168 89300 92170
rect 87781 92112 87786 92168
rect 87842 92112 89300 92168
rect 87781 92110 89300 92112
rect 87781 92107 87847 92110
rect 89294 92108 89300 92110
rect 89364 92108 89370 92172
rect 3062 91968 3378 91969
rect 3062 91904 3068 91968
rect 3132 91904 3148 91968
rect 3212 91904 3228 91968
rect 3292 91904 3308 91968
rect 3372 91904 3378 91968
rect 3062 91903 3378 91904
rect 36946 91968 37262 91969
rect 36946 91904 36952 91968
rect 37016 91904 37032 91968
rect 37096 91904 37112 91968
rect 37176 91904 37192 91968
rect 37256 91904 37262 91968
rect 36946 91903 37262 91904
rect 72946 91968 73262 91969
rect 72946 91904 72952 91968
rect 73016 91904 73032 91968
rect 73096 91904 73112 91968
rect 73176 91904 73192 91968
rect 73256 91904 73262 91968
rect 72946 91903 73262 91904
rect 46749 91626 46815 91629
rect 85205 91626 85271 91629
rect 46749 91624 85271 91626
rect 46749 91568 46754 91624
rect 46810 91568 85210 91624
rect 85266 91568 85271 91624
rect 46749 91566 85271 91568
rect 46749 91563 46815 91566
rect 85205 91563 85271 91566
rect 86677 91626 86743 91629
rect 86902 91626 86908 91628
rect 86677 91624 86908 91626
rect 86677 91568 86682 91624
rect 86738 91568 86908 91624
rect 86677 91566 86908 91568
rect 86677 91563 86743 91566
rect 86902 91564 86908 91566
rect 86972 91564 86978 91628
rect 3798 91424 4114 91425
rect 3798 91360 3804 91424
rect 3868 91360 3884 91424
rect 3948 91360 3964 91424
rect 4028 91360 4044 91424
rect 4108 91360 4114 91424
rect 3798 91359 4114 91360
rect 37606 91424 37922 91425
rect 37606 91360 37612 91424
rect 37676 91360 37692 91424
rect 37756 91360 37772 91424
rect 37836 91360 37852 91424
rect 37916 91360 37922 91424
rect 37606 91359 37922 91360
rect 73606 91424 73922 91425
rect 73606 91360 73612 91424
rect 73676 91360 73692 91424
rect 73756 91360 73772 91424
rect 73836 91360 73852 91424
rect 73916 91360 73922 91424
rect 73606 91359 73922 91360
rect 86401 91356 86467 91357
rect 86350 91354 86356 91356
rect 86310 91294 86356 91354
rect 86420 91352 86467 91356
rect 86462 91296 86467 91352
rect 86350 91292 86356 91294
rect 86420 91292 86467 91296
rect 86401 91291 86467 91292
rect 85941 91218 86007 91221
rect 86718 91218 86724 91220
rect 85941 91216 86724 91218
rect 85941 91160 85946 91216
rect 86002 91160 86724 91216
rect 85941 91158 86724 91160
rect 85941 91155 86007 91158
rect 86718 91156 86724 91158
rect 86788 91156 86794 91220
rect 3062 90880 3378 90881
rect 3062 90816 3068 90880
rect 3132 90816 3148 90880
rect 3212 90816 3228 90880
rect 3292 90816 3308 90880
rect 3372 90816 3378 90880
rect 3062 90815 3378 90816
rect 3798 90336 4114 90337
rect 3798 90272 3804 90336
rect 3868 90272 3884 90336
rect 3948 90272 3964 90336
rect 4028 90272 4044 90336
rect 4108 90272 4114 90336
rect 3798 90271 4114 90272
rect 86033 89858 86099 89861
rect 88374 89858 88380 89860
rect 86033 89856 88380 89858
rect 86033 89800 86038 89856
rect 86094 89800 88380 89856
rect 86033 89798 88380 89800
rect 86033 89795 86099 89798
rect 88374 89796 88380 89798
rect 88444 89796 88450 89860
rect 3062 89792 3378 89793
rect 3062 89728 3068 89792
rect 3132 89728 3148 89792
rect 3212 89728 3228 89792
rect 3292 89728 3308 89792
rect 3372 89728 3378 89792
rect 3062 89727 3378 89728
rect 3798 89248 4114 89249
rect 3798 89184 3804 89248
rect 3868 89184 3884 89248
rect 3948 89184 3964 89248
rect 4028 89184 4044 89248
rect 4108 89184 4114 89248
rect 3798 89183 4114 89184
rect 88425 89178 88491 89181
rect 89200 89178 90000 89208
rect 88425 89176 90000 89178
rect 88425 89120 88430 89176
rect 88486 89120 90000 89176
rect 88425 89118 90000 89120
rect 88425 89115 88491 89118
rect 89200 89088 90000 89118
rect 3062 88704 3378 88705
rect 3062 88640 3068 88704
rect 3132 88640 3148 88704
rect 3212 88640 3228 88704
rect 3292 88640 3308 88704
rect 3372 88640 3378 88704
rect 3062 88639 3378 88640
rect 86493 88498 86559 88501
rect 87270 88498 87276 88500
rect 86493 88496 87276 88498
rect 86493 88440 86498 88496
rect 86554 88440 87276 88496
rect 86493 88438 87276 88440
rect 86493 88435 86559 88438
rect 87270 88436 87276 88438
rect 87340 88436 87346 88500
rect 88333 88498 88399 88501
rect 89200 88498 90000 88528
rect 88333 88496 90000 88498
rect 88333 88440 88338 88496
rect 88394 88440 90000 88496
rect 88333 88438 90000 88440
rect 88333 88435 88399 88438
rect 89200 88408 90000 88438
rect 47301 88362 47367 88365
rect 47710 88362 47716 88364
rect 47301 88360 47716 88362
rect 47301 88304 47306 88360
rect 47362 88304 47716 88360
rect 47301 88302 47716 88304
rect 47301 88299 47367 88302
rect 47710 88300 47716 88302
rect 47780 88300 47786 88364
rect 3798 88160 4114 88161
rect 3798 88096 3804 88160
rect 3868 88096 3884 88160
rect 3948 88096 3964 88160
rect 4028 88096 4044 88160
rect 4108 88096 4114 88160
rect 3798 88095 4114 88096
rect 8518 87892 8524 87956
rect 8588 87892 8594 87956
rect 87137 87954 87203 87957
rect 46828 87894 48116 87954
rect 86940 87952 87203 87954
rect 86940 87896 87142 87952
rect 87198 87896 87203 87952
rect 86940 87894 87203 87896
rect 87137 87891 87203 87894
rect 87321 87818 87387 87821
rect 89200 87818 90000 87848
rect 87321 87816 90000 87818
rect 87321 87760 87326 87816
rect 87382 87760 90000 87816
rect 87321 87758 90000 87760
rect 87321 87755 87387 87758
rect 89200 87728 90000 87758
rect 3062 87616 3378 87617
rect 3062 87552 3068 87616
rect 3132 87552 3148 87616
rect 3212 87552 3228 87616
rect 3292 87552 3308 87616
rect 3372 87552 3378 87616
rect 3062 87551 3378 87552
rect 88333 87410 88399 87413
rect 86542 87408 88399 87410
rect 86542 87352 88338 87408
rect 88394 87352 88399 87408
rect 86542 87350 88399 87352
rect 86542 87276 86602 87350
rect 88333 87347 88399 87350
rect 86534 87212 86540 87276
rect 86604 87212 86610 87276
rect 86769 87274 86835 87277
rect 87597 87274 87663 87277
rect 86769 87272 87663 87274
rect 86769 87216 86774 87272
rect 86830 87216 87602 87272
rect 87658 87216 87663 87272
rect 86769 87214 87663 87216
rect 86769 87211 86835 87214
rect 87597 87211 87663 87214
rect 86902 87076 86908 87140
rect 86972 87138 86978 87140
rect 87137 87138 87203 87141
rect 86972 87136 87203 87138
rect 86972 87080 87142 87136
rect 87198 87080 87203 87136
rect 86972 87078 87203 87080
rect 86972 87076 86978 87078
rect 87137 87075 87203 87078
rect 3798 87072 4114 87073
rect 3798 87008 3804 87072
rect 3868 87008 3884 87072
rect 3948 87008 3964 87072
rect 4028 87008 4044 87072
rect 4108 87008 4114 87072
rect 3798 87007 4114 87008
rect 86718 86940 86724 87004
rect 86788 87002 86794 87004
rect 86953 87002 87019 87005
rect 86788 87000 87019 87002
rect 86788 86944 86958 87000
rect 87014 86944 87019 87000
rect 86788 86942 87019 86944
rect 86788 86940 86794 86942
rect 86953 86939 87019 86942
rect 8293 86730 8359 86733
rect 8293 86728 8402 86730
rect 8293 86672 8298 86728
rect 8354 86672 8402 86728
rect 8293 86667 8402 86672
rect 841 86594 907 86597
rect 798 86592 907 86594
rect 798 86536 846 86592
rect 902 86536 907 86592
rect 8342 86564 8402 86667
rect 87689 86594 87755 86597
rect 798 86531 907 86536
rect 46828 86534 48116 86594
rect 86940 86592 87755 86594
rect 86940 86536 87694 86592
rect 87750 86536 87755 86592
rect 86940 86534 87755 86536
rect 87689 86531 87755 86534
rect 798 86488 858 86531
rect 0 86398 858 86488
rect 3062 86528 3378 86529
rect 3062 86464 3068 86528
rect 3132 86464 3148 86528
rect 3212 86464 3228 86528
rect 3292 86464 3308 86528
rect 3372 86464 3378 86528
rect 3062 86463 3378 86464
rect 88701 86458 88767 86461
rect 89200 86458 90000 86488
rect 88701 86456 90000 86458
rect 88701 86400 88706 86456
rect 88762 86400 90000 86456
rect 88701 86398 90000 86400
rect 0 86368 800 86398
rect 88701 86395 88767 86398
rect 89200 86368 90000 86398
rect 3798 85984 4114 85985
rect 3798 85920 3804 85984
rect 3868 85920 3884 85984
rect 3948 85920 3964 85984
rect 4028 85920 4044 85984
rect 4108 85920 4114 85984
rect 3798 85919 4114 85920
rect 86861 85916 86927 85917
rect 86861 85914 86908 85916
rect 86816 85912 86908 85914
rect 86816 85856 86866 85912
rect 86816 85854 86908 85856
rect 86861 85852 86908 85854
rect 86972 85852 86978 85916
rect 86861 85851 86927 85852
rect 3062 85440 3378 85441
rect 3062 85376 3068 85440
rect 3132 85376 3148 85440
rect 3212 85376 3228 85440
rect 3292 85376 3308 85440
rect 3372 85376 3378 85440
rect 3062 85375 3378 85376
rect 8293 85370 8359 85373
rect 8293 85368 8402 85370
rect 8293 85312 8298 85368
rect 8354 85312 8402 85368
rect 8293 85307 8402 85312
rect 841 85234 907 85237
rect 798 85232 907 85234
rect 798 85176 846 85232
rect 902 85176 907 85232
rect 8342 85204 8402 85307
rect 87505 85234 87571 85237
rect 798 85171 907 85176
rect 46828 85174 48116 85234
rect 86940 85232 87571 85234
rect 86940 85176 87510 85232
rect 87566 85176 87571 85232
rect 86940 85174 87571 85176
rect 87505 85171 87571 85174
rect 798 85128 858 85171
rect 0 85038 858 85128
rect 88517 85098 88583 85101
rect 89200 85098 90000 85128
rect 88517 85096 90000 85098
rect 88517 85040 88522 85096
rect 88578 85040 90000 85096
rect 88517 85038 90000 85040
rect 0 85008 800 85038
rect 88517 85035 88583 85038
rect 89200 85008 90000 85038
rect 3798 84896 4114 84897
rect 3798 84832 3804 84896
rect 3868 84832 3884 84896
rect 3948 84832 3964 84896
rect 4028 84832 4044 84896
rect 4108 84832 4114 84896
rect 3798 84831 4114 84832
rect 3062 84352 3378 84353
rect 3062 84288 3068 84352
rect 3132 84288 3148 84352
rect 3212 84288 3228 84352
rect 3292 84288 3308 84352
rect 3372 84288 3378 84352
rect 3062 84287 3378 84288
rect 8293 84010 8359 84013
rect 8293 84008 8402 84010
rect 8293 83952 8298 84008
rect 8354 83952 8402 84008
rect 8293 83947 8402 83952
rect 841 83874 907 83877
rect 798 83872 907 83874
rect 798 83816 846 83872
rect 902 83816 907 83872
rect 8342 83844 8402 83947
rect 88057 83874 88123 83877
rect 798 83811 907 83816
rect 46828 83814 48116 83874
rect 86940 83872 88123 83874
rect 86940 83816 88062 83872
rect 88118 83816 88123 83872
rect 86940 83814 88123 83816
rect 88057 83811 88123 83814
rect 798 83768 858 83811
rect 0 83678 858 83768
rect 3798 83808 4114 83809
rect 3798 83744 3804 83808
rect 3868 83744 3884 83808
rect 3948 83744 3964 83808
rect 4028 83744 4044 83808
rect 4108 83744 4114 83808
rect 3798 83743 4114 83744
rect 89200 83738 90000 83768
rect 0 83648 800 83678
rect 89164 83648 90000 83738
rect 89164 83466 89224 83648
rect 89529 83466 89595 83469
rect 89164 83464 89595 83466
rect 89164 83408 89534 83464
rect 89590 83408 89595 83464
rect 89164 83406 89595 83408
rect 89529 83403 89595 83406
rect 3062 83264 3378 83265
rect 3062 83200 3068 83264
rect 3132 83200 3148 83264
rect 3212 83200 3228 83264
rect 3292 83200 3308 83264
rect 3372 83200 3378 83264
rect 3062 83199 3378 83200
rect 3798 82720 4114 82721
rect 3798 82656 3804 82720
rect 3868 82656 3884 82720
rect 3948 82656 3964 82720
rect 4028 82656 4044 82720
rect 4108 82656 4114 82720
rect 3798 82655 4114 82656
rect 8293 82650 8359 82653
rect 8293 82648 8402 82650
rect 8293 82592 8298 82648
rect 8354 82592 8402 82648
rect 8293 82587 8402 82592
rect 8342 82484 8402 82587
rect 87965 82514 88031 82517
rect 46828 82454 48116 82514
rect 86940 82512 88031 82514
rect 86940 82456 87970 82512
rect 88026 82456 88031 82512
rect 86940 82454 88031 82456
rect 87965 82451 88031 82454
rect 0 82378 800 82408
rect 88977 82378 89043 82381
rect 89200 82378 90000 82408
rect 0 82288 858 82378
rect 88977 82376 90000 82378
rect 88977 82320 88982 82376
rect 89038 82320 90000 82376
rect 88977 82318 90000 82320
rect 88977 82315 89043 82318
rect 89200 82288 90000 82318
rect 798 82245 858 82288
rect 798 82240 907 82245
rect 798 82184 846 82240
rect 902 82184 907 82240
rect 798 82182 907 82184
rect 841 82179 907 82182
rect 3062 82176 3378 82177
rect 3062 82112 3068 82176
rect 3132 82112 3148 82176
rect 3212 82112 3228 82176
rect 3292 82112 3308 82176
rect 3372 82112 3378 82176
rect 3062 82111 3378 82112
rect 3798 81632 4114 81633
rect 3798 81568 3804 81632
rect 3868 81568 3884 81632
rect 3948 81568 3964 81632
rect 4028 81568 4044 81632
rect 4108 81568 4114 81632
rect 3798 81567 4114 81568
rect 86677 81426 86743 81429
rect 86677 81424 86786 81426
rect 86677 81368 86682 81424
rect 86738 81368 86786 81424
rect 86677 81363 86786 81368
rect 8293 81290 8359 81293
rect 8293 81288 8402 81290
rect 8293 81232 8298 81288
rect 8354 81232 8402 81288
rect 8293 81227 8402 81232
rect 841 81154 907 81157
rect 798 81152 907 81154
rect 798 81096 846 81152
rect 902 81096 907 81152
rect 8342 81124 8402 81227
rect 798 81091 907 81096
rect 46828 81094 48116 81154
rect 86726 81124 86786 81363
rect 798 81048 858 81091
rect 0 80958 858 81048
rect 3062 81088 3378 81089
rect 3062 81024 3068 81088
rect 3132 81024 3148 81088
rect 3212 81024 3228 81088
rect 3292 81024 3308 81088
rect 3372 81024 3378 81088
rect 3062 81023 3378 81024
rect 89069 81018 89135 81021
rect 89200 81018 90000 81048
rect 89069 81016 90000 81018
rect 89069 80960 89074 81016
rect 89130 80960 90000 81016
rect 89069 80958 90000 80960
rect 0 80928 800 80958
rect 89069 80955 89135 80958
rect 89200 80928 90000 80958
rect 3798 80544 4114 80545
rect 3798 80480 3804 80544
rect 3868 80480 3884 80544
rect 3948 80480 3964 80544
rect 4028 80480 4044 80544
rect 4108 80480 4114 80544
rect 3798 80479 4114 80480
rect 3062 80000 3378 80001
rect 3062 79936 3068 80000
rect 3132 79936 3148 80000
rect 3212 79936 3228 80000
rect 3292 79936 3308 80000
rect 3372 79936 3378 80000
rect 3062 79935 3378 79936
rect 8293 79930 8359 79933
rect 89437 79930 89503 79933
rect 8293 79928 8402 79930
rect 8293 79872 8298 79928
rect 8354 79872 8402 79928
rect 8293 79867 8402 79872
rect 8342 79764 8402 79867
rect 89072 79928 89503 79930
rect 89072 79872 89442 79928
rect 89498 79872 89503 79928
rect 89072 79870 89503 79872
rect 88241 79794 88307 79797
rect 46828 79734 48116 79794
rect 86940 79792 88307 79794
rect 86940 79736 88246 79792
rect 88302 79736 88307 79792
rect 86940 79734 88307 79736
rect 88241 79731 88307 79734
rect 0 79658 800 79688
rect 89072 79658 89132 79870
rect 89437 79867 89503 79870
rect 89200 79658 90000 79688
rect 0 79568 858 79658
rect 89072 79598 90000 79658
rect 89200 79568 90000 79598
rect 798 79525 858 79568
rect 798 79520 907 79525
rect 798 79464 846 79520
rect 902 79464 907 79520
rect 798 79462 907 79464
rect 841 79459 907 79462
rect 3798 79456 4114 79457
rect 3798 79392 3804 79456
rect 3868 79392 3884 79456
rect 3948 79392 3964 79456
rect 4028 79392 4044 79456
rect 4108 79392 4114 79456
rect 3798 79391 4114 79392
rect 3062 78912 3378 78913
rect 3062 78848 3068 78912
rect 3132 78848 3148 78912
rect 3212 78848 3228 78912
rect 3292 78848 3308 78912
rect 3372 78848 3378 78912
rect 3062 78847 3378 78848
rect 8293 78570 8359 78573
rect 87045 78570 87111 78573
rect 8293 78568 8402 78570
rect 8293 78512 8298 78568
rect 8354 78512 8402 78568
rect 8293 78507 8402 78512
rect 841 78434 907 78437
rect 798 78432 907 78434
rect 798 78376 846 78432
rect 902 78376 907 78432
rect 8342 78404 8402 78507
rect 86910 78568 87111 78570
rect 86910 78512 87050 78568
rect 87106 78512 87111 78568
rect 86910 78510 87111 78512
rect 798 78371 907 78376
rect 46828 78374 48116 78434
rect 86910 78404 86970 78510
rect 87045 78507 87111 78510
rect 798 78328 858 78371
rect 0 78238 858 78328
rect 3798 78368 4114 78369
rect 3798 78304 3804 78368
rect 3868 78304 3884 78368
rect 3948 78304 3964 78368
rect 4028 78304 4044 78368
rect 4108 78304 4114 78368
rect 3798 78303 4114 78304
rect 89200 78301 90000 78328
rect 89161 78296 90000 78301
rect 89161 78240 89166 78296
rect 89222 78240 90000 78296
rect 0 78208 800 78238
rect 89161 78235 90000 78240
rect 89200 78208 90000 78235
rect 3062 77824 3378 77825
rect 3062 77760 3068 77824
rect 3132 77760 3148 77824
rect 3212 77760 3228 77824
rect 3292 77760 3308 77824
rect 3372 77760 3378 77824
rect 3062 77759 3378 77760
rect 3798 77280 4114 77281
rect 3798 77216 3804 77280
rect 3868 77216 3884 77280
rect 3948 77216 3964 77280
rect 4028 77216 4044 77280
rect 4108 77216 4114 77280
rect 3798 77215 4114 77216
rect 8293 77210 8359 77213
rect 8293 77208 8402 77210
rect 8293 77152 8298 77208
rect 8354 77152 8402 77208
rect 8293 77147 8402 77152
rect 8342 77044 8402 77147
rect 46828 77014 48116 77074
rect 86350 77012 86356 77076
rect 86420 77012 86426 77076
rect 0 76938 800 76968
rect 89200 76941 90000 76968
rect 0 76848 858 76938
rect 89161 76936 90000 76941
rect 89161 76880 89166 76936
rect 89222 76880 90000 76936
rect 89161 76875 90000 76880
rect 89200 76848 90000 76875
rect 798 76805 858 76848
rect 798 76800 907 76805
rect 798 76744 846 76800
rect 902 76744 907 76800
rect 798 76742 907 76744
rect 841 76739 907 76742
rect 3062 76736 3378 76737
rect 3062 76672 3068 76736
rect 3132 76672 3148 76736
rect 3212 76672 3228 76736
rect 3292 76672 3308 76736
rect 3372 76672 3378 76736
rect 3062 76671 3378 76672
rect 3798 76192 4114 76193
rect 3798 76128 3804 76192
rect 3868 76128 3884 76192
rect 3948 76128 3964 76192
rect 4028 76128 4044 76192
rect 4108 76128 4114 76192
rect 3798 76127 4114 76128
rect 841 75714 907 75717
rect 798 75712 907 75714
rect 798 75656 846 75712
rect 902 75656 907 75712
rect 798 75651 907 75656
rect 5533 75714 5599 75717
rect 87413 75714 87479 75717
rect 5533 75712 8188 75714
rect 5533 75656 5538 75712
rect 5594 75656 8188 75712
rect 5533 75654 8188 75656
rect 46828 75654 48116 75714
rect 86940 75712 87479 75714
rect 86940 75656 87418 75712
rect 87474 75656 87479 75712
rect 86940 75654 87479 75656
rect 5533 75651 5599 75654
rect 87413 75651 87479 75654
rect 798 75608 858 75651
rect 0 75518 858 75608
rect 3062 75648 3378 75649
rect 3062 75584 3068 75648
rect 3132 75584 3148 75648
rect 3212 75584 3228 75648
rect 3292 75584 3308 75648
rect 3372 75584 3378 75648
rect 3062 75583 3378 75584
rect 89200 75581 90000 75608
rect 89161 75576 90000 75581
rect 89161 75520 89166 75576
rect 89222 75520 90000 75576
rect 0 75488 800 75518
rect 89161 75515 90000 75520
rect 89200 75488 90000 75515
rect 3798 75104 4114 75105
rect 3798 75040 3804 75104
rect 3868 75040 3884 75104
rect 3948 75040 3964 75104
rect 4028 75040 4044 75104
rect 4108 75040 4114 75104
rect 3798 75039 4114 75040
rect 3062 74560 3378 74561
rect 3062 74496 3068 74560
rect 3132 74496 3148 74560
rect 3212 74496 3228 74560
rect 3292 74496 3308 74560
rect 3372 74496 3378 74560
rect 3062 74495 3378 74496
rect 8293 74490 8359 74493
rect 8293 74488 8402 74490
rect 8293 74432 8298 74488
rect 8354 74432 8402 74488
rect 8293 74427 8402 74432
rect 8342 74324 8402 74427
rect 87505 74354 87571 74357
rect 46828 74294 48116 74354
rect 86940 74352 87571 74354
rect 86940 74296 87510 74352
rect 87566 74296 87571 74352
rect 86940 74294 87571 74296
rect 87505 74291 87571 74294
rect 89110 74292 89116 74356
rect 89180 74354 89186 74356
rect 89180 74292 89224 74354
rect 89164 74248 89224 74292
rect 0 74218 800 74248
rect 0 74128 858 74218
rect 89164 74158 90000 74248
rect 89200 74128 90000 74158
rect 798 74085 858 74128
rect 798 74080 907 74085
rect 798 74024 846 74080
rect 902 74024 907 74080
rect 798 74022 907 74024
rect 841 74019 907 74022
rect 3798 74016 4114 74017
rect 3798 73952 3804 74016
rect 3868 73952 3884 74016
rect 3948 73952 3964 74016
rect 4028 73952 4044 74016
rect 4108 73952 4114 74016
rect 3798 73951 4114 73952
rect 3062 73472 3378 73473
rect 3062 73408 3068 73472
rect 3132 73408 3148 73472
rect 3212 73408 3228 73472
rect 3292 73408 3308 73472
rect 3372 73408 3378 73472
rect 3062 73407 3378 73408
rect 8293 73130 8359 73133
rect 8293 73128 8402 73130
rect 8293 73072 8298 73128
rect 8354 73072 8402 73128
rect 8293 73067 8402 73072
rect 841 72994 907 72997
rect 798 72992 907 72994
rect 798 72936 846 72992
rect 902 72936 907 72992
rect 8342 72964 8402 73067
rect 88425 72994 88491 72997
rect 798 72931 907 72936
rect 46828 72934 48116 72994
rect 86940 72992 88491 72994
rect 86940 72936 88430 72992
rect 88486 72936 88491 72992
rect 86940 72934 88491 72936
rect 88425 72931 88491 72934
rect 798 72888 858 72931
rect 0 72798 858 72888
rect 3798 72928 4114 72929
rect 3798 72864 3804 72928
rect 3868 72864 3884 72928
rect 3948 72864 3964 72928
rect 4028 72864 4044 72928
rect 4108 72864 4114 72928
rect 3798 72863 4114 72864
rect 89200 72860 90000 72888
rect 0 72768 800 72798
rect 89156 72796 89162 72860
rect 89226 72796 90000 72860
rect 89200 72768 90000 72796
rect 3062 72384 3378 72385
rect 3062 72320 3068 72384
rect 3132 72320 3148 72384
rect 3212 72320 3228 72384
rect 3292 72320 3308 72384
rect 3372 72320 3378 72384
rect 3062 72319 3378 72320
rect 3798 71840 4114 71841
rect 3798 71776 3804 71840
rect 3868 71776 3884 71840
rect 3948 71776 3964 71840
rect 4028 71776 4044 71840
rect 4108 71776 4114 71840
rect 3798 71775 4114 71776
rect 8293 71770 8359 71773
rect 8293 71768 8402 71770
rect 8293 71712 8298 71768
rect 8354 71712 8402 71768
rect 8293 71707 8402 71712
rect 8342 71604 8402 71707
rect 87137 71634 87203 71637
rect 46828 71574 48116 71634
rect 86756 71632 87203 71634
rect 86756 71604 87142 71632
rect 86726 71576 87142 71604
rect 87198 71576 87203 71632
rect 86726 71574 87203 71576
rect 0 71498 800 71528
rect 0 71408 858 71498
rect 798 71365 858 71408
rect 86726 71365 86786 71574
rect 87137 71571 87203 71574
rect 89069 71498 89135 71501
rect 89200 71498 90000 71528
rect 89069 71496 90000 71498
rect 89069 71440 89074 71496
rect 89130 71440 90000 71496
rect 89069 71438 90000 71440
rect 89069 71435 89135 71438
rect 89200 71408 90000 71438
rect 798 71360 907 71365
rect 798 71304 846 71360
rect 902 71304 907 71360
rect 798 71302 907 71304
rect 841 71299 907 71302
rect 86677 71360 86786 71365
rect 86677 71304 86682 71360
rect 86738 71304 86786 71360
rect 86677 71302 86786 71304
rect 86677 71299 86743 71302
rect 3062 71296 3378 71297
rect 3062 71232 3068 71296
rect 3132 71232 3148 71296
rect 3212 71232 3228 71296
rect 3292 71232 3308 71296
rect 3372 71232 3378 71296
rect 3062 71231 3378 71232
rect 3798 70752 4114 70753
rect 3798 70688 3804 70752
rect 3868 70688 3884 70752
rect 3948 70688 3964 70752
rect 4028 70688 4044 70752
rect 4108 70688 4114 70752
rect 3798 70687 4114 70688
rect 841 70274 907 70277
rect 798 70272 907 70274
rect 798 70216 846 70272
rect 902 70216 907 70272
rect 798 70211 907 70216
rect 5533 70274 5599 70277
rect 88517 70274 88583 70277
rect 5533 70272 8188 70274
rect 5533 70216 5538 70272
rect 5594 70216 8188 70272
rect 5533 70214 8188 70216
rect 46828 70214 48116 70274
rect 86940 70272 88583 70274
rect 86940 70216 88522 70272
rect 88578 70216 88583 70272
rect 86940 70214 88583 70216
rect 5533 70211 5599 70214
rect 88517 70211 88583 70214
rect 798 70168 858 70211
rect 0 70078 858 70168
rect 3062 70208 3378 70209
rect 3062 70144 3068 70208
rect 3132 70144 3148 70208
rect 3212 70144 3228 70208
rect 3292 70144 3308 70208
rect 3372 70144 3378 70208
rect 3062 70143 3378 70144
rect 89200 70138 90000 70168
rect 89072 70078 90000 70138
rect 0 70048 800 70078
rect 89072 69866 89132 70078
rect 89200 70048 90000 70078
rect 89253 69866 89319 69869
rect 89072 69864 89319 69866
rect 89072 69808 89258 69864
rect 89314 69808 89319 69864
rect 89072 69806 89319 69808
rect 89253 69803 89319 69806
rect 3798 69664 4114 69665
rect 3798 69600 3804 69664
rect 3868 69600 3884 69664
rect 3948 69600 3964 69664
rect 4028 69600 4044 69664
rect 4108 69600 4114 69664
rect 3798 69599 4114 69600
rect 3062 69120 3378 69121
rect 3062 69056 3068 69120
rect 3132 69056 3148 69120
rect 3212 69056 3228 69120
rect 3292 69056 3308 69120
rect 3372 69056 3378 69120
rect 3062 69055 3378 69056
rect 88333 68914 88399 68917
rect 0 68778 800 68808
rect 1209 68778 1275 68781
rect 0 68776 1275 68778
rect 0 68720 1214 68776
rect 1270 68720 1275 68776
rect 0 68718 1275 68720
rect 0 68688 800 68718
rect 1209 68715 1275 68718
rect 8342 68645 8402 68884
rect 46828 68854 48116 68914
rect 86756 68912 88399 68914
rect 86756 68884 88338 68912
rect 86726 68856 88338 68884
rect 88394 68856 88399 68912
rect 86726 68854 88399 68856
rect 8293 68640 8402 68645
rect 8293 68584 8298 68640
rect 8354 68584 8402 68640
rect 8293 68582 8402 68584
rect 8293 68579 8359 68582
rect 3798 68576 4114 68577
rect 3798 68512 3804 68576
rect 3868 68512 3884 68576
rect 3948 68512 3964 68576
rect 4028 68512 4044 68576
rect 4108 68512 4114 68576
rect 3798 68511 4114 68512
rect 86726 68373 86786 68854
rect 88333 68851 88399 68854
rect 88977 68778 89043 68781
rect 89200 68778 90000 68808
rect 88977 68776 90000 68778
rect 88977 68720 88982 68776
rect 89038 68720 90000 68776
rect 88977 68718 90000 68720
rect 88977 68715 89043 68718
rect 89200 68688 90000 68718
rect 86726 68368 86835 68373
rect 86726 68312 86774 68368
rect 86830 68312 86835 68368
rect 86726 68310 86835 68312
rect 86769 68307 86835 68310
rect 3062 68032 3378 68033
rect 3062 67968 3068 68032
rect 3132 67968 3148 68032
rect 3212 67968 3228 68032
rect 3292 67968 3308 68032
rect 3372 67968 3378 68032
rect 3062 67967 3378 67968
rect 5533 67692 5599 67693
rect 5533 67688 5580 67692
rect 5644 67690 5650 67692
rect 5533 67632 5538 67688
rect 5533 67628 5580 67632
rect 5644 67630 5690 67690
rect 5644 67628 5650 67630
rect 5533 67627 5599 67628
rect 5717 67554 5783 67557
rect 88374 67554 88380 67556
rect 5717 67552 8188 67554
rect 5717 67496 5722 67552
rect 5778 67496 8188 67552
rect 5717 67494 8188 67496
rect 46828 67494 48116 67554
rect 86940 67494 88380 67554
rect 5717 67491 5783 67494
rect 88374 67492 88380 67494
rect 88444 67492 88450 67556
rect 3798 67488 4114 67489
rect 0 67418 800 67448
rect 3798 67424 3804 67488
rect 3868 67424 3884 67488
rect 3948 67424 3964 67488
rect 4028 67424 4044 67488
rect 4108 67424 4114 67488
rect 3798 67423 4114 67424
rect 1301 67418 1367 67421
rect 89200 67418 90000 67448
rect 0 67416 1367 67418
rect 0 67360 1306 67416
rect 1362 67360 1367 67416
rect 0 67358 1367 67360
rect 0 67328 800 67358
rect 1301 67355 1367 67358
rect 89072 67358 90000 67418
rect 89072 67146 89132 67358
rect 89200 67328 90000 67358
rect 89345 67146 89411 67149
rect 89072 67144 89411 67146
rect 89072 67088 89350 67144
rect 89406 67088 89411 67144
rect 89072 67086 89411 67088
rect 89345 67083 89411 67086
rect 3062 66944 3378 66945
rect 3062 66880 3068 66944
rect 3132 66880 3148 66944
rect 3212 66880 3228 66944
rect 3292 66880 3308 66944
rect 3372 66880 3378 66944
rect 3062 66879 3378 66880
rect 3798 66400 4114 66401
rect 3798 66336 3804 66400
rect 3868 66336 3884 66400
rect 3948 66336 3964 66400
rect 4028 66336 4044 66400
rect 4108 66336 4114 66400
rect 3798 66335 4114 66336
rect 0 66058 800 66088
rect 1301 66058 1367 66061
rect 0 66056 1367 66058
rect 0 66000 1306 66056
rect 1362 66000 1367 66056
rect 0 65998 1367 66000
rect 0 65968 800 65998
rect 1301 65995 1367 65998
rect 8342 65925 8402 66164
rect 46828 66134 48116 66194
rect 86350 66132 86356 66196
rect 86420 66132 86426 66196
rect 89069 66058 89135 66061
rect 89200 66058 90000 66088
rect 89069 66056 90000 66058
rect 89069 66000 89074 66056
rect 89130 66000 90000 66056
rect 89069 65998 90000 66000
rect 89069 65995 89135 65998
rect 89200 65968 90000 65998
rect 8293 65920 8402 65925
rect 8293 65864 8298 65920
rect 8354 65864 8402 65920
rect 8293 65862 8402 65864
rect 8293 65859 8359 65862
rect 3062 65856 3378 65857
rect 3062 65792 3068 65856
rect 3132 65792 3148 65856
rect 3212 65792 3228 65856
rect 3292 65792 3308 65856
rect 3372 65792 3378 65856
rect 3062 65791 3378 65792
rect 3798 65312 4114 65313
rect 3798 65248 3804 65312
rect 3868 65248 3884 65312
rect 3948 65248 3964 65312
rect 4028 65248 4044 65312
rect 4108 65248 4114 65312
rect 3798 65247 4114 65248
rect 5533 64970 5599 64973
rect 5758 64970 5764 64972
rect 5533 64968 5764 64970
rect 5533 64912 5538 64968
rect 5594 64912 5764 64968
rect 5533 64910 5764 64912
rect 5533 64907 5599 64910
rect 5758 64908 5764 64910
rect 5828 64908 5834 64972
rect 5901 64834 5967 64837
rect 87270 64834 87276 64836
rect 5901 64832 8188 64834
rect 5901 64776 5906 64832
rect 5962 64776 8188 64832
rect 5901 64774 8188 64776
rect 46828 64774 48116 64834
rect 86940 64774 87276 64834
rect 5901 64771 5967 64774
rect 87270 64772 87276 64774
rect 87340 64772 87346 64836
rect 3062 64768 3378 64769
rect 0 64698 800 64728
rect 3062 64704 3068 64768
rect 3132 64704 3148 64768
rect 3212 64704 3228 64768
rect 3292 64704 3308 64768
rect 3372 64704 3378 64768
rect 3062 64703 3378 64704
rect 1301 64698 1367 64701
rect 0 64696 1367 64698
rect 0 64640 1306 64696
rect 1362 64640 1367 64696
rect 0 64638 1367 64640
rect 0 64608 800 64638
rect 1301 64635 1367 64638
rect 87597 64698 87663 64701
rect 89200 64698 90000 64728
rect 87597 64696 90000 64698
rect 87597 64640 87602 64696
rect 87658 64640 90000 64696
rect 87597 64638 90000 64640
rect 87597 64635 87663 64638
rect 89200 64608 90000 64638
rect 3798 64224 4114 64225
rect 3798 64160 3804 64224
rect 3868 64160 3884 64224
rect 3948 64160 3964 64224
rect 4028 64160 4044 64224
rect 4108 64160 4114 64224
rect 3798 64159 4114 64160
rect 3062 63680 3378 63681
rect 3062 63616 3068 63680
rect 3132 63616 3148 63680
rect 3212 63616 3228 63680
rect 3292 63616 3308 63680
rect 3372 63616 3378 63680
rect 3062 63615 3378 63616
rect 0 63338 800 63368
rect 1209 63338 1275 63341
rect 0 63336 1275 63338
rect 0 63280 1214 63336
rect 1270 63280 1275 63336
rect 0 63278 1275 63280
rect 0 63248 800 63278
rect 1209 63275 1275 63278
rect 8342 63205 8402 63444
rect 46828 63414 48116 63474
rect 86534 63412 86540 63476
rect 86604 63412 86610 63476
rect 88885 63338 88951 63341
rect 89200 63338 90000 63368
rect 88885 63336 90000 63338
rect 88885 63280 88890 63336
rect 88946 63280 90000 63336
rect 88885 63278 90000 63280
rect 88885 63275 88951 63278
rect 89200 63248 90000 63278
rect 8293 63200 8402 63205
rect 8293 63144 8298 63200
rect 8354 63144 8402 63200
rect 8293 63142 8402 63144
rect 8293 63139 8359 63142
rect 3798 63136 4114 63137
rect 3798 63072 3804 63136
rect 3868 63072 3884 63136
rect 3948 63072 3964 63136
rect 4028 63072 4044 63136
rect 4108 63072 4114 63136
rect 3798 63071 4114 63072
rect 3062 62592 3378 62593
rect 3062 62528 3068 62592
rect 3132 62528 3148 62592
rect 3212 62528 3228 62592
rect 3292 62528 3308 62592
rect 3372 62528 3378 62592
rect 3062 62527 3378 62528
rect 5901 62252 5967 62253
rect 5901 62248 5948 62252
rect 6012 62250 6018 62252
rect 5901 62192 5906 62248
rect 5901 62188 5948 62192
rect 6012 62190 6058 62250
rect 6012 62188 6018 62190
rect 5901 62187 5967 62188
rect 5533 62114 5599 62117
rect 5533 62112 8188 62114
rect 5533 62056 5538 62112
rect 5594 62056 8188 62112
rect 5533 62054 8188 62056
rect 46828 62054 48116 62114
rect 5533 62051 5599 62054
rect 3798 62048 4114 62049
rect 0 61978 800 62008
rect 3798 61984 3804 62048
rect 3868 61984 3884 62048
rect 3948 61984 3964 62048
rect 4028 61984 4044 62048
rect 4108 61984 4114 62048
rect 3798 61983 4114 61984
rect 1301 61978 1367 61981
rect 0 61976 1367 61978
rect 0 61920 1306 61976
rect 1362 61920 1367 61976
rect 0 61918 1367 61920
rect 0 61888 800 61918
rect 1301 61915 1367 61918
rect 86910 61570 86970 62084
rect 87689 61978 87755 61981
rect 89200 61978 90000 62008
rect 87689 61976 90000 61978
rect 87689 61920 87694 61976
rect 87750 61920 90000 61976
rect 87689 61918 90000 61920
rect 87689 61915 87755 61918
rect 89200 61888 90000 61918
rect 87045 61570 87111 61573
rect 86910 61568 87111 61570
rect 86910 61512 87050 61568
rect 87106 61512 87111 61568
rect 86910 61510 87111 61512
rect 87045 61507 87111 61510
rect 3062 61504 3378 61505
rect 3062 61440 3068 61504
rect 3132 61440 3148 61504
rect 3212 61440 3228 61504
rect 3292 61440 3308 61504
rect 3372 61440 3378 61504
rect 3062 61439 3378 61440
rect 0 61298 800 61328
rect 1301 61298 1367 61301
rect 0 61296 1367 61298
rect 0 61240 1306 61296
rect 1362 61240 1367 61296
rect 0 61238 1367 61240
rect 0 61208 800 61238
rect 1301 61235 1367 61238
rect 8293 61298 8359 61301
rect 8293 61296 8402 61298
rect 8293 61240 8298 61296
rect 8354 61240 8402 61296
rect 8293 61235 8402 61240
rect 3798 60960 4114 60961
rect 3798 60896 3804 60960
rect 3868 60896 3884 60960
rect 3948 60896 3964 60960
rect 4028 60896 4044 60960
rect 4108 60896 4114 60960
rect 3798 60895 4114 60896
rect 8342 60724 8402 61235
rect 46828 60694 48116 60754
rect 86902 60692 86908 60756
rect 86972 60692 86978 60756
rect 0 60618 800 60648
rect 88793 60618 88859 60621
rect 89200 60618 90000 60648
rect 0 60528 858 60618
rect 88793 60616 90000 60618
rect 88793 60560 88798 60616
rect 88854 60560 90000 60616
rect 88793 60558 90000 60560
rect 88793 60555 88859 60558
rect 89200 60528 90000 60558
rect 798 60485 858 60528
rect 798 60480 907 60485
rect 798 60424 846 60480
rect 902 60424 907 60480
rect 798 60422 907 60424
rect 841 60419 907 60422
rect 3062 60416 3378 60417
rect 3062 60352 3068 60416
rect 3132 60352 3148 60416
rect 3212 60352 3228 60416
rect 3292 60352 3308 60416
rect 3372 60352 3378 60416
rect 3062 60351 3378 60352
rect 0 59938 800 59968
rect 1209 59938 1275 59941
rect 0 59936 1275 59938
rect 0 59880 1214 59936
rect 1270 59880 1275 59936
rect 0 59878 1275 59880
rect 0 59848 800 59878
rect 1209 59875 1275 59878
rect 8293 59938 8359 59941
rect 8293 59936 8402 59938
rect 8293 59880 8298 59936
rect 8354 59880 8402 59936
rect 8293 59875 8402 59880
rect 3798 59872 4114 59873
rect 3798 59808 3804 59872
rect 3868 59808 3884 59872
rect 3948 59808 3964 59872
rect 4028 59808 4044 59872
rect 4108 59808 4114 59872
rect 3798 59807 4114 59808
rect 8342 59364 8402 59875
rect 87086 59394 87092 59396
rect 46828 59334 48116 59394
rect 86940 59334 87092 59394
rect 87086 59332 87092 59334
rect 87156 59394 87162 59396
rect 87454 59394 87460 59396
rect 87156 59334 87460 59394
rect 87156 59332 87162 59334
rect 87454 59332 87460 59334
rect 87524 59332 87530 59396
rect 3062 59328 3378 59329
rect 0 59258 800 59288
rect 3062 59264 3068 59328
rect 3132 59264 3148 59328
rect 3212 59264 3228 59328
rect 3292 59264 3308 59328
rect 3372 59264 3378 59328
rect 3062 59263 3378 59264
rect 87781 59258 87847 59261
rect 89200 59258 90000 59288
rect 0 59168 858 59258
rect 87781 59256 90000 59258
rect 87781 59200 87786 59256
rect 87842 59200 90000 59256
rect 87781 59198 90000 59200
rect 87781 59195 87847 59198
rect 89200 59168 90000 59198
rect 798 59125 858 59168
rect 798 59120 907 59125
rect 798 59064 846 59120
rect 902 59064 907 59120
rect 798 59062 907 59064
rect 841 59059 907 59062
rect 3798 58784 4114 58785
rect 3798 58720 3804 58784
rect 3868 58720 3884 58784
rect 3948 58720 3964 58784
rect 4028 58720 4044 58784
rect 4108 58720 4114 58784
rect 3798 58719 4114 58720
rect 0 58578 800 58608
rect 1301 58578 1367 58581
rect 0 58576 1367 58578
rect 0 58520 1306 58576
rect 1362 58520 1367 58576
rect 0 58518 1367 58520
rect 0 58488 800 58518
rect 1301 58515 1367 58518
rect 8293 58578 8359 58581
rect 8293 58576 8402 58578
rect 8293 58520 8298 58576
rect 8354 58520 8402 58576
rect 8293 58515 8402 58520
rect 3062 58240 3378 58241
rect 3062 58176 3068 58240
rect 3132 58176 3148 58240
rect 3212 58176 3228 58240
rect 3292 58176 3308 58240
rect 3372 58176 3378 58240
rect 3062 58175 3378 58176
rect 8342 58004 8402 58515
rect 87137 58034 87203 58037
rect 46828 57974 48116 58034
rect 86940 58032 87203 58034
rect 86940 57976 87142 58032
rect 87198 57976 87203 58032
rect 86940 57974 87203 57976
rect 87137 57971 87203 57974
rect 0 57898 800 57928
rect 88609 57898 88675 57901
rect 89200 57898 90000 57928
rect 0 57808 858 57898
rect 88609 57896 90000 57898
rect 88609 57840 88614 57896
rect 88670 57840 90000 57896
rect 88609 57838 90000 57840
rect 88609 57835 88675 57838
rect 89200 57808 90000 57838
rect 798 57765 858 57808
rect 798 57760 907 57765
rect 798 57704 846 57760
rect 902 57704 907 57760
rect 798 57702 907 57704
rect 841 57699 907 57702
rect 3798 57696 4114 57697
rect 3798 57632 3804 57696
rect 3868 57632 3884 57696
rect 3948 57632 3964 57696
rect 4028 57632 4044 57696
rect 4108 57632 4114 57696
rect 3798 57631 4114 57632
rect 0 57218 800 57248
rect 1301 57218 1367 57221
rect 0 57216 1367 57218
rect 0 57160 1306 57216
rect 1362 57160 1367 57216
rect 0 57158 1367 57160
rect 0 57128 800 57158
rect 1301 57155 1367 57158
rect 8293 57218 8359 57221
rect 86953 57218 87019 57221
rect 8293 57216 8402 57218
rect 8293 57160 8298 57216
rect 8354 57160 8402 57216
rect 8293 57155 8402 57160
rect 3062 57152 3378 57153
rect 3062 57088 3068 57152
rect 3132 57088 3148 57152
rect 3212 57088 3228 57152
rect 3292 57088 3308 57152
rect 3372 57088 3378 57152
rect 3062 57087 3378 57088
rect 8342 56644 8402 57155
rect 86910 57216 87019 57218
rect 86910 57160 86958 57216
rect 87014 57160 87019 57216
rect 86910 57155 87019 57160
rect 86910 56674 86970 57155
rect 87413 56674 87479 56677
rect 46828 56614 48116 56674
rect 86910 56672 87479 56674
rect 86910 56644 87418 56672
rect 86940 56616 87418 56644
rect 87474 56616 87479 56672
rect 86940 56614 87479 56616
rect 87413 56611 87479 56614
rect 3798 56608 4114 56609
rect 0 56538 800 56568
rect 3798 56544 3804 56608
rect 3868 56544 3884 56608
rect 3948 56544 3964 56608
rect 4028 56544 4044 56608
rect 4108 56544 4114 56608
rect 3798 56543 4114 56544
rect 88701 56538 88767 56541
rect 89200 56538 90000 56568
rect 0 56448 858 56538
rect 88701 56536 90000 56538
rect 88701 56480 88706 56536
rect 88762 56480 90000 56536
rect 88701 56478 90000 56480
rect 88701 56475 88767 56478
rect 89200 56448 90000 56478
rect 798 56405 858 56448
rect 798 56400 907 56405
rect 798 56344 846 56400
rect 902 56344 907 56400
rect 798 56342 907 56344
rect 841 56339 907 56342
rect 3062 56064 3378 56065
rect 3062 56000 3068 56064
rect 3132 56000 3148 56064
rect 3212 56000 3228 56064
rect 3292 56000 3308 56064
rect 3372 56000 3378 56064
rect 3062 55999 3378 56000
rect 0 55858 800 55888
rect 1301 55858 1367 55861
rect 0 55856 1367 55858
rect 0 55800 1306 55856
rect 1362 55800 1367 55856
rect 0 55798 1367 55800
rect 0 55768 800 55798
rect 1301 55795 1367 55798
rect 8293 55858 8359 55861
rect 8293 55856 8402 55858
rect 8293 55800 8298 55856
rect 8354 55800 8402 55856
rect 8293 55795 8402 55800
rect 3798 55520 4114 55521
rect 3798 55456 3804 55520
rect 3868 55456 3884 55520
rect 3948 55456 3964 55520
rect 4028 55456 4044 55520
rect 4108 55456 4114 55520
rect 3798 55455 4114 55456
rect 8342 55284 8402 55795
rect 46828 55254 48116 55314
rect 86902 55252 86908 55316
rect 86972 55252 86978 55316
rect 0 55178 800 55208
rect 88517 55178 88583 55181
rect 89200 55178 90000 55208
rect 0 55088 858 55178
rect 88517 55176 90000 55178
rect 88517 55120 88522 55176
rect 88578 55120 90000 55176
rect 88517 55118 90000 55120
rect 88517 55115 88583 55118
rect 89200 55088 90000 55118
rect 798 55045 858 55088
rect 798 55040 907 55045
rect 798 54984 846 55040
rect 902 54984 907 55040
rect 798 54982 907 54984
rect 841 54979 907 54982
rect 3062 54976 3378 54977
rect 3062 54912 3068 54976
rect 3132 54912 3148 54976
rect 3212 54912 3228 54976
rect 3292 54912 3308 54976
rect 3372 54912 3378 54976
rect 3062 54911 3378 54912
rect 0 54498 800 54528
rect 1209 54498 1275 54501
rect 0 54496 1275 54498
rect 0 54440 1214 54496
rect 1270 54440 1275 54496
rect 0 54438 1275 54440
rect 0 54408 800 54438
rect 1209 54435 1275 54438
rect 8293 54498 8359 54501
rect 8293 54496 8402 54498
rect 8293 54440 8298 54496
rect 8354 54440 8402 54496
rect 8293 54435 8402 54440
rect 3798 54432 4114 54433
rect 3798 54368 3804 54432
rect 3868 54368 3884 54432
rect 3948 54368 3964 54432
rect 4028 54368 4044 54432
rect 4108 54368 4114 54432
rect 3798 54367 4114 54368
rect 8342 53924 8402 54435
rect 87321 53954 87387 53957
rect 46828 53894 48116 53954
rect 86940 53952 87387 53954
rect 86940 53896 87326 53952
rect 87382 53896 87387 53952
rect 86940 53894 87387 53896
rect 87321 53891 87387 53894
rect 3062 53888 3378 53889
rect 0 53818 800 53848
rect 3062 53824 3068 53888
rect 3132 53824 3148 53888
rect 3212 53824 3228 53888
rect 3292 53824 3308 53888
rect 3372 53824 3378 53888
rect 3062 53823 3378 53824
rect 88333 53818 88399 53821
rect 89200 53818 90000 53848
rect 0 53728 858 53818
rect 88333 53816 90000 53818
rect 88333 53760 88338 53816
rect 88394 53760 90000 53816
rect 88333 53758 90000 53760
rect 88333 53755 88399 53758
rect 89200 53728 90000 53758
rect 798 53685 858 53728
rect 798 53680 907 53685
rect 798 53624 846 53680
rect 902 53624 907 53680
rect 798 53622 907 53624
rect 841 53619 907 53622
rect 3798 53344 4114 53345
rect 3798 53280 3804 53344
rect 3868 53280 3884 53344
rect 3948 53280 3964 53344
rect 4028 53280 4044 53344
rect 4108 53280 4114 53344
rect 3798 53279 4114 53280
rect 0 53138 800 53168
rect 1301 53138 1367 53141
rect 0 53136 1367 53138
rect 0 53080 1306 53136
rect 1362 53080 1367 53136
rect 0 53078 1367 53080
rect 0 53048 800 53078
rect 1301 53075 1367 53078
rect 8293 53138 8359 53141
rect 8293 53136 8402 53138
rect 8293 53080 8298 53136
rect 8354 53080 8402 53136
rect 8293 53075 8402 53080
rect 3062 52800 3378 52801
rect 3062 52736 3068 52800
rect 3132 52736 3148 52800
rect 3212 52736 3228 52800
rect 3292 52736 3308 52800
rect 3372 52736 3378 52800
rect 3062 52735 3378 52736
rect 8342 52564 8402 53075
rect 87229 52594 87295 52597
rect 46828 52534 48116 52594
rect 86940 52592 87295 52594
rect 86940 52536 87234 52592
rect 87290 52536 87295 52592
rect 86940 52534 87295 52536
rect 87229 52531 87295 52534
rect 0 52458 800 52488
rect 88425 52458 88491 52461
rect 89200 52458 90000 52488
rect 0 52368 858 52458
rect 88425 52456 90000 52458
rect 88425 52400 88430 52456
rect 88486 52400 90000 52456
rect 88425 52398 90000 52400
rect 88425 52395 88491 52398
rect 89200 52368 90000 52398
rect 798 52325 858 52368
rect 798 52320 907 52325
rect 798 52264 846 52320
rect 902 52264 907 52320
rect 798 52262 907 52264
rect 841 52259 907 52262
rect 3798 52256 4114 52257
rect 3798 52192 3804 52256
rect 3868 52192 3884 52256
rect 3948 52192 3964 52256
rect 4028 52192 4044 52256
rect 4108 52192 4114 52256
rect 3798 52191 4114 52192
rect 841 51914 907 51917
rect 798 51912 907 51914
rect 798 51856 846 51912
rect 902 51856 907 51912
rect 798 51851 907 51856
rect 798 51808 858 51851
rect 0 51718 858 51808
rect 0 51688 800 51718
rect 3062 51712 3378 51713
rect 3062 51648 3068 51712
rect 3132 51648 3148 51712
rect 3212 51648 3228 51712
rect 3292 51648 3308 51712
rect 3372 51648 3378 51712
rect 3062 51647 3378 51648
rect 1577 51370 1643 51373
rect 1577 51368 8218 51370
rect 1577 51312 1582 51368
rect 1638 51312 8218 51368
rect 1577 51310 8218 51312
rect 1577 51307 1643 51310
rect 8158 51204 8218 51310
rect 46828 51174 48116 51234
rect 3798 51168 4114 51169
rect 0 51098 800 51128
rect 3798 51104 3804 51168
rect 3868 51104 3884 51168
rect 3948 51104 3964 51168
rect 4028 51104 4044 51168
rect 4108 51104 4114 51168
rect 3798 51103 4114 51104
rect 1025 51098 1091 51101
rect 0 51090 858 51098
rect 982 51096 1091 51098
rect 982 51090 1030 51096
rect 0 51040 1030 51090
rect 1086 51040 1091 51096
rect 0 51035 1091 51040
rect 0 51030 1042 51035
rect 0 51008 800 51030
rect 86910 50962 86970 51204
rect 87137 51098 87203 51101
rect 89200 51098 90000 51128
rect 87137 51096 90000 51098
rect 87137 51040 87142 51096
rect 87198 51040 90000 51096
rect 87137 51038 90000 51040
rect 87137 51035 87203 51038
rect 89200 51008 90000 51038
rect 87137 50962 87203 50965
rect 86910 50960 87203 50962
rect 86910 50904 87142 50960
rect 87198 50904 87203 50960
rect 86910 50902 87203 50904
rect 87137 50899 87203 50902
rect 5758 50764 5764 50828
rect 5828 50826 5834 50828
rect 87597 50826 87663 50829
rect 5828 50824 87663 50826
rect 5828 50768 87602 50824
rect 87658 50768 87663 50824
rect 5828 50766 87663 50768
rect 5828 50764 5834 50766
rect 87597 50763 87663 50766
rect 5574 50628 5580 50692
rect 5644 50690 5650 50692
rect 85246 50690 85252 50692
rect 5644 50630 85252 50690
rect 5644 50628 5650 50630
rect 85246 50628 85252 50630
rect 85316 50628 85322 50692
rect 87045 50690 87111 50693
rect 85438 50688 87111 50690
rect 85438 50632 87050 50688
rect 87106 50632 87111 50688
rect 85438 50630 87111 50632
rect 3062 50624 3378 50625
rect 3062 50560 3068 50624
rect 3132 50560 3148 50624
rect 3212 50560 3228 50624
rect 3292 50560 3308 50624
rect 3372 50560 3378 50624
rect 3062 50559 3378 50560
rect 1393 50554 1459 50557
rect 798 50552 1459 50554
rect 798 50496 1398 50552
rect 1454 50496 1459 50552
rect 798 50494 1459 50496
rect 798 50448 858 50494
rect 1393 50491 1459 50494
rect 5441 50554 5507 50557
rect 46749 50554 46815 50557
rect 85438 50554 85498 50630
rect 87045 50627 87111 50630
rect 5441 50552 85498 50554
rect 5441 50496 5446 50552
rect 5502 50496 46754 50552
rect 46810 50496 85498 50552
rect 5441 50494 85498 50496
rect 85573 50554 85639 50557
rect 86350 50554 86356 50556
rect 85573 50552 86356 50554
rect 85573 50496 85578 50552
rect 85634 50496 86356 50552
rect 85573 50494 86356 50496
rect 5441 50491 5507 50494
rect 46749 50491 46815 50494
rect 85573 50491 85639 50494
rect 86350 50492 86356 50494
rect 86420 50492 86426 50556
rect 0 50358 858 50448
rect 46749 50418 46815 50421
rect 89200 50418 90000 50448
rect 46749 50416 90000 50418
rect 46749 50360 46754 50416
rect 46810 50360 90000 50416
rect 46749 50358 90000 50360
rect 0 50328 800 50358
rect 46749 50355 46815 50358
rect 89200 50328 90000 50358
rect 4797 50282 4863 50285
rect 46841 50282 46907 50285
rect 4797 50280 46907 50282
rect 4797 50224 4802 50280
rect 4858 50224 46846 50280
rect 46902 50224 46907 50280
rect 4797 50222 46907 50224
rect 4797 50219 4863 50222
rect 46841 50219 46907 50222
rect 47710 50220 47716 50284
rect 47780 50282 47786 50284
rect 86953 50282 87019 50285
rect 47780 50280 87019 50282
rect 47780 50224 86958 50280
rect 87014 50224 87019 50280
rect 47780 50222 87019 50224
rect 47780 50220 47786 50222
rect 86953 50219 87019 50222
rect 85246 50084 85252 50148
rect 85316 50146 85322 50148
rect 89345 50146 89411 50149
rect 85316 50144 89411 50146
rect 85316 50088 89350 50144
rect 89406 50088 89411 50144
rect 85316 50086 89411 50088
rect 85316 50084 85322 50086
rect 89345 50083 89411 50086
rect 3798 50080 4114 50081
rect 3798 50016 3804 50080
rect 3868 50016 3884 50080
rect 3948 50016 3964 50080
rect 4028 50016 4044 50080
rect 4108 50016 4114 50080
rect 3798 50015 4114 50016
rect 0 49740 800 49768
rect 0 49676 796 49740
rect 860 49676 866 49740
rect 8385 49738 8451 49741
rect 47209 49738 47275 49741
rect 85573 49738 85639 49741
rect 8385 49736 85639 49738
rect 8385 49680 8390 49736
rect 8446 49680 47214 49736
rect 47270 49680 85578 49736
rect 85634 49680 85639 49736
rect 8385 49678 85639 49680
rect 0 49648 800 49676
rect 8385 49675 8451 49678
rect 47209 49675 47275 49678
rect 85573 49675 85639 49678
rect 4981 49602 5047 49605
rect 87086 49602 87092 49604
rect 4981 49600 87092 49602
rect 4981 49544 4986 49600
rect 5042 49544 87092 49600
rect 4981 49542 87092 49544
rect 4981 49539 5047 49542
rect 87086 49540 87092 49542
rect 87156 49540 87162 49604
rect 3062 49536 3378 49537
rect 3062 49472 3068 49536
rect 3132 49472 3148 49536
rect 3212 49472 3228 49536
rect 3292 49472 3308 49536
rect 3372 49472 3378 49536
rect 3062 49471 3378 49472
rect 790 49404 796 49468
rect 860 49466 866 49468
rect 1393 49466 1459 49469
rect 860 49464 1459 49466
rect 860 49408 1398 49464
rect 1454 49408 1459 49464
rect 860 49406 1459 49408
rect 860 49404 866 49406
rect 1393 49403 1459 49406
rect 5942 49404 5948 49468
rect 6012 49466 6018 49468
rect 87689 49466 87755 49469
rect 6012 49464 87755 49466
rect 6012 49408 87694 49464
rect 87750 49408 87755 49464
rect 6012 49406 87755 49408
rect 6012 49404 6018 49406
rect 87689 49403 87755 49406
rect 790 49268 796 49332
rect 860 49330 866 49332
rect 1393 49330 1459 49333
rect 860 49328 1459 49330
rect 860 49272 1398 49328
rect 1454 49272 1459 49328
rect 860 49270 1459 49272
rect 860 49268 866 49270
rect 1393 49267 1459 49270
rect 4521 49330 4587 49333
rect 40677 49330 40743 49333
rect 4521 49328 40743 49330
rect 4521 49272 4526 49328
rect 4582 49272 40682 49328
rect 40738 49272 40743 49328
rect 4521 49270 40743 49272
rect 4521 49267 4587 49270
rect 40677 49267 40743 49270
rect 48221 49330 48287 49333
rect 87229 49330 87295 49333
rect 48221 49328 87295 49330
rect 48221 49272 48226 49328
rect 48282 49272 87234 49328
rect 87290 49272 87295 49328
rect 48221 49270 87295 49272
rect 48221 49267 48287 49270
rect 87229 49267 87295 49270
rect 4705 49194 4771 49197
rect 48078 49194 48084 49196
rect 4705 49192 48084 49194
rect 4705 49136 4710 49192
rect 4766 49136 48084 49192
rect 4705 49134 48084 49136
rect 4705 49131 4771 49134
rect 48078 49132 48084 49134
rect 48148 49194 48154 49196
rect 86902 49194 86908 49196
rect 48148 49134 86908 49194
rect 48148 49132 48154 49134
rect 86902 49132 86908 49134
rect 86972 49132 86978 49196
rect 0 49060 800 49088
rect 0 48996 796 49060
rect 860 48996 866 49060
rect 5073 49058 5139 49061
rect 47853 49058 47919 49061
rect 87321 49058 87387 49061
rect 5073 49056 87387 49058
rect 5073 49000 5078 49056
rect 5134 49000 47858 49056
rect 47914 49000 87326 49056
rect 87382 49000 87387 49056
rect 5073 48998 87387 49000
rect 0 48968 800 48996
rect 5073 48995 5139 48998
rect 47853 48995 47919 48998
rect 87321 48995 87387 48998
rect 3798 48992 4114 48993
rect 3798 48928 3804 48992
rect 3868 48928 3884 48992
rect 3948 48928 3964 48992
rect 4028 48928 4044 48992
rect 4108 48928 4114 48992
rect 3798 48927 4114 48928
rect 40677 48922 40743 48925
rect 47526 48922 47532 48924
rect 40677 48920 47532 48922
rect 40677 48864 40682 48920
rect 40738 48864 47532 48920
rect 40677 48862 47532 48864
rect 40677 48859 40743 48862
rect 47526 48860 47532 48862
rect 47596 48922 47602 48924
rect 86534 48922 86540 48924
rect 47596 48862 86540 48922
rect 47596 48860 47602 48862
rect 86534 48860 86540 48862
rect 86604 48860 86610 48924
rect 3062 48448 3378 48449
rect 0 48378 800 48408
rect 3062 48384 3068 48448
rect 3132 48384 3148 48448
rect 3212 48384 3228 48448
rect 3292 48384 3308 48448
rect 3372 48384 3378 48448
rect 3062 48383 3378 48384
rect 1301 48378 1367 48381
rect 0 48376 1367 48378
rect 0 48320 1306 48376
rect 1362 48320 1367 48376
rect 0 48318 1367 48320
rect 0 48288 800 48318
rect 1301 48315 1367 48318
rect 4705 48378 4771 48381
rect 48078 48378 48084 48380
rect 4705 48376 48084 48378
rect 4705 48320 4710 48376
rect 4766 48320 48084 48376
rect 4705 48318 48084 48320
rect 4705 48315 4771 48318
rect 48078 48316 48084 48318
rect 48148 48378 48154 48380
rect 87638 48378 87644 48380
rect 48148 48318 87644 48378
rect 48148 48316 48154 48318
rect 87638 48316 87644 48318
rect 87708 48316 87714 48380
rect 4981 48106 5047 48109
rect 47710 48106 47716 48108
rect 4981 48104 47716 48106
rect 4981 48048 4986 48104
rect 5042 48048 47716 48104
rect 4981 48046 47716 48048
rect 4981 48043 5047 48046
rect 47710 48044 47716 48046
rect 47780 48106 47786 48108
rect 48262 48106 48268 48108
rect 47780 48046 48268 48106
rect 47780 48044 47786 48046
rect 48262 48044 48268 48046
rect 48332 48044 48338 48108
rect 790 47908 796 47972
rect 860 47970 866 47972
rect 1393 47970 1459 47973
rect 860 47968 1459 47970
rect 860 47912 1398 47968
rect 1454 47912 1459 47968
rect 860 47910 1459 47912
rect 860 47908 866 47910
rect 1393 47907 1459 47910
rect 4889 47970 4955 47973
rect 88057 47970 88123 47973
rect 4889 47968 88123 47970
rect 4889 47912 4894 47968
rect 4950 47912 88062 47968
rect 88118 47912 88123 47968
rect 4889 47910 88123 47912
rect 4889 47907 4955 47910
rect 88057 47907 88123 47910
rect 3798 47904 4114 47905
rect 3798 47840 3804 47904
rect 3868 47840 3884 47904
rect 3948 47840 3964 47904
rect 4028 47840 4044 47904
rect 4108 47840 4114 47904
rect 3798 47839 4114 47840
rect 4613 47834 4679 47837
rect 47894 47834 47900 47836
rect 4613 47832 47900 47834
rect 4613 47776 4618 47832
rect 4674 47776 47900 47832
rect 4613 47774 47900 47776
rect 4613 47771 4679 47774
rect 47894 47772 47900 47774
rect 47964 47834 47970 47836
rect 87505 47834 87571 47837
rect 47964 47832 87571 47834
rect 47964 47776 87510 47832
rect 87566 47776 87571 47832
rect 47964 47774 87571 47776
rect 47964 47772 47970 47774
rect 87505 47771 87571 47774
rect 0 47700 800 47728
rect 0 47636 796 47700
rect 860 47636 866 47700
rect 6361 47698 6427 47701
rect 6361 47696 26250 47698
rect 6361 47640 6366 47696
rect 6422 47640 26250 47696
rect 6361 47638 26250 47640
rect 0 47608 800 47636
rect 6361 47635 6427 47638
rect 26190 47426 26250 47638
rect 48262 47636 48268 47700
rect 48332 47698 48338 47700
rect 87045 47698 87111 47701
rect 48332 47696 87111 47698
rect 48332 47640 87050 47696
rect 87106 47640 87111 47696
rect 48332 47638 87111 47640
rect 48332 47636 48338 47638
rect 87045 47635 87111 47638
rect 46841 47562 46907 47565
rect 87270 47562 87276 47564
rect 46841 47560 87276 47562
rect 46841 47504 46846 47560
rect 46902 47504 87276 47560
rect 46841 47502 87276 47504
rect 46841 47499 46907 47502
rect 87270 47500 87276 47502
rect 87340 47500 87346 47564
rect 46749 47426 46815 47429
rect 87229 47426 87295 47429
rect 26190 47424 87295 47426
rect 26190 47368 46754 47424
rect 46810 47368 87234 47424
rect 87290 47368 87295 47424
rect 26190 47366 87295 47368
rect 46749 47363 46815 47366
rect 87229 47363 87295 47366
rect 3062 47360 3378 47361
rect 3062 47296 3068 47360
rect 3132 47296 3148 47360
rect 3212 47296 3228 47360
rect 3292 47296 3308 47360
rect 3372 47296 3378 47360
rect 3062 47295 3378 47296
rect 7557 47290 7623 47293
rect 88885 47290 88951 47293
rect 7557 47288 88951 47290
rect 7557 47232 7562 47288
rect 7618 47232 88890 47288
rect 88946 47232 88951 47288
rect 7557 47230 88951 47232
rect 7557 47227 7623 47230
rect 88885 47227 88951 47230
rect 5349 47154 5415 47157
rect 87086 47154 87092 47156
rect 5349 47152 87092 47154
rect 5349 47096 5354 47152
rect 5410 47096 87092 47152
rect 5349 47094 87092 47096
rect 5349 47091 5415 47094
rect 87086 47092 87092 47094
rect 87156 47092 87162 47156
rect 0 47018 800 47048
rect 1393 47018 1459 47021
rect 0 47016 1459 47018
rect 0 46960 1398 47016
rect 1454 46960 1459 47016
rect 0 46958 1459 46960
rect 0 46928 800 46958
rect 1393 46955 1459 46958
rect 5206 46956 5212 47020
rect 5276 47018 5282 47020
rect 11237 47018 11303 47021
rect 5276 47016 11303 47018
rect 5276 46960 11242 47016
rect 11298 46960 11303 47016
rect 5276 46958 11303 46960
rect 5276 46956 5282 46958
rect 11237 46955 11303 46958
rect 3798 46816 4114 46817
rect 3798 46752 3804 46816
rect 3868 46752 3884 46816
rect 3948 46752 3964 46816
rect 4028 46752 4044 46816
rect 4108 46752 4114 46816
rect 3798 46751 4114 46752
rect 47393 46610 47459 46613
rect 51073 46610 51139 46613
rect 87137 46610 87203 46613
rect 47393 46608 51139 46610
rect 47393 46552 47398 46608
rect 47454 46552 51078 46608
rect 51134 46552 51139 46608
rect 47393 46550 51139 46552
rect 47393 46547 47459 46550
rect 51073 46547 51139 46550
rect 64830 46608 87203 46610
rect 64830 46552 87142 46608
rect 87198 46552 87203 46608
rect 64830 46550 87203 46552
rect 5257 46474 5323 46477
rect 64830 46474 64890 46550
rect 87137 46547 87203 46550
rect 5257 46472 64890 46474
rect 5257 46416 5262 46472
rect 5318 46416 64890 46472
rect 5257 46414 64890 46416
rect 85573 46474 85639 46477
rect 85573 46472 86418 46474
rect 85573 46416 85578 46472
rect 85634 46416 86418 46472
rect 85573 46414 86418 46416
rect 5257 46411 5323 46414
rect 85573 46411 85639 46414
rect 0 46338 800 46368
rect 1393 46338 1459 46341
rect 0 46336 1459 46338
rect 0 46280 1398 46336
rect 1454 46280 1459 46336
rect 0 46278 1459 46280
rect 0 46248 800 46278
rect 1393 46275 1459 46278
rect 3062 46272 3378 46273
rect 3062 46208 3068 46272
rect 3132 46208 3148 46272
rect 3212 46208 3228 46272
rect 3292 46208 3308 46272
rect 3372 46208 3378 46272
rect 3062 46207 3378 46208
rect 8293 46066 8359 46069
rect 8293 46064 8402 46066
rect 8293 46008 8298 46064
rect 8354 46008 8402 46064
rect 8293 46003 8402 46008
rect 8342 45900 8402 46003
rect 46828 45870 48116 45930
rect 86358 45900 86418 46414
rect 1485 45794 1551 45797
rect 798 45792 1551 45794
rect 798 45736 1490 45792
rect 1546 45736 1551 45792
rect 798 45734 1551 45736
rect 798 45688 858 45734
rect 1485 45731 1551 45734
rect 0 45598 858 45688
rect 3798 45728 4114 45729
rect 3798 45664 3804 45728
rect 3868 45664 3884 45728
rect 3948 45664 3964 45728
rect 4028 45664 4044 45728
rect 4108 45664 4114 45728
rect 3798 45663 4114 45664
rect 88333 45658 88399 45661
rect 89200 45658 90000 45688
rect 88333 45656 90000 45658
rect 88333 45600 88338 45656
rect 88394 45600 90000 45656
rect 88333 45598 90000 45600
rect 0 45568 800 45598
rect 88333 45595 88399 45598
rect 89200 45568 90000 45598
rect 3062 45184 3378 45185
rect 3062 45120 3068 45184
rect 3132 45120 3148 45184
rect 3212 45120 3228 45184
rect 3292 45120 3308 45184
rect 3372 45120 3378 45184
rect 3062 45119 3378 45120
rect 1393 45114 1459 45117
rect 798 45112 1459 45114
rect 798 45056 1398 45112
rect 1454 45056 1459 45112
rect 798 45054 1459 45056
rect 798 45008 858 45054
rect 1393 45051 1459 45054
rect 0 44918 858 45008
rect 0 44888 800 44918
rect 3798 44640 4114 44641
rect 3798 44576 3804 44640
rect 3868 44576 3884 44640
rect 3948 44576 3964 44640
rect 4028 44576 4044 44640
rect 4108 44576 4114 44640
rect 3798 44575 4114 44576
rect 0 44298 800 44328
rect 8342 44301 8402 44540
rect 46828 44510 48116 44570
rect 1485 44298 1551 44301
rect 0 44296 1551 44298
rect 0 44240 1490 44296
rect 1546 44240 1551 44296
rect 0 44238 1551 44240
rect 0 44208 800 44238
rect 1485 44235 1551 44238
rect 8293 44296 8402 44301
rect 8293 44240 8298 44296
rect 8354 44240 8402 44296
rect 8293 44238 8402 44240
rect 86910 44301 86970 44540
rect 86910 44296 87019 44301
rect 86910 44240 86958 44296
rect 87014 44240 87019 44296
rect 86910 44238 87019 44240
rect 8293 44235 8359 44238
rect 86953 44235 87019 44238
rect 88333 44298 88399 44301
rect 89200 44298 90000 44328
rect 88333 44296 90000 44298
rect 88333 44240 88338 44296
rect 88394 44240 90000 44296
rect 88333 44238 90000 44240
rect 88333 44235 88399 44238
rect 89200 44208 90000 44238
rect 3062 44096 3378 44097
rect 3062 44032 3068 44096
rect 3132 44032 3148 44096
rect 3212 44032 3228 44096
rect 3292 44032 3308 44096
rect 3372 44032 3378 44096
rect 3062 44031 3378 44032
rect 0 43618 800 43648
rect 1209 43618 1275 43621
rect 0 43616 1275 43618
rect 0 43560 1214 43616
rect 1270 43560 1275 43616
rect 0 43558 1275 43560
rect 0 43528 800 43558
rect 1209 43555 1275 43558
rect 3798 43552 4114 43553
rect 3798 43488 3804 43552
rect 3868 43488 3884 43552
rect 3948 43488 3964 43552
rect 4028 43488 4044 43552
rect 4108 43488 4114 43552
rect 3798 43487 4114 43488
rect 8293 43346 8359 43349
rect 86677 43346 86743 43349
rect 8293 43344 8402 43346
rect 8293 43288 8298 43344
rect 8354 43288 8402 43344
rect 8293 43283 8402 43288
rect 86677 43344 86786 43346
rect 86677 43288 86682 43344
rect 86738 43288 86786 43344
rect 86677 43283 86786 43288
rect 8342 43180 8402 43283
rect 86726 43210 86786 43283
rect 87413 43210 87479 43213
rect 46828 43150 48116 43210
rect 86726 43208 87479 43210
rect 86726 43180 87418 43208
rect 86756 43152 87418 43180
rect 87474 43152 87479 43208
rect 86756 43150 87479 43152
rect 87413 43147 87479 43150
rect 1485 43074 1551 43077
rect 798 43072 1551 43074
rect 798 43016 1490 43072
rect 1546 43016 1551 43072
rect 798 43014 1551 43016
rect 798 42968 858 43014
rect 1485 43011 1551 43014
rect 0 42878 858 42968
rect 3062 43008 3378 43009
rect 3062 42944 3068 43008
rect 3132 42944 3148 43008
rect 3212 42944 3228 43008
rect 3292 42944 3308 43008
rect 3372 42944 3378 43008
rect 3062 42943 3378 42944
rect 88517 42938 88583 42941
rect 89200 42938 90000 42968
rect 88517 42936 90000 42938
rect 88517 42880 88522 42936
rect 88578 42880 90000 42936
rect 88517 42878 90000 42880
rect 0 42848 800 42878
rect 88517 42875 88583 42878
rect 89200 42848 90000 42878
rect 3798 42464 4114 42465
rect 3798 42400 3804 42464
rect 3868 42400 3884 42464
rect 3948 42400 3964 42464
rect 4028 42400 4044 42464
rect 4108 42400 4114 42464
rect 3798 42399 4114 42400
rect 86861 41986 86927 41989
rect 86861 41984 86970 41986
rect 86861 41928 86866 41984
rect 86922 41928 86970 41984
rect 86861 41923 86970 41928
rect 3062 41920 3378 41921
rect 3062 41856 3068 41920
rect 3132 41856 3148 41920
rect 3212 41856 3228 41920
rect 3292 41856 3308 41920
rect 3372 41856 3378 41920
rect 3062 41855 3378 41856
rect 86910 41850 86970 41923
rect 88333 41850 88399 41853
rect 0 41578 800 41608
rect 8342 41581 8402 41820
rect 46828 41790 48116 41850
rect 86910 41848 88399 41850
rect 86910 41820 88338 41848
rect 86940 41792 88338 41820
rect 88394 41792 88399 41848
rect 86940 41790 88399 41792
rect 88333 41787 88399 41790
rect 1485 41578 1551 41581
rect 0 41576 1551 41578
rect 0 41520 1490 41576
rect 1546 41520 1551 41576
rect 0 41518 1551 41520
rect 0 41488 800 41518
rect 1485 41515 1551 41518
rect 8293 41576 8402 41581
rect 8293 41520 8298 41576
rect 8354 41520 8402 41576
rect 8293 41518 8402 41520
rect 88701 41578 88767 41581
rect 89200 41578 90000 41608
rect 88701 41576 90000 41578
rect 88701 41520 88706 41576
rect 88762 41520 90000 41576
rect 88701 41518 90000 41520
rect 8293 41515 8359 41518
rect 88701 41515 88767 41518
rect 89200 41488 90000 41518
rect 3798 41376 4114 41377
rect 3798 41312 3804 41376
rect 3868 41312 3884 41376
rect 3948 41312 3964 41376
rect 4028 41312 4044 41376
rect 4108 41312 4114 41376
rect 3798 41311 4114 41312
rect 3062 40832 3378 40833
rect 3062 40768 3068 40832
rect 3132 40768 3148 40832
rect 3212 40768 3228 40832
rect 3292 40768 3308 40832
rect 3372 40768 3378 40832
rect 3062 40767 3378 40768
rect 87270 40700 87276 40764
rect 87340 40762 87346 40764
rect 87873 40762 87939 40765
rect 87340 40760 87939 40762
rect 87340 40704 87878 40760
rect 87934 40704 87939 40760
rect 87340 40702 87939 40704
rect 87340 40700 87346 40702
rect 87873 40699 87939 40702
rect 8293 40626 8359 40629
rect 8293 40624 8402 40626
rect 8293 40568 8298 40624
rect 8354 40568 8402 40624
rect 8293 40563 8402 40568
rect 8342 40460 8402 40563
rect 87270 40490 87276 40492
rect 46828 40430 48116 40490
rect 86940 40430 87276 40490
rect 87270 40428 87276 40430
rect 87340 40428 87346 40492
rect 841 40354 907 40357
rect 798 40352 907 40354
rect 798 40296 846 40352
rect 902 40296 907 40352
rect 798 40291 907 40296
rect 798 40248 858 40291
rect 0 40158 858 40248
rect 3798 40288 4114 40289
rect 3798 40224 3804 40288
rect 3868 40224 3884 40288
rect 3948 40224 3964 40288
rect 4028 40224 4044 40288
rect 4108 40224 4114 40288
rect 3798 40223 4114 40224
rect 88057 40218 88123 40221
rect 89200 40218 90000 40248
rect 88057 40216 90000 40218
rect 88057 40160 88062 40216
rect 88118 40160 90000 40216
rect 88057 40158 90000 40160
rect 0 40128 800 40158
rect 88057 40155 88123 40158
rect 89200 40128 90000 40158
rect 3062 39744 3378 39745
rect 3062 39680 3068 39744
rect 3132 39680 3148 39744
rect 3212 39680 3228 39744
rect 3292 39680 3308 39744
rect 3372 39680 3378 39744
rect 3062 39679 3378 39680
rect 87045 39674 87111 39677
rect 86910 39672 87111 39674
rect 86910 39616 87050 39672
rect 87106 39616 87111 39672
rect 86910 39614 87111 39616
rect 3798 39200 4114 39201
rect 3798 39136 3804 39200
rect 3868 39136 3884 39200
rect 3948 39136 3964 39200
rect 4028 39136 4044 39200
rect 4108 39136 4114 39200
rect 3798 39135 4114 39136
rect 0 38858 800 38888
rect 8342 38861 8402 39100
rect 46828 39070 48116 39130
rect 86910 39100 86970 39614
rect 87045 39611 87111 39614
rect 0 38768 858 38858
rect 8293 38856 8402 38861
rect 8293 38800 8298 38856
rect 8354 38800 8402 38856
rect 8293 38798 8402 38800
rect 88609 38858 88675 38861
rect 89200 38858 90000 38888
rect 88609 38856 90000 38858
rect 88609 38800 88614 38856
rect 88670 38800 90000 38856
rect 88609 38798 90000 38800
rect 8293 38795 8359 38798
rect 88609 38795 88675 38798
rect 89200 38768 90000 38798
rect 798 38725 858 38768
rect 798 38720 907 38725
rect 798 38664 846 38720
rect 902 38664 907 38720
rect 798 38662 907 38664
rect 841 38659 907 38662
rect 3062 38656 3378 38657
rect 3062 38592 3068 38656
rect 3132 38592 3148 38656
rect 3212 38592 3228 38656
rect 3292 38592 3308 38656
rect 3372 38592 3378 38656
rect 3062 38591 3378 38592
rect 3798 38112 4114 38113
rect 3798 38048 3804 38112
rect 3868 38048 3884 38112
rect 3948 38048 3964 38112
rect 4028 38048 4044 38112
rect 4108 38048 4114 38112
rect 3798 38047 4114 38048
rect 8293 37906 8359 37909
rect 8293 37904 8402 37906
rect 8293 37848 8298 37904
rect 8354 37848 8402 37904
rect 8293 37843 8402 37848
rect 8342 37740 8402 37843
rect 87229 37770 87295 37773
rect 46828 37710 48116 37770
rect 86940 37768 87295 37770
rect 86940 37712 87234 37768
rect 87290 37712 87295 37768
rect 86940 37710 87295 37712
rect 87229 37707 87295 37710
rect 841 37634 907 37637
rect 798 37632 907 37634
rect 798 37576 846 37632
rect 902 37576 907 37632
rect 798 37571 907 37576
rect 798 37528 858 37571
rect 0 37438 858 37528
rect 3062 37568 3378 37569
rect 3062 37504 3068 37568
rect 3132 37504 3148 37568
rect 3212 37504 3228 37568
rect 3292 37504 3308 37568
rect 3372 37504 3378 37568
rect 3062 37503 3378 37504
rect 87689 37498 87755 37501
rect 89200 37498 90000 37528
rect 87689 37496 90000 37498
rect 87689 37440 87694 37496
rect 87750 37440 90000 37496
rect 87689 37438 90000 37440
rect 0 37408 800 37438
rect 87689 37435 87755 37438
rect 89200 37408 90000 37438
rect 3798 37024 4114 37025
rect 3798 36960 3804 37024
rect 3868 36960 3884 37024
rect 3948 36960 3964 37024
rect 4028 36960 4044 37024
rect 4108 36960 4114 37024
rect 3798 36959 4114 36960
rect 3062 36480 3378 36481
rect 3062 36416 3068 36480
rect 3132 36416 3148 36480
rect 3212 36416 3228 36480
rect 3292 36416 3308 36480
rect 3372 36416 3378 36480
rect 3062 36415 3378 36416
rect 87505 36410 87571 36413
rect 841 36274 907 36277
rect 798 36272 907 36274
rect 798 36216 846 36272
rect 902 36216 907 36272
rect 798 36211 907 36216
rect 798 36168 858 36211
rect 0 36078 858 36168
rect 8342 36141 8402 36380
rect 46828 36350 48116 36410
rect 86940 36408 87571 36410
rect 86940 36352 87510 36408
rect 87566 36352 87571 36408
rect 86940 36350 87571 36352
rect 87505 36347 87571 36350
rect 8293 36136 8402 36141
rect 8293 36080 8298 36136
rect 8354 36080 8402 36136
rect 8293 36078 8402 36080
rect 88701 36138 88767 36141
rect 89200 36138 90000 36168
rect 88701 36136 90000 36138
rect 88701 36080 88706 36136
rect 88762 36080 90000 36136
rect 88701 36078 90000 36080
rect 0 36048 800 36078
rect 8293 36075 8359 36078
rect 88701 36075 88767 36078
rect 89200 36048 90000 36078
rect 3798 35936 4114 35937
rect 3798 35872 3804 35936
rect 3868 35872 3884 35936
rect 3948 35872 3964 35936
rect 4028 35872 4044 35936
rect 4108 35872 4114 35936
rect 3798 35871 4114 35872
rect 3062 35392 3378 35393
rect 3062 35328 3068 35392
rect 3132 35328 3148 35392
rect 3212 35328 3228 35392
rect 3292 35328 3308 35392
rect 3372 35328 3378 35392
rect 3062 35327 3378 35328
rect 8293 35186 8359 35189
rect 8293 35184 8402 35186
rect 8293 35128 8298 35184
rect 8354 35128 8402 35184
rect 8293 35123 8402 35128
rect 8342 35020 8402 35123
rect 87321 35050 87387 35053
rect 46828 34990 48116 35050
rect 86940 35048 87387 35050
rect 86940 34992 87326 35048
rect 87382 34992 87387 35048
rect 86940 34990 87387 34992
rect 87321 34987 87387 34990
rect 841 34914 907 34917
rect 798 34912 907 34914
rect 798 34856 846 34912
rect 902 34856 907 34912
rect 798 34851 907 34856
rect 798 34808 858 34851
rect 0 34718 858 34808
rect 3798 34848 4114 34849
rect 3798 34784 3804 34848
rect 3868 34784 3884 34848
rect 3948 34784 3964 34848
rect 4028 34784 4044 34848
rect 4108 34784 4114 34848
rect 3798 34783 4114 34784
rect 88793 34778 88859 34781
rect 89200 34778 90000 34808
rect 88793 34776 90000 34778
rect 88793 34720 88798 34776
rect 88854 34720 90000 34776
rect 88793 34718 90000 34720
rect 0 34688 800 34718
rect 88793 34715 88859 34718
rect 89200 34688 90000 34718
rect 3062 34304 3378 34305
rect 3062 34240 3068 34304
rect 3132 34240 3148 34304
rect 3212 34240 3228 34304
rect 3292 34240 3308 34304
rect 3372 34240 3378 34304
rect 3062 34239 3378 34240
rect 3798 33760 4114 33761
rect 3798 33696 3804 33760
rect 3868 33696 3884 33760
rect 3948 33696 3964 33760
rect 4028 33696 4044 33760
rect 4108 33696 4114 33760
rect 3798 33695 4114 33696
rect 0 33418 800 33448
rect 8342 33421 8402 33660
rect 46828 33630 48116 33690
rect 86902 33628 86908 33692
rect 86972 33628 86978 33692
rect 0 33328 858 33418
rect 8293 33416 8402 33421
rect 8293 33360 8298 33416
rect 8354 33360 8402 33416
rect 8293 33358 8402 33360
rect 88977 33418 89043 33421
rect 89200 33418 90000 33448
rect 88977 33416 90000 33418
rect 88977 33360 88982 33416
rect 89038 33360 90000 33416
rect 88977 33358 90000 33360
rect 8293 33355 8359 33358
rect 88977 33355 89043 33358
rect 89200 33328 90000 33358
rect 798 33285 858 33328
rect 798 33280 907 33285
rect 798 33224 846 33280
rect 902 33224 907 33280
rect 798 33222 907 33224
rect 841 33219 907 33222
rect 3062 33216 3378 33217
rect 3062 33152 3068 33216
rect 3132 33152 3148 33216
rect 3212 33152 3228 33216
rect 3292 33152 3308 33216
rect 3372 33152 3378 33216
rect 3062 33151 3378 33152
rect 3798 32672 4114 32673
rect 3798 32608 3804 32672
rect 3868 32608 3884 32672
rect 3948 32608 3964 32672
rect 4028 32608 4044 32672
rect 4108 32608 4114 32672
rect 3798 32607 4114 32608
rect 8293 32466 8359 32469
rect 8293 32464 8402 32466
rect 8293 32408 8298 32464
rect 8354 32408 8402 32464
rect 8293 32403 8402 32408
rect 8342 32300 8402 32403
rect 87086 32330 87092 32332
rect 46828 32270 48116 32330
rect 86940 32270 87092 32330
rect 87086 32268 87092 32270
rect 87156 32268 87162 32332
rect 841 32194 907 32197
rect 798 32192 907 32194
rect 798 32136 846 32192
rect 902 32136 907 32192
rect 798 32131 907 32136
rect 798 32088 858 32131
rect 0 31998 858 32088
rect 3062 32128 3378 32129
rect 3062 32064 3068 32128
rect 3132 32064 3148 32128
rect 3212 32064 3228 32128
rect 3292 32064 3308 32128
rect 3372 32064 3378 32128
rect 3062 32063 3378 32064
rect 88885 32058 88951 32061
rect 89200 32058 90000 32088
rect 88885 32056 90000 32058
rect 88885 32000 88890 32056
rect 88946 32000 90000 32056
rect 88885 31998 90000 32000
rect 0 31968 800 31998
rect 88885 31995 88951 31998
rect 89200 31968 90000 31998
rect 3798 31584 4114 31585
rect 3798 31520 3804 31584
rect 3868 31520 3884 31584
rect 3948 31520 3964 31584
rect 4028 31520 4044 31584
rect 4108 31520 4114 31584
rect 3798 31519 4114 31520
rect 3062 31040 3378 31041
rect 3062 30976 3068 31040
rect 3132 30976 3148 31040
rect 3212 30976 3228 31040
rect 3292 30976 3308 31040
rect 3372 30976 3378 31040
rect 3062 30975 3378 30976
rect 87638 30970 87644 30972
rect 841 30834 907 30837
rect 798 30832 907 30834
rect 798 30776 846 30832
rect 902 30776 907 30832
rect 798 30771 907 30776
rect 798 30728 858 30771
rect 0 30638 858 30728
rect 8342 30701 8402 30940
rect 46828 30910 48116 30970
rect 86940 30910 87644 30970
rect 87638 30908 87644 30910
rect 87708 30908 87714 30972
rect 89200 30701 90000 30728
rect 8293 30696 8402 30701
rect 8293 30640 8298 30696
rect 8354 30640 8402 30696
rect 8293 30638 8402 30640
rect 89161 30696 90000 30701
rect 89161 30640 89166 30696
rect 89222 30640 90000 30696
rect 0 30608 800 30638
rect 8293 30635 8359 30638
rect 89161 30635 90000 30640
rect 89200 30608 90000 30635
rect 3798 30496 4114 30497
rect 3798 30432 3804 30496
rect 3868 30432 3884 30496
rect 3948 30432 3964 30496
rect 4028 30432 4044 30496
rect 4108 30432 4114 30496
rect 3798 30431 4114 30432
rect 3062 29952 3378 29953
rect 3062 29888 3068 29952
rect 3132 29888 3148 29952
rect 3212 29888 3228 29952
rect 3292 29888 3308 29952
rect 3372 29888 3378 29952
rect 3062 29887 3378 29888
rect 8293 29746 8359 29749
rect 8293 29744 8402 29746
rect 8293 29688 8298 29744
rect 8354 29688 8402 29744
rect 8293 29683 8402 29688
rect 8342 29580 8402 29683
rect 87965 29610 88031 29613
rect 46828 29550 48116 29610
rect 86940 29608 88031 29610
rect 86940 29552 87970 29608
rect 88026 29552 88031 29608
rect 86940 29550 88031 29552
rect 87965 29547 88031 29550
rect 841 29474 907 29477
rect 798 29472 907 29474
rect 798 29416 846 29472
rect 902 29416 907 29472
rect 798 29411 907 29416
rect 798 29368 858 29411
rect 0 29278 858 29368
rect 3798 29408 4114 29409
rect 3798 29344 3804 29408
rect 3868 29344 3884 29408
rect 3948 29344 3964 29408
rect 4028 29344 4044 29408
rect 4108 29344 4114 29408
rect 3798 29343 4114 29344
rect 89200 29341 90000 29368
rect 89161 29336 90000 29341
rect 89161 29280 89166 29336
rect 89222 29280 90000 29336
rect 0 29248 800 29278
rect 89161 29275 90000 29280
rect 89200 29248 90000 29275
rect 3062 28864 3378 28865
rect 3062 28800 3068 28864
rect 3132 28800 3148 28864
rect 3212 28800 3228 28864
rect 3292 28800 3308 28864
rect 3372 28800 3378 28864
rect 3062 28799 3378 28800
rect 3798 28320 4114 28321
rect 3798 28256 3804 28320
rect 3868 28256 3884 28320
rect 3948 28256 3964 28320
rect 4028 28256 4044 28320
rect 4108 28256 4114 28320
rect 3798 28255 4114 28256
rect 87137 28250 87203 28253
rect 0 27978 800 28008
rect 8342 27981 8402 28220
rect 46828 28190 48116 28250
rect 86756 28248 87203 28250
rect 86756 28220 87142 28248
rect 86726 28192 87142 28220
rect 87198 28192 87203 28248
rect 86726 28190 87203 28192
rect 86726 27981 86786 28190
rect 87137 28187 87203 28190
rect 0 27888 858 27978
rect 8293 27976 8402 27981
rect 8293 27920 8298 27976
rect 8354 27920 8402 27976
rect 8293 27918 8402 27920
rect 86677 27976 86786 27981
rect 86677 27920 86682 27976
rect 86738 27920 86786 27976
rect 86677 27918 86786 27920
rect 89069 27978 89135 27981
rect 89200 27978 90000 28008
rect 89069 27976 90000 27978
rect 89069 27920 89074 27976
rect 89130 27920 90000 27976
rect 89069 27918 90000 27920
rect 8293 27915 8359 27918
rect 86677 27915 86743 27918
rect 89069 27915 89135 27918
rect 89200 27888 90000 27918
rect 798 27845 858 27888
rect 798 27840 907 27845
rect 798 27784 846 27840
rect 902 27784 907 27840
rect 798 27782 907 27784
rect 841 27779 907 27782
rect 3062 27776 3378 27777
rect 3062 27712 3068 27776
rect 3132 27712 3148 27776
rect 3212 27712 3228 27776
rect 3292 27712 3308 27776
rect 3372 27712 3378 27776
rect 3062 27711 3378 27712
rect 3798 27232 4114 27233
rect 3798 27168 3804 27232
rect 3868 27168 3884 27232
rect 3948 27168 3964 27232
rect 4028 27168 4044 27232
rect 4108 27168 4114 27232
rect 3798 27167 4114 27168
rect 5257 27164 5323 27165
rect 5206 27100 5212 27164
rect 5276 27162 5323 27164
rect 5276 27160 5368 27162
rect 5318 27104 5368 27160
rect 5276 27102 5368 27104
rect 5276 27100 5323 27102
rect 5257 27099 5323 27100
rect 8293 27026 8359 27029
rect 8293 27024 8402 27026
rect 8293 26968 8298 27024
rect 8354 26968 8402 27024
rect 8293 26963 8402 26968
rect 8342 26860 8402 26963
rect 87873 26890 87939 26893
rect 46828 26830 48116 26890
rect 86940 26888 87939 26890
rect 86940 26832 87878 26888
rect 87934 26832 87939 26888
rect 86940 26830 87939 26832
rect 87873 26827 87939 26830
rect 3062 26688 3378 26689
rect 0 26618 800 26648
rect 3062 26624 3068 26688
rect 3132 26624 3148 26688
rect 3212 26624 3228 26688
rect 3292 26624 3308 26688
rect 3372 26624 3378 26688
rect 3062 26623 3378 26624
rect 1301 26618 1367 26621
rect 0 26616 1367 26618
rect 0 26560 1306 26616
rect 1362 26560 1367 26616
rect 0 26558 1367 26560
rect 0 26528 800 26558
rect 1301 26555 1367 26558
rect 87597 26618 87663 26621
rect 89200 26618 90000 26648
rect 87597 26616 90000 26618
rect 87597 26560 87602 26616
rect 87658 26560 90000 26616
rect 87597 26558 90000 26560
rect 87597 26555 87663 26558
rect 89200 26528 90000 26558
rect 3798 26144 4114 26145
rect 3798 26080 3804 26144
rect 3868 26080 3884 26144
rect 3948 26080 3964 26144
rect 4028 26080 4044 26144
rect 4108 26080 4114 26144
rect 3798 26079 4114 26080
rect 8293 25666 8359 25669
rect 8293 25664 8402 25666
rect 8293 25608 8298 25664
rect 8354 25608 8402 25664
rect 8293 25603 8402 25608
rect 3062 25600 3378 25601
rect 3062 25536 3068 25600
rect 3132 25536 3148 25600
rect 3212 25536 3228 25600
rect 3292 25536 3308 25600
rect 3372 25536 3378 25600
rect 3062 25535 3378 25536
rect 8342 25500 8402 25603
rect 87229 25530 87295 25533
rect 46828 25470 48116 25530
rect 86940 25528 87295 25530
rect 86940 25472 87234 25528
rect 87290 25472 87295 25528
rect 86940 25470 87295 25472
rect 87229 25467 87295 25470
rect 0 25258 800 25288
rect 89200 25261 90000 25288
rect 1209 25258 1275 25261
rect 0 25256 1275 25258
rect 0 25200 1214 25256
rect 1270 25200 1275 25256
rect 0 25198 1275 25200
rect 0 25168 800 25198
rect 1209 25195 1275 25198
rect 89161 25256 90000 25261
rect 89161 25200 89166 25256
rect 89222 25200 90000 25256
rect 89161 25195 90000 25200
rect 89200 25168 90000 25195
rect 3798 25056 4114 25057
rect 3798 24992 3804 25056
rect 3868 24992 3884 25056
rect 3948 24992 3964 25056
rect 4028 24992 4044 25056
rect 4108 24992 4114 25056
rect 3798 24991 4114 24992
rect 3062 24512 3378 24513
rect 3062 24448 3068 24512
rect 3132 24448 3148 24512
rect 3212 24448 3228 24512
rect 3292 24448 3308 24512
rect 3372 24448 3378 24512
rect 3062 24447 3378 24448
rect 8293 24306 8359 24309
rect 8293 24304 8402 24306
rect 8293 24248 8298 24304
rect 8354 24248 8402 24304
rect 8293 24243 8402 24248
rect 8342 24140 8402 24243
rect 88742 24170 88748 24172
rect 46828 24110 48116 24170
rect 86940 24110 88748 24170
rect 88742 24108 88748 24110
rect 88812 24108 88818 24172
rect 3798 23968 4114 23969
rect 0 23898 800 23928
rect 3798 23904 3804 23968
rect 3868 23904 3884 23968
rect 3948 23904 3964 23968
rect 4028 23904 4044 23968
rect 4108 23904 4114 23968
rect 3798 23903 4114 23904
rect 1301 23898 1367 23901
rect 0 23896 1367 23898
rect 0 23840 1306 23896
rect 1362 23840 1367 23896
rect 0 23838 1367 23840
rect 0 23808 800 23838
rect 1301 23835 1367 23838
rect 88558 23836 88564 23900
rect 88628 23898 88634 23900
rect 89200 23898 90000 23928
rect 88628 23838 90000 23898
rect 88628 23836 88634 23838
rect 89200 23808 90000 23838
rect 3062 23424 3378 23425
rect 3062 23360 3068 23424
rect 3132 23360 3148 23424
rect 3212 23360 3228 23424
rect 3292 23360 3308 23424
rect 3372 23360 3378 23424
rect 3062 23359 3378 23360
rect 3798 22880 4114 22881
rect 3798 22816 3804 22880
rect 3868 22816 3884 22880
rect 3948 22816 3964 22880
rect 4028 22816 4044 22880
rect 4108 22816 4114 22880
rect 3798 22815 4114 22816
rect 0 22538 800 22568
rect 8342 22541 8402 22780
rect 46828 22750 48116 22810
rect 86350 22748 86356 22812
rect 86420 22748 86426 22812
rect 1301 22538 1367 22541
rect 0 22536 1367 22538
rect 0 22480 1306 22536
rect 1362 22480 1367 22536
rect 0 22478 1367 22480
rect 0 22448 800 22478
rect 1301 22475 1367 22478
rect 8293 22536 8402 22541
rect 8293 22480 8298 22536
rect 8354 22480 8402 22536
rect 8293 22478 8402 22480
rect 89069 22538 89135 22541
rect 89200 22538 90000 22568
rect 89069 22536 90000 22538
rect 89069 22480 89074 22536
rect 89130 22480 90000 22536
rect 89069 22478 90000 22480
rect 8293 22475 8359 22478
rect 89069 22475 89135 22478
rect 89200 22448 90000 22478
rect 3062 22336 3378 22337
rect 3062 22272 3068 22336
rect 3132 22272 3148 22336
rect 3212 22272 3228 22336
rect 3292 22272 3308 22336
rect 3372 22272 3378 22336
rect 3062 22271 3378 22272
rect 3798 21792 4114 21793
rect 3798 21728 3804 21792
rect 3868 21728 3884 21792
rect 3948 21728 3964 21792
rect 4028 21728 4044 21792
rect 4108 21728 4114 21792
rect 3798 21727 4114 21728
rect 8293 21586 8359 21589
rect 8293 21584 8402 21586
rect 8293 21528 8298 21584
rect 8354 21528 8402 21584
rect 8293 21523 8402 21528
rect 8342 21420 8402 21523
rect 88190 21450 88196 21452
rect 46828 21390 48116 21450
rect 86940 21390 88196 21450
rect 88190 21388 88196 21390
rect 88260 21388 88266 21452
rect 3062 21248 3378 21249
rect 0 21178 800 21208
rect 3062 21184 3068 21248
rect 3132 21184 3148 21248
rect 3212 21184 3228 21248
rect 3292 21184 3308 21248
rect 3372 21184 3378 21248
rect 3062 21183 3378 21184
rect 1301 21178 1367 21181
rect 0 21176 1367 21178
rect 0 21120 1306 21176
rect 1362 21120 1367 21176
rect 0 21118 1367 21120
rect 0 21088 800 21118
rect 1301 21115 1367 21118
rect 88425 21178 88491 21181
rect 89200 21178 90000 21208
rect 88425 21176 90000 21178
rect 88425 21120 88430 21176
rect 88486 21120 90000 21176
rect 88425 21118 90000 21120
rect 88425 21115 88491 21118
rect 89200 21088 90000 21118
rect 3798 20704 4114 20705
rect 3798 20640 3804 20704
rect 3868 20640 3884 20704
rect 3948 20640 3964 20704
rect 4028 20640 4044 20704
rect 4108 20640 4114 20704
rect 3798 20639 4114 20640
rect 8293 20226 8359 20229
rect 8293 20224 8402 20226
rect 8293 20168 8298 20224
rect 8354 20168 8402 20224
rect 8293 20163 8402 20168
rect 3062 20160 3378 20161
rect 3062 20096 3068 20160
rect 3132 20096 3148 20160
rect 3212 20096 3228 20160
rect 3292 20096 3308 20160
rect 3372 20096 3378 20160
rect 3062 20095 3378 20096
rect 8342 20060 8402 20163
rect 87505 20090 87571 20093
rect 46828 20030 48116 20090
rect 86940 20088 87571 20090
rect 86940 20032 87510 20088
rect 87566 20032 87571 20088
rect 86940 20030 87571 20032
rect 87505 20027 87571 20030
rect 0 19818 800 19848
rect 1209 19818 1275 19821
rect 89200 19818 90000 19848
rect 0 19816 1275 19818
rect 0 19760 1214 19816
rect 1270 19760 1275 19816
rect 0 19758 1275 19760
rect 0 19728 800 19758
rect 1209 19755 1275 19758
rect 89072 19758 90000 19818
rect 3798 19616 4114 19617
rect 3798 19552 3804 19616
rect 3868 19552 3884 19616
rect 3948 19552 3964 19616
rect 4028 19552 4044 19616
rect 4108 19552 4114 19616
rect 3798 19551 4114 19552
rect 89072 19546 89132 19758
rect 89200 19728 90000 19758
rect 89253 19546 89319 19549
rect 89072 19544 89319 19546
rect 89072 19488 89258 19544
rect 89314 19488 89319 19544
rect 89072 19486 89319 19488
rect 89253 19483 89319 19486
rect 3062 19072 3378 19073
rect 3062 19008 3068 19072
rect 3132 19008 3148 19072
rect 3212 19008 3228 19072
rect 3292 19008 3308 19072
rect 3372 19008 3378 19072
rect 3062 19007 3378 19008
rect 8293 18866 8359 18869
rect 8293 18864 8402 18866
rect 8293 18808 8298 18864
rect 8354 18808 8402 18864
rect 8293 18803 8402 18808
rect 8342 18700 8402 18803
rect 87873 18730 87939 18733
rect 46828 18670 48116 18730
rect 86940 18728 87939 18730
rect 86940 18672 87878 18728
rect 87934 18672 87939 18728
rect 86940 18670 87939 18672
rect 87873 18667 87939 18670
rect 3798 18528 4114 18529
rect 0 18458 800 18488
rect 3798 18464 3804 18528
rect 3868 18464 3884 18528
rect 3948 18464 3964 18528
rect 4028 18464 4044 18528
rect 4108 18464 4114 18528
rect 3798 18463 4114 18464
rect 1301 18458 1367 18461
rect 89200 18458 90000 18488
rect 0 18456 1367 18458
rect 0 18400 1306 18456
rect 1362 18400 1367 18456
rect 0 18398 1367 18400
rect 0 18368 800 18398
rect 1301 18395 1367 18398
rect 89072 18398 90000 18458
rect 89072 18186 89132 18398
rect 89200 18368 90000 18398
rect 89345 18186 89411 18189
rect 89072 18184 89411 18186
rect 89072 18128 89350 18184
rect 89406 18128 89411 18184
rect 89072 18126 89411 18128
rect 89345 18123 89411 18126
rect 3062 17984 3378 17985
rect 3062 17920 3068 17984
rect 3132 17920 3148 17984
rect 3212 17920 3228 17984
rect 3292 17920 3308 17984
rect 3372 17920 3378 17984
rect 3062 17919 3378 17920
rect 3798 17440 4114 17441
rect 3798 17376 3804 17440
rect 3868 17376 3884 17440
rect 3948 17376 3964 17440
rect 4028 17376 4044 17440
rect 4108 17376 4114 17440
rect 3798 17375 4114 17376
rect 87137 17370 87203 17373
rect 0 17098 800 17128
rect 8342 17101 8402 17340
rect 46828 17310 48116 17370
rect 86940 17368 87203 17370
rect 86940 17312 87142 17368
rect 87198 17312 87203 17368
rect 86940 17310 87203 17312
rect 87137 17307 87203 17310
rect 1301 17098 1367 17101
rect 0 17096 1367 17098
rect 0 17040 1306 17096
rect 1362 17040 1367 17096
rect 0 17038 1367 17040
rect 0 17008 800 17038
rect 1301 17035 1367 17038
rect 8293 17096 8402 17101
rect 8293 17040 8298 17096
rect 8354 17040 8402 17096
rect 8293 17038 8402 17040
rect 89069 17098 89135 17101
rect 89200 17098 90000 17128
rect 89069 17096 90000 17098
rect 89069 17040 89074 17096
rect 89130 17040 90000 17096
rect 89069 17038 90000 17040
rect 8293 17035 8359 17038
rect 89069 17035 89135 17038
rect 89200 17008 90000 17038
rect 3062 16896 3378 16897
rect 3062 16832 3068 16896
rect 3132 16832 3148 16896
rect 3212 16832 3228 16896
rect 3292 16832 3308 16896
rect 3372 16832 3378 16896
rect 3062 16831 3378 16832
rect 3798 16352 4114 16353
rect 3798 16288 3804 16352
rect 3868 16288 3884 16352
rect 3948 16288 3964 16352
rect 4028 16288 4044 16352
rect 4108 16288 4114 16352
rect 3798 16287 4114 16288
rect 8293 16146 8359 16149
rect 8293 16144 8402 16146
rect 8293 16088 8298 16144
rect 8354 16088 8402 16144
rect 8293 16083 8402 16088
rect 8342 15980 8402 16083
rect 46828 15950 48116 16010
rect 3062 15808 3378 15809
rect 0 15738 800 15768
rect 3062 15744 3068 15808
rect 3132 15744 3148 15808
rect 3212 15744 3228 15808
rect 3292 15744 3308 15808
rect 3372 15744 3378 15808
rect 3062 15743 3378 15744
rect 1301 15738 1367 15741
rect 0 15736 1367 15738
rect 0 15680 1306 15736
rect 1362 15680 1367 15736
rect 0 15678 1367 15680
rect 0 15648 800 15678
rect 1301 15675 1367 15678
rect 86910 15466 86970 15980
rect 88977 15738 89043 15741
rect 89200 15738 90000 15768
rect 88977 15736 90000 15738
rect 88977 15680 88982 15736
rect 89038 15680 90000 15736
rect 88977 15678 90000 15680
rect 88977 15675 89043 15678
rect 89200 15648 90000 15678
rect 87045 15466 87111 15469
rect 86910 15464 87111 15466
rect 86910 15408 87050 15464
rect 87106 15408 87111 15464
rect 86910 15406 87111 15408
rect 87045 15403 87111 15406
rect 3798 15264 4114 15265
rect 3798 15200 3804 15264
rect 3868 15200 3884 15264
rect 3948 15200 3964 15264
rect 4028 15200 4044 15264
rect 4108 15200 4114 15264
rect 3798 15199 4114 15200
rect 8293 14786 8359 14789
rect 8293 14784 8402 14786
rect 8293 14728 8298 14784
rect 8354 14728 8402 14784
rect 8293 14723 8402 14728
rect 3062 14720 3378 14721
rect 3062 14656 3068 14720
rect 3132 14656 3148 14720
rect 3212 14656 3228 14720
rect 3292 14656 3308 14720
rect 3372 14656 3378 14720
rect 3062 14655 3378 14656
rect 8342 14620 8402 14723
rect 88609 14650 88675 14653
rect 46828 14590 48116 14650
rect 86940 14648 88675 14650
rect 86940 14592 88614 14648
rect 88670 14592 88675 14648
rect 86940 14590 88675 14592
rect 88609 14587 88675 14590
rect 0 14378 800 14408
rect 1209 14378 1275 14381
rect 89200 14378 90000 14408
rect 0 14376 1275 14378
rect 0 14320 1214 14376
rect 1270 14320 1275 14376
rect 0 14318 1275 14320
rect 0 14288 800 14318
rect 1209 14315 1275 14318
rect 89072 14318 90000 14378
rect 3798 14176 4114 14177
rect 3798 14112 3804 14176
rect 3868 14112 3884 14176
rect 3948 14112 3964 14176
rect 4028 14112 4044 14176
rect 4108 14112 4114 14176
rect 3798 14111 4114 14112
rect 89072 14106 89132 14318
rect 89200 14288 90000 14318
rect 89437 14106 89503 14109
rect 89072 14104 89503 14106
rect 89072 14048 89442 14104
rect 89498 14048 89503 14104
rect 89072 14046 89503 14048
rect 89437 14043 89503 14046
rect 86350 13636 86356 13700
rect 86420 13698 86426 13700
rect 86585 13698 86651 13701
rect 86420 13696 86651 13698
rect 86420 13640 86590 13696
rect 86646 13640 86651 13696
rect 86420 13638 86651 13640
rect 86420 13636 86426 13638
rect 86585 13635 86651 13638
rect 3062 13632 3378 13633
rect 3062 13568 3068 13632
rect 3132 13568 3148 13632
rect 3212 13568 3228 13632
rect 3292 13568 3308 13632
rect 3372 13568 3378 13632
rect 3062 13567 3378 13568
rect 8293 13426 8359 13429
rect 8293 13424 8402 13426
rect 8293 13368 8298 13424
rect 8354 13368 8402 13424
rect 8293 13363 8402 13368
rect 8342 13260 8402 13363
rect 87413 13290 87479 13293
rect 46828 13230 48116 13290
rect 86940 13288 87479 13290
rect 86940 13232 87418 13288
rect 87474 13232 87479 13288
rect 86940 13230 87479 13232
rect 87413 13227 87479 13230
rect 3798 13088 4114 13089
rect 0 13018 800 13048
rect 3798 13024 3804 13088
rect 3868 13024 3884 13088
rect 3948 13024 3964 13088
rect 4028 13024 4044 13088
rect 4108 13024 4114 13088
rect 3798 13023 4114 13024
rect 1301 13018 1367 13021
rect 0 13016 1367 13018
rect 0 12960 1306 13016
rect 1362 12960 1367 13016
rect 0 12958 1367 12960
rect 0 12928 800 12958
rect 1301 12955 1367 12958
rect 88885 13018 88951 13021
rect 89200 13018 90000 13048
rect 88885 13016 90000 13018
rect 88885 12960 88890 13016
rect 88946 12960 90000 13016
rect 88885 12958 90000 12960
rect 88885 12955 88951 12958
rect 89200 12928 90000 12958
rect 86534 12548 86540 12612
rect 86604 12610 86610 12612
rect 87321 12610 87387 12613
rect 86604 12608 87387 12610
rect 86604 12552 87326 12608
rect 87382 12552 87387 12608
rect 86604 12550 87387 12552
rect 86604 12548 86610 12550
rect 87321 12547 87387 12550
rect 3062 12544 3378 12545
rect 3062 12480 3068 12544
rect 3132 12480 3148 12544
rect 3212 12480 3228 12544
rect 3292 12480 3308 12544
rect 3372 12480 3378 12544
rect 3062 12479 3378 12480
rect 3798 12000 4114 12001
rect 3798 11936 3804 12000
rect 3868 11936 3884 12000
rect 3948 11936 3964 12000
rect 4028 11936 4044 12000
rect 4108 11936 4114 12000
rect 3798 11935 4114 11936
rect 87781 11930 87847 11933
rect 0 11658 800 11688
rect 8342 11661 8402 11900
rect 46828 11870 48116 11930
rect 86940 11928 87847 11930
rect 86940 11872 87786 11928
rect 87842 11872 87847 11928
rect 86940 11870 87847 11872
rect 87781 11867 87847 11870
rect 1301 11658 1367 11661
rect 0 11656 1367 11658
rect 0 11600 1306 11656
rect 1362 11600 1367 11656
rect 0 11598 1367 11600
rect 0 11568 800 11598
rect 1301 11595 1367 11598
rect 8293 11656 8402 11661
rect 8293 11600 8298 11656
rect 8354 11600 8402 11656
rect 8293 11598 8402 11600
rect 88793 11658 88859 11661
rect 89200 11658 90000 11688
rect 88793 11656 90000 11658
rect 88793 11600 88798 11656
rect 88854 11600 90000 11656
rect 88793 11598 90000 11600
rect 8293 11595 8359 11598
rect 88793 11595 88859 11598
rect 89200 11568 90000 11598
rect 3062 11456 3378 11457
rect 3062 11392 3068 11456
rect 3132 11392 3148 11456
rect 3212 11392 3228 11456
rect 3292 11392 3308 11456
rect 3372 11392 3378 11456
rect 3062 11391 3378 11392
rect 87965 11114 88031 11117
rect 88374 11114 88380 11116
rect 87965 11112 88380 11114
rect 87965 11056 87970 11112
rect 88026 11056 88380 11112
rect 87965 11054 88380 11056
rect 87965 11051 88031 11054
rect 88374 11052 88380 11054
rect 88444 11052 88450 11116
rect 3798 10912 4114 10913
rect 3798 10848 3804 10912
rect 3868 10848 3884 10912
rect 3948 10848 3964 10912
rect 4028 10848 4044 10912
rect 4108 10848 4114 10912
rect 3798 10847 4114 10848
rect 87965 10570 88031 10573
rect 3062 10368 3378 10369
rect 3062 10304 3068 10368
rect 3132 10304 3148 10368
rect 3212 10304 3228 10368
rect 3292 10304 3308 10368
rect 3372 10304 3378 10368
rect 3062 10303 3378 10304
rect 8158 10029 8218 10540
rect 46828 10510 48116 10570
rect 86940 10568 88031 10570
rect 86940 10512 87970 10568
rect 88026 10512 88031 10568
rect 86940 10510 88031 10512
rect 87965 10507 88031 10510
rect 88701 10298 88767 10301
rect 89200 10298 90000 10328
rect 88701 10296 90000 10298
rect 88701 10240 88706 10296
rect 88762 10240 90000 10296
rect 88701 10238 90000 10240
rect 88701 10235 88767 10238
rect 89200 10208 90000 10238
rect 8109 10024 8218 10029
rect 8109 9968 8114 10024
rect 8170 9968 8218 10024
rect 8109 9966 8218 9968
rect 8109 9963 8175 9966
rect 3798 9824 4114 9825
rect 3798 9760 3804 9824
rect 3868 9760 3884 9824
rect 3948 9760 3964 9824
rect 4028 9760 4044 9824
rect 4108 9760 4114 9824
rect 3798 9759 4114 9760
rect 88241 9618 88307 9621
rect 88742 9618 88748 9620
rect 88241 9616 88748 9618
rect 88241 9560 88246 9616
rect 88302 9560 88748 9616
rect 88241 9558 88748 9560
rect 88241 9555 88307 9558
rect 88742 9556 88748 9558
rect 88812 9556 88818 9620
rect 89200 9618 90000 9648
rect 88934 9558 90000 9618
rect 88934 9346 88994 9558
rect 89200 9528 90000 9558
rect 87094 9286 88994 9346
rect 3062 9280 3378 9281
rect 3062 9216 3068 9280
rect 3132 9216 3148 9280
rect 3212 9216 3228 9280
rect 3292 9216 3308 9280
rect 3372 9216 3378 9280
rect 3062 9215 3378 9216
rect 3798 8736 4114 8737
rect 3798 8672 3804 8736
rect 3868 8672 3884 8736
rect 3948 8672 3964 8736
rect 4028 8672 4044 8736
rect 4108 8672 4114 8736
rect 3798 8671 4114 8672
rect 8342 8669 8402 9180
rect 46828 9150 48116 9210
rect 8293 8664 8402 8669
rect 8293 8608 8298 8664
rect 8354 8608 8402 8664
rect 8293 8606 8402 8608
rect 86358 8669 86418 9180
rect 86358 8664 86467 8669
rect 86358 8608 86406 8664
rect 86462 8608 86467 8664
rect 86358 8606 86467 8608
rect 8293 8603 8359 8606
rect 86401 8603 86467 8606
rect 86585 8530 86651 8533
rect 87094 8530 87154 9286
rect 88333 8938 88399 8941
rect 89200 8938 90000 8968
rect 88333 8936 90000 8938
rect 88333 8880 88338 8936
rect 88394 8880 90000 8936
rect 88333 8878 90000 8880
rect 88333 8875 88399 8878
rect 89200 8848 90000 8878
rect 86585 8528 87154 8530
rect 86585 8472 86590 8528
rect 86646 8472 87154 8528
rect 86585 8470 87154 8472
rect 86585 8467 86651 8470
rect 86033 8394 86099 8397
rect 88374 8394 88380 8396
rect 86033 8392 88380 8394
rect 86033 8336 86038 8392
rect 86094 8336 88380 8392
rect 86033 8334 88380 8336
rect 86033 8331 86099 8334
rect 88374 8332 88380 8334
rect 88444 8332 88450 8396
rect 85665 8258 85731 8261
rect 86902 8258 86908 8260
rect 85665 8256 86908 8258
rect 85665 8200 85670 8256
rect 85726 8200 86908 8256
rect 85665 8198 86908 8200
rect 85665 8195 85731 8198
rect 86902 8196 86908 8198
rect 86972 8196 86978 8260
rect 89200 8258 90000 8288
rect 87830 8198 90000 8258
rect 3062 8192 3378 8193
rect 3062 8128 3068 8192
rect 3132 8128 3148 8192
rect 3212 8128 3228 8192
rect 3292 8128 3308 8192
rect 3372 8128 3378 8192
rect 3062 8127 3378 8128
rect 86309 8122 86375 8125
rect 87830 8122 87890 8198
rect 89200 8168 90000 8198
rect 86309 8120 87890 8122
rect 86309 8064 86314 8120
rect 86370 8064 87890 8120
rect 86309 8062 87890 8064
rect 86309 8059 86375 8062
rect 85757 7986 85823 7989
rect 87086 7986 87092 7988
rect 85757 7984 87092 7986
rect 85757 7928 85762 7984
rect 85818 7928 87092 7984
rect 85757 7926 87092 7928
rect 85757 7923 85823 7926
rect 87086 7924 87092 7926
rect 87156 7924 87162 7988
rect 3798 7648 4114 7649
rect 3798 7584 3804 7648
rect 3868 7584 3884 7648
rect 3948 7584 3964 7648
rect 4028 7584 4044 7648
rect 4108 7584 4114 7648
rect 3798 7583 4114 7584
rect 3062 7104 3378 7105
rect 3062 7040 3068 7104
rect 3132 7040 3148 7104
rect 3212 7040 3228 7104
rect 3292 7040 3308 7104
rect 3372 7040 3378 7104
rect 3062 7039 3378 7040
rect 3798 6560 4114 6561
rect 3798 6496 3804 6560
rect 3868 6496 3884 6560
rect 3948 6496 3964 6560
rect 4028 6496 4044 6560
rect 4108 6496 4114 6560
rect 3798 6495 4114 6496
rect 3062 6016 3378 6017
rect 3062 5952 3068 6016
rect 3132 5952 3148 6016
rect 3212 5952 3228 6016
rect 3292 5952 3308 6016
rect 3372 5952 3378 6016
rect 3062 5951 3378 5952
rect 72946 6016 73262 6017
rect 72946 5952 72952 6016
rect 73016 5952 73032 6016
rect 73096 5952 73112 6016
rect 73176 5952 73192 6016
rect 73256 5952 73262 6016
rect 72946 5951 73262 5952
rect 88517 5948 88583 5949
rect 88517 5946 88564 5948
rect 88472 5944 88564 5946
rect 88472 5888 88522 5944
rect 88472 5886 88564 5888
rect 88517 5884 88564 5886
rect 88628 5884 88634 5948
rect 88517 5883 88583 5884
rect 47710 5748 47716 5812
rect 47780 5810 47786 5812
rect 85113 5810 85179 5813
rect 47780 5808 85179 5810
rect 47780 5752 85118 5808
rect 85174 5752 85179 5808
rect 47780 5750 85179 5752
rect 47780 5748 47786 5750
rect 85113 5747 85179 5750
rect 48078 5612 48084 5676
rect 48148 5674 48154 5676
rect 85573 5674 85639 5677
rect 48148 5672 85639 5674
rect 48148 5616 85578 5672
rect 85634 5616 85639 5672
rect 48148 5614 85639 5616
rect 48148 5612 48154 5614
rect 85573 5611 85639 5614
rect 88241 5540 88307 5541
rect 88190 5538 88196 5540
rect 88150 5478 88196 5538
rect 88260 5536 88307 5540
rect 88302 5480 88307 5536
rect 88190 5476 88196 5478
rect 88260 5476 88307 5480
rect 88241 5475 88307 5476
rect 3798 5472 4114 5473
rect 3798 5408 3804 5472
rect 3868 5408 3884 5472
rect 3948 5408 3964 5472
rect 4028 5408 4044 5472
rect 4108 5408 4114 5472
rect 3798 5407 4114 5408
rect 37606 5472 37922 5473
rect 37606 5408 37612 5472
rect 37676 5408 37692 5472
rect 37756 5408 37772 5472
rect 37836 5408 37852 5472
rect 37916 5408 37922 5472
rect 37606 5407 37922 5408
rect 73606 5472 73922 5473
rect 73606 5408 73612 5472
rect 73676 5408 73692 5472
rect 73756 5408 73772 5472
rect 73836 5408 73852 5472
rect 73916 5408 73922 5472
rect 73606 5407 73922 5408
rect 86493 5404 86559 5405
rect 86493 5402 86540 5404
rect 86448 5400 86540 5402
rect 86448 5344 86498 5400
rect 86448 5342 86540 5344
rect 86493 5340 86540 5342
rect 86604 5340 86610 5404
rect 86493 5339 86559 5340
rect 36946 4928 37262 4929
rect 36946 4864 36952 4928
rect 37016 4864 37032 4928
rect 37096 4864 37112 4928
rect 37176 4864 37192 4928
rect 37256 4864 37262 4928
rect 36946 4863 37262 4864
rect 72946 4928 73262 4929
rect 72946 4864 72952 4928
rect 73016 4864 73032 4928
rect 73096 4864 73112 4928
rect 73176 4864 73192 4928
rect 73256 4864 73262 4928
rect 72946 4863 73262 4864
rect 87229 4860 87295 4861
rect 87229 4858 87276 4860
rect 87184 4856 87276 4858
rect 87184 4800 87234 4856
rect 87184 4798 87276 4800
rect 87229 4796 87276 4798
rect 87340 4796 87346 4860
rect 87229 4795 87295 4796
rect 47894 4524 47900 4588
rect 47964 4586 47970 4588
rect 86953 4586 87019 4589
rect 47964 4584 87019 4586
rect 47964 4528 86958 4584
rect 87014 4528 87019 4584
rect 47964 4526 87019 4528
rect 47964 4524 47970 4526
rect 86953 4523 87019 4526
rect 37606 4384 37922 4385
rect 37606 4320 37612 4384
rect 37676 4320 37692 4384
rect 37756 4320 37772 4384
rect 37836 4320 37852 4384
rect 37916 4320 37922 4384
rect 37606 4319 37922 4320
rect 73606 4384 73922 4385
rect 73606 4320 73612 4384
rect 73676 4320 73692 4384
rect 73756 4320 73772 4384
rect 73836 4320 73852 4384
rect 73916 4320 73922 4384
rect 73606 4319 73922 4320
rect 36946 3840 37262 3841
rect 36946 3776 36952 3840
rect 37016 3776 37032 3840
rect 37096 3776 37112 3840
rect 37176 3776 37192 3840
rect 37256 3776 37262 3840
rect 36946 3775 37262 3776
rect 72946 3840 73262 3841
rect 72946 3776 72952 3840
rect 73016 3776 73032 3840
rect 73096 3776 73112 3840
rect 73176 3776 73192 3840
rect 73256 3776 73262 3840
rect 72946 3775 73262 3776
rect 37606 3296 37922 3297
rect 37606 3232 37612 3296
rect 37676 3232 37692 3296
rect 37756 3232 37772 3296
rect 37836 3232 37852 3296
rect 37916 3232 37922 3296
rect 37606 3231 37922 3232
rect 73606 3296 73922 3297
rect 73606 3232 73612 3296
rect 73676 3232 73692 3296
rect 73756 3232 73772 3296
rect 73836 3232 73852 3296
rect 73916 3232 73922 3296
rect 73606 3231 73922 3232
rect 36946 2752 37262 2753
rect 36946 2688 36952 2752
rect 37016 2688 37032 2752
rect 37096 2688 37112 2752
rect 37176 2688 37192 2752
rect 37256 2688 37262 2752
rect 36946 2687 37262 2688
rect 72946 2752 73262 2753
rect 72946 2688 72952 2752
rect 73016 2688 73032 2752
rect 73096 2688 73112 2752
rect 73176 2688 73192 2752
rect 73256 2688 73262 2752
rect 72946 2687 73262 2688
rect 37606 2208 37922 2209
rect 37606 2144 37612 2208
rect 37676 2144 37692 2208
rect 37756 2144 37772 2208
rect 37836 2144 37852 2208
rect 37916 2144 37922 2208
rect 37606 2143 37922 2144
rect 73606 2208 73922 2209
rect 73606 2144 73612 2208
rect 73676 2144 73692 2208
rect 73756 2144 73772 2208
rect 73836 2144 73852 2208
rect 73916 2144 73922 2208
rect 73606 2143 73922 2144
<< via3 >>
rect 37612 95772 37676 95776
rect 37612 95716 37616 95772
rect 37616 95716 37672 95772
rect 37672 95716 37676 95772
rect 37612 95712 37676 95716
rect 37692 95772 37756 95776
rect 37692 95716 37696 95772
rect 37696 95716 37752 95772
rect 37752 95716 37756 95772
rect 37692 95712 37756 95716
rect 37772 95772 37836 95776
rect 37772 95716 37776 95772
rect 37776 95716 37832 95772
rect 37832 95716 37836 95772
rect 37772 95712 37836 95716
rect 37852 95772 37916 95776
rect 37852 95716 37856 95772
rect 37856 95716 37912 95772
rect 37912 95716 37916 95772
rect 37852 95712 37916 95716
rect 73612 95772 73676 95776
rect 73612 95716 73616 95772
rect 73616 95716 73672 95772
rect 73672 95716 73676 95772
rect 73612 95712 73676 95716
rect 73692 95772 73756 95776
rect 73692 95716 73696 95772
rect 73696 95716 73752 95772
rect 73752 95716 73756 95772
rect 73692 95712 73756 95716
rect 73772 95772 73836 95776
rect 73772 95716 73776 95772
rect 73776 95716 73832 95772
rect 73832 95716 73836 95772
rect 73772 95712 73836 95716
rect 73852 95772 73916 95776
rect 73852 95716 73856 95772
rect 73856 95716 73912 95772
rect 73912 95716 73916 95772
rect 73852 95712 73916 95716
rect 8524 95296 8588 95300
rect 8524 95240 8538 95296
rect 8538 95240 8588 95296
rect 8524 95236 8588 95240
rect 36952 95228 37016 95232
rect 36952 95172 36956 95228
rect 36956 95172 37012 95228
rect 37012 95172 37016 95228
rect 36952 95168 37016 95172
rect 37032 95228 37096 95232
rect 37032 95172 37036 95228
rect 37036 95172 37092 95228
rect 37092 95172 37096 95228
rect 37032 95168 37096 95172
rect 37112 95228 37176 95232
rect 37112 95172 37116 95228
rect 37116 95172 37172 95228
rect 37172 95172 37176 95228
rect 37112 95168 37176 95172
rect 37192 95228 37256 95232
rect 37192 95172 37196 95228
rect 37196 95172 37252 95228
rect 37252 95172 37256 95228
rect 37192 95168 37256 95172
rect 72952 95228 73016 95232
rect 72952 95172 72956 95228
rect 72956 95172 73012 95228
rect 73012 95172 73016 95228
rect 72952 95168 73016 95172
rect 73032 95228 73096 95232
rect 73032 95172 73036 95228
rect 73036 95172 73092 95228
rect 73092 95172 73096 95228
rect 73032 95168 73096 95172
rect 73112 95228 73176 95232
rect 73112 95172 73116 95228
rect 73116 95172 73172 95228
rect 73172 95172 73176 95228
rect 73112 95168 73176 95172
rect 73192 95228 73256 95232
rect 73192 95172 73196 95228
rect 73196 95172 73252 95228
rect 73252 95172 73256 95228
rect 73192 95168 73256 95172
rect 37612 94684 37676 94688
rect 37612 94628 37616 94684
rect 37616 94628 37672 94684
rect 37672 94628 37676 94684
rect 37612 94624 37676 94628
rect 37692 94684 37756 94688
rect 37692 94628 37696 94684
rect 37696 94628 37752 94684
rect 37752 94628 37756 94684
rect 37692 94624 37756 94628
rect 37772 94684 37836 94688
rect 37772 94628 37776 94684
rect 37776 94628 37832 94684
rect 37832 94628 37836 94684
rect 37772 94624 37836 94628
rect 37852 94684 37916 94688
rect 37852 94628 37856 94684
rect 37856 94628 37912 94684
rect 37912 94628 37916 94684
rect 37852 94624 37916 94628
rect 73612 94684 73676 94688
rect 73612 94628 73616 94684
rect 73616 94628 73672 94684
rect 73672 94628 73676 94684
rect 73612 94624 73676 94628
rect 73692 94684 73756 94688
rect 73692 94628 73696 94684
rect 73696 94628 73752 94684
rect 73752 94628 73756 94684
rect 73692 94624 73756 94628
rect 73772 94684 73836 94688
rect 73772 94628 73776 94684
rect 73776 94628 73832 94684
rect 73832 94628 73836 94684
rect 73772 94624 73836 94628
rect 73852 94684 73916 94688
rect 73852 94628 73856 94684
rect 73856 94628 73912 94684
rect 73912 94628 73916 94684
rect 73852 94624 73916 94628
rect 36952 94140 37016 94144
rect 36952 94084 36956 94140
rect 36956 94084 37012 94140
rect 37012 94084 37016 94140
rect 36952 94080 37016 94084
rect 37032 94140 37096 94144
rect 37032 94084 37036 94140
rect 37036 94084 37092 94140
rect 37092 94084 37096 94140
rect 37032 94080 37096 94084
rect 37112 94140 37176 94144
rect 37112 94084 37116 94140
rect 37116 94084 37172 94140
rect 37172 94084 37176 94140
rect 37112 94080 37176 94084
rect 37192 94140 37256 94144
rect 37192 94084 37196 94140
rect 37196 94084 37252 94140
rect 37252 94084 37256 94140
rect 37192 94080 37256 94084
rect 72952 94140 73016 94144
rect 72952 94084 72956 94140
rect 72956 94084 73012 94140
rect 73012 94084 73016 94140
rect 72952 94080 73016 94084
rect 73032 94140 73096 94144
rect 73032 94084 73036 94140
rect 73036 94084 73092 94140
rect 73092 94084 73096 94140
rect 73032 94080 73096 94084
rect 73112 94140 73176 94144
rect 73112 94084 73116 94140
rect 73116 94084 73172 94140
rect 73172 94084 73176 94140
rect 73112 94080 73176 94084
rect 73192 94140 73256 94144
rect 73192 94084 73196 94140
rect 73196 94084 73252 94140
rect 73252 94084 73256 94140
rect 73192 94080 73256 94084
rect 37612 93596 37676 93600
rect 37612 93540 37616 93596
rect 37616 93540 37672 93596
rect 37672 93540 37676 93596
rect 37612 93536 37676 93540
rect 37692 93596 37756 93600
rect 37692 93540 37696 93596
rect 37696 93540 37752 93596
rect 37752 93540 37756 93596
rect 37692 93536 37756 93540
rect 37772 93596 37836 93600
rect 37772 93540 37776 93596
rect 37776 93540 37832 93596
rect 37832 93540 37836 93596
rect 37772 93536 37836 93540
rect 37852 93596 37916 93600
rect 37852 93540 37856 93596
rect 37856 93540 37912 93596
rect 37912 93540 37916 93596
rect 37852 93536 37916 93540
rect 73612 93596 73676 93600
rect 73612 93540 73616 93596
rect 73616 93540 73672 93596
rect 73672 93540 73676 93596
rect 73612 93536 73676 93540
rect 73692 93596 73756 93600
rect 73692 93540 73696 93596
rect 73696 93540 73752 93596
rect 73752 93540 73756 93596
rect 73692 93536 73756 93540
rect 73772 93596 73836 93600
rect 73772 93540 73776 93596
rect 73776 93540 73832 93596
rect 73832 93540 73836 93596
rect 73772 93536 73836 93540
rect 73852 93596 73916 93600
rect 73852 93540 73856 93596
rect 73856 93540 73912 93596
rect 73912 93540 73916 93596
rect 73852 93536 73916 93540
rect 36952 93052 37016 93056
rect 36952 92996 36956 93052
rect 36956 92996 37012 93052
rect 37012 92996 37016 93052
rect 36952 92992 37016 92996
rect 37032 93052 37096 93056
rect 37032 92996 37036 93052
rect 37036 92996 37092 93052
rect 37092 92996 37096 93052
rect 37032 92992 37096 92996
rect 37112 93052 37176 93056
rect 37112 92996 37116 93052
rect 37116 92996 37172 93052
rect 37172 92996 37176 93052
rect 37112 92992 37176 92996
rect 37192 93052 37256 93056
rect 37192 92996 37196 93052
rect 37196 92996 37252 93052
rect 37252 92996 37256 93052
rect 37192 92992 37256 92996
rect 72952 93052 73016 93056
rect 72952 92996 72956 93052
rect 72956 92996 73012 93052
rect 73012 92996 73016 93052
rect 72952 92992 73016 92996
rect 73032 93052 73096 93056
rect 73032 92996 73036 93052
rect 73036 92996 73092 93052
rect 73092 92996 73096 93052
rect 73032 92992 73096 92996
rect 73112 93052 73176 93056
rect 73112 92996 73116 93052
rect 73116 92996 73172 93052
rect 73172 92996 73176 93052
rect 73112 92992 73176 92996
rect 73192 93052 73256 93056
rect 73192 92996 73196 93052
rect 73196 92996 73252 93052
rect 73252 92996 73256 93052
rect 73192 92992 73256 92996
rect 48084 92788 48148 92852
rect 47532 92652 47596 92716
rect 89116 92652 89180 92716
rect 86540 92576 86604 92580
rect 86540 92520 86590 92576
rect 86590 92520 86604 92576
rect 86540 92516 86604 92520
rect 87092 92576 87156 92580
rect 87092 92520 87106 92576
rect 87106 92520 87156 92576
rect 87092 92516 87156 92520
rect 37612 92508 37676 92512
rect 37612 92452 37616 92508
rect 37616 92452 37672 92508
rect 37672 92452 37676 92508
rect 37612 92448 37676 92452
rect 37692 92508 37756 92512
rect 37692 92452 37696 92508
rect 37696 92452 37752 92508
rect 37752 92452 37756 92508
rect 37692 92448 37756 92452
rect 37772 92508 37836 92512
rect 37772 92452 37776 92508
rect 37776 92452 37832 92508
rect 37832 92452 37836 92508
rect 37772 92448 37836 92452
rect 37852 92508 37916 92512
rect 37852 92452 37856 92508
rect 37856 92452 37912 92508
rect 37912 92452 37916 92508
rect 37852 92448 37916 92452
rect 73612 92508 73676 92512
rect 73612 92452 73616 92508
rect 73616 92452 73672 92508
rect 73672 92452 73676 92508
rect 73612 92448 73676 92452
rect 73692 92508 73756 92512
rect 73692 92452 73696 92508
rect 73696 92452 73752 92508
rect 73752 92452 73756 92508
rect 73692 92448 73756 92452
rect 73772 92508 73836 92512
rect 73772 92452 73776 92508
rect 73776 92452 73832 92508
rect 73832 92452 73836 92508
rect 73772 92448 73836 92452
rect 73852 92508 73916 92512
rect 73852 92452 73856 92508
rect 73856 92452 73912 92508
rect 73912 92452 73916 92508
rect 73852 92448 73916 92452
rect 89300 92108 89364 92172
rect 3068 91964 3132 91968
rect 3068 91908 3072 91964
rect 3072 91908 3128 91964
rect 3128 91908 3132 91964
rect 3068 91904 3132 91908
rect 3148 91964 3212 91968
rect 3148 91908 3152 91964
rect 3152 91908 3208 91964
rect 3208 91908 3212 91964
rect 3148 91904 3212 91908
rect 3228 91964 3292 91968
rect 3228 91908 3232 91964
rect 3232 91908 3288 91964
rect 3288 91908 3292 91964
rect 3228 91904 3292 91908
rect 3308 91964 3372 91968
rect 3308 91908 3312 91964
rect 3312 91908 3368 91964
rect 3368 91908 3372 91964
rect 3308 91904 3372 91908
rect 36952 91964 37016 91968
rect 36952 91908 36956 91964
rect 36956 91908 37012 91964
rect 37012 91908 37016 91964
rect 36952 91904 37016 91908
rect 37032 91964 37096 91968
rect 37032 91908 37036 91964
rect 37036 91908 37092 91964
rect 37092 91908 37096 91964
rect 37032 91904 37096 91908
rect 37112 91964 37176 91968
rect 37112 91908 37116 91964
rect 37116 91908 37172 91964
rect 37172 91908 37176 91964
rect 37112 91904 37176 91908
rect 37192 91964 37256 91968
rect 37192 91908 37196 91964
rect 37196 91908 37252 91964
rect 37252 91908 37256 91964
rect 37192 91904 37256 91908
rect 72952 91964 73016 91968
rect 72952 91908 72956 91964
rect 72956 91908 73012 91964
rect 73012 91908 73016 91964
rect 72952 91904 73016 91908
rect 73032 91964 73096 91968
rect 73032 91908 73036 91964
rect 73036 91908 73092 91964
rect 73092 91908 73096 91964
rect 73032 91904 73096 91908
rect 73112 91964 73176 91968
rect 73112 91908 73116 91964
rect 73116 91908 73172 91964
rect 73172 91908 73176 91964
rect 73112 91904 73176 91908
rect 73192 91964 73256 91968
rect 73192 91908 73196 91964
rect 73196 91908 73252 91964
rect 73252 91908 73256 91964
rect 73192 91904 73256 91908
rect 86908 91564 86972 91628
rect 3804 91420 3868 91424
rect 3804 91364 3808 91420
rect 3808 91364 3864 91420
rect 3864 91364 3868 91420
rect 3804 91360 3868 91364
rect 3884 91420 3948 91424
rect 3884 91364 3888 91420
rect 3888 91364 3944 91420
rect 3944 91364 3948 91420
rect 3884 91360 3948 91364
rect 3964 91420 4028 91424
rect 3964 91364 3968 91420
rect 3968 91364 4024 91420
rect 4024 91364 4028 91420
rect 3964 91360 4028 91364
rect 4044 91420 4108 91424
rect 4044 91364 4048 91420
rect 4048 91364 4104 91420
rect 4104 91364 4108 91420
rect 4044 91360 4108 91364
rect 37612 91420 37676 91424
rect 37612 91364 37616 91420
rect 37616 91364 37672 91420
rect 37672 91364 37676 91420
rect 37612 91360 37676 91364
rect 37692 91420 37756 91424
rect 37692 91364 37696 91420
rect 37696 91364 37752 91420
rect 37752 91364 37756 91420
rect 37692 91360 37756 91364
rect 37772 91420 37836 91424
rect 37772 91364 37776 91420
rect 37776 91364 37832 91420
rect 37832 91364 37836 91420
rect 37772 91360 37836 91364
rect 37852 91420 37916 91424
rect 37852 91364 37856 91420
rect 37856 91364 37912 91420
rect 37912 91364 37916 91420
rect 37852 91360 37916 91364
rect 73612 91420 73676 91424
rect 73612 91364 73616 91420
rect 73616 91364 73672 91420
rect 73672 91364 73676 91420
rect 73612 91360 73676 91364
rect 73692 91420 73756 91424
rect 73692 91364 73696 91420
rect 73696 91364 73752 91420
rect 73752 91364 73756 91420
rect 73692 91360 73756 91364
rect 73772 91420 73836 91424
rect 73772 91364 73776 91420
rect 73776 91364 73832 91420
rect 73832 91364 73836 91420
rect 73772 91360 73836 91364
rect 73852 91420 73916 91424
rect 73852 91364 73856 91420
rect 73856 91364 73912 91420
rect 73912 91364 73916 91420
rect 73852 91360 73916 91364
rect 86356 91352 86420 91356
rect 86356 91296 86406 91352
rect 86406 91296 86420 91352
rect 86356 91292 86420 91296
rect 86724 91156 86788 91220
rect 3068 90876 3132 90880
rect 3068 90820 3072 90876
rect 3072 90820 3128 90876
rect 3128 90820 3132 90876
rect 3068 90816 3132 90820
rect 3148 90876 3212 90880
rect 3148 90820 3152 90876
rect 3152 90820 3208 90876
rect 3208 90820 3212 90876
rect 3148 90816 3212 90820
rect 3228 90876 3292 90880
rect 3228 90820 3232 90876
rect 3232 90820 3288 90876
rect 3288 90820 3292 90876
rect 3228 90816 3292 90820
rect 3308 90876 3372 90880
rect 3308 90820 3312 90876
rect 3312 90820 3368 90876
rect 3368 90820 3372 90876
rect 3308 90816 3372 90820
rect 3804 90332 3868 90336
rect 3804 90276 3808 90332
rect 3808 90276 3864 90332
rect 3864 90276 3868 90332
rect 3804 90272 3868 90276
rect 3884 90332 3948 90336
rect 3884 90276 3888 90332
rect 3888 90276 3944 90332
rect 3944 90276 3948 90332
rect 3884 90272 3948 90276
rect 3964 90332 4028 90336
rect 3964 90276 3968 90332
rect 3968 90276 4024 90332
rect 4024 90276 4028 90332
rect 3964 90272 4028 90276
rect 4044 90332 4108 90336
rect 4044 90276 4048 90332
rect 4048 90276 4104 90332
rect 4104 90276 4108 90332
rect 4044 90272 4108 90276
rect 88380 89796 88444 89860
rect 3068 89788 3132 89792
rect 3068 89732 3072 89788
rect 3072 89732 3128 89788
rect 3128 89732 3132 89788
rect 3068 89728 3132 89732
rect 3148 89788 3212 89792
rect 3148 89732 3152 89788
rect 3152 89732 3208 89788
rect 3208 89732 3212 89788
rect 3148 89728 3212 89732
rect 3228 89788 3292 89792
rect 3228 89732 3232 89788
rect 3232 89732 3288 89788
rect 3288 89732 3292 89788
rect 3228 89728 3292 89732
rect 3308 89788 3372 89792
rect 3308 89732 3312 89788
rect 3312 89732 3368 89788
rect 3368 89732 3372 89788
rect 3308 89728 3372 89732
rect 3804 89244 3868 89248
rect 3804 89188 3808 89244
rect 3808 89188 3864 89244
rect 3864 89188 3868 89244
rect 3804 89184 3868 89188
rect 3884 89244 3948 89248
rect 3884 89188 3888 89244
rect 3888 89188 3944 89244
rect 3944 89188 3948 89244
rect 3884 89184 3948 89188
rect 3964 89244 4028 89248
rect 3964 89188 3968 89244
rect 3968 89188 4024 89244
rect 4024 89188 4028 89244
rect 3964 89184 4028 89188
rect 4044 89244 4108 89248
rect 4044 89188 4048 89244
rect 4048 89188 4104 89244
rect 4104 89188 4108 89244
rect 4044 89184 4108 89188
rect 3068 88700 3132 88704
rect 3068 88644 3072 88700
rect 3072 88644 3128 88700
rect 3128 88644 3132 88700
rect 3068 88640 3132 88644
rect 3148 88700 3212 88704
rect 3148 88644 3152 88700
rect 3152 88644 3208 88700
rect 3208 88644 3212 88700
rect 3148 88640 3212 88644
rect 3228 88700 3292 88704
rect 3228 88644 3232 88700
rect 3232 88644 3288 88700
rect 3288 88644 3292 88700
rect 3228 88640 3292 88644
rect 3308 88700 3372 88704
rect 3308 88644 3312 88700
rect 3312 88644 3368 88700
rect 3368 88644 3372 88700
rect 3308 88640 3372 88644
rect 87276 88436 87340 88500
rect 47716 88300 47780 88364
rect 3804 88156 3868 88160
rect 3804 88100 3808 88156
rect 3808 88100 3864 88156
rect 3864 88100 3868 88156
rect 3804 88096 3868 88100
rect 3884 88156 3948 88160
rect 3884 88100 3888 88156
rect 3888 88100 3944 88156
rect 3944 88100 3948 88156
rect 3884 88096 3948 88100
rect 3964 88156 4028 88160
rect 3964 88100 3968 88156
rect 3968 88100 4024 88156
rect 4024 88100 4028 88156
rect 3964 88096 4028 88100
rect 4044 88156 4108 88160
rect 4044 88100 4048 88156
rect 4048 88100 4104 88156
rect 4104 88100 4108 88156
rect 4044 88096 4108 88100
rect 8524 87892 8588 87956
rect 3068 87612 3132 87616
rect 3068 87556 3072 87612
rect 3072 87556 3128 87612
rect 3128 87556 3132 87612
rect 3068 87552 3132 87556
rect 3148 87612 3212 87616
rect 3148 87556 3152 87612
rect 3152 87556 3208 87612
rect 3208 87556 3212 87612
rect 3148 87552 3212 87556
rect 3228 87612 3292 87616
rect 3228 87556 3232 87612
rect 3232 87556 3288 87612
rect 3288 87556 3292 87612
rect 3228 87552 3292 87556
rect 3308 87612 3372 87616
rect 3308 87556 3312 87612
rect 3312 87556 3368 87612
rect 3368 87556 3372 87612
rect 3308 87552 3372 87556
rect 86540 87212 86604 87276
rect 86908 87076 86972 87140
rect 3804 87068 3868 87072
rect 3804 87012 3808 87068
rect 3808 87012 3864 87068
rect 3864 87012 3868 87068
rect 3804 87008 3868 87012
rect 3884 87068 3948 87072
rect 3884 87012 3888 87068
rect 3888 87012 3944 87068
rect 3944 87012 3948 87068
rect 3884 87008 3948 87012
rect 3964 87068 4028 87072
rect 3964 87012 3968 87068
rect 3968 87012 4024 87068
rect 4024 87012 4028 87068
rect 3964 87008 4028 87012
rect 4044 87068 4108 87072
rect 4044 87012 4048 87068
rect 4048 87012 4104 87068
rect 4104 87012 4108 87068
rect 4044 87008 4108 87012
rect 86724 86940 86788 87004
rect 3068 86524 3132 86528
rect 3068 86468 3072 86524
rect 3072 86468 3128 86524
rect 3128 86468 3132 86524
rect 3068 86464 3132 86468
rect 3148 86524 3212 86528
rect 3148 86468 3152 86524
rect 3152 86468 3208 86524
rect 3208 86468 3212 86524
rect 3148 86464 3212 86468
rect 3228 86524 3292 86528
rect 3228 86468 3232 86524
rect 3232 86468 3288 86524
rect 3288 86468 3292 86524
rect 3228 86464 3292 86468
rect 3308 86524 3372 86528
rect 3308 86468 3312 86524
rect 3312 86468 3368 86524
rect 3368 86468 3372 86524
rect 3308 86464 3372 86468
rect 3804 85980 3868 85984
rect 3804 85924 3808 85980
rect 3808 85924 3864 85980
rect 3864 85924 3868 85980
rect 3804 85920 3868 85924
rect 3884 85980 3948 85984
rect 3884 85924 3888 85980
rect 3888 85924 3944 85980
rect 3944 85924 3948 85980
rect 3884 85920 3948 85924
rect 3964 85980 4028 85984
rect 3964 85924 3968 85980
rect 3968 85924 4024 85980
rect 4024 85924 4028 85980
rect 3964 85920 4028 85924
rect 4044 85980 4108 85984
rect 4044 85924 4048 85980
rect 4048 85924 4104 85980
rect 4104 85924 4108 85980
rect 4044 85920 4108 85924
rect 86908 85912 86972 85916
rect 86908 85856 86922 85912
rect 86922 85856 86972 85912
rect 86908 85852 86972 85856
rect 3068 85436 3132 85440
rect 3068 85380 3072 85436
rect 3072 85380 3128 85436
rect 3128 85380 3132 85436
rect 3068 85376 3132 85380
rect 3148 85436 3212 85440
rect 3148 85380 3152 85436
rect 3152 85380 3208 85436
rect 3208 85380 3212 85436
rect 3148 85376 3212 85380
rect 3228 85436 3292 85440
rect 3228 85380 3232 85436
rect 3232 85380 3288 85436
rect 3288 85380 3292 85436
rect 3228 85376 3292 85380
rect 3308 85436 3372 85440
rect 3308 85380 3312 85436
rect 3312 85380 3368 85436
rect 3368 85380 3372 85436
rect 3308 85376 3372 85380
rect 3804 84892 3868 84896
rect 3804 84836 3808 84892
rect 3808 84836 3864 84892
rect 3864 84836 3868 84892
rect 3804 84832 3868 84836
rect 3884 84892 3948 84896
rect 3884 84836 3888 84892
rect 3888 84836 3944 84892
rect 3944 84836 3948 84892
rect 3884 84832 3948 84836
rect 3964 84892 4028 84896
rect 3964 84836 3968 84892
rect 3968 84836 4024 84892
rect 4024 84836 4028 84892
rect 3964 84832 4028 84836
rect 4044 84892 4108 84896
rect 4044 84836 4048 84892
rect 4048 84836 4104 84892
rect 4104 84836 4108 84892
rect 4044 84832 4108 84836
rect 3068 84348 3132 84352
rect 3068 84292 3072 84348
rect 3072 84292 3128 84348
rect 3128 84292 3132 84348
rect 3068 84288 3132 84292
rect 3148 84348 3212 84352
rect 3148 84292 3152 84348
rect 3152 84292 3208 84348
rect 3208 84292 3212 84348
rect 3148 84288 3212 84292
rect 3228 84348 3292 84352
rect 3228 84292 3232 84348
rect 3232 84292 3288 84348
rect 3288 84292 3292 84348
rect 3228 84288 3292 84292
rect 3308 84348 3372 84352
rect 3308 84292 3312 84348
rect 3312 84292 3368 84348
rect 3368 84292 3372 84348
rect 3308 84288 3372 84292
rect 3804 83804 3868 83808
rect 3804 83748 3808 83804
rect 3808 83748 3864 83804
rect 3864 83748 3868 83804
rect 3804 83744 3868 83748
rect 3884 83804 3948 83808
rect 3884 83748 3888 83804
rect 3888 83748 3944 83804
rect 3944 83748 3948 83804
rect 3884 83744 3948 83748
rect 3964 83804 4028 83808
rect 3964 83748 3968 83804
rect 3968 83748 4024 83804
rect 4024 83748 4028 83804
rect 3964 83744 4028 83748
rect 4044 83804 4108 83808
rect 4044 83748 4048 83804
rect 4048 83748 4104 83804
rect 4104 83748 4108 83804
rect 4044 83744 4108 83748
rect 3068 83260 3132 83264
rect 3068 83204 3072 83260
rect 3072 83204 3128 83260
rect 3128 83204 3132 83260
rect 3068 83200 3132 83204
rect 3148 83260 3212 83264
rect 3148 83204 3152 83260
rect 3152 83204 3208 83260
rect 3208 83204 3212 83260
rect 3148 83200 3212 83204
rect 3228 83260 3292 83264
rect 3228 83204 3232 83260
rect 3232 83204 3288 83260
rect 3288 83204 3292 83260
rect 3228 83200 3292 83204
rect 3308 83260 3372 83264
rect 3308 83204 3312 83260
rect 3312 83204 3368 83260
rect 3368 83204 3372 83260
rect 3308 83200 3372 83204
rect 3804 82716 3868 82720
rect 3804 82660 3808 82716
rect 3808 82660 3864 82716
rect 3864 82660 3868 82716
rect 3804 82656 3868 82660
rect 3884 82716 3948 82720
rect 3884 82660 3888 82716
rect 3888 82660 3944 82716
rect 3944 82660 3948 82716
rect 3884 82656 3948 82660
rect 3964 82716 4028 82720
rect 3964 82660 3968 82716
rect 3968 82660 4024 82716
rect 4024 82660 4028 82716
rect 3964 82656 4028 82660
rect 4044 82716 4108 82720
rect 4044 82660 4048 82716
rect 4048 82660 4104 82716
rect 4104 82660 4108 82716
rect 4044 82656 4108 82660
rect 3068 82172 3132 82176
rect 3068 82116 3072 82172
rect 3072 82116 3128 82172
rect 3128 82116 3132 82172
rect 3068 82112 3132 82116
rect 3148 82172 3212 82176
rect 3148 82116 3152 82172
rect 3152 82116 3208 82172
rect 3208 82116 3212 82172
rect 3148 82112 3212 82116
rect 3228 82172 3292 82176
rect 3228 82116 3232 82172
rect 3232 82116 3288 82172
rect 3288 82116 3292 82172
rect 3228 82112 3292 82116
rect 3308 82172 3372 82176
rect 3308 82116 3312 82172
rect 3312 82116 3368 82172
rect 3368 82116 3372 82172
rect 3308 82112 3372 82116
rect 3804 81628 3868 81632
rect 3804 81572 3808 81628
rect 3808 81572 3864 81628
rect 3864 81572 3868 81628
rect 3804 81568 3868 81572
rect 3884 81628 3948 81632
rect 3884 81572 3888 81628
rect 3888 81572 3944 81628
rect 3944 81572 3948 81628
rect 3884 81568 3948 81572
rect 3964 81628 4028 81632
rect 3964 81572 3968 81628
rect 3968 81572 4024 81628
rect 4024 81572 4028 81628
rect 3964 81568 4028 81572
rect 4044 81628 4108 81632
rect 4044 81572 4048 81628
rect 4048 81572 4104 81628
rect 4104 81572 4108 81628
rect 4044 81568 4108 81572
rect 3068 81084 3132 81088
rect 3068 81028 3072 81084
rect 3072 81028 3128 81084
rect 3128 81028 3132 81084
rect 3068 81024 3132 81028
rect 3148 81084 3212 81088
rect 3148 81028 3152 81084
rect 3152 81028 3208 81084
rect 3208 81028 3212 81084
rect 3148 81024 3212 81028
rect 3228 81084 3292 81088
rect 3228 81028 3232 81084
rect 3232 81028 3288 81084
rect 3288 81028 3292 81084
rect 3228 81024 3292 81028
rect 3308 81084 3372 81088
rect 3308 81028 3312 81084
rect 3312 81028 3368 81084
rect 3368 81028 3372 81084
rect 3308 81024 3372 81028
rect 3804 80540 3868 80544
rect 3804 80484 3808 80540
rect 3808 80484 3864 80540
rect 3864 80484 3868 80540
rect 3804 80480 3868 80484
rect 3884 80540 3948 80544
rect 3884 80484 3888 80540
rect 3888 80484 3944 80540
rect 3944 80484 3948 80540
rect 3884 80480 3948 80484
rect 3964 80540 4028 80544
rect 3964 80484 3968 80540
rect 3968 80484 4024 80540
rect 4024 80484 4028 80540
rect 3964 80480 4028 80484
rect 4044 80540 4108 80544
rect 4044 80484 4048 80540
rect 4048 80484 4104 80540
rect 4104 80484 4108 80540
rect 4044 80480 4108 80484
rect 3068 79996 3132 80000
rect 3068 79940 3072 79996
rect 3072 79940 3128 79996
rect 3128 79940 3132 79996
rect 3068 79936 3132 79940
rect 3148 79996 3212 80000
rect 3148 79940 3152 79996
rect 3152 79940 3208 79996
rect 3208 79940 3212 79996
rect 3148 79936 3212 79940
rect 3228 79996 3292 80000
rect 3228 79940 3232 79996
rect 3232 79940 3288 79996
rect 3288 79940 3292 79996
rect 3228 79936 3292 79940
rect 3308 79996 3372 80000
rect 3308 79940 3312 79996
rect 3312 79940 3368 79996
rect 3368 79940 3372 79996
rect 3308 79936 3372 79940
rect 3804 79452 3868 79456
rect 3804 79396 3808 79452
rect 3808 79396 3864 79452
rect 3864 79396 3868 79452
rect 3804 79392 3868 79396
rect 3884 79452 3948 79456
rect 3884 79396 3888 79452
rect 3888 79396 3944 79452
rect 3944 79396 3948 79452
rect 3884 79392 3948 79396
rect 3964 79452 4028 79456
rect 3964 79396 3968 79452
rect 3968 79396 4024 79452
rect 4024 79396 4028 79452
rect 3964 79392 4028 79396
rect 4044 79452 4108 79456
rect 4044 79396 4048 79452
rect 4048 79396 4104 79452
rect 4104 79396 4108 79452
rect 4044 79392 4108 79396
rect 3068 78908 3132 78912
rect 3068 78852 3072 78908
rect 3072 78852 3128 78908
rect 3128 78852 3132 78908
rect 3068 78848 3132 78852
rect 3148 78908 3212 78912
rect 3148 78852 3152 78908
rect 3152 78852 3208 78908
rect 3208 78852 3212 78908
rect 3148 78848 3212 78852
rect 3228 78908 3292 78912
rect 3228 78852 3232 78908
rect 3232 78852 3288 78908
rect 3288 78852 3292 78908
rect 3228 78848 3292 78852
rect 3308 78908 3372 78912
rect 3308 78852 3312 78908
rect 3312 78852 3368 78908
rect 3368 78852 3372 78908
rect 3308 78848 3372 78852
rect 3804 78364 3868 78368
rect 3804 78308 3808 78364
rect 3808 78308 3864 78364
rect 3864 78308 3868 78364
rect 3804 78304 3868 78308
rect 3884 78364 3948 78368
rect 3884 78308 3888 78364
rect 3888 78308 3944 78364
rect 3944 78308 3948 78364
rect 3884 78304 3948 78308
rect 3964 78364 4028 78368
rect 3964 78308 3968 78364
rect 3968 78308 4024 78364
rect 4024 78308 4028 78364
rect 3964 78304 4028 78308
rect 4044 78364 4108 78368
rect 4044 78308 4048 78364
rect 4048 78308 4104 78364
rect 4104 78308 4108 78364
rect 4044 78304 4108 78308
rect 3068 77820 3132 77824
rect 3068 77764 3072 77820
rect 3072 77764 3128 77820
rect 3128 77764 3132 77820
rect 3068 77760 3132 77764
rect 3148 77820 3212 77824
rect 3148 77764 3152 77820
rect 3152 77764 3208 77820
rect 3208 77764 3212 77820
rect 3148 77760 3212 77764
rect 3228 77820 3292 77824
rect 3228 77764 3232 77820
rect 3232 77764 3288 77820
rect 3288 77764 3292 77820
rect 3228 77760 3292 77764
rect 3308 77820 3372 77824
rect 3308 77764 3312 77820
rect 3312 77764 3368 77820
rect 3368 77764 3372 77820
rect 3308 77760 3372 77764
rect 3804 77276 3868 77280
rect 3804 77220 3808 77276
rect 3808 77220 3864 77276
rect 3864 77220 3868 77276
rect 3804 77216 3868 77220
rect 3884 77276 3948 77280
rect 3884 77220 3888 77276
rect 3888 77220 3944 77276
rect 3944 77220 3948 77276
rect 3884 77216 3948 77220
rect 3964 77276 4028 77280
rect 3964 77220 3968 77276
rect 3968 77220 4024 77276
rect 4024 77220 4028 77276
rect 3964 77216 4028 77220
rect 4044 77276 4108 77280
rect 4044 77220 4048 77276
rect 4048 77220 4104 77276
rect 4104 77220 4108 77276
rect 4044 77216 4108 77220
rect 86356 77012 86420 77076
rect 3068 76732 3132 76736
rect 3068 76676 3072 76732
rect 3072 76676 3128 76732
rect 3128 76676 3132 76732
rect 3068 76672 3132 76676
rect 3148 76732 3212 76736
rect 3148 76676 3152 76732
rect 3152 76676 3208 76732
rect 3208 76676 3212 76732
rect 3148 76672 3212 76676
rect 3228 76732 3292 76736
rect 3228 76676 3232 76732
rect 3232 76676 3288 76732
rect 3288 76676 3292 76732
rect 3228 76672 3292 76676
rect 3308 76732 3372 76736
rect 3308 76676 3312 76732
rect 3312 76676 3368 76732
rect 3368 76676 3372 76732
rect 3308 76672 3372 76676
rect 3804 76188 3868 76192
rect 3804 76132 3808 76188
rect 3808 76132 3864 76188
rect 3864 76132 3868 76188
rect 3804 76128 3868 76132
rect 3884 76188 3948 76192
rect 3884 76132 3888 76188
rect 3888 76132 3944 76188
rect 3944 76132 3948 76188
rect 3884 76128 3948 76132
rect 3964 76188 4028 76192
rect 3964 76132 3968 76188
rect 3968 76132 4024 76188
rect 4024 76132 4028 76188
rect 3964 76128 4028 76132
rect 4044 76188 4108 76192
rect 4044 76132 4048 76188
rect 4048 76132 4104 76188
rect 4104 76132 4108 76188
rect 4044 76128 4108 76132
rect 3068 75644 3132 75648
rect 3068 75588 3072 75644
rect 3072 75588 3128 75644
rect 3128 75588 3132 75644
rect 3068 75584 3132 75588
rect 3148 75644 3212 75648
rect 3148 75588 3152 75644
rect 3152 75588 3208 75644
rect 3208 75588 3212 75644
rect 3148 75584 3212 75588
rect 3228 75644 3292 75648
rect 3228 75588 3232 75644
rect 3232 75588 3288 75644
rect 3288 75588 3292 75644
rect 3228 75584 3292 75588
rect 3308 75644 3372 75648
rect 3308 75588 3312 75644
rect 3312 75588 3368 75644
rect 3368 75588 3372 75644
rect 3308 75584 3372 75588
rect 3804 75100 3868 75104
rect 3804 75044 3808 75100
rect 3808 75044 3864 75100
rect 3864 75044 3868 75100
rect 3804 75040 3868 75044
rect 3884 75100 3948 75104
rect 3884 75044 3888 75100
rect 3888 75044 3944 75100
rect 3944 75044 3948 75100
rect 3884 75040 3948 75044
rect 3964 75100 4028 75104
rect 3964 75044 3968 75100
rect 3968 75044 4024 75100
rect 4024 75044 4028 75100
rect 3964 75040 4028 75044
rect 4044 75100 4108 75104
rect 4044 75044 4048 75100
rect 4048 75044 4104 75100
rect 4104 75044 4108 75100
rect 4044 75040 4108 75044
rect 3068 74556 3132 74560
rect 3068 74500 3072 74556
rect 3072 74500 3128 74556
rect 3128 74500 3132 74556
rect 3068 74496 3132 74500
rect 3148 74556 3212 74560
rect 3148 74500 3152 74556
rect 3152 74500 3208 74556
rect 3208 74500 3212 74556
rect 3148 74496 3212 74500
rect 3228 74556 3292 74560
rect 3228 74500 3232 74556
rect 3232 74500 3288 74556
rect 3288 74500 3292 74556
rect 3228 74496 3292 74500
rect 3308 74556 3372 74560
rect 3308 74500 3312 74556
rect 3312 74500 3368 74556
rect 3368 74500 3372 74556
rect 3308 74496 3372 74500
rect 89116 74292 89180 74356
rect 3804 74012 3868 74016
rect 3804 73956 3808 74012
rect 3808 73956 3864 74012
rect 3864 73956 3868 74012
rect 3804 73952 3868 73956
rect 3884 74012 3948 74016
rect 3884 73956 3888 74012
rect 3888 73956 3944 74012
rect 3944 73956 3948 74012
rect 3884 73952 3948 73956
rect 3964 74012 4028 74016
rect 3964 73956 3968 74012
rect 3968 73956 4024 74012
rect 4024 73956 4028 74012
rect 3964 73952 4028 73956
rect 4044 74012 4108 74016
rect 4044 73956 4048 74012
rect 4048 73956 4104 74012
rect 4104 73956 4108 74012
rect 4044 73952 4108 73956
rect 3068 73468 3132 73472
rect 3068 73412 3072 73468
rect 3072 73412 3128 73468
rect 3128 73412 3132 73468
rect 3068 73408 3132 73412
rect 3148 73468 3212 73472
rect 3148 73412 3152 73468
rect 3152 73412 3208 73468
rect 3208 73412 3212 73468
rect 3148 73408 3212 73412
rect 3228 73468 3292 73472
rect 3228 73412 3232 73468
rect 3232 73412 3288 73468
rect 3288 73412 3292 73468
rect 3228 73408 3292 73412
rect 3308 73468 3372 73472
rect 3308 73412 3312 73468
rect 3312 73412 3368 73468
rect 3368 73412 3372 73468
rect 3308 73408 3372 73412
rect 3804 72924 3868 72928
rect 3804 72868 3808 72924
rect 3808 72868 3864 72924
rect 3864 72868 3868 72924
rect 3804 72864 3868 72868
rect 3884 72924 3948 72928
rect 3884 72868 3888 72924
rect 3888 72868 3944 72924
rect 3944 72868 3948 72924
rect 3884 72864 3948 72868
rect 3964 72924 4028 72928
rect 3964 72868 3968 72924
rect 3968 72868 4024 72924
rect 4024 72868 4028 72924
rect 3964 72864 4028 72868
rect 4044 72924 4108 72928
rect 4044 72868 4048 72924
rect 4048 72868 4104 72924
rect 4104 72868 4108 72924
rect 4044 72864 4108 72868
rect 89162 72796 89226 72860
rect 3068 72380 3132 72384
rect 3068 72324 3072 72380
rect 3072 72324 3128 72380
rect 3128 72324 3132 72380
rect 3068 72320 3132 72324
rect 3148 72380 3212 72384
rect 3148 72324 3152 72380
rect 3152 72324 3208 72380
rect 3208 72324 3212 72380
rect 3148 72320 3212 72324
rect 3228 72380 3292 72384
rect 3228 72324 3232 72380
rect 3232 72324 3288 72380
rect 3288 72324 3292 72380
rect 3228 72320 3292 72324
rect 3308 72380 3372 72384
rect 3308 72324 3312 72380
rect 3312 72324 3368 72380
rect 3368 72324 3372 72380
rect 3308 72320 3372 72324
rect 3804 71836 3868 71840
rect 3804 71780 3808 71836
rect 3808 71780 3864 71836
rect 3864 71780 3868 71836
rect 3804 71776 3868 71780
rect 3884 71836 3948 71840
rect 3884 71780 3888 71836
rect 3888 71780 3944 71836
rect 3944 71780 3948 71836
rect 3884 71776 3948 71780
rect 3964 71836 4028 71840
rect 3964 71780 3968 71836
rect 3968 71780 4024 71836
rect 4024 71780 4028 71836
rect 3964 71776 4028 71780
rect 4044 71836 4108 71840
rect 4044 71780 4048 71836
rect 4048 71780 4104 71836
rect 4104 71780 4108 71836
rect 4044 71776 4108 71780
rect 3068 71292 3132 71296
rect 3068 71236 3072 71292
rect 3072 71236 3128 71292
rect 3128 71236 3132 71292
rect 3068 71232 3132 71236
rect 3148 71292 3212 71296
rect 3148 71236 3152 71292
rect 3152 71236 3208 71292
rect 3208 71236 3212 71292
rect 3148 71232 3212 71236
rect 3228 71292 3292 71296
rect 3228 71236 3232 71292
rect 3232 71236 3288 71292
rect 3288 71236 3292 71292
rect 3228 71232 3292 71236
rect 3308 71292 3372 71296
rect 3308 71236 3312 71292
rect 3312 71236 3368 71292
rect 3368 71236 3372 71292
rect 3308 71232 3372 71236
rect 3804 70748 3868 70752
rect 3804 70692 3808 70748
rect 3808 70692 3864 70748
rect 3864 70692 3868 70748
rect 3804 70688 3868 70692
rect 3884 70748 3948 70752
rect 3884 70692 3888 70748
rect 3888 70692 3944 70748
rect 3944 70692 3948 70748
rect 3884 70688 3948 70692
rect 3964 70748 4028 70752
rect 3964 70692 3968 70748
rect 3968 70692 4024 70748
rect 4024 70692 4028 70748
rect 3964 70688 4028 70692
rect 4044 70748 4108 70752
rect 4044 70692 4048 70748
rect 4048 70692 4104 70748
rect 4104 70692 4108 70748
rect 4044 70688 4108 70692
rect 3068 70204 3132 70208
rect 3068 70148 3072 70204
rect 3072 70148 3128 70204
rect 3128 70148 3132 70204
rect 3068 70144 3132 70148
rect 3148 70204 3212 70208
rect 3148 70148 3152 70204
rect 3152 70148 3208 70204
rect 3208 70148 3212 70204
rect 3148 70144 3212 70148
rect 3228 70204 3292 70208
rect 3228 70148 3232 70204
rect 3232 70148 3288 70204
rect 3288 70148 3292 70204
rect 3228 70144 3292 70148
rect 3308 70204 3372 70208
rect 3308 70148 3312 70204
rect 3312 70148 3368 70204
rect 3368 70148 3372 70204
rect 3308 70144 3372 70148
rect 3804 69660 3868 69664
rect 3804 69604 3808 69660
rect 3808 69604 3864 69660
rect 3864 69604 3868 69660
rect 3804 69600 3868 69604
rect 3884 69660 3948 69664
rect 3884 69604 3888 69660
rect 3888 69604 3944 69660
rect 3944 69604 3948 69660
rect 3884 69600 3948 69604
rect 3964 69660 4028 69664
rect 3964 69604 3968 69660
rect 3968 69604 4024 69660
rect 4024 69604 4028 69660
rect 3964 69600 4028 69604
rect 4044 69660 4108 69664
rect 4044 69604 4048 69660
rect 4048 69604 4104 69660
rect 4104 69604 4108 69660
rect 4044 69600 4108 69604
rect 3068 69116 3132 69120
rect 3068 69060 3072 69116
rect 3072 69060 3128 69116
rect 3128 69060 3132 69116
rect 3068 69056 3132 69060
rect 3148 69116 3212 69120
rect 3148 69060 3152 69116
rect 3152 69060 3208 69116
rect 3208 69060 3212 69116
rect 3148 69056 3212 69060
rect 3228 69116 3292 69120
rect 3228 69060 3232 69116
rect 3232 69060 3288 69116
rect 3288 69060 3292 69116
rect 3228 69056 3292 69060
rect 3308 69116 3372 69120
rect 3308 69060 3312 69116
rect 3312 69060 3368 69116
rect 3368 69060 3372 69116
rect 3308 69056 3372 69060
rect 3804 68572 3868 68576
rect 3804 68516 3808 68572
rect 3808 68516 3864 68572
rect 3864 68516 3868 68572
rect 3804 68512 3868 68516
rect 3884 68572 3948 68576
rect 3884 68516 3888 68572
rect 3888 68516 3944 68572
rect 3944 68516 3948 68572
rect 3884 68512 3948 68516
rect 3964 68572 4028 68576
rect 3964 68516 3968 68572
rect 3968 68516 4024 68572
rect 4024 68516 4028 68572
rect 3964 68512 4028 68516
rect 4044 68572 4108 68576
rect 4044 68516 4048 68572
rect 4048 68516 4104 68572
rect 4104 68516 4108 68572
rect 4044 68512 4108 68516
rect 3068 68028 3132 68032
rect 3068 67972 3072 68028
rect 3072 67972 3128 68028
rect 3128 67972 3132 68028
rect 3068 67968 3132 67972
rect 3148 68028 3212 68032
rect 3148 67972 3152 68028
rect 3152 67972 3208 68028
rect 3208 67972 3212 68028
rect 3148 67968 3212 67972
rect 3228 68028 3292 68032
rect 3228 67972 3232 68028
rect 3232 67972 3288 68028
rect 3288 67972 3292 68028
rect 3228 67968 3292 67972
rect 3308 68028 3372 68032
rect 3308 67972 3312 68028
rect 3312 67972 3368 68028
rect 3368 67972 3372 68028
rect 3308 67968 3372 67972
rect 5580 67688 5644 67692
rect 5580 67632 5594 67688
rect 5594 67632 5644 67688
rect 5580 67628 5644 67632
rect 88380 67492 88444 67556
rect 3804 67484 3868 67488
rect 3804 67428 3808 67484
rect 3808 67428 3864 67484
rect 3864 67428 3868 67484
rect 3804 67424 3868 67428
rect 3884 67484 3948 67488
rect 3884 67428 3888 67484
rect 3888 67428 3944 67484
rect 3944 67428 3948 67484
rect 3884 67424 3948 67428
rect 3964 67484 4028 67488
rect 3964 67428 3968 67484
rect 3968 67428 4024 67484
rect 4024 67428 4028 67484
rect 3964 67424 4028 67428
rect 4044 67484 4108 67488
rect 4044 67428 4048 67484
rect 4048 67428 4104 67484
rect 4104 67428 4108 67484
rect 4044 67424 4108 67428
rect 3068 66940 3132 66944
rect 3068 66884 3072 66940
rect 3072 66884 3128 66940
rect 3128 66884 3132 66940
rect 3068 66880 3132 66884
rect 3148 66940 3212 66944
rect 3148 66884 3152 66940
rect 3152 66884 3208 66940
rect 3208 66884 3212 66940
rect 3148 66880 3212 66884
rect 3228 66940 3292 66944
rect 3228 66884 3232 66940
rect 3232 66884 3288 66940
rect 3288 66884 3292 66940
rect 3228 66880 3292 66884
rect 3308 66940 3372 66944
rect 3308 66884 3312 66940
rect 3312 66884 3368 66940
rect 3368 66884 3372 66940
rect 3308 66880 3372 66884
rect 3804 66396 3868 66400
rect 3804 66340 3808 66396
rect 3808 66340 3864 66396
rect 3864 66340 3868 66396
rect 3804 66336 3868 66340
rect 3884 66396 3948 66400
rect 3884 66340 3888 66396
rect 3888 66340 3944 66396
rect 3944 66340 3948 66396
rect 3884 66336 3948 66340
rect 3964 66396 4028 66400
rect 3964 66340 3968 66396
rect 3968 66340 4024 66396
rect 4024 66340 4028 66396
rect 3964 66336 4028 66340
rect 4044 66396 4108 66400
rect 4044 66340 4048 66396
rect 4048 66340 4104 66396
rect 4104 66340 4108 66396
rect 4044 66336 4108 66340
rect 86356 66132 86420 66196
rect 3068 65852 3132 65856
rect 3068 65796 3072 65852
rect 3072 65796 3128 65852
rect 3128 65796 3132 65852
rect 3068 65792 3132 65796
rect 3148 65852 3212 65856
rect 3148 65796 3152 65852
rect 3152 65796 3208 65852
rect 3208 65796 3212 65852
rect 3148 65792 3212 65796
rect 3228 65852 3292 65856
rect 3228 65796 3232 65852
rect 3232 65796 3288 65852
rect 3288 65796 3292 65852
rect 3228 65792 3292 65796
rect 3308 65852 3372 65856
rect 3308 65796 3312 65852
rect 3312 65796 3368 65852
rect 3368 65796 3372 65852
rect 3308 65792 3372 65796
rect 3804 65308 3868 65312
rect 3804 65252 3808 65308
rect 3808 65252 3864 65308
rect 3864 65252 3868 65308
rect 3804 65248 3868 65252
rect 3884 65308 3948 65312
rect 3884 65252 3888 65308
rect 3888 65252 3944 65308
rect 3944 65252 3948 65308
rect 3884 65248 3948 65252
rect 3964 65308 4028 65312
rect 3964 65252 3968 65308
rect 3968 65252 4024 65308
rect 4024 65252 4028 65308
rect 3964 65248 4028 65252
rect 4044 65308 4108 65312
rect 4044 65252 4048 65308
rect 4048 65252 4104 65308
rect 4104 65252 4108 65308
rect 4044 65248 4108 65252
rect 5764 64908 5828 64972
rect 87276 64772 87340 64836
rect 3068 64764 3132 64768
rect 3068 64708 3072 64764
rect 3072 64708 3128 64764
rect 3128 64708 3132 64764
rect 3068 64704 3132 64708
rect 3148 64764 3212 64768
rect 3148 64708 3152 64764
rect 3152 64708 3208 64764
rect 3208 64708 3212 64764
rect 3148 64704 3212 64708
rect 3228 64764 3292 64768
rect 3228 64708 3232 64764
rect 3232 64708 3288 64764
rect 3288 64708 3292 64764
rect 3228 64704 3292 64708
rect 3308 64764 3372 64768
rect 3308 64708 3312 64764
rect 3312 64708 3368 64764
rect 3368 64708 3372 64764
rect 3308 64704 3372 64708
rect 3804 64220 3868 64224
rect 3804 64164 3808 64220
rect 3808 64164 3864 64220
rect 3864 64164 3868 64220
rect 3804 64160 3868 64164
rect 3884 64220 3948 64224
rect 3884 64164 3888 64220
rect 3888 64164 3944 64220
rect 3944 64164 3948 64220
rect 3884 64160 3948 64164
rect 3964 64220 4028 64224
rect 3964 64164 3968 64220
rect 3968 64164 4024 64220
rect 4024 64164 4028 64220
rect 3964 64160 4028 64164
rect 4044 64220 4108 64224
rect 4044 64164 4048 64220
rect 4048 64164 4104 64220
rect 4104 64164 4108 64220
rect 4044 64160 4108 64164
rect 3068 63676 3132 63680
rect 3068 63620 3072 63676
rect 3072 63620 3128 63676
rect 3128 63620 3132 63676
rect 3068 63616 3132 63620
rect 3148 63676 3212 63680
rect 3148 63620 3152 63676
rect 3152 63620 3208 63676
rect 3208 63620 3212 63676
rect 3148 63616 3212 63620
rect 3228 63676 3292 63680
rect 3228 63620 3232 63676
rect 3232 63620 3288 63676
rect 3288 63620 3292 63676
rect 3228 63616 3292 63620
rect 3308 63676 3372 63680
rect 3308 63620 3312 63676
rect 3312 63620 3368 63676
rect 3368 63620 3372 63676
rect 3308 63616 3372 63620
rect 86540 63412 86604 63476
rect 3804 63132 3868 63136
rect 3804 63076 3808 63132
rect 3808 63076 3864 63132
rect 3864 63076 3868 63132
rect 3804 63072 3868 63076
rect 3884 63132 3948 63136
rect 3884 63076 3888 63132
rect 3888 63076 3944 63132
rect 3944 63076 3948 63132
rect 3884 63072 3948 63076
rect 3964 63132 4028 63136
rect 3964 63076 3968 63132
rect 3968 63076 4024 63132
rect 4024 63076 4028 63132
rect 3964 63072 4028 63076
rect 4044 63132 4108 63136
rect 4044 63076 4048 63132
rect 4048 63076 4104 63132
rect 4104 63076 4108 63132
rect 4044 63072 4108 63076
rect 3068 62588 3132 62592
rect 3068 62532 3072 62588
rect 3072 62532 3128 62588
rect 3128 62532 3132 62588
rect 3068 62528 3132 62532
rect 3148 62588 3212 62592
rect 3148 62532 3152 62588
rect 3152 62532 3208 62588
rect 3208 62532 3212 62588
rect 3148 62528 3212 62532
rect 3228 62588 3292 62592
rect 3228 62532 3232 62588
rect 3232 62532 3288 62588
rect 3288 62532 3292 62588
rect 3228 62528 3292 62532
rect 3308 62588 3372 62592
rect 3308 62532 3312 62588
rect 3312 62532 3368 62588
rect 3368 62532 3372 62588
rect 3308 62528 3372 62532
rect 5948 62248 6012 62252
rect 5948 62192 5962 62248
rect 5962 62192 6012 62248
rect 5948 62188 6012 62192
rect 3804 62044 3868 62048
rect 3804 61988 3808 62044
rect 3808 61988 3864 62044
rect 3864 61988 3868 62044
rect 3804 61984 3868 61988
rect 3884 62044 3948 62048
rect 3884 61988 3888 62044
rect 3888 61988 3944 62044
rect 3944 61988 3948 62044
rect 3884 61984 3948 61988
rect 3964 62044 4028 62048
rect 3964 61988 3968 62044
rect 3968 61988 4024 62044
rect 4024 61988 4028 62044
rect 3964 61984 4028 61988
rect 4044 62044 4108 62048
rect 4044 61988 4048 62044
rect 4048 61988 4104 62044
rect 4104 61988 4108 62044
rect 4044 61984 4108 61988
rect 3068 61500 3132 61504
rect 3068 61444 3072 61500
rect 3072 61444 3128 61500
rect 3128 61444 3132 61500
rect 3068 61440 3132 61444
rect 3148 61500 3212 61504
rect 3148 61444 3152 61500
rect 3152 61444 3208 61500
rect 3208 61444 3212 61500
rect 3148 61440 3212 61444
rect 3228 61500 3292 61504
rect 3228 61444 3232 61500
rect 3232 61444 3288 61500
rect 3288 61444 3292 61500
rect 3228 61440 3292 61444
rect 3308 61500 3372 61504
rect 3308 61444 3312 61500
rect 3312 61444 3368 61500
rect 3368 61444 3372 61500
rect 3308 61440 3372 61444
rect 3804 60956 3868 60960
rect 3804 60900 3808 60956
rect 3808 60900 3864 60956
rect 3864 60900 3868 60956
rect 3804 60896 3868 60900
rect 3884 60956 3948 60960
rect 3884 60900 3888 60956
rect 3888 60900 3944 60956
rect 3944 60900 3948 60956
rect 3884 60896 3948 60900
rect 3964 60956 4028 60960
rect 3964 60900 3968 60956
rect 3968 60900 4024 60956
rect 4024 60900 4028 60956
rect 3964 60896 4028 60900
rect 4044 60956 4108 60960
rect 4044 60900 4048 60956
rect 4048 60900 4104 60956
rect 4104 60900 4108 60956
rect 4044 60896 4108 60900
rect 86908 60692 86972 60756
rect 3068 60412 3132 60416
rect 3068 60356 3072 60412
rect 3072 60356 3128 60412
rect 3128 60356 3132 60412
rect 3068 60352 3132 60356
rect 3148 60412 3212 60416
rect 3148 60356 3152 60412
rect 3152 60356 3208 60412
rect 3208 60356 3212 60412
rect 3148 60352 3212 60356
rect 3228 60412 3292 60416
rect 3228 60356 3232 60412
rect 3232 60356 3288 60412
rect 3288 60356 3292 60412
rect 3228 60352 3292 60356
rect 3308 60412 3372 60416
rect 3308 60356 3312 60412
rect 3312 60356 3368 60412
rect 3368 60356 3372 60412
rect 3308 60352 3372 60356
rect 3804 59868 3868 59872
rect 3804 59812 3808 59868
rect 3808 59812 3864 59868
rect 3864 59812 3868 59868
rect 3804 59808 3868 59812
rect 3884 59868 3948 59872
rect 3884 59812 3888 59868
rect 3888 59812 3944 59868
rect 3944 59812 3948 59868
rect 3884 59808 3948 59812
rect 3964 59868 4028 59872
rect 3964 59812 3968 59868
rect 3968 59812 4024 59868
rect 4024 59812 4028 59868
rect 3964 59808 4028 59812
rect 4044 59868 4108 59872
rect 4044 59812 4048 59868
rect 4048 59812 4104 59868
rect 4104 59812 4108 59868
rect 4044 59808 4108 59812
rect 87092 59332 87156 59396
rect 87460 59332 87524 59396
rect 3068 59324 3132 59328
rect 3068 59268 3072 59324
rect 3072 59268 3128 59324
rect 3128 59268 3132 59324
rect 3068 59264 3132 59268
rect 3148 59324 3212 59328
rect 3148 59268 3152 59324
rect 3152 59268 3208 59324
rect 3208 59268 3212 59324
rect 3148 59264 3212 59268
rect 3228 59324 3292 59328
rect 3228 59268 3232 59324
rect 3232 59268 3288 59324
rect 3288 59268 3292 59324
rect 3228 59264 3292 59268
rect 3308 59324 3372 59328
rect 3308 59268 3312 59324
rect 3312 59268 3368 59324
rect 3368 59268 3372 59324
rect 3308 59264 3372 59268
rect 3804 58780 3868 58784
rect 3804 58724 3808 58780
rect 3808 58724 3864 58780
rect 3864 58724 3868 58780
rect 3804 58720 3868 58724
rect 3884 58780 3948 58784
rect 3884 58724 3888 58780
rect 3888 58724 3944 58780
rect 3944 58724 3948 58780
rect 3884 58720 3948 58724
rect 3964 58780 4028 58784
rect 3964 58724 3968 58780
rect 3968 58724 4024 58780
rect 4024 58724 4028 58780
rect 3964 58720 4028 58724
rect 4044 58780 4108 58784
rect 4044 58724 4048 58780
rect 4048 58724 4104 58780
rect 4104 58724 4108 58780
rect 4044 58720 4108 58724
rect 3068 58236 3132 58240
rect 3068 58180 3072 58236
rect 3072 58180 3128 58236
rect 3128 58180 3132 58236
rect 3068 58176 3132 58180
rect 3148 58236 3212 58240
rect 3148 58180 3152 58236
rect 3152 58180 3208 58236
rect 3208 58180 3212 58236
rect 3148 58176 3212 58180
rect 3228 58236 3292 58240
rect 3228 58180 3232 58236
rect 3232 58180 3288 58236
rect 3288 58180 3292 58236
rect 3228 58176 3292 58180
rect 3308 58236 3372 58240
rect 3308 58180 3312 58236
rect 3312 58180 3368 58236
rect 3368 58180 3372 58236
rect 3308 58176 3372 58180
rect 3804 57692 3868 57696
rect 3804 57636 3808 57692
rect 3808 57636 3864 57692
rect 3864 57636 3868 57692
rect 3804 57632 3868 57636
rect 3884 57692 3948 57696
rect 3884 57636 3888 57692
rect 3888 57636 3944 57692
rect 3944 57636 3948 57692
rect 3884 57632 3948 57636
rect 3964 57692 4028 57696
rect 3964 57636 3968 57692
rect 3968 57636 4024 57692
rect 4024 57636 4028 57692
rect 3964 57632 4028 57636
rect 4044 57692 4108 57696
rect 4044 57636 4048 57692
rect 4048 57636 4104 57692
rect 4104 57636 4108 57692
rect 4044 57632 4108 57636
rect 3068 57148 3132 57152
rect 3068 57092 3072 57148
rect 3072 57092 3128 57148
rect 3128 57092 3132 57148
rect 3068 57088 3132 57092
rect 3148 57148 3212 57152
rect 3148 57092 3152 57148
rect 3152 57092 3208 57148
rect 3208 57092 3212 57148
rect 3148 57088 3212 57092
rect 3228 57148 3292 57152
rect 3228 57092 3232 57148
rect 3232 57092 3288 57148
rect 3288 57092 3292 57148
rect 3228 57088 3292 57092
rect 3308 57148 3372 57152
rect 3308 57092 3312 57148
rect 3312 57092 3368 57148
rect 3368 57092 3372 57148
rect 3308 57088 3372 57092
rect 3804 56604 3868 56608
rect 3804 56548 3808 56604
rect 3808 56548 3864 56604
rect 3864 56548 3868 56604
rect 3804 56544 3868 56548
rect 3884 56604 3948 56608
rect 3884 56548 3888 56604
rect 3888 56548 3944 56604
rect 3944 56548 3948 56604
rect 3884 56544 3948 56548
rect 3964 56604 4028 56608
rect 3964 56548 3968 56604
rect 3968 56548 4024 56604
rect 4024 56548 4028 56604
rect 3964 56544 4028 56548
rect 4044 56604 4108 56608
rect 4044 56548 4048 56604
rect 4048 56548 4104 56604
rect 4104 56548 4108 56604
rect 4044 56544 4108 56548
rect 3068 56060 3132 56064
rect 3068 56004 3072 56060
rect 3072 56004 3128 56060
rect 3128 56004 3132 56060
rect 3068 56000 3132 56004
rect 3148 56060 3212 56064
rect 3148 56004 3152 56060
rect 3152 56004 3208 56060
rect 3208 56004 3212 56060
rect 3148 56000 3212 56004
rect 3228 56060 3292 56064
rect 3228 56004 3232 56060
rect 3232 56004 3288 56060
rect 3288 56004 3292 56060
rect 3228 56000 3292 56004
rect 3308 56060 3372 56064
rect 3308 56004 3312 56060
rect 3312 56004 3368 56060
rect 3368 56004 3372 56060
rect 3308 56000 3372 56004
rect 3804 55516 3868 55520
rect 3804 55460 3808 55516
rect 3808 55460 3864 55516
rect 3864 55460 3868 55516
rect 3804 55456 3868 55460
rect 3884 55516 3948 55520
rect 3884 55460 3888 55516
rect 3888 55460 3944 55516
rect 3944 55460 3948 55516
rect 3884 55456 3948 55460
rect 3964 55516 4028 55520
rect 3964 55460 3968 55516
rect 3968 55460 4024 55516
rect 4024 55460 4028 55516
rect 3964 55456 4028 55460
rect 4044 55516 4108 55520
rect 4044 55460 4048 55516
rect 4048 55460 4104 55516
rect 4104 55460 4108 55516
rect 4044 55456 4108 55460
rect 86908 55252 86972 55316
rect 3068 54972 3132 54976
rect 3068 54916 3072 54972
rect 3072 54916 3128 54972
rect 3128 54916 3132 54972
rect 3068 54912 3132 54916
rect 3148 54972 3212 54976
rect 3148 54916 3152 54972
rect 3152 54916 3208 54972
rect 3208 54916 3212 54972
rect 3148 54912 3212 54916
rect 3228 54972 3292 54976
rect 3228 54916 3232 54972
rect 3232 54916 3288 54972
rect 3288 54916 3292 54972
rect 3228 54912 3292 54916
rect 3308 54972 3372 54976
rect 3308 54916 3312 54972
rect 3312 54916 3368 54972
rect 3368 54916 3372 54972
rect 3308 54912 3372 54916
rect 3804 54428 3868 54432
rect 3804 54372 3808 54428
rect 3808 54372 3864 54428
rect 3864 54372 3868 54428
rect 3804 54368 3868 54372
rect 3884 54428 3948 54432
rect 3884 54372 3888 54428
rect 3888 54372 3944 54428
rect 3944 54372 3948 54428
rect 3884 54368 3948 54372
rect 3964 54428 4028 54432
rect 3964 54372 3968 54428
rect 3968 54372 4024 54428
rect 4024 54372 4028 54428
rect 3964 54368 4028 54372
rect 4044 54428 4108 54432
rect 4044 54372 4048 54428
rect 4048 54372 4104 54428
rect 4104 54372 4108 54428
rect 4044 54368 4108 54372
rect 3068 53884 3132 53888
rect 3068 53828 3072 53884
rect 3072 53828 3128 53884
rect 3128 53828 3132 53884
rect 3068 53824 3132 53828
rect 3148 53884 3212 53888
rect 3148 53828 3152 53884
rect 3152 53828 3208 53884
rect 3208 53828 3212 53884
rect 3148 53824 3212 53828
rect 3228 53884 3292 53888
rect 3228 53828 3232 53884
rect 3232 53828 3288 53884
rect 3288 53828 3292 53884
rect 3228 53824 3292 53828
rect 3308 53884 3372 53888
rect 3308 53828 3312 53884
rect 3312 53828 3368 53884
rect 3368 53828 3372 53884
rect 3308 53824 3372 53828
rect 3804 53340 3868 53344
rect 3804 53284 3808 53340
rect 3808 53284 3864 53340
rect 3864 53284 3868 53340
rect 3804 53280 3868 53284
rect 3884 53340 3948 53344
rect 3884 53284 3888 53340
rect 3888 53284 3944 53340
rect 3944 53284 3948 53340
rect 3884 53280 3948 53284
rect 3964 53340 4028 53344
rect 3964 53284 3968 53340
rect 3968 53284 4024 53340
rect 4024 53284 4028 53340
rect 3964 53280 4028 53284
rect 4044 53340 4108 53344
rect 4044 53284 4048 53340
rect 4048 53284 4104 53340
rect 4104 53284 4108 53340
rect 4044 53280 4108 53284
rect 3068 52796 3132 52800
rect 3068 52740 3072 52796
rect 3072 52740 3128 52796
rect 3128 52740 3132 52796
rect 3068 52736 3132 52740
rect 3148 52796 3212 52800
rect 3148 52740 3152 52796
rect 3152 52740 3208 52796
rect 3208 52740 3212 52796
rect 3148 52736 3212 52740
rect 3228 52796 3292 52800
rect 3228 52740 3232 52796
rect 3232 52740 3288 52796
rect 3288 52740 3292 52796
rect 3228 52736 3292 52740
rect 3308 52796 3372 52800
rect 3308 52740 3312 52796
rect 3312 52740 3368 52796
rect 3368 52740 3372 52796
rect 3308 52736 3372 52740
rect 3804 52252 3868 52256
rect 3804 52196 3808 52252
rect 3808 52196 3864 52252
rect 3864 52196 3868 52252
rect 3804 52192 3868 52196
rect 3884 52252 3948 52256
rect 3884 52196 3888 52252
rect 3888 52196 3944 52252
rect 3944 52196 3948 52252
rect 3884 52192 3948 52196
rect 3964 52252 4028 52256
rect 3964 52196 3968 52252
rect 3968 52196 4024 52252
rect 4024 52196 4028 52252
rect 3964 52192 4028 52196
rect 4044 52252 4108 52256
rect 4044 52196 4048 52252
rect 4048 52196 4104 52252
rect 4104 52196 4108 52252
rect 4044 52192 4108 52196
rect 3068 51708 3132 51712
rect 3068 51652 3072 51708
rect 3072 51652 3128 51708
rect 3128 51652 3132 51708
rect 3068 51648 3132 51652
rect 3148 51708 3212 51712
rect 3148 51652 3152 51708
rect 3152 51652 3208 51708
rect 3208 51652 3212 51708
rect 3148 51648 3212 51652
rect 3228 51708 3292 51712
rect 3228 51652 3232 51708
rect 3232 51652 3288 51708
rect 3288 51652 3292 51708
rect 3228 51648 3292 51652
rect 3308 51708 3372 51712
rect 3308 51652 3312 51708
rect 3312 51652 3368 51708
rect 3368 51652 3372 51708
rect 3308 51648 3372 51652
rect 3804 51164 3868 51168
rect 3804 51108 3808 51164
rect 3808 51108 3864 51164
rect 3864 51108 3868 51164
rect 3804 51104 3868 51108
rect 3884 51164 3948 51168
rect 3884 51108 3888 51164
rect 3888 51108 3944 51164
rect 3944 51108 3948 51164
rect 3884 51104 3948 51108
rect 3964 51164 4028 51168
rect 3964 51108 3968 51164
rect 3968 51108 4024 51164
rect 4024 51108 4028 51164
rect 3964 51104 4028 51108
rect 4044 51164 4108 51168
rect 4044 51108 4048 51164
rect 4048 51108 4104 51164
rect 4104 51108 4108 51164
rect 4044 51104 4108 51108
rect 5764 50764 5828 50828
rect 5580 50628 5644 50692
rect 85252 50628 85316 50692
rect 3068 50620 3132 50624
rect 3068 50564 3072 50620
rect 3072 50564 3128 50620
rect 3128 50564 3132 50620
rect 3068 50560 3132 50564
rect 3148 50620 3212 50624
rect 3148 50564 3152 50620
rect 3152 50564 3208 50620
rect 3208 50564 3212 50620
rect 3148 50560 3212 50564
rect 3228 50620 3292 50624
rect 3228 50564 3232 50620
rect 3232 50564 3288 50620
rect 3288 50564 3292 50620
rect 3228 50560 3292 50564
rect 3308 50620 3372 50624
rect 3308 50564 3312 50620
rect 3312 50564 3368 50620
rect 3368 50564 3372 50620
rect 3308 50560 3372 50564
rect 86356 50492 86420 50556
rect 47716 50220 47780 50284
rect 85252 50084 85316 50148
rect 3804 50076 3868 50080
rect 3804 50020 3808 50076
rect 3808 50020 3864 50076
rect 3864 50020 3868 50076
rect 3804 50016 3868 50020
rect 3884 50076 3948 50080
rect 3884 50020 3888 50076
rect 3888 50020 3944 50076
rect 3944 50020 3948 50076
rect 3884 50016 3948 50020
rect 3964 50076 4028 50080
rect 3964 50020 3968 50076
rect 3968 50020 4024 50076
rect 4024 50020 4028 50076
rect 3964 50016 4028 50020
rect 4044 50076 4108 50080
rect 4044 50020 4048 50076
rect 4048 50020 4104 50076
rect 4104 50020 4108 50076
rect 4044 50016 4108 50020
rect 796 49676 860 49740
rect 87092 49540 87156 49604
rect 3068 49532 3132 49536
rect 3068 49476 3072 49532
rect 3072 49476 3128 49532
rect 3128 49476 3132 49532
rect 3068 49472 3132 49476
rect 3148 49532 3212 49536
rect 3148 49476 3152 49532
rect 3152 49476 3208 49532
rect 3208 49476 3212 49532
rect 3148 49472 3212 49476
rect 3228 49532 3292 49536
rect 3228 49476 3232 49532
rect 3232 49476 3288 49532
rect 3288 49476 3292 49532
rect 3228 49472 3292 49476
rect 3308 49532 3372 49536
rect 3308 49476 3312 49532
rect 3312 49476 3368 49532
rect 3368 49476 3372 49532
rect 3308 49472 3372 49476
rect 796 49404 860 49468
rect 5948 49404 6012 49468
rect 796 49268 860 49332
rect 48084 49132 48148 49196
rect 86908 49132 86972 49196
rect 796 48996 860 49060
rect 3804 48988 3868 48992
rect 3804 48932 3808 48988
rect 3808 48932 3864 48988
rect 3864 48932 3868 48988
rect 3804 48928 3868 48932
rect 3884 48988 3948 48992
rect 3884 48932 3888 48988
rect 3888 48932 3944 48988
rect 3944 48932 3948 48988
rect 3884 48928 3948 48932
rect 3964 48988 4028 48992
rect 3964 48932 3968 48988
rect 3968 48932 4024 48988
rect 4024 48932 4028 48988
rect 3964 48928 4028 48932
rect 4044 48988 4108 48992
rect 4044 48932 4048 48988
rect 4048 48932 4104 48988
rect 4104 48932 4108 48988
rect 4044 48928 4108 48932
rect 47532 48860 47596 48924
rect 86540 48860 86604 48924
rect 3068 48444 3132 48448
rect 3068 48388 3072 48444
rect 3072 48388 3128 48444
rect 3128 48388 3132 48444
rect 3068 48384 3132 48388
rect 3148 48444 3212 48448
rect 3148 48388 3152 48444
rect 3152 48388 3208 48444
rect 3208 48388 3212 48444
rect 3148 48384 3212 48388
rect 3228 48444 3292 48448
rect 3228 48388 3232 48444
rect 3232 48388 3288 48444
rect 3288 48388 3292 48444
rect 3228 48384 3292 48388
rect 3308 48444 3372 48448
rect 3308 48388 3312 48444
rect 3312 48388 3368 48444
rect 3368 48388 3372 48444
rect 3308 48384 3372 48388
rect 48084 48316 48148 48380
rect 87644 48316 87708 48380
rect 47716 48044 47780 48108
rect 48268 48044 48332 48108
rect 796 47908 860 47972
rect 3804 47900 3868 47904
rect 3804 47844 3808 47900
rect 3808 47844 3864 47900
rect 3864 47844 3868 47900
rect 3804 47840 3868 47844
rect 3884 47900 3948 47904
rect 3884 47844 3888 47900
rect 3888 47844 3944 47900
rect 3944 47844 3948 47900
rect 3884 47840 3948 47844
rect 3964 47900 4028 47904
rect 3964 47844 3968 47900
rect 3968 47844 4024 47900
rect 4024 47844 4028 47900
rect 3964 47840 4028 47844
rect 4044 47900 4108 47904
rect 4044 47844 4048 47900
rect 4048 47844 4104 47900
rect 4104 47844 4108 47900
rect 4044 47840 4108 47844
rect 47900 47772 47964 47836
rect 796 47636 860 47700
rect 48268 47636 48332 47700
rect 87276 47500 87340 47564
rect 3068 47356 3132 47360
rect 3068 47300 3072 47356
rect 3072 47300 3128 47356
rect 3128 47300 3132 47356
rect 3068 47296 3132 47300
rect 3148 47356 3212 47360
rect 3148 47300 3152 47356
rect 3152 47300 3208 47356
rect 3208 47300 3212 47356
rect 3148 47296 3212 47300
rect 3228 47356 3292 47360
rect 3228 47300 3232 47356
rect 3232 47300 3288 47356
rect 3288 47300 3292 47356
rect 3228 47296 3292 47300
rect 3308 47356 3372 47360
rect 3308 47300 3312 47356
rect 3312 47300 3368 47356
rect 3368 47300 3372 47356
rect 3308 47296 3372 47300
rect 87092 47092 87156 47156
rect 5212 46956 5276 47020
rect 3804 46812 3868 46816
rect 3804 46756 3808 46812
rect 3808 46756 3864 46812
rect 3864 46756 3868 46812
rect 3804 46752 3868 46756
rect 3884 46812 3948 46816
rect 3884 46756 3888 46812
rect 3888 46756 3944 46812
rect 3944 46756 3948 46812
rect 3884 46752 3948 46756
rect 3964 46812 4028 46816
rect 3964 46756 3968 46812
rect 3968 46756 4024 46812
rect 4024 46756 4028 46812
rect 3964 46752 4028 46756
rect 4044 46812 4108 46816
rect 4044 46756 4048 46812
rect 4048 46756 4104 46812
rect 4104 46756 4108 46812
rect 4044 46752 4108 46756
rect 3068 46268 3132 46272
rect 3068 46212 3072 46268
rect 3072 46212 3128 46268
rect 3128 46212 3132 46268
rect 3068 46208 3132 46212
rect 3148 46268 3212 46272
rect 3148 46212 3152 46268
rect 3152 46212 3208 46268
rect 3208 46212 3212 46268
rect 3148 46208 3212 46212
rect 3228 46268 3292 46272
rect 3228 46212 3232 46268
rect 3232 46212 3288 46268
rect 3288 46212 3292 46268
rect 3228 46208 3292 46212
rect 3308 46268 3372 46272
rect 3308 46212 3312 46268
rect 3312 46212 3368 46268
rect 3368 46212 3372 46268
rect 3308 46208 3372 46212
rect 3804 45724 3868 45728
rect 3804 45668 3808 45724
rect 3808 45668 3864 45724
rect 3864 45668 3868 45724
rect 3804 45664 3868 45668
rect 3884 45724 3948 45728
rect 3884 45668 3888 45724
rect 3888 45668 3944 45724
rect 3944 45668 3948 45724
rect 3884 45664 3948 45668
rect 3964 45724 4028 45728
rect 3964 45668 3968 45724
rect 3968 45668 4024 45724
rect 4024 45668 4028 45724
rect 3964 45664 4028 45668
rect 4044 45724 4108 45728
rect 4044 45668 4048 45724
rect 4048 45668 4104 45724
rect 4104 45668 4108 45724
rect 4044 45664 4108 45668
rect 3068 45180 3132 45184
rect 3068 45124 3072 45180
rect 3072 45124 3128 45180
rect 3128 45124 3132 45180
rect 3068 45120 3132 45124
rect 3148 45180 3212 45184
rect 3148 45124 3152 45180
rect 3152 45124 3208 45180
rect 3208 45124 3212 45180
rect 3148 45120 3212 45124
rect 3228 45180 3292 45184
rect 3228 45124 3232 45180
rect 3232 45124 3288 45180
rect 3288 45124 3292 45180
rect 3228 45120 3292 45124
rect 3308 45180 3372 45184
rect 3308 45124 3312 45180
rect 3312 45124 3368 45180
rect 3368 45124 3372 45180
rect 3308 45120 3372 45124
rect 3804 44636 3868 44640
rect 3804 44580 3808 44636
rect 3808 44580 3864 44636
rect 3864 44580 3868 44636
rect 3804 44576 3868 44580
rect 3884 44636 3948 44640
rect 3884 44580 3888 44636
rect 3888 44580 3944 44636
rect 3944 44580 3948 44636
rect 3884 44576 3948 44580
rect 3964 44636 4028 44640
rect 3964 44580 3968 44636
rect 3968 44580 4024 44636
rect 4024 44580 4028 44636
rect 3964 44576 4028 44580
rect 4044 44636 4108 44640
rect 4044 44580 4048 44636
rect 4048 44580 4104 44636
rect 4104 44580 4108 44636
rect 4044 44576 4108 44580
rect 3068 44092 3132 44096
rect 3068 44036 3072 44092
rect 3072 44036 3128 44092
rect 3128 44036 3132 44092
rect 3068 44032 3132 44036
rect 3148 44092 3212 44096
rect 3148 44036 3152 44092
rect 3152 44036 3208 44092
rect 3208 44036 3212 44092
rect 3148 44032 3212 44036
rect 3228 44092 3292 44096
rect 3228 44036 3232 44092
rect 3232 44036 3288 44092
rect 3288 44036 3292 44092
rect 3228 44032 3292 44036
rect 3308 44092 3372 44096
rect 3308 44036 3312 44092
rect 3312 44036 3368 44092
rect 3368 44036 3372 44092
rect 3308 44032 3372 44036
rect 3804 43548 3868 43552
rect 3804 43492 3808 43548
rect 3808 43492 3864 43548
rect 3864 43492 3868 43548
rect 3804 43488 3868 43492
rect 3884 43548 3948 43552
rect 3884 43492 3888 43548
rect 3888 43492 3944 43548
rect 3944 43492 3948 43548
rect 3884 43488 3948 43492
rect 3964 43548 4028 43552
rect 3964 43492 3968 43548
rect 3968 43492 4024 43548
rect 4024 43492 4028 43548
rect 3964 43488 4028 43492
rect 4044 43548 4108 43552
rect 4044 43492 4048 43548
rect 4048 43492 4104 43548
rect 4104 43492 4108 43548
rect 4044 43488 4108 43492
rect 3068 43004 3132 43008
rect 3068 42948 3072 43004
rect 3072 42948 3128 43004
rect 3128 42948 3132 43004
rect 3068 42944 3132 42948
rect 3148 43004 3212 43008
rect 3148 42948 3152 43004
rect 3152 42948 3208 43004
rect 3208 42948 3212 43004
rect 3148 42944 3212 42948
rect 3228 43004 3292 43008
rect 3228 42948 3232 43004
rect 3232 42948 3288 43004
rect 3288 42948 3292 43004
rect 3228 42944 3292 42948
rect 3308 43004 3372 43008
rect 3308 42948 3312 43004
rect 3312 42948 3368 43004
rect 3368 42948 3372 43004
rect 3308 42944 3372 42948
rect 3804 42460 3868 42464
rect 3804 42404 3808 42460
rect 3808 42404 3864 42460
rect 3864 42404 3868 42460
rect 3804 42400 3868 42404
rect 3884 42460 3948 42464
rect 3884 42404 3888 42460
rect 3888 42404 3944 42460
rect 3944 42404 3948 42460
rect 3884 42400 3948 42404
rect 3964 42460 4028 42464
rect 3964 42404 3968 42460
rect 3968 42404 4024 42460
rect 4024 42404 4028 42460
rect 3964 42400 4028 42404
rect 4044 42460 4108 42464
rect 4044 42404 4048 42460
rect 4048 42404 4104 42460
rect 4104 42404 4108 42460
rect 4044 42400 4108 42404
rect 3068 41916 3132 41920
rect 3068 41860 3072 41916
rect 3072 41860 3128 41916
rect 3128 41860 3132 41916
rect 3068 41856 3132 41860
rect 3148 41916 3212 41920
rect 3148 41860 3152 41916
rect 3152 41860 3208 41916
rect 3208 41860 3212 41916
rect 3148 41856 3212 41860
rect 3228 41916 3292 41920
rect 3228 41860 3232 41916
rect 3232 41860 3288 41916
rect 3288 41860 3292 41916
rect 3228 41856 3292 41860
rect 3308 41916 3372 41920
rect 3308 41860 3312 41916
rect 3312 41860 3368 41916
rect 3368 41860 3372 41916
rect 3308 41856 3372 41860
rect 3804 41372 3868 41376
rect 3804 41316 3808 41372
rect 3808 41316 3864 41372
rect 3864 41316 3868 41372
rect 3804 41312 3868 41316
rect 3884 41372 3948 41376
rect 3884 41316 3888 41372
rect 3888 41316 3944 41372
rect 3944 41316 3948 41372
rect 3884 41312 3948 41316
rect 3964 41372 4028 41376
rect 3964 41316 3968 41372
rect 3968 41316 4024 41372
rect 4024 41316 4028 41372
rect 3964 41312 4028 41316
rect 4044 41372 4108 41376
rect 4044 41316 4048 41372
rect 4048 41316 4104 41372
rect 4104 41316 4108 41372
rect 4044 41312 4108 41316
rect 3068 40828 3132 40832
rect 3068 40772 3072 40828
rect 3072 40772 3128 40828
rect 3128 40772 3132 40828
rect 3068 40768 3132 40772
rect 3148 40828 3212 40832
rect 3148 40772 3152 40828
rect 3152 40772 3208 40828
rect 3208 40772 3212 40828
rect 3148 40768 3212 40772
rect 3228 40828 3292 40832
rect 3228 40772 3232 40828
rect 3232 40772 3288 40828
rect 3288 40772 3292 40828
rect 3228 40768 3292 40772
rect 3308 40828 3372 40832
rect 3308 40772 3312 40828
rect 3312 40772 3368 40828
rect 3368 40772 3372 40828
rect 3308 40768 3372 40772
rect 87276 40700 87340 40764
rect 87276 40428 87340 40492
rect 3804 40284 3868 40288
rect 3804 40228 3808 40284
rect 3808 40228 3864 40284
rect 3864 40228 3868 40284
rect 3804 40224 3868 40228
rect 3884 40284 3948 40288
rect 3884 40228 3888 40284
rect 3888 40228 3944 40284
rect 3944 40228 3948 40284
rect 3884 40224 3948 40228
rect 3964 40284 4028 40288
rect 3964 40228 3968 40284
rect 3968 40228 4024 40284
rect 4024 40228 4028 40284
rect 3964 40224 4028 40228
rect 4044 40284 4108 40288
rect 4044 40228 4048 40284
rect 4048 40228 4104 40284
rect 4104 40228 4108 40284
rect 4044 40224 4108 40228
rect 3068 39740 3132 39744
rect 3068 39684 3072 39740
rect 3072 39684 3128 39740
rect 3128 39684 3132 39740
rect 3068 39680 3132 39684
rect 3148 39740 3212 39744
rect 3148 39684 3152 39740
rect 3152 39684 3208 39740
rect 3208 39684 3212 39740
rect 3148 39680 3212 39684
rect 3228 39740 3292 39744
rect 3228 39684 3232 39740
rect 3232 39684 3288 39740
rect 3288 39684 3292 39740
rect 3228 39680 3292 39684
rect 3308 39740 3372 39744
rect 3308 39684 3312 39740
rect 3312 39684 3368 39740
rect 3368 39684 3372 39740
rect 3308 39680 3372 39684
rect 3804 39196 3868 39200
rect 3804 39140 3808 39196
rect 3808 39140 3864 39196
rect 3864 39140 3868 39196
rect 3804 39136 3868 39140
rect 3884 39196 3948 39200
rect 3884 39140 3888 39196
rect 3888 39140 3944 39196
rect 3944 39140 3948 39196
rect 3884 39136 3948 39140
rect 3964 39196 4028 39200
rect 3964 39140 3968 39196
rect 3968 39140 4024 39196
rect 4024 39140 4028 39196
rect 3964 39136 4028 39140
rect 4044 39196 4108 39200
rect 4044 39140 4048 39196
rect 4048 39140 4104 39196
rect 4104 39140 4108 39196
rect 4044 39136 4108 39140
rect 3068 38652 3132 38656
rect 3068 38596 3072 38652
rect 3072 38596 3128 38652
rect 3128 38596 3132 38652
rect 3068 38592 3132 38596
rect 3148 38652 3212 38656
rect 3148 38596 3152 38652
rect 3152 38596 3208 38652
rect 3208 38596 3212 38652
rect 3148 38592 3212 38596
rect 3228 38652 3292 38656
rect 3228 38596 3232 38652
rect 3232 38596 3288 38652
rect 3288 38596 3292 38652
rect 3228 38592 3292 38596
rect 3308 38652 3372 38656
rect 3308 38596 3312 38652
rect 3312 38596 3368 38652
rect 3368 38596 3372 38652
rect 3308 38592 3372 38596
rect 3804 38108 3868 38112
rect 3804 38052 3808 38108
rect 3808 38052 3864 38108
rect 3864 38052 3868 38108
rect 3804 38048 3868 38052
rect 3884 38108 3948 38112
rect 3884 38052 3888 38108
rect 3888 38052 3944 38108
rect 3944 38052 3948 38108
rect 3884 38048 3948 38052
rect 3964 38108 4028 38112
rect 3964 38052 3968 38108
rect 3968 38052 4024 38108
rect 4024 38052 4028 38108
rect 3964 38048 4028 38052
rect 4044 38108 4108 38112
rect 4044 38052 4048 38108
rect 4048 38052 4104 38108
rect 4104 38052 4108 38108
rect 4044 38048 4108 38052
rect 3068 37564 3132 37568
rect 3068 37508 3072 37564
rect 3072 37508 3128 37564
rect 3128 37508 3132 37564
rect 3068 37504 3132 37508
rect 3148 37564 3212 37568
rect 3148 37508 3152 37564
rect 3152 37508 3208 37564
rect 3208 37508 3212 37564
rect 3148 37504 3212 37508
rect 3228 37564 3292 37568
rect 3228 37508 3232 37564
rect 3232 37508 3288 37564
rect 3288 37508 3292 37564
rect 3228 37504 3292 37508
rect 3308 37564 3372 37568
rect 3308 37508 3312 37564
rect 3312 37508 3368 37564
rect 3368 37508 3372 37564
rect 3308 37504 3372 37508
rect 3804 37020 3868 37024
rect 3804 36964 3808 37020
rect 3808 36964 3864 37020
rect 3864 36964 3868 37020
rect 3804 36960 3868 36964
rect 3884 37020 3948 37024
rect 3884 36964 3888 37020
rect 3888 36964 3944 37020
rect 3944 36964 3948 37020
rect 3884 36960 3948 36964
rect 3964 37020 4028 37024
rect 3964 36964 3968 37020
rect 3968 36964 4024 37020
rect 4024 36964 4028 37020
rect 3964 36960 4028 36964
rect 4044 37020 4108 37024
rect 4044 36964 4048 37020
rect 4048 36964 4104 37020
rect 4104 36964 4108 37020
rect 4044 36960 4108 36964
rect 3068 36476 3132 36480
rect 3068 36420 3072 36476
rect 3072 36420 3128 36476
rect 3128 36420 3132 36476
rect 3068 36416 3132 36420
rect 3148 36476 3212 36480
rect 3148 36420 3152 36476
rect 3152 36420 3208 36476
rect 3208 36420 3212 36476
rect 3148 36416 3212 36420
rect 3228 36476 3292 36480
rect 3228 36420 3232 36476
rect 3232 36420 3288 36476
rect 3288 36420 3292 36476
rect 3228 36416 3292 36420
rect 3308 36476 3372 36480
rect 3308 36420 3312 36476
rect 3312 36420 3368 36476
rect 3368 36420 3372 36476
rect 3308 36416 3372 36420
rect 3804 35932 3868 35936
rect 3804 35876 3808 35932
rect 3808 35876 3864 35932
rect 3864 35876 3868 35932
rect 3804 35872 3868 35876
rect 3884 35932 3948 35936
rect 3884 35876 3888 35932
rect 3888 35876 3944 35932
rect 3944 35876 3948 35932
rect 3884 35872 3948 35876
rect 3964 35932 4028 35936
rect 3964 35876 3968 35932
rect 3968 35876 4024 35932
rect 4024 35876 4028 35932
rect 3964 35872 4028 35876
rect 4044 35932 4108 35936
rect 4044 35876 4048 35932
rect 4048 35876 4104 35932
rect 4104 35876 4108 35932
rect 4044 35872 4108 35876
rect 3068 35388 3132 35392
rect 3068 35332 3072 35388
rect 3072 35332 3128 35388
rect 3128 35332 3132 35388
rect 3068 35328 3132 35332
rect 3148 35388 3212 35392
rect 3148 35332 3152 35388
rect 3152 35332 3208 35388
rect 3208 35332 3212 35388
rect 3148 35328 3212 35332
rect 3228 35388 3292 35392
rect 3228 35332 3232 35388
rect 3232 35332 3288 35388
rect 3288 35332 3292 35388
rect 3228 35328 3292 35332
rect 3308 35388 3372 35392
rect 3308 35332 3312 35388
rect 3312 35332 3368 35388
rect 3368 35332 3372 35388
rect 3308 35328 3372 35332
rect 3804 34844 3868 34848
rect 3804 34788 3808 34844
rect 3808 34788 3864 34844
rect 3864 34788 3868 34844
rect 3804 34784 3868 34788
rect 3884 34844 3948 34848
rect 3884 34788 3888 34844
rect 3888 34788 3944 34844
rect 3944 34788 3948 34844
rect 3884 34784 3948 34788
rect 3964 34844 4028 34848
rect 3964 34788 3968 34844
rect 3968 34788 4024 34844
rect 4024 34788 4028 34844
rect 3964 34784 4028 34788
rect 4044 34844 4108 34848
rect 4044 34788 4048 34844
rect 4048 34788 4104 34844
rect 4104 34788 4108 34844
rect 4044 34784 4108 34788
rect 3068 34300 3132 34304
rect 3068 34244 3072 34300
rect 3072 34244 3128 34300
rect 3128 34244 3132 34300
rect 3068 34240 3132 34244
rect 3148 34300 3212 34304
rect 3148 34244 3152 34300
rect 3152 34244 3208 34300
rect 3208 34244 3212 34300
rect 3148 34240 3212 34244
rect 3228 34300 3292 34304
rect 3228 34244 3232 34300
rect 3232 34244 3288 34300
rect 3288 34244 3292 34300
rect 3228 34240 3292 34244
rect 3308 34300 3372 34304
rect 3308 34244 3312 34300
rect 3312 34244 3368 34300
rect 3368 34244 3372 34300
rect 3308 34240 3372 34244
rect 3804 33756 3868 33760
rect 3804 33700 3808 33756
rect 3808 33700 3864 33756
rect 3864 33700 3868 33756
rect 3804 33696 3868 33700
rect 3884 33756 3948 33760
rect 3884 33700 3888 33756
rect 3888 33700 3944 33756
rect 3944 33700 3948 33756
rect 3884 33696 3948 33700
rect 3964 33756 4028 33760
rect 3964 33700 3968 33756
rect 3968 33700 4024 33756
rect 4024 33700 4028 33756
rect 3964 33696 4028 33700
rect 4044 33756 4108 33760
rect 4044 33700 4048 33756
rect 4048 33700 4104 33756
rect 4104 33700 4108 33756
rect 4044 33696 4108 33700
rect 86908 33628 86972 33692
rect 3068 33212 3132 33216
rect 3068 33156 3072 33212
rect 3072 33156 3128 33212
rect 3128 33156 3132 33212
rect 3068 33152 3132 33156
rect 3148 33212 3212 33216
rect 3148 33156 3152 33212
rect 3152 33156 3208 33212
rect 3208 33156 3212 33212
rect 3148 33152 3212 33156
rect 3228 33212 3292 33216
rect 3228 33156 3232 33212
rect 3232 33156 3288 33212
rect 3288 33156 3292 33212
rect 3228 33152 3292 33156
rect 3308 33212 3372 33216
rect 3308 33156 3312 33212
rect 3312 33156 3368 33212
rect 3368 33156 3372 33212
rect 3308 33152 3372 33156
rect 3804 32668 3868 32672
rect 3804 32612 3808 32668
rect 3808 32612 3864 32668
rect 3864 32612 3868 32668
rect 3804 32608 3868 32612
rect 3884 32668 3948 32672
rect 3884 32612 3888 32668
rect 3888 32612 3944 32668
rect 3944 32612 3948 32668
rect 3884 32608 3948 32612
rect 3964 32668 4028 32672
rect 3964 32612 3968 32668
rect 3968 32612 4024 32668
rect 4024 32612 4028 32668
rect 3964 32608 4028 32612
rect 4044 32668 4108 32672
rect 4044 32612 4048 32668
rect 4048 32612 4104 32668
rect 4104 32612 4108 32668
rect 4044 32608 4108 32612
rect 87092 32268 87156 32332
rect 3068 32124 3132 32128
rect 3068 32068 3072 32124
rect 3072 32068 3128 32124
rect 3128 32068 3132 32124
rect 3068 32064 3132 32068
rect 3148 32124 3212 32128
rect 3148 32068 3152 32124
rect 3152 32068 3208 32124
rect 3208 32068 3212 32124
rect 3148 32064 3212 32068
rect 3228 32124 3292 32128
rect 3228 32068 3232 32124
rect 3232 32068 3288 32124
rect 3288 32068 3292 32124
rect 3228 32064 3292 32068
rect 3308 32124 3372 32128
rect 3308 32068 3312 32124
rect 3312 32068 3368 32124
rect 3368 32068 3372 32124
rect 3308 32064 3372 32068
rect 3804 31580 3868 31584
rect 3804 31524 3808 31580
rect 3808 31524 3864 31580
rect 3864 31524 3868 31580
rect 3804 31520 3868 31524
rect 3884 31580 3948 31584
rect 3884 31524 3888 31580
rect 3888 31524 3944 31580
rect 3944 31524 3948 31580
rect 3884 31520 3948 31524
rect 3964 31580 4028 31584
rect 3964 31524 3968 31580
rect 3968 31524 4024 31580
rect 4024 31524 4028 31580
rect 3964 31520 4028 31524
rect 4044 31580 4108 31584
rect 4044 31524 4048 31580
rect 4048 31524 4104 31580
rect 4104 31524 4108 31580
rect 4044 31520 4108 31524
rect 3068 31036 3132 31040
rect 3068 30980 3072 31036
rect 3072 30980 3128 31036
rect 3128 30980 3132 31036
rect 3068 30976 3132 30980
rect 3148 31036 3212 31040
rect 3148 30980 3152 31036
rect 3152 30980 3208 31036
rect 3208 30980 3212 31036
rect 3148 30976 3212 30980
rect 3228 31036 3292 31040
rect 3228 30980 3232 31036
rect 3232 30980 3288 31036
rect 3288 30980 3292 31036
rect 3228 30976 3292 30980
rect 3308 31036 3372 31040
rect 3308 30980 3312 31036
rect 3312 30980 3368 31036
rect 3368 30980 3372 31036
rect 3308 30976 3372 30980
rect 87644 30908 87708 30972
rect 3804 30492 3868 30496
rect 3804 30436 3808 30492
rect 3808 30436 3864 30492
rect 3864 30436 3868 30492
rect 3804 30432 3868 30436
rect 3884 30492 3948 30496
rect 3884 30436 3888 30492
rect 3888 30436 3944 30492
rect 3944 30436 3948 30492
rect 3884 30432 3948 30436
rect 3964 30492 4028 30496
rect 3964 30436 3968 30492
rect 3968 30436 4024 30492
rect 4024 30436 4028 30492
rect 3964 30432 4028 30436
rect 4044 30492 4108 30496
rect 4044 30436 4048 30492
rect 4048 30436 4104 30492
rect 4104 30436 4108 30492
rect 4044 30432 4108 30436
rect 3068 29948 3132 29952
rect 3068 29892 3072 29948
rect 3072 29892 3128 29948
rect 3128 29892 3132 29948
rect 3068 29888 3132 29892
rect 3148 29948 3212 29952
rect 3148 29892 3152 29948
rect 3152 29892 3208 29948
rect 3208 29892 3212 29948
rect 3148 29888 3212 29892
rect 3228 29948 3292 29952
rect 3228 29892 3232 29948
rect 3232 29892 3288 29948
rect 3288 29892 3292 29948
rect 3228 29888 3292 29892
rect 3308 29948 3372 29952
rect 3308 29892 3312 29948
rect 3312 29892 3368 29948
rect 3368 29892 3372 29948
rect 3308 29888 3372 29892
rect 3804 29404 3868 29408
rect 3804 29348 3808 29404
rect 3808 29348 3864 29404
rect 3864 29348 3868 29404
rect 3804 29344 3868 29348
rect 3884 29404 3948 29408
rect 3884 29348 3888 29404
rect 3888 29348 3944 29404
rect 3944 29348 3948 29404
rect 3884 29344 3948 29348
rect 3964 29404 4028 29408
rect 3964 29348 3968 29404
rect 3968 29348 4024 29404
rect 4024 29348 4028 29404
rect 3964 29344 4028 29348
rect 4044 29404 4108 29408
rect 4044 29348 4048 29404
rect 4048 29348 4104 29404
rect 4104 29348 4108 29404
rect 4044 29344 4108 29348
rect 3068 28860 3132 28864
rect 3068 28804 3072 28860
rect 3072 28804 3128 28860
rect 3128 28804 3132 28860
rect 3068 28800 3132 28804
rect 3148 28860 3212 28864
rect 3148 28804 3152 28860
rect 3152 28804 3208 28860
rect 3208 28804 3212 28860
rect 3148 28800 3212 28804
rect 3228 28860 3292 28864
rect 3228 28804 3232 28860
rect 3232 28804 3288 28860
rect 3288 28804 3292 28860
rect 3228 28800 3292 28804
rect 3308 28860 3372 28864
rect 3308 28804 3312 28860
rect 3312 28804 3368 28860
rect 3368 28804 3372 28860
rect 3308 28800 3372 28804
rect 3804 28316 3868 28320
rect 3804 28260 3808 28316
rect 3808 28260 3864 28316
rect 3864 28260 3868 28316
rect 3804 28256 3868 28260
rect 3884 28316 3948 28320
rect 3884 28260 3888 28316
rect 3888 28260 3944 28316
rect 3944 28260 3948 28316
rect 3884 28256 3948 28260
rect 3964 28316 4028 28320
rect 3964 28260 3968 28316
rect 3968 28260 4024 28316
rect 4024 28260 4028 28316
rect 3964 28256 4028 28260
rect 4044 28316 4108 28320
rect 4044 28260 4048 28316
rect 4048 28260 4104 28316
rect 4104 28260 4108 28316
rect 4044 28256 4108 28260
rect 3068 27772 3132 27776
rect 3068 27716 3072 27772
rect 3072 27716 3128 27772
rect 3128 27716 3132 27772
rect 3068 27712 3132 27716
rect 3148 27772 3212 27776
rect 3148 27716 3152 27772
rect 3152 27716 3208 27772
rect 3208 27716 3212 27772
rect 3148 27712 3212 27716
rect 3228 27772 3292 27776
rect 3228 27716 3232 27772
rect 3232 27716 3288 27772
rect 3288 27716 3292 27772
rect 3228 27712 3292 27716
rect 3308 27772 3372 27776
rect 3308 27716 3312 27772
rect 3312 27716 3368 27772
rect 3368 27716 3372 27772
rect 3308 27712 3372 27716
rect 3804 27228 3868 27232
rect 3804 27172 3808 27228
rect 3808 27172 3864 27228
rect 3864 27172 3868 27228
rect 3804 27168 3868 27172
rect 3884 27228 3948 27232
rect 3884 27172 3888 27228
rect 3888 27172 3944 27228
rect 3944 27172 3948 27228
rect 3884 27168 3948 27172
rect 3964 27228 4028 27232
rect 3964 27172 3968 27228
rect 3968 27172 4024 27228
rect 4024 27172 4028 27228
rect 3964 27168 4028 27172
rect 4044 27228 4108 27232
rect 4044 27172 4048 27228
rect 4048 27172 4104 27228
rect 4104 27172 4108 27228
rect 4044 27168 4108 27172
rect 5212 27160 5276 27164
rect 5212 27104 5262 27160
rect 5262 27104 5276 27160
rect 5212 27100 5276 27104
rect 3068 26684 3132 26688
rect 3068 26628 3072 26684
rect 3072 26628 3128 26684
rect 3128 26628 3132 26684
rect 3068 26624 3132 26628
rect 3148 26684 3212 26688
rect 3148 26628 3152 26684
rect 3152 26628 3208 26684
rect 3208 26628 3212 26684
rect 3148 26624 3212 26628
rect 3228 26684 3292 26688
rect 3228 26628 3232 26684
rect 3232 26628 3288 26684
rect 3288 26628 3292 26684
rect 3228 26624 3292 26628
rect 3308 26684 3372 26688
rect 3308 26628 3312 26684
rect 3312 26628 3368 26684
rect 3368 26628 3372 26684
rect 3308 26624 3372 26628
rect 3804 26140 3868 26144
rect 3804 26084 3808 26140
rect 3808 26084 3864 26140
rect 3864 26084 3868 26140
rect 3804 26080 3868 26084
rect 3884 26140 3948 26144
rect 3884 26084 3888 26140
rect 3888 26084 3944 26140
rect 3944 26084 3948 26140
rect 3884 26080 3948 26084
rect 3964 26140 4028 26144
rect 3964 26084 3968 26140
rect 3968 26084 4024 26140
rect 4024 26084 4028 26140
rect 3964 26080 4028 26084
rect 4044 26140 4108 26144
rect 4044 26084 4048 26140
rect 4048 26084 4104 26140
rect 4104 26084 4108 26140
rect 4044 26080 4108 26084
rect 3068 25596 3132 25600
rect 3068 25540 3072 25596
rect 3072 25540 3128 25596
rect 3128 25540 3132 25596
rect 3068 25536 3132 25540
rect 3148 25596 3212 25600
rect 3148 25540 3152 25596
rect 3152 25540 3208 25596
rect 3208 25540 3212 25596
rect 3148 25536 3212 25540
rect 3228 25596 3292 25600
rect 3228 25540 3232 25596
rect 3232 25540 3288 25596
rect 3288 25540 3292 25596
rect 3228 25536 3292 25540
rect 3308 25596 3372 25600
rect 3308 25540 3312 25596
rect 3312 25540 3368 25596
rect 3368 25540 3372 25596
rect 3308 25536 3372 25540
rect 3804 25052 3868 25056
rect 3804 24996 3808 25052
rect 3808 24996 3864 25052
rect 3864 24996 3868 25052
rect 3804 24992 3868 24996
rect 3884 25052 3948 25056
rect 3884 24996 3888 25052
rect 3888 24996 3944 25052
rect 3944 24996 3948 25052
rect 3884 24992 3948 24996
rect 3964 25052 4028 25056
rect 3964 24996 3968 25052
rect 3968 24996 4024 25052
rect 4024 24996 4028 25052
rect 3964 24992 4028 24996
rect 4044 25052 4108 25056
rect 4044 24996 4048 25052
rect 4048 24996 4104 25052
rect 4104 24996 4108 25052
rect 4044 24992 4108 24996
rect 3068 24508 3132 24512
rect 3068 24452 3072 24508
rect 3072 24452 3128 24508
rect 3128 24452 3132 24508
rect 3068 24448 3132 24452
rect 3148 24508 3212 24512
rect 3148 24452 3152 24508
rect 3152 24452 3208 24508
rect 3208 24452 3212 24508
rect 3148 24448 3212 24452
rect 3228 24508 3292 24512
rect 3228 24452 3232 24508
rect 3232 24452 3288 24508
rect 3288 24452 3292 24508
rect 3228 24448 3292 24452
rect 3308 24508 3372 24512
rect 3308 24452 3312 24508
rect 3312 24452 3368 24508
rect 3368 24452 3372 24508
rect 3308 24448 3372 24452
rect 88748 24108 88812 24172
rect 3804 23964 3868 23968
rect 3804 23908 3808 23964
rect 3808 23908 3864 23964
rect 3864 23908 3868 23964
rect 3804 23904 3868 23908
rect 3884 23964 3948 23968
rect 3884 23908 3888 23964
rect 3888 23908 3944 23964
rect 3944 23908 3948 23964
rect 3884 23904 3948 23908
rect 3964 23964 4028 23968
rect 3964 23908 3968 23964
rect 3968 23908 4024 23964
rect 4024 23908 4028 23964
rect 3964 23904 4028 23908
rect 4044 23964 4108 23968
rect 4044 23908 4048 23964
rect 4048 23908 4104 23964
rect 4104 23908 4108 23964
rect 4044 23904 4108 23908
rect 88564 23836 88628 23900
rect 3068 23420 3132 23424
rect 3068 23364 3072 23420
rect 3072 23364 3128 23420
rect 3128 23364 3132 23420
rect 3068 23360 3132 23364
rect 3148 23420 3212 23424
rect 3148 23364 3152 23420
rect 3152 23364 3208 23420
rect 3208 23364 3212 23420
rect 3148 23360 3212 23364
rect 3228 23420 3292 23424
rect 3228 23364 3232 23420
rect 3232 23364 3288 23420
rect 3288 23364 3292 23420
rect 3228 23360 3292 23364
rect 3308 23420 3372 23424
rect 3308 23364 3312 23420
rect 3312 23364 3368 23420
rect 3368 23364 3372 23420
rect 3308 23360 3372 23364
rect 3804 22876 3868 22880
rect 3804 22820 3808 22876
rect 3808 22820 3864 22876
rect 3864 22820 3868 22876
rect 3804 22816 3868 22820
rect 3884 22876 3948 22880
rect 3884 22820 3888 22876
rect 3888 22820 3944 22876
rect 3944 22820 3948 22876
rect 3884 22816 3948 22820
rect 3964 22876 4028 22880
rect 3964 22820 3968 22876
rect 3968 22820 4024 22876
rect 4024 22820 4028 22876
rect 3964 22816 4028 22820
rect 4044 22876 4108 22880
rect 4044 22820 4048 22876
rect 4048 22820 4104 22876
rect 4104 22820 4108 22876
rect 4044 22816 4108 22820
rect 86356 22748 86420 22812
rect 3068 22332 3132 22336
rect 3068 22276 3072 22332
rect 3072 22276 3128 22332
rect 3128 22276 3132 22332
rect 3068 22272 3132 22276
rect 3148 22332 3212 22336
rect 3148 22276 3152 22332
rect 3152 22276 3208 22332
rect 3208 22276 3212 22332
rect 3148 22272 3212 22276
rect 3228 22332 3292 22336
rect 3228 22276 3232 22332
rect 3232 22276 3288 22332
rect 3288 22276 3292 22332
rect 3228 22272 3292 22276
rect 3308 22332 3372 22336
rect 3308 22276 3312 22332
rect 3312 22276 3368 22332
rect 3368 22276 3372 22332
rect 3308 22272 3372 22276
rect 3804 21788 3868 21792
rect 3804 21732 3808 21788
rect 3808 21732 3864 21788
rect 3864 21732 3868 21788
rect 3804 21728 3868 21732
rect 3884 21788 3948 21792
rect 3884 21732 3888 21788
rect 3888 21732 3944 21788
rect 3944 21732 3948 21788
rect 3884 21728 3948 21732
rect 3964 21788 4028 21792
rect 3964 21732 3968 21788
rect 3968 21732 4024 21788
rect 4024 21732 4028 21788
rect 3964 21728 4028 21732
rect 4044 21788 4108 21792
rect 4044 21732 4048 21788
rect 4048 21732 4104 21788
rect 4104 21732 4108 21788
rect 4044 21728 4108 21732
rect 88196 21388 88260 21452
rect 3068 21244 3132 21248
rect 3068 21188 3072 21244
rect 3072 21188 3128 21244
rect 3128 21188 3132 21244
rect 3068 21184 3132 21188
rect 3148 21244 3212 21248
rect 3148 21188 3152 21244
rect 3152 21188 3208 21244
rect 3208 21188 3212 21244
rect 3148 21184 3212 21188
rect 3228 21244 3292 21248
rect 3228 21188 3232 21244
rect 3232 21188 3288 21244
rect 3288 21188 3292 21244
rect 3228 21184 3292 21188
rect 3308 21244 3372 21248
rect 3308 21188 3312 21244
rect 3312 21188 3368 21244
rect 3368 21188 3372 21244
rect 3308 21184 3372 21188
rect 3804 20700 3868 20704
rect 3804 20644 3808 20700
rect 3808 20644 3864 20700
rect 3864 20644 3868 20700
rect 3804 20640 3868 20644
rect 3884 20700 3948 20704
rect 3884 20644 3888 20700
rect 3888 20644 3944 20700
rect 3944 20644 3948 20700
rect 3884 20640 3948 20644
rect 3964 20700 4028 20704
rect 3964 20644 3968 20700
rect 3968 20644 4024 20700
rect 4024 20644 4028 20700
rect 3964 20640 4028 20644
rect 4044 20700 4108 20704
rect 4044 20644 4048 20700
rect 4048 20644 4104 20700
rect 4104 20644 4108 20700
rect 4044 20640 4108 20644
rect 3068 20156 3132 20160
rect 3068 20100 3072 20156
rect 3072 20100 3128 20156
rect 3128 20100 3132 20156
rect 3068 20096 3132 20100
rect 3148 20156 3212 20160
rect 3148 20100 3152 20156
rect 3152 20100 3208 20156
rect 3208 20100 3212 20156
rect 3148 20096 3212 20100
rect 3228 20156 3292 20160
rect 3228 20100 3232 20156
rect 3232 20100 3288 20156
rect 3288 20100 3292 20156
rect 3228 20096 3292 20100
rect 3308 20156 3372 20160
rect 3308 20100 3312 20156
rect 3312 20100 3368 20156
rect 3368 20100 3372 20156
rect 3308 20096 3372 20100
rect 3804 19612 3868 19616
rect 3804 19556 3808 19612
rect 3808 19556 3864 19612
rect 3864 19556 3868 19612
rect 3804 19552 3868 19556
rect 3884 19612 3948 19616
rect 3884 19556 3888 19612
rect 3888 19556 3944 19612
rect 3944 19556 3948 19612
rect 3884 19552 3948 19556
rect 3964 19612 4028 19616
rect 3964 19556 3968 19612
rect 3968 19556 4024 19612
rect 4024 19556 4028 19612
rect 3964 19552 4028 19556
rect 4044 19612 4108 19616
rect 4044 19556 4048 19612
rect 4048 19556 4104 19612
rect 4104 19556 4108 19612
rect 4044 19552 4108 19556
rect 3068 19068 3132 19072
rect 3068 19012 3072 19068
rect 3072 19012 3128 19068
rect 3128 19012 3132 19068
rect 3068 19008 3132 19012
rect 3148 19068 3212 19072
rect 3148 19012 3152 19068
rect 3152 19012 3208 19068
rect 3208 19012 3212 19068
rect 3148 19008 3212 19012
rect 3228 19068 3292 19072
rect 3228 19012 3232 19068
rect 3232 19012 3288 19068
rect 3288 19012 3292 19068
rect 3228 19008 3292 19012
rect 3308 19068 3372 19072
rect 3308 19012 3312 19068
rect 3312 19012 3368 19068
rect 3368 19012 3372 19068
rect 3308 19008 3372 19012
rect 3804 18524 3868 18528
rect 3804 18468 3808 18524
rect 3808 18468 3864 18524
rect 3864 18468 3868 18524
rect 3804 18464 3868 18468
rect 3884 18524 3948 18528
rect 3884 18468 3888 18524
rect 3888 18468 3944 18524
rect 3944 18468 3948 18524
rect 3884 18464 3948 18468
rect 3964 18524 4028 18528
rect 3964 18468 3968 18524
rect 3968 18468 4024 18524
rect 4024 18468 4028 18524
rect 3964 18464 4028 18468
rect 4044 18524 4108 18528
rect 4044 18468 4048 18524
rect 4048 18468 4104 18524
rect 4104 18468 4108 18524
rect 4044 18464 4108 18468
rect 3068 17980 3132 17984
rect 3068 17924 3072 17980
rect 3072 17924 3128 17980
rect 3128 17924 3132 17980
rect 3068 17920 3132 17924
rect 3148 17980 3212 17984
rect 3148 17924 3152 17980
rect 3152 17924 3208 17980
rect 3208 17924 3212 17980
rect 3148 17920 3212 17924
rect 3228 17980 3292 17984
rect 3228 17924 3232 17980
rect 3232 17924 3288 17980
rect 3288 17924 3292 17980
rect 3228 17920 3292 17924
rect 3308 17980 3372 17984
rect 3308 17924 3312 17980
rect 3312 17924 3368 17980
rect 3368 17924 3372 17980
rect 3308 17920 3372 17924
rect 3804 17436 3868 17440
rect 3804 17380 3808 17436
rect 3808 17380 3864 17436
rect 3864 17380 3868 17436
rect 3804 17376 3868 17380
rect 3884 17436 3948 17440
rect 3884 17380 3888 17436
rect 3888 17380 3944 17436
rect 3944 17380 3948 17436
rect 3884 17376 3948 17380
rect 3964 17436 4028 17440
rect 3964 17380 3968 17436
rect 3968 17380 4024 17436
rect 4024 17380 4028 17436
rect 3964 17376 4028 17380
rect 4044 17436 4108 17440
rect 4044 17380 4048 17436
rect 4048 17380 4104 17436
rect 4104 17380 4108 17436
rect 4044 17376 4108 17380
rect 3068 16892 3132 16896
rect 3068 16836 3072 16892
rect 3072 16836 3128 16892
rect 3128 16836 3132 16892
rect 3068 16832 3132 16836
rect 3148 16892 3212 16896
rect 3148 16836 3152 16892
rect 3152 16836 3208 16892
rect 3208 16836 3212 16892
rect 3148 16832 3212 16836
rect 3228 16892 3292 16896
rect 3228 16836 3232 16892
rect 3232 16836 3288 16892
rect 3288 16836 3292 16892
rect 3228 16832 3292 16836
rect 3308 16892 3372 16896
rect 3308 16836 3312 16892
rect 3312 16836 3368 16892
rect 3368 16836 3372 16892
rect 3308 16832 3372 16836
rect 3804 16348 3868 16352
rect 3804 16292 3808 16348
rect 3808 16292 3864 16348
rect 3864 16292 3868 16348
rect 3804 16288 3868 16292
rect 3884 16348 3948 16352
rect 3884 16292 3888 16348
rect 3888 16292 3944 16348
rect 3944 16292 3948 16348
rect 3884 16288 3948 16292
rect 3964 16348 4028 16352
rect 3964 16292 3968 16348
rect 3968 16292 4024 16348
rect 4024 16292 4028 16348
rect 3964 16288 4028 16292
rect 4044 16348 4108 16352
rect 4044 16292 4048 16348
rect 4048 16292 4104 16348
rect 4104 16292 4108 16348
rect 4044 16288 4108 16292
rect 3068 15804 3132 15808
rect 3068 15748 3072 15804
rect 3072 15748 3128 15804
rect 3128 15748 3132 15804
rect 3068 15744 3132 15748
rect 3148 15804 3212 15808
rect 3148 15748 3152 15804
rect 3152 15748 3208 15804
rect 3208 15748 3212 15804
rect 3148 15744 3212 15748
rect 3228 15804 3292 15808
rect 3228 15748 3232 15804
rect 3232 15748 3288 15804
rect 3288 15748 3292 15804
rect 3228 15744 3292 15748
rect 3308 15804 3372 15808
rect 3308 15748 3312 15804
rect 3312 15748 3368 15804
rect 3368 15748 3372 15804
rect 3308 15744 3372 15748
rect 3804 15260 3868 15264
rect 3804 15204 3808 15260
rect 3808 15204 3864 15260
rect 3864 15204 3868 15260
rect 3804 15200 3868 15204
rect 3884 15260 3948 15264
rect 3884 15204 3888 15260
rect 3888 15204 3944 15260
rect 3944 15204 3948 15260
rect 3884 15200 3948 15204
rect 3964 15260 4028 15264
rect 3964 15204 3968 15260
rect 3968 15204 4024 15260
rect 4024 15204 4028 15260
rect 3964 15200 4028 15204
rect 4044 15260 4108 15264
rect 4044 15204 4048 15260
rect 4048 15204 4104 15260
rect 4104 15204 4108 15260
rect 4044 15200 4108 15204
rect 3068 14716 3132 14720
rect 3068 14660 3072 14716
rect 3072 14660 3128 14716
rect 3128 14660 3132 14716
rect 3068 14656 3132 14660
rect 3148 14716 3212 14720
rect 3148 14660 3152 14716
rect 3152 14660 3208 14716
rect 3208 14660 3212 14716
rect 3148 14656 3212 14660
rect 3228 14716 3292 14720
rect 3228 14660 3232 14716
rect 3232 14660 3288 14716
rect 3288 14660 3292 14716
rect 3228 14656 3292 14660
rect 3308 14716 3372 14720
rect 3308 14660 3312 14716
rect 3312 14660 3368 14716
rect 3368 14660 3372 14716
rect 3308 14656 3372 14660
rect 3804 14172 3868 14176
rect 3804 14116 3808 14172
rect 3808 14116 3864 14172
rect 3864 14116 3868 14172
rect 3804 14112 3868 14116
rect 3884 14172 3948 14176
rect 3884 14116 3888 14172
rect 3888 14116 3944 14172
rect 3944 14116 3948 14172
rect 3884 14112 3948 14116
rect 3964 14172 4028 14176
rect 3964 14116 3968 14172
rect 3968 14116 4024 14172
rect 4024 14116 4028 14172
rect 3964 14112 4028 14116
rect 4044 14172 4108 14176
rect 4044 14116 4048 14172
rect 4048 14116 4104 14172
rect 4104 14116 4108 14172
rect 4044 14112 4108 14116
rect 86356 13636 86420 13700
rect 3068 13628 3132 13632
rect 3068 13572 3072 13628
rect 3072 13572 3128 13628
rect 3128 13572 3132 13628
rect 3068 13568 3132 13572
rect 3148 13628 3212 13632
rect 3148 13572 3152 13628
rect 3152 13572 3208 13628
rect 3208 13572 3212 13628
rect 3148 13568 3212 13572
rect 3228 13628 3292 13632
rect 3228 13572 3232 13628
rect 3232 13572 3288 13628
rect 3288 13572 3292 13628
rect 3228 13568 3292 13572
rect 3308 13628 3372 13632
rect 3308 13572 3312 13628
rect 3312 13572 3368 13628
rect 3368 13572 3372 13628
rect 3308 13568 3372 13572
rect 3804 13084 3868 13088
rect 3804 13028 3808 13084
rect 3808 13028 3864 13084
rect 3864 13028 3868 13084
rect 3804 13024 3868 13028
rect 3884 13084 3948 13088
rect 3884 13028 3888 13084
rect 3888 13028 3944 13084
rect 3944 13028 3948 13084
rect 3884 13024 3948 13028
rect 3964 13084 4028 13088
rect 3964 13028 3968 13084
rect 3968 13028 4024 13084
rect 4024 13028 4028 13084
rect 3964 13024 4028 13028
rect 4044 13084 4108 13088
rect 4044 13028 4048 13084
rect 4048 13028 4104 13084
rect 4104 13028 4108 13084
rect 4044 13024 4108 13028
rect 86540 12548 86604 12612
rect 3068 12540 3132 12544
rect 3068 12484 3072 12540
rect 3072 12484 3128 12540
rect 3128 12484 3132 12540
rect 3068 12480 3132 12484
rect 3148 12540 3212 12544
rect 3148 12484 3152 12540
rect 3152 12484 3208 12540
rect 3208 12484 3212 12540
rect 3148 12480 3212 12484
rect 3228 12540 3292 12544
rect 3228 12484 3232 12540
rect 3232 12484 3288 12540
rect 3288 12484 3292 12540
rect 3228 12480 3292 12484
rect 3308 12540 3372 12544
rect 3308 12484 3312 12540
rect 3312 12484 3368 12540
rect 3368 12484 3372 12540
rect 3308 12480 3372 12484
rect 3804 11996 3868 12000
rect 3804 11940 3808 11996
rect 3808 11940 3864 11996
rect 3864 11940 3868 11996
rect 3804 11936 3868 11940
rect 3884 11996 3948 12000
rect 3884 11940 3888 11996
rect 3888 11940 3944 11996
rect 3944 11940 3948 11996
rect 3884 11936 3948 11940
rect 3964 11996 4028 12000
rect 3964 11940 3968 11996
rect 3968 11940 4024 11996
rect 4024 11940 4028 11996
rect 3964 11936 4028 11940
rect 4044 11996 4108 12000
rect 4044 11940 4048 11996
rect 4048 11940 4104 11996
rect 4104 11940 4108 11996
rect 4044 11936 4108 11940
rect 3068 11452 3132 11456
rect 3068 11396 3072 11452
rect 3072 11396 3128 11452
rect 3128 11396 3132 11452
rect 3068 11392 3132 11396
rect 3148 11452 3212 11456
rect 3148 11396 3152 11452
rect 3152 11396 3208 11452
rect 3208 11396 3212 11452
rect 3148 11392 3212 11396
rect 3228 11452 3292 11456
rect 3228 11396 3232 11452
rect 3232 11396 3288 11452
rect 3288 11396 3292 11452
rect 3228 11392 3292 11396
rect 3308 11452 3372 11456
rect 3308 11396 3312 11452
rect 3312 11396 3368 11452
rect 3368 11396 3372 11452
rect 3308 11392 3372 11396
rect 88380 11052 88444 11116
rect 3804 10908 3868 10912
rect 3804 10852 3808 10908
rect 3808 10852 3864 10908
rect 3864 10852 3868 10908
rect 3804 10848 3868 10852
rect 3884 10908 3948 10912
rect 3884 10852 3888 10908
rect 3888 10852 3944 10908
rect 3944 10852 3948 10908
rect 3884 10848 3948 10852
rect 3964 10908 4028 10912
rect 3964 10852 3968 10908
rect 3968 10852 4024 10908
rect 4024 10852 4028 10908
rect 3964 10848 4028 10852
rect 4044 10908 4108 10912
rect 4044 10852 4048 10908
rect 4048 10852 4104 10908
rect 4104 10852 4108 10908
rect 4044 10848 4108 10852
rect 3068 10364 3132 10368
rect 3068 10308 3072 10364
rect 3072 10308 3128 10364
rect 3128 10308 3132 10364
rect 3068 10304 3132 10308
rect 3148 10364 3212 10368
rect 3148 10308 3152 10364
rect 3152 10308 3208 10364
rect 3208 10308 3212 10364
rect 3148 10304 3212 10308
rect 3228 10364 3292 10368
rect 3228 10308 3232 10364
rect 3232 10308 3288 10364
rect 3288 10308 3292 10364
rect 3228 10304 3292 10308
rect 3308 10364 3372 10368
rect 3308 10308 3312 10364
rect 3312 10308 3368 10364
rect 3368 10308 3372 10364
rect 3308 10304 3372 10308
rect 3804 9820 3868 9824
rect 3804 9764 3808 9820
rect 3808 9764 3864 9820
rect 3864 9764 3868 9820
rect 3804 9760 3868 9764
rect 3884 9820 3948 9824
rect 3884 9764 3888 9820
rect 3888 9764 3944 9820
rect 3944 9764 3948 9820
rect 3884 9760 3948 9764
rect 3964 9820 4028 9824
rect 3964 9764 3968 9820
rect 3968 9764 4024 9820
rect 4024 9764 4028 9820
rect 3964 9760 4028 9764
rect 4044 9820 4108 9824
rect 4044 9764 4048 9820
rect 4048 9764 4104 9820
rect 4104 9764 4108 9820
rect 4044 9760 4108 9764
rect 88748 9556 88812 9620
rect 3068 9276 3132 9280
rect 3068 9220 3072 9276
rect 3072 9220 3128 9276
rect 3128 9220 3132 9276
rect 3068 9216 3132 9220
rect 3148 9276 3212 9280
rect 3148 9220 3152 9276
rect 3152 9220 3208 9276
rect 3208 9220 3212 9276
rect 3148 9216 3212 9220
rect 3228 9276 3292 9280
rect 3228 9220 3232 9276
rect 3232 9220 3288 9276
rect 3288 9220 3292 9276
rect 3228 9216 3292 9220
rect 3308 9276 3372 9280
rect 3308 9220 3312 9276
rect 3312 9220 3368 9276
rect 3368 9220 3372 9276
rect 3308 9216 3372 9220
rect 3804 8732 3868 8736
rect 3804 8676 3808 8732
rect 3808 8676 3864 8732
rect 3864 8676 3868 8732
rect 3804 8672 3868 8676
rect 3884 8732 3948 8736
rect 3884 8676 3888 8732
rect 3888 8676 3944 8732
rect 3944 8676 3948 8732
rect 3884 8672 3948 8676
rect 3964 8732 4028 8736
rect 3964 8676 3968 8732
rect 3968 8676 4024 8732
rect 4024 8676 4028 8732
rect 3964 8672 4028 8676
rect 4044 8732 4108 8736
rect 4044 8676 4048 8732
rect 4048 8676 4104 8732
rect 4104 8676 4108 8732
rect 4044 8672 4108 8676
rect 88380 8332 88444 8396
rect 86908 8196 86972 8260
rect 3068 8188 3132 8192
rect 3068 8132 3072 8188
rect 3072 8132 3128 8188
rect 3128 8132 3132 8188
rect 3068 8128 3132 8132
rect 3148 8188 3212 8192
rect 3148 8132 3152 8188
rect 3152 8132 3208 8188
rect 3208 8132 3212 8188
rect 3148 8128 3212 8132
rect 3228 8188 3292 8192
rect 3228 8132 3232 8188
rect 3232 8132 3288 8188
rect 3288 8132 3292 8188
rect 3228 8128 3292 8132
rect 3308 8188 3372 8192
rect 3308 8132 3312 8188
rect 3312 8132 3368 8188
rect 3368 8132 3372 8188
rect 3308 8128 3372 8132
rect 87092 7924 87156 7988
rect 3804 7644 3868 7648
rect 3804 7588 3808 7644
rect 3808 7588 3864 7644
rect 3864 7588 3868 7644
rect 3804 7584 3868 7588
rect 3884 7644 3948 7648
rect 3884 7588 3888 7644
rect 3888 7588 3944 7644
rect 3944 7588 3948 7644
rect 3884 7584 3948 7588
rect 3964 7644 4028 7648
rect 3964 7588 3968 7644
rect 3968 7588 4024 7644
rect 4024 7588 4028 7644
rect 3964 7584 4028 7588
rect 4044 7644 4108 7648
rect 4044 7588 4048 7644
rect 4048 7588 4104 7644
rect 4104 7588 4108 7644
rect 4044 7584 4108 7588
rect 3068 7100 3132 7104
rect 3068 7044 3072 7100
rect 3072 7044 3128 7100
rect 3128 7044 3132 7100
rect 3068 7040 3132 7044
rect 3148 7100 3212 7104
rect 3148 7044 3152 7100
rect 3152 7044 3208 7100
rect 3208 7044 3212 7100
rect 3148 7040 3212 7044
rect 3228 7100 3292 7104
rect 3228 7044 3232 7100
rect 3232 7044 3288 7100
rect 3288 7044 3292 7100
rect 3228 7040 3292 7044
rect 3308 7100 3372 7104
rect 3308 7044 3312 7100
rect 3312 7044 3368 7100
rect 3368 7044 3372 7100
rect 3308 7040 3372 7044
rect 3804 6556 3868 6560
rect 3804 6500 3808 6556
rect 3808 6500 3864 6556
rect 3864 6500 3868 6556
rect 3804 6496 3868 6500
rect 3884 6556 3948 6560
rect 3884 6500 3888 6556
rect 3888 6500 3944 6556
rect 3944 6500 3948 6556
rect 3884 6496 3948 6500
rect 3964 6556 4028 6560
rect 3964 6500 3968 6556
rect 3968 6500 4024 6556
rect 4024 6500 4028 6556
rect 3964 6496 4028 6500
rect 4044 6556 4108 6560
rect 4044 6500 4048 6556
rect 4048 6500 4104 6556
rect 4104 6500 4108 6556
rect 4044 6496 4108 6500
rect 3068 6012 3132 6016
rect 3068 5956 3072 6012
rect 3072 5956 3128 6012
rect 3128 5956 3132 6012
rect 3068 5952 3132 5956
rect 3148 6012 3212 6016
rect 3148 5956 3152 6012
rect 3152 5956 3208 6012
rect 3208 5956 3212 6012
rect 3148 5952 3212 5956
rect 3228 6012 3292 6016
rect 3228 5956 3232 6012
rect 3232 5956 3288 6012
rect 3288 5956 3292 6012
rect 3228 5952 3292 5956
rect 3308 6012 3372 6016
rect 3308 5956 3312 6012
rect 3312 5956 3368 6012
rect 3368 5956 3372 6012
rect 3308 5952 3372 5956
rect 72952 6012 73016 6016
rect 72952 5956 72956 6012
rect 72956 5956 73012 6012
rect 73012 5956 73016 6012
rect 72952 5952 73016 5956
rect 73032 6012 73096 6016
rect 73032 5956 73036 6012
rect 73036 5956 73092 6012
rect 73092 5956 73096 6012
rect 73032 5952 73096 5956
rect 73112 6012 73176 6016
rect 73112 5956 73116 6012
rect 73116 5956 73172 6012
rect 73172 5956 73176 6012
rect 73112 5952 73176 5956
rect 73192 6012 73256 6016
rect 73192 5956 73196 6012
rect 73196 5956 73252 6012
rect 73252 5956 73256 6012
rect 73192 5952 73256 5956
rect 88564 5944 88628 5948
rect 88564 5888 88578 5944
rect 88578 5888 88628 5944
rect 88564 5884 88628 5888
rect 47716 5748 47780 5812
rect 48084 5612 48148 5676
rect 88196 5536 88260 5540
rect 88196 5480 88246 5536
rect 88246 5480 88260 5536
rect 88196 5476 88260 5480
rect 3804 5468 3868 5472
rect 3804 5412 3808 5468
rect 3808 5412 3864 5468
rect 3864 5412 3868 5468
rect 3804 5408 3868 5412
rect 3884 5468 3948 5472
rect 3884 5412 3888 5468
rect 3888 5412 3944 5468
rect 3944 5412 3948 5468
rect 3884 5408 3948 5412
rect 3964 5468 4028 5472
rect 3964 5412 3968 5468
rect 3968 5412 4024 5468
rect 4024 5412 4028 5468
rect 3964 5408 4028 5412
rect 4044 5468 4108 5472
rect 4044 5412 4048 5468
rect 4048 5412 4104 5468
rect 4104 5412 4108 5468
rect 4044 5408 4108 5412
rect 37612 5468 37676 5472
rect 37612 5412 37616 5468
rect 37616 5412 37672 5468
rect 37672 5412 37676 5468
rect 37612 5408 37676 5412
rect 37692 5468 37756 5472
rect 37692 5412 37696 5468
rect 37696 5412 37752 5468
rect 37752 5412 37756 5468
rect 37692 5408 37756 5412
rect 37772 5468 37836 5472
rect 37772 5412 37776 5468
rect 37776 5412 37832 5468
rect 37832 5412 37836 5468
rect 37772 5408 37836 5412
rect 37852 5468 37916 5472
rect 37852 5412 37856 5468
rect 37856 5412 37912 5468
rect 37912 5412 37916 5468
rect 37852 5408 37916 5412
rect 73612 5468 73676 5472
rect 73612 5412 73616 5468
rect 73616 5412 73672 5468
rect 73672 5412 73676 5468
rect 73612 5408 73676 5412
rect 73692 5468 73756 5472
rect 73692 5412 73696 5468
rect 73696 5412 73752 5468
rect 73752 5412 73756 5468
rect 73692 5408 73756 5412
rect 73772 5468 73836 5472
rect 73772 5412 73776 5468
rect 73776 5412 73832 5468
rect 73832 5412 73836 5468
rect 73772 5408 73836 5412
rect 73852 5468 73916 5472
rect 73852 5412 73856 5468
rect 73856 5412 73912 5468
rect 73912 5412 73916 5468
rect 73852 5408 73916 5412
rect 86540 5400 86604 5404
rect 86540 5344 86554 5400
rect 86554 5344 86604 5400
rect 86540 5340 86604 5344
rect 36952 4924 37016 4928
rect 36952 4868 36956 4924
rect 36956 4868 37012 4924
rect 37012 4868 37016 4924
rect 36952 4864 37016 4868
rect 37032 4924 37096 4928
rect 37032 4868 37036 4924
rect 37036 4868 37092 4924
rect 37092 4868 37096 4924
rect 37032 4864 37096 4868
rect 37112 4924 37176 4928
rect 37112 4868 37116 4924
rect 37116 4868 37172 4924
rect 37172 4868 37176 4924
rect 37112 4864 37176 4868
rect 37192 4924 37256 4928
rect 37192 4868 37196 4924
rect 37196 4868 37252 4924
rect 37252 4868 37256 4924
rect 37192 4864 37256 4868
rect 72952 4924 73016 4928
rect 72952 4868 72956 4924
rect 72956 4868 73012 4924
rect 73012 4868 73016 4924
rect 72952 4864 73016 4868
rect 73032 4924 73096 4928
rect 73032 4868 73036 4924
rect 73036 4868 73092 4924
rect 73092 4868 73096 4924
rect 73032 4864 73096 4868
rect 73112 4924 73176 4928
rect 73112 4868 73116 4924
rect 73116 4868 73172 4924
rect 73172 4868 73176 4924
rect 73112 4864 73176 4868
rect 73192 4924 73256 4928
rect 73192 4868 73196 4924
rect 73196 4868 73252 4924
rect 73252 4868 73256 4924
rect 73192 4864 73256 4868
rect 87276 4856 87340 4860
rect 87276 4800 87290 4856
rect 87290 4800 87340 4856
rect 87276 4796 87340 4800
rect 47900 4524 47964 4588
rect 37612 4380 37676 4384
rect 37612 4324 37616 4380
rect 37616 4324 37672 4380
rect 37672 4324 37676 4380
rect 37612 4320 37676 4324
rect 37692 4380 37756 4384
rect 37692 4324 37696 4380
rect 37696 4324 37752 4380
rect 37752 4324 37756 4380
rect 37692 4320 37756 4324
rect 37772 4380 37836 4384
rect 37772 4324 37776 4380
rect 37776 4324 37832 4380
rect 37832 4324 37836 4380
rect 37772 4320 37836 4324
rect 37852 4380 37916 4384
rect 37852 4324 37856 4380
rect 37856 4324 37912 4380
rect 37912 4324 37916 4380
rect 37852 4320 37916 4324
rect 73612 4380 73676 4384
rect 73612 4324 73616 4380
rect 73616 4324 73672 4380
rect 73672 4324 73676 4380
rect 73612 4320 73676 4324
rect 73692 4380 73756 4384
rect 73692 4324 73696 4380
rect 73696 4324 73752 4380
rect 73752 4324 73756 4380
rect 73692 4320 73756 4324
rect 73772 4380 73836 4384
rect 73772 4324 73776 4380
rect 73776 4324 73832 4380
rect 73832 4324 73836 4380
rect 73772 4320 73836 4324
rect 73852 4380 73916 4384
rect 73852 4324 73856 4380
rect 73856 4324 73912 4380
rect 73912 4324 73916 4380
rect 73852 4320 73916 4324
rect 36952 3836 37016 3840
rect 36952 3780 36956 3836
rect 36956 3780 37012 3836
rect 37012 3780 37016 3836
rect 36952 3776 37016 3780
rect 37032 3836 37096 3840
rect 37032 3780 37036 3836
rect 37036 3780 37092 3836
rect 37092 3780 37096 3836
rect 37032 3776 37096 3780
rect 37112 3836 37176 3840
rect 37112 3780 37116 3836
rect 37116 3780 37172 3836
rect 37172 3780 37176 3836
rect 37112 3776 37176 3780
rect 37192 3836 37256 3840
rect 37192 3780 37196 3836
rect 37196 3780 37252 3836
rect 37252 3780 37256 3836
rect 37192 3776 37256 3780
rect 72952 3836 73016 3840
rect 72952 3780 72956 3836
rect 72956 3780 73012 3836
rect 73012 3780 73016 3836
rect 72952 3776 73016 3780
rect 73032 3836 73096 3840
rect 73032 3780 73036 3836
rect 73036 3780 73092 3836
rect 73092 3780 73096 3836
rect 73032 3776 73096 3780
rect 73112 3836 73176 3840
rect 73112 3780 73116 3836
rect 73116 3780 73172 3836
rect 73172 3780 73176 3836
rect 73112 3776 73176 3780
rect 73192 3836 73256 3840
rect 73192 3780 73196 3836
rect 73196 3780 73252 3836
rect 73252 3780 73256 3836
rect 73192 3776 73256 3780
rect 37612 3292 37676 3296
rect 37612 3236 37616 3292
rect 37616 3236 37672 3292
rect 37672 3236 37676 3292
rect 37612 3232 37676 3236
rect 37692 3292 37756 3296
rect 37692 3236 37696 3292
rect 37696 3236 37752 3292
rect 37752 3236 37756 3292
rect 37692 3232 37756 3236
rect 37772 3292 37836 3296
rect 37772 3236 37776 3292
rect 37776 3236 37832 3292
rect 37832 3236 37836 3292
rect 37772 3232 37836 3236
rect 37852 3292 37916 3296
rect 37852 3236 37856 3292
rect 37856 3236 37912 3292
rect 37912 3236 37916 3292
rect 37852 3232 37916 3236
rect 73612 3292 73676 3296
rect 73612 3236 73616 3292
rect 73616 3236 73672 3292
rect 73672 3236 73676 3292
rect 73612 3232 73676 3236
rect 73692 3292 73756 3296
rect 73692 3236 73696 3292
rect 73696 3236 73752 3292
rect 73752 3236 73756 3292
rect 73692 3232 73756 3236
rect 73772 3292 73836 3296
rect 73772 3236 73776 3292
rect 73776 3236 73832 3292
rect 73832 3236 73836 3292
rect 73772 3232 73836 3236
rect 73852 3292 73916 3296
rect 73852 3236 73856 3292
rect 73856 3236 73912 3292
rect 73912 3236 73916 3292
rect 73852 3232 73916 3236
rect 36952 2748 37016 2752
rect 36952 2692 36956 2748
rect 36956 2692 37012 2748
rect 37012 2692 37016 2748
rect 36952 2688 37016 2692
rect 37032 2748 37096 2752
rect 37032 2692 37036 2748
rect 37036 2692 37092 2748
rect 37092 2692 37096 2748
rect 37032 2688 37096 2692
rect 37112 2748 37176 2752
rect 37112 2692 37116 2748
rect 37116 2692 37172 2748
rect 37172 2692 37176 2748
rect 37112 2688 37176 2692
rect 37192 2748 37256 2752
rect 37192 2692 37196 2748
rect 37196 2692 37252 2748
rect 37252 2692 37256 2748
rect 37192 2688 37256 2692
rect 72952 2748 73016 2752
rect 72952 2692 72956 2748
rect 72956 2692 73012 2748
rect 73012 2692 73016 2748
rect 72952 2688 73016 2692
rect 73032 2748 73096 2752
rect 73032 2692 73036 2748
rect 73036 2692 73092 2748
rect 73092 2692 73096 2748
rect 73032 2688 73096 2692
rect 73112 2748 73176 2752
rect 73112 2692 73116 2748
rect 73116 2692 73172 2748
rect 73172 2692 73176 2748
rect 73112 2688 73176 2692
rect 73192 2748 73256 2752
rect 73192 2692 73196 2748
rect 73196 2692 73252 2748
rect 73252 2692 73256 2748
rect 73192 2688 73256 2692
rect 37612 2204 37676 2208
rect 37612 2148 37616 2204
rect 37616 2148 37672 2204
rect 37672 2148 37676 2204
rect 37612 2144 37676 2148
rect 37692 2204 37756 2208
rect 37692 2148 37696 2204
rect 37696 2148 37752 2204
rect 37752 2148 37756 2204
rect 37692 2144 37756 2148
rect 37772 2204 37836 2208
rect 37772 2148 37776 2204
rect 37776 2148 37832 2204
rect 37832 2148 37836 2204
rect 37772 2144 37836 2148
rect 37852 2204 37916 2208
rect 37852 2148 37856 2204
rect 37856 2148 37912 2204
rect 37912 2148 37916 2204
rect 37852 2144 37916 2148
rect 73612 2204 73676 2208
rect 73612 2148 73616 2204
rect 73616 2148 73672 2204
rect 73672 2148 73676 2204
rect 73612 2144 73676 2148
rect 73692 2204 73756 2208
rect 73692 2148 73696 2204
rect 73696 2148 73752 2204
rect 73752 2148 73756 2204
rect 73692 2144 73756 2148
rect 73772 2204 73836 2208
rect 73772 2148 73776 2204
rect 73776 2148 73832 2204
rect 73832 2148 73836 2204
rect 73772 2144 73836 2148
rect 73852 2204 73916 2208
rect 73852 2148 73856 2204
rect 73856 2148 73912 2204
rect 73912 2148 73916 2204
rect 73852 2144 73916 2148
<< metal4 >>
rect -1076 97882 -756 97924
rect -1076 97646 -1034 97882
rect -798 97646 -756 97882
rect -1076 69754 -756 97646
rect -1076 69518 -1034 69754
rect -798 69518 -756 69754
rect -1076 36354 -756 69518
rect -1076 36118 -1034 36354
rect -798 36118 -756 36354
rect -1076 274 -756 36118
rect -416 97222 -96 97264
rect -416 96986 -374 97222
rect -138 96986 -96 97222
rect -416 69094 -96 96986
rect 36944 97222 37264 97924
rect 36944 96986 36986 97222
rect 37222 96986 37264 97222
rect 8523 95300 8589 95301
rect 8523 95236 8524 95300
rect 8588 95236 8589 95300
rect 8523 95235 8589 95236
rect -416 68858 -374 69094
rect -138 68858 -96 69094
rect -416 35694 -96 68858
rect 3060 91968 3380 91984
rect 3060 91904 3068 91968
rect 3132 91904 3148 91968
rect 3212 91904 3228 91968
rect 3292 91904 3308 91968
rect 3372 91904 3380 91968
rect 3060 90880 3380 91904
rect 3060 90816 3068 90880
rect 3132 90816 3148 90880
rect 3212 90816 3228 90880
rect 3292 90816 3308 90880
rect 3372 90816 3380 90880
rect 3060 89792 3380 90816
rect 3060 89728 3068 89792
rect 3132 89728 3148 89792
rect 3212 89728 3228 89792
rect 3292 89728 3308 89792
rect 3372 89728 3380 89792
rect 3060 88704 3380 89728
rect 3060 88640 3068 88704
rect 3132 88640 3148 88704
rect 3212 88640 3228 88704
rect 3292 88640 3308 88704
rect 3372 88640 3380 88704
rect 3060 87616 3380 88640
rect 3060 87552 3068 87616
rect 3132 87552 3148 87616
rect 3212 87552 3228 87616
rect 3292 87552 3308 87616
rect 3372 87552 3380 87616
rect 3060 86528 3380 87552
rect 3060 86464 3068 86528
rect 3132 86464 3148 86528
rect 3212 86464 3228 86528
rect 3292 86464 3308 86528
rect 3372 86464 3380 86528
rect 3060 85440 3380 86464
rect 3060 85376 3068 85440
rect 3132 85376 3148 85440
rect 3212 85376 3228 85440
rect 3292 85376 3308 85440
rect 3372 85376 3380 85440
rect 3060 84352 3380 85376
rect 3060 84288 3068 84352
rect 3132 84288 3148 84352
rect 3212 84288 3228 84352
rect 3292 84288 3308 84352
rect 3372 84288 3380 84352
rect 3060 83264 3380 84288
rect 3060 83200 3068 83264
rect 3132 83200 3148 83264
rect 3212 83200 3228 83264
rect 3292 83200 3308 83264
rect 3372 83200 3380 83264
rect 3060 82176 3380 83200
rect 3060 82112 3068 82176
rect 3132 82112 3148 82176
rect 3212 82112 3228 82176
rect 3292 82112 3308 82176
rect 3372 82112 3380 82176
rect 3060 81088 3380 82112
rect 3060 81024 3068 81088
rect 3132 81024 3148 81088
rect 3212 81024 3228 81088
rect 3292 81024 3308 81088
rect 3372 81024 3380 81088
rect 3060 80000 3380 81024
rect 3060 79936 3068 80000
rect 3132 79936 3148 80000
rect 3212 79936 3228 80000
rect 3292 79936 3308 80000
rect 3372 79936 3380 80000
rect 3060 78912 3380 79936
rect 3060 78848 3068 78912
rect 3132 78848 3148 78912
rect 3212 78848 3228 78912
rect 3292 78848 3308 78912
rect 3372 78848 3380 78912
rect 3060 77824 3380 78848
rect 3060 77760 3068 77824
rect 3132 77760 3148 77824
rect 3212 77760 3228 77824
rect 3292 77760 3308 77824
rect 3372 77760 3380 77824
rect 3060 76736 3380 77760
rect 3060 76672 3068 76736
rect 3132 76672 3148 76736
rect 3212 76672 3228 76736
rect 3292 76672 3308 76736
rect 3372 76672 3380 76736
rect 3060 75648 3380 76672
rect 3060 75584 3068 75648
rect 3132 75584 3148 75648
rect 3212 75584 3228 75648
rect 3292 75584 3308 75648
rect 3372 75584 3380 75648
rect 3060 74560 3380 75584
rect 3060 74496 3068 74560
rect 3132 74496 3148 74560
rect 3212 74496 3228 74560
rect 3292 74496 3308 74560
rect 3372 74496 3380 74560
rect 3060 73472 3380 74496
rect 3060 73408 3068 73472
rect 3132 73408 3148 73472
rect 3212 73408 3228 73472
rect 3292 73408 3308 73472
rect 3372 73408 3380 73472
rect 3060 72384 3380 73408
rect 3060 72320 3068 72384
rect 3132 72320 3148 72384
rect 3212 72320 3228 72384
rect 3292 72320 3308 72384
rect 3372 72320 3380 72384
rect 3060 71296 3380 72320
rect 3060 71232 3068 71296
rect 3132 71232 3148 71296
rect 3212 71232 3228 71296
rect 3292 71232 3308 71296
rect 3372 71232 3380 71296
rect 3060 70208 3380 71232
rect 3060 70144 3068 70208
rect 3132 70144 3148 70208
rect 3212 70144 3228 70208
rect 3292 70144 3308 70208
rect 3372 70144 3380 70208
rect 3060 69120 3380 70144
rect 3060 69056 3068 69120
rect 3132 69094 3148 69120
rect 3212 69094 3228 69120
rect 3292 69094 3308 69120
rect 3372 69056 3380 69120
rect 3060 68858 3102 69056
rect 3338 68858 3380 69056
rect 3060 68032 3380 68858
rect 3060 67968 3068 68032
rect 3132 67968 3148 68032
rect 3212 67968 3228 68032
rect 3292 67968 3308 68032
rect 3372 67968 3380 68032
rect 3060 66944 3380 67968
rect 3060 66880 3068 66944
rect 3132 66880 3148 66944
rect 3212 66880 3228 66944
rect 3292 66880 3308 66944
rect 3372 66880 3380 66944
rect 3060 65856 3380 66880
rect 3060 65792 3068 65856
rect 3132 65792 3148 65856
rect 3212 65792 3228 65856
rect 3292 65792 3308 65856
rect 3372 65792 3380 65856
rect 3060 64768 3380 65792
rect 3060 64704 3068 64768
rect 3132 64704 3148 64768
rect 3212 64704 3228 64768
rect 3292 64704 3308 64768
rect 3372 64704 3380 64768
rect 3060 63680 3380 64704
rect 3060 63616 3068 63680
rect 3132 63616 3148 63680
rect 3212 63616 3228 63680
rect 3292 63616 3308 63680
rect 3372 63616 3380 63680
rect 3060 62592 3380 63616
rect 3060 62528 3068 62592
rect 3132 62528 3148 62592
rect 3212 62528 3228 62592
rect 3292 62528 3308 62592
rect 3372 62528 3380 62592
rect 3060 61504 3380 62528
rect 3060 61440 3068 61504
rect 3132 61440 3148 61504
rect 3212 61440 3228 61504
rect 3292 61440 3308 61504
rect 3372 61440 3380 61504
rect 3060 60416 3380 61440
rect 3060 60352 3068 60416
rect 3132 60352 3148 60416
rect 3212 60352 3228 60416
rect 3292 60352 3308 60416
rect 3372 60352 3380 60416
rect 3060 59328 3380 60352
rect 3060 59264 3068 59328
rect 3132 59264 3148 59328
rect 3212 59264 3228 59328
rect 3292 59264 3308 59328
rect 3372 59264 3380 59328
rect 3060 58240 3380 59264
rect 3060 58176 3068 58240
rect 3132 58176 3148 58240
rect 3212 58176 3228 58240
rect 3292 58176 3308 58240
rect 3372 58176 3380 58240
rect 3060 57152 3380 58176
rect 3060 57088 3068 57152
rect 3132 57088 3148 57152
rect 3212 57088 3228 57152
rect 3292 57088 3308 57152
rect 3372 57088 3380 57152
rect 3060 56064 3380 57088
rect 3060 56000 3068 56064
rect 3132 56000 3148 56064
rect 3212 56000 3228 56064
rect 3292 56000 3308 56064
rect 3372 56000 3380 56064
rect 3060 54976 3380 56000
rect 3060 54912 3068 54976
rect 3132 54912 3148 54976
rect 3212 54912 3228 54976
rect 3292 54912 3308 54976
rect 3372 54912 3380 54976
rect 3060 53888 3380 54912
rect 3060 53824 3068 53888
rect 3132 53824 3148 53888
rect 3212 53824 3228 53888
rect 3292 53824 3308 53888
rect 3372 53824 3380 53888
rect 3060 52800 3380 53824
rect 3060 52736 3068 52800
rect 3132 52736 3148 52800
rect 3212 52736 3228 52800
rect 3292 52736 3308 52800
rect 3372 52736 3380 52800
rect 3060 51712 3380 52736
rect 3060 51648 3068 51712
rect 3132 51648 3148 51712
rect 3212 51648 3228 51712
rect 3292 51648 3308 51712
rect 3372 51648 3380 51712
rect 3060 50624 3380 51648
rect 3060 50560 3068 50624
rect 3132 50560 3148 50624
rect 3212 50560 3228 50624
rect 3292 50560 3308 50624
rect 3372 50560 3380 50624
rect 795 49740 861 49741
rect 795 49676 796 49740
rect 860 49676 861 49740
rect 795 49675 861 49676
rect 798 49469 858 49675
rect 3060 49536 3380 50560
rect 3060 49472 3068 49536
rect 3132 49472 3148 49536
rect 3212 49472 3228 49536
rect 3292 49472 3308 49536
rect 3372 49472 3380 49536
rect 795 49468 861 49469
rect 795 49404 796 49468
rect 860 49404 861 49468
rect 795 49403 861 49404
rect 795 49332 861 49333
rect 795 49268 796 49332
rect 860 49268 861 49332
rect 795 49267 861 49268
rect 798 49061 858 49267
rect 795 49060 861 49061
rect 795 48996 796 49060
rect 860 48996 861 49060
rect 795 48995 861 48996
rect 3060 48448 3380 49472
rect 3060 48384 3068 48448
rect 3132 48384 3148 48448
rect 3212 48384 3228 48448
rect 3292 48384 3308 48448
rect 3372 48384 3380 48448
rect 795 47972 861 47973
rect 795 47908 796 47972
rect 860 47908 861 47972
rect 795 47907 861 47908
rect 798 47701 858 47907
rect 795 47700 861 47701
rect 795 47636 796 47700
rect 860 47636 861 47700
rect 795 47635 861 47636
rect -416 35458 -374 35694
rect -138 35458 -96 35694
rect -416 934 -96 35458
rect 3060 47360 3380 48384
rect 3060 47296 3068 47360
rect 3132 47296 3148 47360
rect 3212 47296 3228 47360
rect 3292 47296 3308 47360
rect 3372 47296 3380 47360
rect 3060 46272 3380 47296
rect 3060 46208 3068 46272
rect 3132 46208 3148 46272
rect 3212 46208 3228 46272
rect 3292 46208 3308 46272
rect 3372 46208 3380 46272
rect 3060 45184 3380 46208
rect 3060 45120 3068 45184
rect 3132 45120 3148 45184
rect 3212 45120 3228 45184
rect 3292 45120 3308 45184
rect 3372 45120 3380 45184
rect 3060 44096 3380 45120
rect 3060 44032 3068 44096
rect 3132 44032 3148 44096
rect 3212 44032 3228 44096
rect 3292 44032 3308 44096
rect 3372 44032 3380 44096
rect 3060 43008 3380 44032
rect 3060 42944 3068 43008
rect 3132 42944 3148 43008
rect 3212 42944 3228 43008
rect 3292 42944 3308 43008
rect 3372 42944 3380 43008
rect 3060 41920 3380 42944
rect 3060 41856 3068 41920
rect 3132 41856 3148 41920
rect 3212 41856 3228 41920
rect 3292 41856 3308 41920
rect 3372 41856 3380 41920
rect 3060 40832 3380 41856
rect 3060 40768 3068 40832
rect 3132 40768 3148 40832
rect 3212 40768 3228 40832
rect 3292 40768 3308 40832
rect 3372 40768 3380 40832
rect 3060 39744 3380 40768
rect 3060 39680 3068 39744
rect 3132 39680 3148 39744
rect 3212 39680 3228 39744
rect 3292 39680 3308 39744
rect 3372 39680 3380 39744
rect 3060 38656 3380 39680
rect 3060 38592 3068 38656
rect 3132 38592 3148 38656
rect 3212 38592 3228 38656
rect 3292 38592 3308 38656
rect 3372 38592 3380 38656
rect 3060 37568 3380 38592
rect 3060 37504 3068 37568
rect 3132 37504 3148 37568
rect 3212 37504 3228 37568
rect 3292 37504 3308 37568
rect 3372 37504 3380 37568
rect 3060 36480 3380 37504
rect 3060 36416 3068 36480
rect 3132 36416 3148 36480
rect 3212 36416 3228 36480
rect 3292 36416 3308 36480
rect 3372 36416 3380 36480
rect 3060 35694 3380 36416
rect 3060 35458 3102 35694
rect 3338 35458 3380 35694
rect 3060 35392 3380 35458
rect 3060 35328 3068 35392
rect 3132 35328 3148 35392
rect 3212 35328 3228 35392
rect 3292 35328 3308 35392
rect 3372 35328 3380 35392
rect 3060 34304 3380 35328
rect 3060 34240 3068 34304
rect 3132 34240 3148 34304
rect 3212 34240 3228 34304
rect 3292 34240 3308 34304
rect 3372 34240 3380 34304
rect 3060 33216 3380 34240
rect 3060 33152 3068 33216
rect 3132 33152 3148 33216
rect 3212 33152 3228 33216
rect 3292 33152 3308 33216
rect 3372 33152 3380 33216
rect 3060 32128 3380 33152
rect 3060 32064 3068 32128
rect 3132 32064 3148 32128
rect 3212 32064 3228 32128
rect 3292 32064 3308 32128
rect 3372 32064 3380 32128
rect 3060 31040 3380 32064
rect 3060 30976 3068 31040
rect 3132 30976 3148 31040
rect 3212 30976 3228 31040
rect 3292 30976 3308 31040
rect 3372 30976 3380 31040
rect 3060 29952 3380 30976
rect 3060 29888 3068 29952
rect 3132 29888 3148 29952
rect 3212 29888 3228 29952
rect 3292 29888 3308 29952
rect 3372 29888 3380 29952
rect 3060 28864 3380 29888
rect 3060 28800 3068 28864
rect 3132 28800 3148 28864
rect 3212 28800 3228 28864
rect 3292 28800 3308 28864
rect 3372 28800 3380 28864
rect 3060 27776 3380 28800
rect 3060 27712 3068 27776
rect 3132 27712 3148 27776
rect 3212 27712 3228 27776
rect 3292 27712 3308 27776
rect 3372 27712 3380 27776
rect 3060 26688 3380 27712
rect 3060 26624 3068 26688
rect 3132 26624 3148 26688
rect 3212 26624 3228 26688
rect 3292 26624 3308 26688
rect 3372 26624 3380 26688
rect 3060 25600 3380 26624
rect 3060 25536 3068 25600
rect 3132 25536 3148 25600
rect 3212 25536 3228 25600
rect 3292 25536 3308 25600
rect 3372 25536 3380 25600
rect 3060 24512 3380 25536
rect 3060 24448 3068 24512
rect 3132 24448 3148 24512
rect 3212 24448 3228 24512
rect 3292 24448 3308 24512
rect 3372 24448 3380 24512
rect 3060 23424 3380 24448
rect 3060 23360 3068 23424
rect 3132 23360 3148 23424
rect 3212 23360 3228 23424
rect 3292 23360 3308 23424
rect 3372 23360 3380 23424
rect 3060 22336 3380 23360
rect 3060 22272 3068 22336
rect 3132 22272 3148 22336
rect 3212 22272 3228 22336
rect 3292 22272 3308 22336
rect 3372 22272 3380 22336
rect 3060 21248 3380 22272
rect 3060 21184 3068 21248
rect 3132 21184 3148 21248
rect 3212 21184 3228 21248
rect 3292 21184 3308 21248
rect 3372 21184 3380 21248
rect 3060 20160 3380 21184
rect 3060 20096 3068 20160
rect 3132 20096 3148 20160
rect 3212 20096 3228 20160
rect 3292 20096 3308 20160
rect 3372 20096 3380 20160
rect 3060 19072 3380 20096
rect 3060 19008 3068 19072
rect 3132 19008 3148 19072
rect 3212 19008 3228 19072
rect 3292 19008 3308 19072
rect 3372 19008 3380 19072
rect 3060 17984 3380 19008
rect 3060 17920 3068 17984
rect 3132 17920 3148 17984
rect 3212 17920 3228 17984
rect 3292 17920 3308 17984
rect 3372 17920 3380 17984
rect 3060 16896 3380 17920
rect 3060 16832 3068 16896
rect 3132 16832 3148 16896
rect 3212 16832 3228 16896
rect 3292 16832 3308 16896
rect 3372 16832 3380 16896
rect 3060 15808 3380 16832
rect 3060 15744 3068 15808
rect 3132 15744 3148 15808
rect 3212 15744 3228 15808
rect 3292 15744 3308 15808
rect 3372 15744 3380 15808
rect 3060 14720 3380 15744
rect 3060 14656 3068 14720
rect 3132 14656 3148 14720
rect 3212 14656 3228 14720
rect 3292 14656 3308 14720
rect 3372 14656 3380 14720
rect 3060 13632 3380 14656
rect 3060 13568 3068 13632
rect 3132 13568 3148 13632
rect 3212 13568 3228 13632
rect 3292 13568 3308 13632
rect 3372 13568 3380 13632
rect 3060 12544 3380 13568
rect 3060 12480 3068 12544
rect 3132 12480 3148 12544
rect 3212 12480 3228 12544
rect 3292 12480 3308 12544
rect 3372 12480 3380 12544
rect 3060 11456 3380 12480
rect 3060 11392 3068 11456
rect 3132 11392 3148 11456
rect 3212 11392 3228 11456
rect 3292 11392 3308 11456
rect 3372 11392 3380 11456
rect 3060 10368 3380 11392
rect 3060 10304 3068 10368
rect 3132 10304 3148 10368
rect 3212 10304 3228 10368
rect 3292 10304 3308 10368
rect 3372 10304 3380 10368
rect 3060 9280 3380 10304
rect 3060 9216 3068 9280
rect 3132 9216 3148 9280
rect 3212 9216 3228 9280
rect 3292 9216 3308 9280
rect 3372 9216 3380 9280
rect 3060 8192 3380 9216
rect 3060 8128 3068 8192
rect 3132 8128 3148 8192
rect 3212 8128 3228 8192
rect 3292 8128 3308 8192
rect 3372 8128 3380 8192
rect 3060 7104 3380 8128
rect 3060 7040 3068 7104
rect 3132 7040 3148 7104
rect 3212 7040 3228 7104
rect 3292 7040 3308 7104
rect 3372 7040 3380 7104
rect 3060 6016 3380 7040
rect 3060 5952 3068 6016
rect 3132 5952 3148 6016
rect 3212 5952 3228 6016
rect 3292 5952 3308 6016
rect 3372 5952 3380 6016
rect 3060 5392 3380 5952
rect 3796 91424 4116 91984
rect 3796 91360 3804 91424
rect 3868 91360 3884 91424
rect 3948 91360 3964 91424
rect 4028 91360 4044 91424
rect 4108 91360 4116 91424
rect 3796 90336 4116 91360
rect 3796 90272 3804 90336
rect 3868 90272 3884 90336
rect 3948 90272 3964 90336
rect 4028 90272 4044 90336
rect 4108 90272 4116 90336
rect 3796 89248 4116 90272
rect 3796 89184 3804 89248
rect 3868 89184 3884 89248
rect 3948 89184 3964 89248
rect 4028 89184 4044 89248
rect 4108 89184 4116 89248
rect 3796 88160 4116 89184
rect 3796 88096 3804 88160
rect 3868 88096 3884 88160
rect 3948 88096 3964 88160
rect 4028 88096 4044 88160
rect 4108 88096 4116 88160
rect 3796 87072 4116 88096
rect 8526 87957 8586 95235
rect 36944 95232 37264 96986
rect 36944 95168 36952 95232
rect 37016 95168 37032 95232
rect 37096 95168 37112 95232
rect 37176 95168 37192 95232
rect 37256 95168 37264 95232
rect 36944 94144 37264 95168
rect 36944 94080 36952 94144
rect 37016 94080 37032 94144
rect 37096 94080 37112 94144
rect 37176 94080 37192 94144
rect 37256 94080 37264 94144
rect 36944 93056 37264 94080
rect 36944 92992 36952 93056
rect 37016 92992 37032 93056
rect 37096 92992 37112 93056
rect 37176 92992 37192 93056
rect 37256 92992 37264 93056
rect 36944 91968 37264 92992
rect 36944 91904 36952 91968
rect 37016 91904 37032 91968
rect 37096 91904 37112 91968
rect 37176 91904 37192 91968
rect 37256 91904 37264 91968
rect 36944 90377 37264 91904
rect 37604 97882 37924 97924
rect 37604 97646 37646 97882
rect 37882 97646 37924 97882
rect 37604 95776 37924 97646
rect 37604 95712 37612 95776
rect 37676 95712 37692 95776
rect 37756 95712 37772 95776
rect 37836 95712 37852 95776
rect 37916 95712 37924 95776
rect 37604 94688 37924 95712
rect 37604 94624 37612 94688
rect 37676 94624 37692 94688
rect 37756 94624 37772 94688
rect 37836 94624 37852 94688
rect 37916 94624 37924 94688
rect 37604 93600 37924 94624
rect 37604 93536 37612 93600
rect 37676 93536 37692 93600
rect 37756 93536 37772 93600
rect 37836 93536 37852 93600
rect 37916 93536 37924 93600
rect 37604 92512 37924 93536
rect 72944 97222 73264 97924
rect 72944 96986 72986 97222
rect 73222 96986 73264 97222
rect 72944 95232 73264 96986
rect 72944 95168 72952 95232
rect 73016 95168 73032 95232
rect 73096 95168 73112 95232
rect 73176 95168 73192 95232
rect 73256 95168 73264 95232
rect 72944 94144 73264 95168
rect 72944 94080 72952 94144
rect 73016 94080 73032 94144
rect 73096 94080 73112 94144
rect 73176 94080 73192 94144
rect 73256 94080 73264 94144
rect 72944 93056 73264 94080
rect 72944 92992 72952 93056
rect 73016 92992 73032 93056
rect 73096 92992 73112 93056
rect 73176 92992 73192 93056
rect 73256 92992 73264 93056
rect 48083 92852 48149 92853
rect 48083 92788 48084 92852
rect 48148 92788 48149 92852
rect 48083 92787 48149 92788
rect 47531 92716 47597 92717
rect 47531 92652 47532 92716
rect 47596 92652 47597 92716
rect 47531 92651 47597 92652
rect 37604 92448 37612 92512
rect 37676 92448 37692 92512
rect 37756 92448 37772 92512
rect 37836 92448 37852 92512
rect 37916 92448 37924 92512
rect 37604 91424 37924 92448
rect 37604 91360 37612 91424
rect 37676 91360 37692 91424
rect 37756 91360 37772 91424
rect 37836 91360 37852 91424
rect 37916 91360 37924 91424
rect 37604 90377 37924 91360
rect 8523 87956 8589 87957
rect 8523 87892 8524 87956
rect 8588 87892 8589 87956
rect 8523 87891 8589 87892
rect 3796 87008 3804 87072
rect 3868 87008 3884 87072
rect 3948 87008 3964 87072
rect 4028 87008 4044 87072
rect 4108 87008 4116 87072
rect 3796 85984 4116 87008
rect 9604 86118 9646 86354
rect 9882 86118 9924 86354
rect 45604 86118 45646 86354
rect 45882 86118 45924 86354
rect 3796 85920 3804 85984
rect 3868 85920 3884 85984
rect 3948 85920 3964 85984
rect 4028 85920 4044 85984
rect 4108 85920 4116 85984
rect 3796 84896 4116 85920
rect 8944 85458 8986 85694
rect 9222 85458 9264 85694
rect 44944 85458 44986 85694
rect 45222 85458 45264 85694
rect 3796 84832 3804 84896
rect 3868 84832 3884 84896
rect 3948 84832 3964 84896
rect 4028 84832 4044 84896
rect 4108 84832 4116 84896
rect 3796 83808 4116 84832
rect 3796 83744 3804 83808
rect 3868 83744 3884 83808
rect 3948 83744 3964 83808
rect 4028 83744 4044 83808
rect 4108 83744 4116 83808
rect 3796 82720 4116 83744
rect 3796 82656 3804 82720
rect 3868 82656 3884 82720
rect 3948 82656 3964 82720
rect 4028 82656 4044 82720
rect 4108 82656 4116 82720
rect 3796 81632 4116 82656
rect 3796 81568 3804 81632
rect 3868 81568 3884 81632
rect 3948 81568 3964 81632
rect 4028 81568 4044 81632
rect 4108 81568 4116 81632
rect 3796 80544 4116 81568
rect 3796 80480 3804 80544
rect 3868 80480 3884 80544
rect 3948 80480 3964 80544
rect 4028 80480 4044 80544
rect 4108 80480 4116 80544
rect 3796 79456 4116 80480
rect 3796 79392 3804 79456
rect 3868 79392 3884 79456
rect 3948 79392 3964 79456
rect 4028 79392 4044 79456
rect 4108 79392 4116 79456
rect 3796 78368 4116 79392
rect 3796 78304 3804 78368
rect 3868 78304 3884 78368
rect 3948 78304 3964 78368
rect 4028 78304 4044 78368
rect 4108 78304 4116 78368
rect 3796 77280 4116 78304
rect 3796 77216 3804 77280
rect 3868 77216 3884 77280
rect 3948 77216 3964 77280
rect 4028 77216 4044 77280
rect 4108 77216 4116 77280
rect 3796 76192 4116 77216
rect 3796 76128 3804 76192
rect 3868 76128 3884 76192
rect 3948 76128 3964 76192
rect 4028 76128 4044 76192
rect 4108 76128 4116 76192
rect 3796 75104 4116 76128
rect 3796 75040 3804 75104
rect 3868 75040 3884 75104
rect 3948 75040 3964 75104
rect 4028 75040 4044 75104
rect 4108 75040 4116 75104
rect 3796 74016 4116 75040
rect 3796 73952 3804 74016
rect 3868 73952 3884 74016
rect 3948 73952 3964 74016
rect 4028 73952 4044 74016
rect 4108 73952 4116 74016
rect 3796 72928 4116 73952
rect 3796 72864 3804 72928
rect 3868 72864 3884 72928
rect 3948 72864 3964 72928
rect 4028 72864 4044 72928
rect 4108 72864 4116 72928
rect 3796 71840 4116 72864
rect 3796 71776 3804 71840
rect 3868 71776 3884 71840
rect 3948 71776 3964 71840
rect 4028 71776 4044 71840
rect 4108 71776 4116 71840
rect 3796 70752 4116 71776
rect 3796 70688 3804 70752
rect 3868 70688 3884 70752
rect 3948 70688 3964 70752
rect 4028 70688 4044 70752
rect 4108 70688 4116 70752
rect 3796 69754 4116 70688
rect 3796 69664 3838 69754
rect 4074 69664 4116 69754
rect 3796 69600 3804 69664
rect 4108 69600 4116 69664
rect 3796 69518 3838 69600
rect 4074 69518 4116 69600
rect 9604 69518 9646 69754
rect 9882 69518 9924 69754
rect 45604 69518 45646 69754
rect 45882 69518 45924 69754
rect 3796 68576 4116 69518
rect 8944 68858 8986 69094
rect 9222 68858 9264 69094
rect 44944 68858 44986 69094
rect 45222 68858 45264 69094
rect 3796 68512 3804 68576
rect 3868 68512 3884 68576
rect 3948 68512 3964 68576
rect 4028 68512 4044 68576
rect 4108 68512 4116 68576
rect 3796 67488 4116 68512
rect 5579 67692 5645 67693
rect 5579 67628 5580 67692
rect 5644 67628 5645 67692
rect 5579 67627 5645 67628
rect 3796 67424 3804 67488
rect 3868 67424 3884 67488
rect 3948 67424 3964 67488
rect 4028 67424 4044 67488
rect 4108 67424 4116 67488
rect 3796 66400 4116 67424
rect 3796 66336 3804 66400
rect 3868 66336 3884 66400
rect 3948 66336 3964 66400
rect 4028 66336 4044 66400
rect 4108 66336 4116 66400
rect 3796 65312 4116 66336
rect 3796 65248 3804 65312
rect 3868 65248 3884 65312
rect 3948 65248 3964 65312
rect 4028 65248 4044 65312
rect 4108 65248 4116 65312
rect 3796 64224 4116 65248
rect 3796 64160 3804 64224
rect 3868 64160 3884 64224
rect 3948 64160 3964 64224
rect 4028 64160 4044 64224
rect 4108 64160 4116 64224
rect 3796 63136 4116 64160
rect 3796 63072 3804 63136
rect 3868 63072 3884 63136
rect 3948 63072 3964 63136
rect 4028 63072 4044 63136
rect 4108 63072 4116 63136
rect 3796 62048 4116 63072
rect 3796 61984 3804 62048
rect 3868 61984 3884 62048
rect 3948 61984 3964 62048
rect 4028 61984 4044 62048
rect 4108 61984 4116 62048
rect 3796 60960 4116 61984
rect 3796 60896 3804 60960
rect 3868 60896 3884 60960
rect 3948 60896 3964 60960
rect 4028 60896 4044 60960
rect 4108 60896 4116 60960
rect 3796 59872 4116 60896
rect 3796 59808 3804 59872
rect 3868 59808 3884 59872
rect 3948 59808 3964 59872
rect 4028 59808 4044 59872
rect 4108 59808 4116 59872
rect 3796 58784 4116 59808
rect 3796 58720 3804 58784
rect 3868 58720 3884 58784
rect 3948 58720 3964 58784
rect 4028 58720 4044 58784
rect 4108 58720 4116 58784
rect 3796 57696 4116 58720
rect 3796 57632 3804 57696
rect 3868 57632 3884 57696
rect 3948 57632 3964 57696
rect 4028 57632 4044 57696
rect 4108 57632 4116 57696
rect 3796 56608 4116 57632
rect 3796 56544 3804 56608
rect 3868 56544 3884 56608
rect 3948 56544 3964 56608
rect 4028 56544 4044 56608
rect 4108 56544 4116 56608
rect 3796 55520 4116 56544
rect 3796 55456 3804 55520
rect 3868 55456 3884 55520
rect 3948 55456 3964 55520
rect 4028 55456 4044 55520
rect 4108 55456 4116 55520
rect 3796 54432 4116 55456
rect 3796 54368 3804 54432
rect 3868 54368 3884 54432
rect 3948 54368 3964 54432
rect 4028 54368 4044 54432
rect 4108 54368 4116 54432
rect 3796 53344 4116 54368
rect 3796 53280 3804 53344
rect 3868 53280 3884 53344
rect 3948 53280 3964 53344
rect 4028 53280 4044 53344
rect 4108 53280 4116 53344
rect 3796 52256 4116 53280
rect 3796 52192 3804 52256
rect 3868 52192 3884 52256
rect 3948 52192 3964 52256
rect 4028 52192 4044 52256
rect 4108 52192 4116 52256
rect 3796 51168 4116 52192
rect 3796 51104 3804 51168
rect 3868 51104 3884 51168
rect 3948 51104 3964 51168
rect 4028 51104 4044 51168
rect 4108 51104 4116 51168
rect 3796 50080 4116 51104
rect 5582 50693 5642 67627
rect 5763 64972 5829 64973
rect 5763 64908 5764 64972
rect 5828 64908 5829 64972
rect 5763 64907 5829 64908
rect 5766 50829 5826 64907
rect 5947 62252 6013 62253
rect 5947 62188 5948 62252
rect 6012 62188 6013 62252
rect 5947 62187 6013 62188
rect 5763 50828 5829 50829
rect 5763 50764 5764 50828
rect 5828 50764 5829 50828
rect 5763 50763 5829 50764
rect 5579 50692 5645 50693
rect 5579 50628 5580 50692
rect 5644 50628 5645 50692
rect 5579 50627 5645 50628
rect 3796 50016 3804 50080
rect 3868 50016 3884 50080
rect 3948 50016 3964 50080
rect 4028 50016 4044 50080
rect 4108 50016 4116 50080
rect 3796 48992 4116 50016
rect 5950 49469 6010 62187
rect 9604 52718 9646 52954
rect 9882 52718 9924 52954
rect 45604 52718 45646 52954
rect 45882 52718 45924 52954
rect 8944 52058 8986 52294
rect 9222 52058 9264 52294
rect 44944 52058 44986 52294
rect 45222 52058 45264 52294
rect 5947 49468 6013 49469
rect 5947 49404 5948 49468
rect 6012 49404 6013 49468
rect 5947 49403 6013 49404
rect 3796 48928 3804 48992
rect 3868 48928 3884 48992
rect 3948 48928 3964 48992
rect 4028 48928 4044 48992
rect 4108 48928 4116 48992
rect 3796 47904 4116 48928
rect 47534 48925 47594 92651
rect 47715 88364 47781 88365
rect 47715 88300 47716 88364
rect 47780 88300 47781 88364
rect 47715 88299 47781 88300
rect 47718 50285 47778 88299
rect 47715 50284 47781 50285
rect 47715 50220 47716 50284
rect 47780 50220 47781 50284
rect 47715 50219 47781 50220
rect 48086 49197 48146 92787
rect 72944 91968 73264 92992
rect 72944 91904 72952 91968
rect 73016 91904 73032 91968
rect 73096 91904 73112 91968
rect 73176 91904 73192 91968
rect 73256 91904 73264 91968
rect 72944 90377 73264 91904
rect 73604 97882 73924 97924
rect 73604 97646 73646 97882
rect 73882 97646 73924 97882
rect 73604 95776 73924 97646
rect 90732 97882 91052 97924
rect 90732 97646 90774 97882
rect 91010 97646 91052 97882
rect 73604 95712 73612 95776
rect 73676 95712 73692 95776
rect 73756 95712 73772 95776
rect 73836 95712 73852 95776
rect 73916 95712 73924 95776
rect 73604 94688 73924 95712
rect 73604 94624 73612 94688
rect 73676 94624 73692 94688
rect 73756 94624 73772 94688
rect 73836 94624 73852 94688
rect 73916 94624 73924 94688
rect 73604 93600 73924 94624
rect 73604 93536 73612 93600
rect 73676 93536 73692 93600
rect 73756 93536 73772 93600
rect 73836 93536 73852 93600
rect 73916 93536 73924 93600
rect 73604 92512 73924 93536
rect 90072 97222 90392 97264
rect 90072 96986 90114 97222
rect 90350 96986 90392 97222
rect 89115 92716 89181 92717
rect 89115 92652 89116 92716
rect 89180 92652 89181 92716
rect 89115 92651 89181 92652
rect 86539 92580 86605 92581
rect 86539 92516 86540 92580
rect 86604 92516 86605 92580
rect 86539 92515 86605 92516
rect 87091 92580 87157 92581
rect 87091 92516 87092 92580
rect 87156 92516 87157 92580
rect 87091 92515 87157 92516
rect 73604 92448 73612 92512
rect 73676 92448 73692 92512
rect 73756 92448 73772 92512
rect 73836 92448 73852 92512
rect 73916 92448 73924 92512
rect 73604 91424 73924 92448
rect 73604 91360 73612 91424
rect 73676 91360 73692 91424
rect 73756 91360 73772 91424
rect 73836 91360 73852 91424
rect 73916 91360 73924 91424
rect 73604 90377 73924 91360
rect 86355 91356 86421 91357
rect 86355 91292 86356 91356
rect 86420 91292 86421 91356
rect 86355 91291 86421 91292
rect 49604 86118 49646 86354
rect 49882 86118 49924 86354
rect 85604 86118 85646 86354
rect 85882 86118 85924 86354
rect 48944 85458 48986 85694
rect 49222 85458 49264 85694
rect 84944 85458 84986 85694
rect 85222 85458 85264 85694
rect 86358 77077 86418 91291
rect 86542 87277 86602 92515
rect 86907 91628 86973 91629
rect 86907 91564 86908 91628
rect 86972 91564 86973 91628
rect 86907 91563 86973 91564
rect 86723 91220 86789 91221
rect 86723 91156 86724 91220
rect 86788 91156 86789 91220
rect 86723 91155 86789 91156
rect 86539 87276 86605 87277
rect 86539 87212 86540 87276
rect 86604 87212 86605 87276
rect 86539 87211 86605 87212
rect 86726 87005 86786 91155
rect 86910 87141 86970 91563
rect 86907 87140 86973 87141
rect 86907 87076 86908 87140
rect 86972 87076 86973 87140
rect 86907 87075 86973 87076
rect 86723 87004 86789 87005
rect 86723 86940 86724 87004
rect 86788 86940 86789 87004
rect 86723 86939 86789 86940
rect 86907 85916 86973 85917
rect 86907 85852 86908 85916
rect 86972 85852 86973 85916
rect 86907 85851 86973 85852
rect 86355 77076 86421 77077
rect 86355 77012 86356 77076
rect 86420 77012 86421 77076
rect 86355 77011 86421 77012
rect 49604 69518 49646 69754
rect 49882 69518 49924 69754
rect 85604 69518 85646 69754
rect 85882 69518 85924 69754
rect 48944 68858 48986 69094
rect 49222 68858 49264 69094
rect 84944 68858 84986 69094
rect 85222 68858 85264 69094
rect 86355 66196 86421 66197
rect 86355 66132 86356 66196
rect 86420 66132 86421 66196
rect 86355 66131 86421 66132
rect 49604 52718 49646 52954
rect 49882 52718 49924 52954
rect 85604 52718 85646 52954
rect 85882 52718 85924 52954
rect 48944 52058 48986 52294
rect 49222 52058 49264 52294
rect 84944 52058 84986 52294
rect 85222 52058 85264 52294
rect 85251 50692 85317 50693
rect 85251 50628 85252 50692
rect 85316 50628 85317 50692
rect 85251 50627 85317 50628
rect 85254 50149 85314 50627
rect 86358 50557 86418 66131
rect 86539 63476 86605 63477
rect 86539 63412 86540 63476
rect 86604 63412 86605 63476
rect 86539 63411 86605 63412
rect 86355 50556 86421 50557
rect 86355 50492 86356 50556
rect 86420 50492 86421 50556
rect 86355 50491 86421 50492
rect 85251 50148 85317 50149
rect 85251 50084 85252 50148
rect 85316 50084 85317 50148
rect 85251 50083 85317 50084
rect 48083 49196 48149 49197
rect 48083 49132 48084 49196
rect 48148 49132 48149 49196
rect 48083 49131 48149 49132
rect 86542 48925 86602 63411
rect 86910 60757 86970 85851
rect 86907 60756 86973 60757
rect 86907 60692 86908 60756
rect 86972 60692 86973 60756
rect 86907 60691 86973 60692
rect 87094 60750 87154 92515
rect 88379 89860 88445 89861
rect 88379 89796 88380 89860
rect 88444 89796 88445 89860
rect 88379 89795 88445 89796
rect 87275 88500 87341 88501
rect 87275 88436 87276 88500
rect 87340 88436 87341 88500
rect 87275 88435 87341 88436
rect 87278 64837 87338 88435
rect 88382 67557 88442 89795
rect 89118 74357 89178 92651
rect 89299 92172 89365 92173
rect 89299 92108 89300 92172
rect 89364 92108 89365 92172
rect 89299 92107 89365 92108
rect 89115 74356 89181 74357
rect 89115 74292 89116 74356
rect 89180 74292 89181 74356
rect 89115 74291 89181 74292
rect 89302 73130 89362 92107
rect 89164 73070 89362 73130
rect 89164 72861 89224 73070
rect 89161 72860 89227 72861
rect 89161 72796 89162 72860
rect 89226 72796 89227 72860
rect 89161 72795 89227 72796
rect 90072 69094 90392 96986
rect 90072 68858 90114 69094
rect 90350 68858 90392 69094
rect 88379 67556 88445 67557
rect 88379 67492 88380 67556
rect 88444 67492 88445 67556
rect 88379 67491 88445 67492
rect 87275 64836 87341 64837
rect 87275 64772 87276 64836
rect 87340 64772 87341 64836
rect 87275 64771 87341 64772
rect 87094 60690 87522 60750
rect 87462 59397 87522 60690
rect 87091 59396 87157 59397
rect 87091 59332 87092 59396
rect 87156 59332 87157 59396
rect 87091 59331 87157 59332
rect 87459 59396 87525 59397
rect 87459 59332 87460 59396
rect 87524 59332 87525 59396
rect 87459 59331 87525 59332
rect 86907 55316 86973 55317
rect 86907 55252 86908 55316
rect 86972 55252 86973 55316
rect 86907 55251 86973 55252
rect 86910 49197 86970 55251
rect 87094 49605 87154 59331
rect 87091 49604 87157 49605
rect 87091 49540 87092 49604
rect 87156 49540 87157 49604
rect 87091 49539 87157 49540
rect 86907 49196 86973 49197
rect 86907 49132 86908 49196
rect 86972 49132 86973 49196
rect 86907 49131 86973 49132
rect 47531 48924 47597 48925
rect 47531 48860 47532 48924
rect 47596 48860 47597 48924
rect 47531 48859 47597 48860
rect 86539 48924 86605 48925
rect 86539 48860 86540 48924
rect 86604 48860 86605 48924
rect 86539 48859 86605 48860
rect 48083 48380 48149 48381
rect 48083 48316 48084 48380
rect 48148 48316 48149 48380
rect 48083 48315 48149 48316
rect 87643 48380 87709 48381
rect 87643 48316 87644 48380
rect 87708 48316 87709 48380
rect 87643 48315 87709 48316
rect 47715 48108 47781 48109
rect 47715 48044 47716 48108
rect 47780 48044 47781 48108
rect 47715 48043 47781 48044
rect 3796 47840 3804 47904
rect 3868 47840 3884 47904
rect 3948 47840 3964 47904
rect 4028 47840 4044 47904
rect 4108 47840 4116 47904
rect 3796 46816 4116 47840
rect 5211 47020 5277 47021
rect 5211 46956 5212 47020
rect 5276 46956 5277 47020
rect 5211 46955 5277 46956
rect 3796 46752 3804 46816
rect 3868 46752 3884 46816
rect 3948 46752 3964 46816
rect 4028 46752 4044 46816
rect 4108 46752 4116 46816
rect 3796 45728 4116 46752
rect 3796 45664 3804 45728
rect 3868 45664 3884 45728
rect 3948 45664 3964 45728
rect 4028 45664 4044 45728
rect 4108 45664 4116 45728
rect 3796 44640 4116 45664
rect 3796 44576 3804 44640
rect 3868 44576 3884 44640
rect 3948 44576 3964 44640
rect 4028 44576 4044 44640
rect 4108 44576 4116 44640
rect 3796 43552 4116 44576
rect 3796 43488 3804 43552
rect 3868 43488 3884 43552
rect 3948 43488 3964 43552
rect 4028 43488 4044 43552
rect 4108 43488 4116 43552
rect 3796 42464 4116 43488
rect 3796 42400 3804 42464
rect 3868 42400 3884 42464
rect 3948 42400 3964 42464
rect 4028 42400 4044 42464
rect 4108 42400 4116 42464
rect 3796 41376 4116 42400
rect 3796 41312 3804 41376
rect 3868 41312 3884 41376
rect 3948 41312 3964 41376
rect 4028 41312 4044 41376
rect 4108 41312 4116 41376
rect 3796 40288 4116 41312
rect 3796 40224 3804 40288
rect 3868 40224 3884 40288
rect 3948 40224 3964 40288
rect 4028 40224 4044 40288
rect 4108 40224 4116 40288
rect 3796 39200 4116 40224
rect 3796 39136 3804 39200
rect 3868 39136 3884 39200
rect 3948 39136 3964 39200
rect 4028 39136 4044 39200
rect 4108 39136 4116 39200
rect 3796 38112 4116 39136
rect 3796 38048 3804 38112
rect 3868 38048 3884 38112
rect 3948 38048 3964 38112
rect 4028 38048 4044 38112
rect 4108 38048 4116 38112
rect 3796 37024 4116 38048
rect 3796 36960 3804 37024
rect 3868 36960 3884 37024
rect 3948 36960 3964 37024
rect 4028 36960 4044 37024
rect 4108 36960 4116 37024
rect 3796 36354 4116 36960
rect 3796 36118 3838 36354
rect 4074 36118 4116 36354
rect 3796 35936 4116 36118
rect 3796 35872 3804 35936
rect 3868 35872 3884 35936
rect 3948 35872 3964 35936
rect 4028 35872 4044 35936
rect 4108 35872 4116 35936
rect 3796 34848 4116 35872
rect 3796 34784 3804 34848
rect 3868 34784 3884 34848
rect 3948 34784 3964 34848
rect 4028 34784 4044 34848
rect 4108 34784 4116 34848
rect 3796 33760 4116 34784
rect 3796 33696 3804 33760
rect 3868 33696 3884 33760
rect 3948 33696 3964 33760
rect 4028 33696 4044 33760
rect 4108 33696 4116 33760
rect 3796 32672 4116 33696
rect 3796 32608 3804 32672
rect 3868 32608 3884 32672
rect 3948 32608 3964 32672
rect 4028 32608 4044 32672
rect 4108 32608 4116 32672
rect 3796 31584 4116 32608
rect 3796 31520 3804 31584
rect 3868 31520 3884 31584
rect 3948 31520 3964 31584
rect 4028 31520 4044 31584
rect 4108 31520 4116 31584
rect 3796 30496 4116 31520
rect 3796 30432 3804 30496
rect 3868 30432 3884 30496
rect 3948 30432 3964 30496
rect 4028 30432 4044 30496
rect 4108 30432 4116 30496
rect 3796 29408 4116 30432
rect 3796 29344 3804 29408
rect 3868 29344 3884 29408
rect 3948 29344 3964 29408
rect 4028 29344 4044 29408
rect 4108 29344 4116 29408
rect 3796 28320 4116 29344
rect 3796 28256 3804 28320
rect 3868 28256 3884 28320
rect 3948 28256 3964 28320
rect 4028 28256 4044 28320
rect 4108 28256 4116 28320
rect 3796 27232 4116 28256
rect 3796 27168 3804 27232
rect 3868 27168 3884 27232
rect 3948 27168 3964 27232
rect 4028 27168 4044 27232
rect 4108 27168 4116 27232
rect 3796 26144 4116 27168
rect 5214 27165 5274 46955
rect 9604 44118 9646 44354
rect 9882 44118 9924 44354
rect 45604 44118 45646 44354
rect 45882 44118 45924 44354
rect 8944 43458 8986 43694
rect 9222 43458 9264 43694
rect 44944 43458 44986 43694
rect 45222 43458 45264 43694
rect 9604 36118 9646 36354
rect 9882 36118 9924 36354
rect 45604 36118 45646 36354
rect 45882 36118 45924 36354
rect 8944 35458 8986 35694
rect 9222 35458 9264 35694
rect 44944 35458 44986 35694
rect 45222 35458 45264 35694
rect 5211 27164 5277 27165
rect 5211 27100 5212 27164
rect 5276 27100 5277 27164
rect 5211 27099 5277 27100
rect 3796 26080 3804 26144
rect 3868 26080 3884 26144
rect 3948 26080 3964 26144
rect 4028 26080 4044 26144
rect 4108 26080 4116 26144
rect 3796 25056 4116 26080
rect 3796 24992 3804 25056
rect 3868 24992 3884 25056
rect 3948 24992 3964 25056
rect 4028 24992 4044 25056
rect 4108 24992 4116 25056
rect 3796 23968 4116 24992
rect 3796 23904 3804 23968
rect 3868 23904 3884 23968
rect 3948 23904 3964 23968
rect 4028 23904 4044 23968
rect 4108 23904 4116 23968
rect 3796 22880 4116 23904
rect 3796 22816 3804 22880
rect 3868 22816 3884 22880
rect 3948 22816 3964 22880
rect 4028 22816 4044 22880
rect 4108 22816 4116 22880
rect 3796 21792 4116 22816
rect 3796 21728 3804 21792
rect 3868 21728 3884 21792
rect 3948 21728 3964 21792
rect 4028 21728 4044 21792
rect 4108 21728 4116 21792
rect 3796 20704 4116 21728
rect 3796 20640 3804 20704
rect 3868 20640 3884 20704
rect 3948 20640 3964 20704
rect 4028 20640 4044 20704
rect 4108 20640 4116 20704
rect 3796 19616 4116 20640
rect 3796 19552 3804 19616
rect 3868 19552 3884 19616
rect 3948 19552 3964 19616
rect 4028 19552 4044 19616
rect 4108 19552 4116 19616
rect 3796 18528 4116 19552
rect 3796 18464 3804 18528
rect 3868 18464 3884 18528
rect 3948 18464 3964 18528
rect 4028 18464 4044 18528
rect 4108 18464 4116 18528
rect 3796 17440 4116 18464
rect 3796 17376 3804 17440
rect 3868 17376 3884 17440
rect 3948 17376 3964 17440
rect 4028 17376 4044 17440
rect 4108 17376 4116 17440
rect 3796 16352 4116 17376
rect 3796 16288 3804 16352
rect 3868 16288 3884 16352
rect 3948 16288 3964 16352
rect 4028 16288 4044 16352
rect 4108 16288 4116 16352
rect 3796 15264 4116 16288
rect 3796 15200 3804 15264
rect 3868 15200 3884 15264
rect 3948 15200 3964 15264
rect 4028 15200 4044 15264
rect 4108 15200 4116 15264
rect 3796 14176 4116 15200
rect 3796 14112 3804 14176
rect 3868 14112 3884 14176
rect 3948 14112 3964 14176
rect 4028 14112 4044 14176
rect 4108 14112 4116 14176
rect 3796 13088 4116 14112
rect 3796 13024 3804 13088
rect 3868 13024 3884 13088
rect 3948 13024 3964 13088
rect 4028 13024 4044 13088
rect 4108 13024 4116 13088
rect 3796 12000 4116 13024
rect 3796 11936 3804 12000
rect 3868 11936 3884 12000
rect 3948 11936 3964 12000
rect 4028 11936 4044 12000
rect 4108 11936 4116 12000
rect 3796 10912 4116 11936
rect 3796 10848 3804 10912
rect 3868 10848 3884 10912
rect 3948 10848 3964 10912
rect 4028 10848 4044 10912
rect 4108 10848 4116 10912
rect 3796 9824 4116 10848
rect 9604 10718 9646 10954
rect 9882 10718 9924 10954
rect 45604 10718 45646 10954
rect 45882 10718 45924 10954
rect 8944 10058 8986 10294
rect 9222 10058 9264 10294
rect 44944 10058 44986 10294
rect 45222 10058 45264 10294
rect 3796 9760 3804 9824
rect 3868 9760 3884 9824
rect 3948 9760 3964 9824
rect 4028 9760 4044 9824
rect 4108 9760 4116 9824
rect 3796 8736 4116 9760
rect 3796 8672 3804 8736
rect 3868 8672 3884 8736
rect 3948 8672 3964 8736
rect 4028 8672 4044 8736
rect 4108 8672 4116 8736
rect 3796 7648 4116 8672
rect 3796 7584 3804 7648
rect 3868 7584 3884 7648
rect 3948 7584 3964 7648
rect 4028 7584 4044 7648
rect 4108 7584 4116 7648
rect 3796 6560 4116 7584
rect 3796 6496 3804 6560
rect 3868 6496 3884 6560
rect 3948 6496 3964 6560
rect 4028 6496 4044 6560
rect 4108 6496 4116 6560
rect 3796 5472 4116 6496
rect 3796 5408 3804 5472
rect 3868 5408 3884 5472
rect 3948 5408 3964 5472
rect 4028 5408 4044 5472
rect 4108 5408 4116 5472
rect 3796 5392 4116 5408
rect -416 698 -374 934
rect -138 698 -96 934
rect -416 656 -96 698
rect 36944 4928 37264 8559
rect 36944 4864 36952 4928
rect 37016 4864 37032 4928
rect 37096 4864 37112 4928
rect 37176 4864 37192 4928
rect 37256 4864 37264 4928
rect 36944 3840 37264 4864
rect 36944 3776 36952 3840
rect 37016 3776 37032 3840
rect 37096 3776 37112 3840
rect 37176 3776 37192 3840
rect 37256 3776 37264 3840
rect 36944 2752 37264 3776
rect 36944 2688 36952 2752
rect 37016 2688 37032 2752
rect 37096 2688 37112 2752
rect 37176 2688 37192 2752
rect 37256 2688 37264 2752
rect 36944 934 37264 2688
rect 36944 698 36986 934
rect 37222 698 37264 934
rect -1076 38 -1034 274
rect -798 38 -756 274
rect -1076 -4 -756 38
rect 36944 -4 37264 698
rect 37604 5472 37924 8559
rect 47718 5813 47778 48043
rect 47899 47836 47965 47837
rect 47899 47772 47900 47836
rect 47964 47772 47965 47836
rect 47899 47771 47965 47772
rect 47715 5812 47781 5813
rect 47715 5748 47716 5812
rect 47780 5748 47781 5812
rect 47715 5747 47781 5748
rect 37604 5408 37612 5472
rect 37676 5408 37692 5472
rect 37756 5408 37772 5472
rect 37836 5408 37852 5472
rect 37916 5408 37924 5472
rect 37604 4384 37924 5408
rect 47902 4589 47962 47771
rect 48086 5677 48146 48315
rect 48267 48108 48333 48109
rect 48267 48044 48268 48108
rect 48332 48044 48333 48108
rect 48267 48043 48333 48044
rect 48270 47701 48330 48043
rect 48267 47700 48333 47701
rect 48267 47636 48268 47700
rect 48332 47636 48333 47700
rect 48267 47635 48333 47636
rect 87275 47564 87341 47565
rect 87275 47500 87276 47564
rect 87340 47500 87341 47564
rect 87275 47499 87341 47500
rect 87091 47156 87157 47157
rect 87091 47092 87092 47156
rect 87156 47092 87157 47156
rect 87091 47091 87157 47092
rect 49604 44118 49646 44354
rect 49882 44118 49924 44354
rect 85604 44118 85646 44354
rect 85882 44118 85924 44354
rect 48944 43458 48986 43694
rect 49222 43458 49264 43694
rect 84944 43458 84986 43694
rect 85222 43458 85264 43694
rect 87094 40490 87154 47091
rect 87278 40765 87338 47499
rect 87275 40764 87341 40765
rect 87275 40700 87276 40764
rect 87340 40700 87341 40764
rect 87275 40699 87341 40700
rect 87275 40492 87341 40493
rect 87275 40490 87276 40492
rect 87094 40430 87276 40490
rect 87275 40428 87276 40430
rect 87340 40428 87341 40492
rect 87275 40427 87341 40428
rect 49604 36118 49646 36354
rect 49882 36118 49924 36354
rect 85604 36118 85646 36354
rect 85882 36118 85924 36354
rect 48944 35458 48986 35694
rect 49222 35458 49264 35694
rect 84944 35458 84986 35694
rect 85222 35458 85264 35694
rect 86907 33692 86973 33693
rect 86907 33628 86908 33692
rect 86972 33628 86973 33692
rect 86907 33627 86973 33628
rect 86355 22812 86421 22813
rect 86355 22748 86356 22812
rect 86420 22748 86421 22812
rect 86355 22747 86421 22748
rect 86358 13701 86418 22747
rect 86355 13700 86421 13701
rect 86355 13636 86356 13700
rect 86420 13636 86421 13700
rect 86355 13635 86421 13636
rect 86539 12612 86605 12613
rect 86539 12548 86540 12612
rect 86604 12548 86605 12612
rect 86539 12547 86605 12548
rect 49604 10718 49646 10954
rect 49882 10718 49924 10954
rect 85604 10718 85646 10954
rect 85882 10718 85924 10954
rect 48944 10058 48986 10294
rect 49222 10058 49264 10294
rect 84944 10058 84986 10294
rect 85222 10058 85264 10294
rect 72944 6016 73264 8559
rect 72944 5952 72952 6016
rect 73016 5952 73032 6016
rect 73096 5952 73112 6016
rect 73176 5952 73192 6016
rect 73256 5952 73264 6016
rect 48083 5676 48149 5677
rect 48083 5612 48084 5676
rect 48148 5612 48149 5676
rect 48083 5611 48149 5612
rect 72944 4928 73264 5952
rect 72944 4864 72952 4928
rect 73016 4864 73032 4928
rect 73096 4864 73112 4928
rect 73176 4864 73192 4928
rect 73256 4864 73264 4928
rect 47899 4588 47965 4589
rect 47899 4524 47900 4588
rect 47964 4524 47965 4588
rect 47899 4523 47965 4524
rect 37604 4320 37612 4384
rect 37676 4320 37692 4384
rect 37756 4320 37772 4384
rect 37836 4320 37852 4384
rect 37916 4320 37924 4384
rect 37604 3296 37924 4320
rect 37604 3232 37612 3296
rect 37676 3232 37692 3296
rect 37756 3232 37772 3296
rect 37836 3232 37852 3296
rect 37916 3232 37924 3296
rect 37604 2208 37924 3232
rect 37604 2144 37612 2208
rect 37676 2144 37692 2208
rect 37756 2144 37772 2208
rect 37836 2144 37852 2208
rect 37916 2144 37924 2208
rect 37604 274 37924 2144
rect 37604 38 37646 274
rect 37882 38 37924 274
rect 37604 -4 37924 38
rect 72944 3840 73264 4864
rect 72944 3776 72952 3840
rect 73016 3776 73032 3840
rect 73096 3776 73112 3840
rect 73176 3776 73192 3840
rect 73256 3776 73264 3840
rect 72944 2752 73264 3776
rect 72944 2688 72952 2752
rect 73016 2688 73032 2752
rect 73096 2688 73112 2752
rect 73176 2688 73192 2752
rect 73256 2688 73264 2752
rect 72944 934 73264 2688
rect 72944 698 72986 934
rect 73222 698 73264 934
rect 72944 -4 73264 698
rect 73604 5472 73924 8559
rect 73604 5408 73612 5472
rect 73676 5408 73692 5472
rect 73756 5408 73772 5472
rect 73836 5408 73852 5472
rect 73916 5408 73924 5472
rect 73604 4384 73924 5408
rect 86542 5405 86602 12547
rect 86910 8261 86970 33627
rect 87091 32332 87157 32333
rect 87091 32268 87092 32332
rect 87156 32268 87157 32332
rect 87091 32267 87157 32268
rect 86907 8260 86973 8261
rect 86907 8196 86908 8260
rect 86972 8196 86973 8260
rect 86907 8195 86973 8196
rect 87094 7989 87154 32267
rect 87091 7988 87157 7989
rect 87091 7924 87092 7988
rect 87156 7924 87157 7988
rect 87091 7923 87157 7924
rect 86539 5404 86605 5405
rect 86539 5340 86540 5404
rect 86604 5340 86605 5404
rect 86539 5339 86605 5340
rect 87278 4861 87338 40427
rect 87646 30973 87706 48315
rect 90072 35694 90392 68858
rect 90072 35458 90114 35694
rect 90350 35458 90392 35694
rect 87643 30972 87709 30973
rect 87643 30908 87644 30972
rect 87708 30908 87709 30972
rect 87643 30907 87709 30908
rect 88747 24172 88813 24173
rect 88747 24108 88748 24172
rect 88812 24108 88813 24172
rect 88747 24107 88813 24108
rect 88563 23900 88629 23901
rect 88563 23836 88564 23900
rect 88628 23836 88629 23900
rect 88563 23835 88629 23836
rect 88195 21452 88261 21453
rect 88195 21388 88196 21452
rect 88260 21388 88261 21452
rect 88195 21387 88261 21388
rect 88198 5541 88258 21387
rect 88379 11116 88445 11117
rect 88379 11052 88380 11116
rect 88444 11052 88445 11116
rect 88379 11051 88445 11052
rect 88382 8397 88442 11051
rect 88379 8396 88445 8397
rect 88379 8332 88380 8396
rect 88444 8332 88445 8396
rect 88379 8331 88445 8332
rect 88566 5949 88626 23835
rect 88750 9621 88810 24107
rect 88747 9620 88813 9621
rect 88747 9556 88748 9620
rect 88812 9556 88813 9620
rect 88747 9555 88813 9556
rect 88563 5948 88629 5949
rect 88563 5884 88564 5948
rect 88628 5884 88629 5948
rect 88563 5883 88629 5884
rect 88195 5540 88261 5541
rect 88195 5476 88196 5540
rect 88260 5476 88261 5540
rect 88195 5475 88261 5476
rect 87275 4860 87341 4861
rect 87275 4796 87276 4860
rect 87340 4796 87341 4860
rect 87275 4795 87341 4796
rect 73604 4320 73612 4384
rect 73676 4320 73692 4384
rect 73756 4320 73772 4384
rect 73836 4320 73852 4384
rect 73916 4320 73924 4384
rect 73604 3296 73924 4320
rect 73604 3232 73612 3296
rect 73676 3232 73692 3296
rect 73756 3232 73772 3296
rect 73836 3232 73852 3296
rect 73916 3232 73924 3296
rect 73604 2208 73924 3232
rect 73604 2144 73612 2208
rect 73676 2144 73692 2208
rect 73756 2144 73772 2208
rect 73836 2144 73852 2208
rect 73916 2144 73924 2208
rect 73604 274 73924 2144
rect 90072 934 90392 35458
rect 90072 698 90114 934
rect 90350 698 90392 934
rect 90072 656 90392 698
rect 90732 69754 91052 97646
rect 90732 69518 90774 69754
rect 91010 69518 91052 69754
rect 90732 36354 91052 69518
rect 90732 36118 90774 36354
rect 91010 36118 91052 36354
rect 73604 38 73646 274
rect 73882 38 73924 274
rect 73604 -4 73924 38
rect 90732 274 91052 36118
rect 90732 38 90774 274
rect 91010 38 91052 274
rect 90732 -4 91052 38
<< via4 >>
rect -1034 97646 -798 97882
rect -1034 69518 -798 69754
rect -1034 36118 -798 36354
rect -374 96986 -138 97222
rect 36986 96986 37222 97222
rect -374 68858 -138 69094
rect 3102 69056 3132 69094
rect 3132 69056 3148 69094
rect 3148 69056 3212 69094
rect 3212 69056 3228 69094
rect 3228 69056 3292 69094
rect 3292 69056 3308 69094
rect 3308 69056 3338 69094
rect 3102 68858 3338 69056
rect -374 35458 -138 35694
rect 3102 35458 3338 35694
rect 37646 97646 37882 97882
rect 72986 96986 73222 97222
rect 9646 86118 9882 86354
rect 45646 86118 45882 86354
rect 8986 85458 9222 85694
rect 44986 85458 45222 85694
rect 3838 69664 4074 69754
rect 3838 69600 3868 69664
rect 3868 69600 3884 69664
rect 3884 69600 3948 69664
rect 3948 69600 3964 69664
rect 3964 69600 4028 69664
rect 4028 69600 4044 69664
rect 4044 69600 4074 69664
rect 3838 69518 4074 69600
rect 9646 69518 9882 69754
rect 45646 69518 45882 69754
rect 8986 68858 9222 69094
rect 44986 68858 45222 69094
rect 9646 52718 9882 52954
rect 45646 52718 45882 52954
rect 8986 52058 9222 52294
rect 44986 52058 45222 52294
rect 73646 97646 73882 97882
rect 90774 97646 91010 97882
rect 90114 96986 90350 97222
rect 49646 86118 49882 86354
rect 85646 86118 85882 86354
rect 48986 85458 49222 85694
rect 84986 85458 85222 85694
rect 49646 69518 49882 69754
rect 85646 69518 85882 69754
rect 48986 68858 49222 69094
rect 84986 68858 85222 69094
rect 49646 52718 49882 52954
rect 85646 52718 85882 52954
rect 48986 52058 49222 52294
rect 84986 52058 85222 52294
rect 90114 68858 90350 69094
rect 3838 36118 4074 36354
rect 9646 44118 9882 44354
rect 45646 44118 45882 44354
rect 8986 43458 9222 43694
rect 44986 43458 45222 43694
rect 9646 36118 9882 36354
rect 45646 36118 45882 36354
rect 8986 35458 9222 35694
rect 44986 35458 45222 35694
rect 9646 10718 9882 10954
rect 45646 10718 45882 10954
rect 8986 10058 9222 10294
rect 44986 10058 45222 10294
rect -374 698 -138 934
rect 36986 698 37222 934
rect -1034 38 -798 274
rect 49646 44118 49882 44354
rect 85646 44118 85882 44354
rect 48986 43458 49222 43694
rect 84986 43458 85222 43694
rect 49646 36118 49882 36354
rect 85646 36118 85882 36354
rect 48986 35458 49222 35694
rect 84986 35458 85222 35694
rect 49646 10718 49882 10954
rect 85646 10718 85882 10954
rect 48986 10058 49222 10294
rect 84986 10058 85222 10294
rect 37646 38 37882 274
rect 72986 698 73222 934
rect 90114 35458 90350 35694
rect 90114 698 90350 934
rect 90774 69518 91010 69754
rect 90774 36118 91010 36354
rect 73646 38 73882 274
rect 90774 38 91010 274
<< metal5 >>
rect -1076 97882 91052 97924
rect -1076 97646 -1034 97882
rect -798 97646 37646 97882
rect 37882 97646 73646 97882
rect 73882 97646 90774 97882
rect 91010 97646 91052 97882
rect -1076 97604 91052 97646
rect -416 97222 90392 97264
rect -416 96986 -374 97222
rect -138 96986 36986 97222
rect 37222 96986 72986 97222
rect 73222 96986 90114 97222
rect 90350 96986 90392 97222
rect -416 96944 90392 96986
rect 9622 86354 9906 86396
rect 9622 86118 9646 86354
rect 9882 86118 9906 86354
rect 9622 86076 9906 86118
rect 45622 86354 45906 86396
rect 45622 86118 45646 86354
rect 45882 86118 45906 86354
rect 45622 86076 45906 86118
rect 49622 86354 49906 86396
rect 49622 86118 49646 86354
rect 49882 86118 49906 86354
rect 49622 86076 49906 86118
rect 85622 86354 85906 86396
rect 85622 86118 85646 86354
rect 85882 86118 85906 86354
rect 85622 86076 85906 86118
rect 8962 85694 9246 85736
rect 8962 85458 8986 85694
rect 9222 85458 9246 85694
rect 8962 85416 9246 85458
rect 44962 85694 45246 85736
rect 44962 85458 44986 85694
rect 45222 85458 45246 85694
rect 44962 85416 45246 85458
rect 48962 85694 49246 85736
rect 48962 85458 48986 85694
rect 49222 85458 49246 85694
rect 48962 85416 49246 85458
rect 84962 85694 85246 85736
rect 84962 85458 84986 85694
rect 85222 85458 85246 85694
rect 84962 85416 85246 85458
rect -1076 69754 91052 69796
rect -1076 69518 -1034 69754
rect -798 69518 3838 69754
rect 4074 69518 9646 69754
rect 9882 69518 45646 69754
rect 45882 69518 49646 69754
rect 49882 69518 85646 69754
rect 85882 69518 90774 69754
rect 91010 69518 91052 69754
rect -1076 69476 91052 69518
rect -1076 69094 91052 69136
rect -1076 68858 -374 69094
rect -138 68858 3102 69094
rect 3338 68858 8986 69094
rect 9222 68858 44986 69094
rect 45222 68858 48986 69094
rect 49222 68858 84986 69094
rect 85222 68858 90114 69094
rect 90350 68858 91052 69094
rect -1076 68816 91052 68858
rect 9622 52954 9906 52996
rect 9622 52718 9646 52954
rect 9882 52718 9906 52954
rect 9622 52676 9906 52718
rect 45622 52954 45906 52996
rect 45622 52718 45646 52954
rect 45882 52718 45906 52954
rect 45622 52676 45906 52718
rect 49622 52954 49906 52996
rect 49622 52718 49646 52954
rect 49882 52718 49906 52954
rect 49622 52676 49906 52718
rect 85622 52954 85906 52996
rect 85622 52718 85646 52954
rect 85882 52718 85906 52954
rect 85622 52676 85906 52718
rect 8962 52294 9246 52336
rect 8962 52058 8986 52294
rect 9222 52058 9246 52294
rect 8962 52016 9246 52058
rect 44962 52294 45246 52336
rect 44962 52058 44986 52294
rect 45222 52058 45246 52294
rect 44962 52016 45246 52058
rect 48962 52294 49246 52336
rect 48962 52058 48986 52294
rect 49222 52058 49246 52294
rect 48962 52016 49246 52058
rect 84962 52294 85246 52336
rect 84962 52058 84986 52294
rect 85222 52058 85246 52294
rect 84962 52016 85246 52058
rect 9622 44354 9906 44396
rect 9622 44118 9646 44354
rect 9882 44118 9906 44354
rect 9622 44076 9906 44118
rect 45622 44354 45906 44396
rect 45622 44118 45646 44354
rect 45882 44118 45906 44354
rect 45622 44076 45906 44118
rect 49622 44354 49906 44396
rect 49622 44118 49646 44354
rect 49882 44118 49906 44354
rect 49622 44076 49906 44118
rect 85622 44354 85906 44396
rect 85622 44118 85646 44354
rect 85882 44118 85906 44354
rect 85622 44076 85906 44118
rect 8962 43694 9246 43736
rect 8962 43458 8986 43694
rect 9222 43458 9246 43694
rect 8962 43416 9246 43458
rect 44962 43694 45246 43736
rect 44962 43458 44986 43694
rect 45222 43458 45246 43694
rect 44962 43416 45246 43458
rect 48962 43694 49246 43736
rect 48962 43458 48986 43694
rect 49222 43458 49246 43694
rect 48962 43416 49246 43458
rect 84962 43694 85246 43736
rect 84962 43458 84986 43694
rect 85222 43458 85246 43694
rect 84962 43416 85246 43458
rect -1076 36354 91052 36396
rect -1076 36118 -1034 36354
rect -798 36118 3838 36354
rect 4074 36118 9646 36354
rect 9882 36118 45646 36354
rect 45882 36118 49646 36354
rect 49882 36118 85646 36354
rect 85882 36118 90774 36354
rect 91010 36118 91052 36354
rect -1076 36076 91052 36118
rect -1076 35694 91052 35736
rect -1076 35458 -374 35694
rect -138 35458 3102 35694
rect 3338 35458 8986 35694
rect 9222 35458 44986 35694
rect 45222 35458 48986 35694
rect 49222 35458 84986 35694
rect 85222 35458 90114 35694
rect 90350 35458 91052 35694
rect -1076 35416 91052 35458
rect 9622 10954 9906 10996
rect 9622 10718 9646 10954
rect 9882 10718 9906 10954
rect 9622 10676 9906 10718
rect 45622 10954 45906 10996
rect 45622 10718 45646 10954
rect 45882 10718 45906 10954
rect 45622 10676 45906 10718
rect 49622 10954 49906 10996
rect 49622 10718 49646 10954
rect 49882 10718 49906 10954
rect 49622 10676 49906 10718
rect 85622 10954 85906 10996
rect 85622 10718 85646 10954
rect 85882 10718 85906 10954
rect 85622 10676 85906 10718
rect 8962 10294 9246 10336
rect 8962 10058 8986 10294
rect 9222 10058 9246 10294
rect 8962 10016 9246 10058
rect 44962 10294 45246 10336
rect 44962 10058 44986 10294
rect 45222 10058 45246 10294
rect 44962 10016 45246 10058
rect 48962 10294 49246 10336
rect 48962 10058 48986 10294
rect 49222 10058 49246 10294
rect 48962 10016 49246 10058
rect 84962 10294 85246 10336
rect 84962 10058 84986 10294
rect 85222 10058 85246 10294
rect 84962 10016 85246 10058
rect -416 934 90392 976
rect -416 698 -374 934
rect -138 698 36986 934
rect 37222 698 72986 934
rect 73222 698 90114 934
rect 90350 698 90392 934
rect -416 656 90392 698
rect -1076 274 91052 316
rect -1076 38 -1034 274
rect -798 38 37646 274
rect 37882 38 73646 274
rect 73882 38 90774 274
rect 91010 38 91052 274
rect -1076 -4 91052 38
use sky130_fd_sc_hd__diode_2  ANTENNA_cell0_clk
timestamp 18001
transform 1 0 5520 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell0_config_data_out
timestamp 18001
transform -1 0 9844 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell0_config_en
timestamp 18001
transform -1 0 5520 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell0_le_clk
timestamp 18001
transform 1 0 10764 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell0_le_en
timestamp 18001
transform 1 0 11868 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell0_le_nrst
timestamp 18001
transform 1 0 12972 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell0_nrst
timestamp 18001
transform -1 0 5336 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell1_CBeast_in[0]
timestamp 18001
transform -1 0 86756 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell1_CBeast_in[1]
timestamp 18001
transform -1 0 86204 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell1_CBeast_in[2]
timestamp 18001
transform -1 0 85652 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell1_CBeast_in[3]
timestamp 18001
transform -1 0 86940 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell1_CBeast_in[4]
timestamp 18001
transform -1 0 86020 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell1_CBeast_in[5]
timestamp 18001
transform -1 0 85468 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell1_CBeast_in[6]
timestamp 18001
transform -1 0 87124 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell1_CBeast_in[7]
timestamp 18001
transform -1 0 85836 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell1_CBeast_in[8]
timestamp 18001
transform -1 0 85284 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell1_CBeast_in[9]
timestamp 18001
transform -1 0 87308 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell1_CBeast_in[10]
timestamp 18001
transform -1 0 85836 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell1_CBeast_in[11]
timestamp 18001
transform -1 0 86572 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell1_CBeast_in[12]
timestamp 18001
transform -1 0 86388 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell1_CBeast_in[13]
timestamp 18001
transform -1 0 86756 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell1_CBeast_out[10]
timestamp 18001
transform -1 0 85100 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell1_CBeast_out[11]
timestamp 18001
transform 1 0 87308 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell1_CBeast_out[12]
timestamp 18001
transform -1 0 84916 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell1_CBeast_out[13]
timestamp 18001
transform -1 0 86572 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell1_clk
timestamp 18001
transform -1 0 50416 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell1_config_data_in
timestamp 18001
transform -1 0 53728 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell1_config_data_out
timestamp 18001
transform -1 0 49864 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell1_config_en
timestamp 18001
transform -1 0 52624 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell1_le_clk
timestamp 18001
transform -1 0 50968 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell1_le_en
timestamp 18001
transform -1 0 52072 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell1_le_nrst
timestamp 18001
transform 1 0 52992 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell1_nrst
timestamp 18001
transform -1 0 51520 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell2_clk
timestamp 18001
transform 1 0 10212 0 1 91392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell2_config_data_in
timestamp 18001
transform -1 0 13708 0 1 91392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell2_config_data_out
timestamp 18001
transform -1 0 5336 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell2_config_en
timestamp 18001
transform 1 0 12420 0 1 91392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell2_le_clk
timestamp 18001
transform -1 0 5704 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell2_le_en
timestamp 18001
transform -1 0 5152 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell2_le_nrst
timestamp 18001
transform -1 0 5520 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell2_nrst
timestamp 18001
transform 1 0 11500 0 1 91392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell3_CBeast_in[0]
timestamp 18001
transform -1 0 86480 0 1 91392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell3_CBeast_in[1]
timestamp 18001
transform -1 0 86756 0 -1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell3_CBeast_in[2]
timestamp 18001
transform -1 0 86112 0 1 91392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell3_CBeast_in[3]
timestamp 18001
transform 1 0 86756 0 -1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell3_CBeast_out[0]
timestamp 18001
transform -1 0 85928 0 1 91392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell3_CBeast_out[1]
timestamp 18001
transform -1 0 86204 0 -1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell3_CBeast_out[2]
timestamp 18001
transform -1 0 85560 0 1 91392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell3_CBeast_out[3]
timestamp 18001
transform -1 0 86940 0 1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell3_CBeast_out[4]
timestamp 18001
transform -1 0 86020 0 -1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell3_CBeast_out[5]
timestamp 18001
transform -1 0 85376 0 1 91392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell3_CBeast_out[6]
timestamp 18001
transform -1 0 87124 0 1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell3_CBeast_out[7]
timestamp 18001
transform -1 0 85836 0 -1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell3_CBeast_out[8]
timestamp 18001
transform -1 0 85192 0 1 91392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell3_CBeast_out[9]
timestamp 18001
transform -1 0 87308 0 1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell3_CBeast_out[10]
timestamp 18001
transform -1 0 86572 0 -1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell3_CBeast_out[11]
timestamp 18001
transform -1 0 86388 0 -1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell3_CBeast_out[12]
timestamp 18001
transform -1 0 85744 0 1 91392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell3_CBeast_out[13]
timestamp 18001
transform -1 0 86756 0 1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell3_clk
timestamp 18001
transform -1 0 50416 0 1 91392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell3_config_data_in
timestamp 18001
transform -1 0 54372 0 1 91392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell3_config_data_out
timestamp 18001
transform -1 0 49864 0 1 91392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell3_config_en
timestamp 18001
transform 1 0 52440 0 -1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell3_le_clk
timestamp 18001
transform -1 0 50968 0 1 91392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell3_le_en
timestamp 18001
transform -1 0 52072 0 -1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell3_le_nrst
timestamp 18001
transform -1 0 53268 0 -1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell3_nrst
timestamp 18001
transform 1 0 50968 0 1 91392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 18001
transform 1 0 32384 0 1 91392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_X
timestamp 18001
transform 1 0 32200 0 1 91392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0__f_clk_A
timestamp 18001
transform 1 0 5336 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0__f_clk_X
timestamp 18001
transform -1 0 5704 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1__f_clk_A
timestamp 18001
transform -1 0 32568 0 -1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1__f_clk_X
timestamp 18001
transform 1 0 32200 0 -1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 18001
transform -1 0 2116 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 18001
transform -1 0 52716 0 1 94656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_X
timestamp 18001
transform 1 0 54188 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 18001
transform -1 0 5244 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_X
timestamp 18001
transform -1 0 5428 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 18001
transform -1 0 5152 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_X
timestamp 18001
transform -1 0 5336 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 18001
transform -1 0 5152 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_X
timestamp 18001
transform -1 0 5336 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 18001
transform -1 0 5152 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_X
timestamp 18001
transform -1 0 5336 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 18001
transform -1 0 5152 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_X
timestamp 18001
transform -1 0 5336 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 18001
transform -1 0 5244 0 -1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_X
timestamp 18001
transform -1 0 5428 0 -1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 18001
transform -1 0 5244 0 -1 71808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_X
timestamp 18001
transform -1 0 5428 0 -1 71808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 18001
transform -1 0 88228 0 -1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_X
timestamp 18001
transform -1 0 88596 0 -1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 18001
transform -1 0 86572 0 1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_X
timestamp 18001
transform -1 0 88596 0 -1 94656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 18001
transform -1 0 5244 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_X
timestamp 18001
transform -1 0 5428 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 18001
transform -1 0 87768 0 -1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 18001
transform -1 0 88136 0 1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 18001
transform -1 0 87492 0 -1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 18001
transform -1 0 88596 0 1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 18001
transform -1 0 87492 0 1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 18001
transform -1 0 88412 0 -1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 18001
transform -1 0 87952 0 1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 18001
transform -1 0 88044 0 -1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 18001
transform -1 0 88412 0 1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 18001
transform -1 0 87676 0 1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 18001
transform -1 0 5244 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_X
timestamp 18001
transform -1 0 5428 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 18001
transform -1 0 5244 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_X
timestamp 18001
transform -1 0 5428 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 18001
transform -1 0 5244 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_X
timestamp 18001
transform -1 0 5428 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 18001
transform -1 0 5244 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_X
timestamp 18001
transform -1 0 5428 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 18001
transform -1 0 5244 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_X
timestamp 18001
transform -1 0 5428 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 18001
transform -1 0 5152 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_X
timestamp 18001
transform -1 0 5336 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 18001
transform -1 0 5244 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_X
timestamp 18001
transform -1 0 5428 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 18001
transform -1 0 5152 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_X
timestamp 18001
transform -1 0 5336 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 18001
transform -1 0 14904 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 18001
transform -1 0 25852 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 18001
transform -1 0 27140 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 18001
transform -1 0 27784 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 18001
transform -1 0 29072 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 18001
transform -1 0 56028 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 18001
transform -1 0 56672 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 18001
transform -1 0 57316 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 18001
transform -1 0 58052 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 18001
transform -1 0 16100 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 18001
transform -1 0 59340 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 18001
transform -1 0 60628 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 18001
transform -1 0 61272 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 18001
transform -1 0 62560 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 18001
transform -1 0 63848 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 18001
transform -1 0 65320 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 18001
transform -1 0 65780 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 18001
transform -1 0 67068 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 18001
transform -1 0 67712 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 18001
transform -1 0 69000 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 18001
transform -1 0 16836 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 18001
transform -1 0 18124 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 18001
transform -1 0 19412 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 18001
transform -1 0 20608 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 18001
transform -1 0 21344 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 18001
transform -1 0 22632 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 18001
transform -1 0 23276 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 18001
transform -1 0 24564 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 18001
transform -1 0 31004 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 18001
transform -1 0 41952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 18001
transform -1 0 42596 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 18001
transform -1 0 43884 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 18001
transform -1 0 45172 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 18001
transform -1 0 70932 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 18001
transform -1 0 71576 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 18001
transform -1 0 72864 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 18001
transform -1 0 74152 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 18001
transform -1 0 31648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 18001
transform -1 0 75440 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 18001
transform -1 0 76084 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 18001
transform -1 0 77372 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 18001
transform -1 0 78660 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 18001
transform -1 0 80132 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 18001
transform -1 0 80592 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 18001
transform -1 0 81880 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 18001
transform -1 0 83168 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input77_A
timestamp 18001
transform -1 0 87676 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input78_A
timestamp 18001
transform 1 0 86204 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 18001
transform -1 0 32936 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 18001
transform -1 0 34224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input81_A
timestamp 18001
transform -1 0 34868 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input82_A
timestamp 18001
transform -1 0 36156 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input83_A
timestamp 18001
transform -1 0 37444 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input84_A
timestamp 18001
transform -1 0 38732 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input85_A
timestamp 18001
transform -1 0 40388 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input86_A
timestamp 18001
transform -1 0 40664 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input87_A
timestamp 18001
transform -1 0 7820 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input88_A
timestamp 18001
transform -1 0 1840 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input89_A
timestamp 18001
transform -1 0 1840 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input90_A
timestamp 18001
transform -1 0 1840 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input91_A
timestamp 18001
transform -1 0 1840 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input92_A
timestamp 18001
transform -1 0 1840 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input93_A
timestamp 18001
transform -1 0 1840 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input94_A
timestamp 18001
transform -1 0 1840 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input95_A
timestamp 18001
transform -1 0 1840 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input96_A
timestamp 18001
transform -1 0 8464 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input97_A
timestamp 18001
transform -1 0 1840 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input98_A
timestamp 18001
transform -1 0 1840 0 1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input99_A
timestamp 18001
transform -1 0 1840 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input100_A
timestamp 18001
transform -1 0 1840 0 -1 62016
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input101_A
timestamp 18001
transform -1 0 1840 0 1 62016
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input102_A
timestamp 18001
transform -1 0 1840 0 1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input103_A
timestamp 18001
transform -1 0 1840 0 -1 65280
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input104_A
timestamp 18001
transform -1 0 1840 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input105_A
timestamp 18001
transform -1 0 1840 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input106_A
timestamp 18001
transform -1 0 1840 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input107_A
timestamp 18001
transform -1 0 1840 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input108_A
timestamp 18001
transform -1 0 1840 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input109_A
timestamp 18001
transform -1 0 1840 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input110_A
timestamp 18001
transform -1 0 1840 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input111_A
timestamp 18001
transform -1 0 1840 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input112_A
timestamp 18001
transform -1 0 1840 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input113_A
timestamp 18001
transform -1 0 1840 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input114_A
timestamp 18001
transform -1 0 1840 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input115_A
timestamp 18001
transform -1 0 11960 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input115_X
timestamp 18001
transform 1 0 11592 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input116_A
timestamp 18001
transform -1 0 12328 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input116_X
timestamp 18001
transform 1 0 13340 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input117_A
timestamp 18001
transform -1 0 13984 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input117_X
timestamp 18001
transform 1 0 15088 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input118_A
timestamp 18001
transform -1 0 50968 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input118_X
timestamp 18001
transform 1 0 52440 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_max_cap232_A
timestamp 18001
transform -1 0 54556 0 1 91392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_max_cap232_X
timestamp 18001
transform -1 0 54740 0 1 91392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_max_cap233_A
timestamp 18001
transform -1 0 52900 0 -1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_max_cap233_X
timestamp 18001
transform -1 0 53084 0 -1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output119_A
timestamp 18001
transform -1 0 4968 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output121_A
timestamp 18001
transform -1 0 87860 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output122_A
timestamp 18001
transform -1 0 88228 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output123_A
timestamp 18001
transform -1 0 5336 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output124_A
timestamp 18001
transform -1 0 5336 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output125_A
timestamp 18001
transform -1 0 5336 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output126_A
timestamp 18001
transform -1 0 5336 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output127_A
timestamp 18001
transform -1 0 5336 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output128_A
timestamp 18001
transform -1 0 5336 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output130_A
timestamp 18001
transform -1 0 5336 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output131_A
timestamp 18001
transform -1 0 5336 0 1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output132_A
timestamp 18001
transform -1 0 5336 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output133_A
timestamp 18001
transform -1 0 5336 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output134_A
timestamp 18001
transform -1 0 5336 0 1 62016
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output135_A
timestamp 18001
transform -1 0 5336 0 1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output136_A
timestamp 18001
transform -1 0 5336 0 -1 65280
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output137_A
timestamp 18001
transform -1 0 5336 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output138_A
timestamp 18001
transform -1 0 5336 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output139_A
timestamp 18001
transform -1 0 5336 0 1 68544
box -38 -48 222 592
use fpgacell  cell0
timestamp 0
transform 1 0 8000 0 1 8000
box 0 0 39000 39000
use fpgacell  cell1
timestamp 0
transform 1 0 48000 0 1 8000
box 0 0 39000 39000
use fpgacell  cell2
timestamp 0
transform 1 0 8000 0 1 50000
box 0 0 39000 39000
use fpgacell  cell3
timestamp 0
transform 1 0 48000 0 1 50000
box 0 0 39000 39000
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 18001
transform -1 0 32016 0 1 91392
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 18001
transform -1 0 5704 0 1 56576
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 18001
transform -1 0 32016 0 -1 92480
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3
timestamp 1636986456
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1636986456
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp 18001
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1636986456
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1636986456
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp 18001
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1636986456
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_69
timestamp 18001
transform 1 0 7452 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76
timestamp 18001
transform 1 0 8096 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 18001
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1636986456
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_97
timestamp 18001
transform 1 0 10028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113
timestamp 18001
transform 1 0 11500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_118
timestamp 18001
transform 1 0 11960 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_135
timestamp 18001
transform 1 0 13524 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_154
timestamp 18001
transform 1 0 15272 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_161
timestamp 18001
transform 1 0 15916 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_169
timestamp 18001
transform 1 0 16652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_177
timestamp 18001
transform 1 0 17388 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_182
timestamp 18001
transform 1 0 17848 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_190
timestamp 18001
transform 1 0 18584 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 18001
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_203
timestamp 18001
transform 1 0 19780 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_211
timestamp 18001
transform 1 0 20516 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_217
timestamp 18001
transform 1 0 21068 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 18001
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 18001
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_231
timestamp 18001
transform 1 0 22356 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_239
timestamp 18001
transform 1 0 23092 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_245
timestamp 18001
transform 1 0 23644 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_253
timestamp 18001
transform 1 0 24380 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_261
timestamp 18001
transform 1 0 25116 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_266
timestamp 18001
transform 1 0 25576 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_274
timestamp 18001
transform 1 0 26312 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 18001
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_287
timestamp 18001
transform 1 0 27508 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_295
timestamp 18001
transform 1 0 28244 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_301
timestamp 18001
transform 1 0 28796 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 18001
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 18001
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_315
timestamp 18001
transform 1 0 30084 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_328
timestamp 18001
transform 1 0 31280 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_335
timestamp 18001
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_337
timestamp 18001
transform 1 0 32108 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_343
timestamp 18001
transform 1 0 32660 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_349
timestamp 18001
transform 1 0 33212 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_357
timestamp 18001
transform 1 0 33948 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 18001
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_370
timestamp 18001
transform 1 0 35144 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_378
timestamp 18001
transform 1 0 35880 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_384
timestamp 18001
transform 1 0 36432 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_398
timestamp 18001
transform 1 0 37720 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_406
timestamp 18001
transform 1 0 38456 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_419
timestamp 18001
transform 1 0 39652 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_427
timestamp 18001
transform 1 0 40388 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_434
timestamp 18001
transform 1 0 41032 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_455
timestamp 18001
transform 1 0 42964 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_469
timestamp 18001
transform 1 0 44252 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_475
timestamp 18001
transform 1 0 44804 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_482
timestamp 1636986456
transform 1 0 45448 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_494
timestamp 18001
transform 1 0 46552 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_502
timestamp 18001
transform 1 0 47288 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_505
timestamp 1636986456
transform 1 0 47564 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_517
timestamp 1636986456
transform 1 0 48668 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_529
timestamp 18001
transform 1 0 49772 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_533
timestamp 1636986456
transform 1 0 50140 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_545
timestamp 1636986456
transform 1 0 51244 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_557
timestamp 18001
transform 1 0 52348 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_561
timestamp 1636986456
transform 1 0 52716 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_573
timestamp 1636986456
transform 1 0 53820 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_585
timestamp 18001
transform 1 0 54924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_589
timestamp 18001
transform 1 0 55292 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_595
timestamp 18001
transform 1 0 55844 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_602
timestamp 18001
transform 1 0 56488 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_610
timestamp 18001
transform 1 0 57224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_617
timestamp 18001
transform 1 0 57868 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_625
timestamp 18001
transform 1 0 58604 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_630
timestamp 18001
transform 1 0 59064 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_638
timestamp 18001
transform 1 0 59800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_645
timestamp 18001
transform 1 0 60444 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_651
timestamp 18001
transform 1 0 60996 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_659
timestamp 18001
transform 1 0 61732 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_665
timestamp 18001
transform 1 0 62284 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_671
timestamp 18001
transform 1 0 62836 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_673
timestamp 18001
transform 1 0 63020 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_679
timestamp 18001
transform 1 0 63572 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_686
timestamp 18001
transform 1 0 64216 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_694
timestamp 18001
transform 1 0 64952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_701
timestamp 18001
transform 1 0 65596 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_709
timestamp 18001
transform 1 0 66332 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_714
timestamp 18001
transform 1 0 66792 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_722
timestamp 18001
transform 1 0 67528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_729
timestamp 18001
transform 1 0 68172 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_735
timestamp 18001
transform 1 0 68724 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_743
timestamp 18001
transform 1 0 69460 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_749
timestamp 18001
transform 1 0 70012 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_755
timestamp 18001
transform 1 0 70564 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_762
timestamp 18001
transform 1 0 71208 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_769
timestamp 18001
transform 1 0 71852 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_777
timestamp 18001
transform 1 0 72588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_783
timestamp 18001
transform 1 0 73140 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_785
timestamp 18001
transform 1 0 73324 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_791
timestamp 18001
transform 1 0 73876 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_797
timestamp 18001
transform 1 0 74428 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_805
timestamp 18001
transform 1 0 75164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_811
timestamp 18001
transform 1 0 75716 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_818
timestamp 18001
transform 1 0 76360 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_826
timestamp 18001
transform 1 0 77096 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_832
timestamp 18001
transform 1 0 77648 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_859
timestamp 18001
transform 1 0 80132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_869
timestamp 18001
transform 1 0 81052 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_875
timestamp 18001
transform 1 0 81604 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_882
timestamp 18001
transform 1 0 82248 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_897
timestamp 1636986456
transform 1 0 83628 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_909
timestamp 1636986456
transform 1 0 84732 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_921
timestamp 18001
transform 1 0 85836 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_925
timestamp 1636986456
transform 1 0 86204 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_937
timestamp 1636986456
transform 1 0 87308 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_949
timestamp 18001
transform 1 0 88412 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1636986456
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1636986456
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1636986456
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1636986456
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 18001
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 18001
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1636986456
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1636986456
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1636986456
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1636986456
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 18001
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 18001
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1636986456
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1636986456
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1636986456
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1636986456
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 18001
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 18001
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1636986456
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1636986456
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1636986456
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1636986456
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 18001
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 18001
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1636986456
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1636986456
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1636986456
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1636986456
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 18001
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 18001
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1636986456
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1636986456
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1636986456
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1636986456
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 18001
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 18001
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1636986456
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1636986456
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1636986456
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1636986456
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 18001
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 18001
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1636986456
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_405
timestamp 1636986456
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_417
timestamp 1636986456
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_429
timestamp 1636986456
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 18001
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 18001
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_449
timestamp 1636986456
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_461
timestamp 1636986456
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_473
timestamp 1636986456
transform 1 0 44620 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_485
timestamp 1636986456
transform 1 0 45724 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_497
timestamp 18001
transform 1 0 46828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 18001
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_505
timestamp 1636986456
transform 1 0 47564 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_517
timestamp 1636986456
transform 1 0 48668 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_529
timestamp 1636986456
transform 1 0 49772 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_541
timestamp 1636986456
transform 1 0 50876 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_553
timestamp 18001
transform 1 0 51980 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_559
timestamp 18001
transform 1 0 52532 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_561
timestamp 1636986456
transform 1 0 52716 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_573
timestamp 1636986456
transform 1 0 53820 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_585
timestamp 1636986456
transform 1 0 54924 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_597
timestamp 1636986456
transform 1 0 56028 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_609
timestamp 18001
transform 1 0 57132 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_615
timestamp 18001
transform 1 0 57684 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_617
timestamp 1636986456
transform 1 0 57868 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_629
timestamp 1636986456
transform 1 0 58972 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_641
timestamp 1636986456
transform 1 0 60076 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_653
timestamp 1636986456
transform 1 0 61180 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_665
timestamp 18001
transform 1 0 62284 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_671
timestamp 18001
transform 1 0 62836 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_673
timestamp 1636986456
transform 1 0 63020 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_685
timestamp 1636986456
transform 1 0 64124 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_697
timestamp 1636986456
transform 1 0 65228 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_709
timestamp 1636986456
transform 1 0 66332 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_721
timestamp 18001
transform 1 0 67436 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_727
timestamp 18001
transform 1 0 67988 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_729
timestamp 1636986456
transform 1 0 68172 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_741
timestamp 1636986456
transform 1 0 69276 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_753
timestamp 1636986456
transform 1 0 70380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_765
timestamp 1636986456
transform 1 0 71484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_777
timestamp 18001
transform 1 0 72588 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_783
timestamp 18001
transform 1 0 73140 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_785
timestamp 1636986456
transform 1 0 73324 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_797
timestamp 1636986456
transform 1 0 74428 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_809
timestamp 1636986456
transform 1 0 75532 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_821
timestamp 1636986456
transform 1 0 76636 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_833
timestamp 18001
transform 1 0 77740 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_839
timestamp 18001
transform 1 0 78292 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_841
timestamp 1636986456
transform 1 0 78476 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_853
timestamp 1636986456
transform 1 0 79580 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_865
timestamp 1636986456
transform 1 0 80684 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_877
timestamp 1636986456
transform 1 0 81788 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_889
timestamp 18001
transform 1 0 82892 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_895
timestamp 18001
transform 1 0 83444 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_897
timestamp 1636986456
transform 1 0 83628 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_909
timestamp 1636986456
transform 1 0 84732 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_921
timestamp 1636986456
transform 1 0 85836 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_933
timestamp 1636986456
transform 1 0 86940 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_945
timestamp 18001
transform 1 0 88044 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1636986456
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1636986456
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 18001
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1636986456
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1636986456
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1636986456
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1636986456
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 18001
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 18001
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1636986456
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1636986456
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1636986456
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1636986456
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 18001
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 18001
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1636986456
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1636986456
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1636986456
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1636986456
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 18001
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 18001
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1636986456
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1636986456
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1636986456
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1636986456
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 18001
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 18001
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1636986456
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1636986456
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1636986456
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1636986456
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 18001
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 18001
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1636986456
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1636986456
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1636986456
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1636986456
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 18001
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 18001
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1636986456
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1636986456
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1636986456
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1636986456
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 18001
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 18001
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1636986456
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1636986456
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 1636986456
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_457
timestamp 1636986456
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 18001
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 18001
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_477
timestamp 1636986456
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_489
timestamp 1636986456
transform 1 0 46092 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_501
timestamp 1636986456
transform 1 0 47196 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_513
timestamp 1636986456
transform 1 0 48300 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_525
timestamp 18001
transform 1 0 49404 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 18001
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_533
timestamp 1636986456
transform 1 0 50140 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_545
timestamp 1636986456
transform 1 0 51244 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_557
timestamp 1636986456
transform 1 0 52348 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_569
timestamp 1636986456
transform 1 0 53452 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_581
timestamp 18001
transform 1 0 54556 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 18001
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_589
timestamp 1636986456
transform 1 0 55292 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_601
timestamp 1636986456
transform 1 0 56396 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_613
timestamp 1636986456
transform 1 0 57500 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_625
timestamp 1636986456
transform 1 0 58604 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_637
timestamp 18001
transform 1 0 59708 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_643
timestamp 18001
transform 1 0 60260 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_645
timestamp 1636986456
transform 1 0 60444 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_657
timestamp 1636986456
transform 1 0 61548 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_669
timestamp 1636986456
transform 1 0 62652 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_681
timestamp 1636986456
transform 1 0 63756 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_693
timestamp 18001
transform 1 0 64860 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_699
timestamp 18001
transform 1 0 65412 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_701
timestamp 1636986456
transform 1 0 65596 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_713
timestamp 1636986456
transform 1 0 66700 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_725
timestamp 1636986456
transform 1 0 67804 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_737
timestamp 1636986456
transform 1 0 68908 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_749
timestamp 18001
transform 1 0 70012 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_755
timestamp 18001
transform 1 0 70564 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_757
timestamp 1636986456
transform 1 0 70748 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_769
timestamp 1636986456
transform 1 0 71852 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_781
timestamp 1636986456
transform 1 0 72956 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_793
timestamp 1636986456
transform 1 0 74060 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_805
timestamp 18001
transform 1 0 75164 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_811
timestamp 18001
transform 1 0 75716 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_813
timestamp 1636986456
transform 1 0 75900 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_825
timestamp 1636986456
transform 1 0 77004 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_837
timestamp 1636986456
transform 1 0 78108 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_849
timestamp 1636986456
transform 1 0 79212 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_861
timestamp 18001
transform 1 0 80316 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_867
timestamp 18001
transform 1 0 80868 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_869
timestamp 1636986456
transform 1 0 81052 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_881
timestamp 1636986456
transform 1 0 82156 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_893
timestamp 1636986456
transform 1 0 83260 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_905
timestamp 1636986456
transform 1 0 84364 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_917
timestamp 18001
transform 1 0 85468 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_923
timestamp 18001
transform 1 0 86020 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_925
timestamp 1636986456
transform 1 0 86204 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_937
timestamp 1636986456
transform 1 0 87308 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_949
timestamp 18001
transform 1 0 88412 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1636986456
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1636986456
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1636986456
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1636986456
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 18001
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 18001
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1636986456
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1636986456
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1636986456
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1636986456
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 18001
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 18001
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1636986456
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1636986456
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1636986456
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1636986456
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 18001
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 18001
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1636986456
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1636986456
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1636986456
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1636986456
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 18001
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 18001
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1636986456
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1636986456
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1636986456
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1636986456
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 18001
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 18001
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1636986456
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1636986456
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1636986456
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1636986456
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 18001
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 18001
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1636986456
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1636986456
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1636986456
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1636986456
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 18001
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 18001
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1636986456
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1636986456
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1636986456
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1636986456
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 18001
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 18001
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1636986456
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1636986456
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1636986456
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1636986456
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 18001
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 18001
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_505
timestamp 1636986456
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_517
timestamp 1636986456
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_529
timestamp 1636986456
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_541
timestamp 1636986456
transform 1 0 50876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_553
timestamp 18001
transform 1 0 51980 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 18001
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_561
timestamp 1636986456
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_573
timestamp 1636986456
transform 1 0 53820 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_585
timestamp 1636986456
transform 1 0 54924 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_597
timestamp 1636986456
transform 1 0 56028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_609
timestamp 18001
transform 1 0 57132 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 18001
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_617
timestamp 1636986456
transform 1 0 57868 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_629
timestamp 1636986456
transform 1 0 58972 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_641
timestamp 1636986456
transform 1 0 60076 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_653
timestamp 1636986456
transform 1 0 61180 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_665
timestamp 18001
transform 1 0 62284 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_671
timestamp 18001
transform 1 0 62836 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_673
timestamp 1636986456
transform 1 0 63020 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_685
timestamp 1636986456
transform 1 0 64124 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_697
timestamp 1636986456
transform 1 0 65228 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_709
timestamp 1636986456
transform 1 0 66332 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_721
timestamp 18001
transform 1 0 67436 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_727
timestamp 18001
transform 1 0 67988 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_729
timestamp 1636986456
transform 1 0 68172 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_741
timestamp 1636986456
transform 1 0 69276 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_753
timestamp 1636986456
transform 1 0 70380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_765
timestamp 1636986456
transform 1 0 71484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_777
timestamp 18001
transform 1 0 72588 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_783
timestamp 18001
transform 1 0 73140 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_785
timestamp 1636986456
transform 1 0 73324 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_797
timestamp 1636986456
transform 1 0 74428 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_809
timestamp 1636986456
transform 1 0 75532 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_821
timestamp 1636986456
transform 1 0 76636 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_833
timestamp 18001
transform 1 0 77740 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_839
timestamp 18001
transform 1 0 78292 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_841
timestamp 1636986456
transform 1 0 78476 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_853
timestamp 1636986456
transform 1 0 79580 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_865
timestamp 1636986456
transform 1 0 80684 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_877
timestamp 1636986456
transform 1 0 81788 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_889
timestamp 18001
transform 1 0 82892 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_895
timestamp 18001
transform 1 0 83444 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_897
timestamp 1636986456
transform 1 0 83628 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_909
timestamp 1636986456
transform 1 0 84732 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_921
timestamp 1636986456
transform 1 0 85836 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_933
timestamp 1636986456
transform 1 0 86940 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_947
timestamp 18001
transform 1 0 88228 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1636986456
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1636986456
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 18001
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1636986456
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1636986456
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1636986456
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1636986456
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 18001
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 18001
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1636986456
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1636986456
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1636986456
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1636986456
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 18001
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 18001
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1636986456
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1636986456
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1636986456
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1636986456
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 18001
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 18001
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1636986456
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1636986456
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1636986456
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1636986456
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 18001
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 18001
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1636986456
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1636986456
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1636986456
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1636986456
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 18001
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 18001
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1636986456
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1636986456
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1636986456
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1636986456
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 18001
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 18001
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1636986456
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1636986456
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1636986456
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1636986456
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 18001
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 18001
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1636986456
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1636986456
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1636986456
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1636986456
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 18001
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 18001
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1636986456
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1636986456
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_501
timestamp 1636986456
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_513
timestamp 1636986456
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_525
timestamp 18001
transform 1 0 49404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 18001
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_533
timestamp 1636986456
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_545
timestamp 1636986456
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_557
timestamp 1636986456
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_569
timestamp 1636986456
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_581
timestamp 18001
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 18001
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_589
timestamp 1636986456
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_601
timestamp 1636986456
transform 1 0 56396 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_613
timestamp 1636986456
transform 1 0 57500 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_625
timestamp 1636986456
transform 1 0 58604 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_637
timestamp 18001
transform 1 0 59708 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_643
timestamp 18001
transform 1 0 60260 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_645
timestamp 1636986456
transform 1 0 60444 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_657
timestamp 1636986456
transform 1 0 61548 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_669
timestamp 1636986456
transform 1 0 62652 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_681
timestamp 1636986456
transform 1 0 63756 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_693
timestamp 18001
transform 1 0 64860 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_699
timestamp 18001
transform 1 0 65412 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_701
timestamp 1636986456
transform 1 0 65596 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_713
timestamp 1636986456
transform 1 0 66700 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_725
timestamp 1636986456
transform 1 0 67804 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_737
timestamp 1636986456
transform 1 0 68908 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_749
timestamp 18001
transform 1 0 70012 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_755
timestamp 18001
transform 1 0 70564 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_757
timestamp 1636986456
transform 1 0 70748 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_769
timestamp 1636986456
transform 1 0 71852 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_781
timestamp 1636986456
transform 1 0 72956 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_793
timestamp 1636986456
transform 1 0 74060 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_805
timestamp 18001
transform 1 0 75164 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_811
timestamp 18001
transform 1 0 75716 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_813
timestamp 1636986456
transform 1 0 75900 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_825
timestamp 1636986456
transform 1 0 77004 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_837
timestamp 1636986456
transform 1 0 78108 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_849
timestamp 1636986456
transform 1 0 79212 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_861
timestamp 18001
transform 1 0 80316 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_867
timestamp 18001
transform 1 0 80868 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_869
timestamp 1636986456
transform 1 0 81052 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_881
timestamp 1636986456
transform 1 0 82156 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_893
timestamp 1636986456
transform 1 0 83260 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_905
timestamp 1636986456
transform 1 0 84364 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_917
timestamp 18001
transform 1 0 85468 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_923
timestamp 18001
transform 1 0 86020 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_925
timestamp 18001
transform 1 0 86204 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1636986456
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1636986456
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1636986456
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1636986456
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 18001
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 18001
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1636986456
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1636986456
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1636986456
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1636986456
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 18001
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 18001
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1636986456
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1636986456
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1636986456
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1636986456
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 18001
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 18001
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1636986456
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1636986456
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1636986456
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1636986456
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 18001
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 18001
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1636986456
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1636986456
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1636986456
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1636986456
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 18001
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 18001
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1636986456
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1636986456
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1636986456
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1636986456
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 18001
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 18001
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1636986456
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1636986456
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1636986456
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1636986456
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 18001
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 18001
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1636986456
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1636986456
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1636986456
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1636986456
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 18001
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 18001
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1636986456
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1636986456
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1636986456
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1636986456
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 18001
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 18001
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1636986456
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_517
timestamp 1636986456
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_529
timestamp 1636986456
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_541
timestamp 1636986456
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 18001
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 18001
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_561
timestamp 1636986456
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_573
timestamp 1636986456
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_585
timestamp 1636986456
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_597
timestamp 1636986456
transform 1 0 56028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_609
timestamp 18001
transform 1 0 57132 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_615
timestamp 18001
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_617
timestamp 1636986456
transform 1 0 57868 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_629
timestamp 1636986456
transform 1 0 58972 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_641
timestamp 1636986456
transform 1 0 60076 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_653
timestamp 1636986456
transform 1 0 61180 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_665
timestamp 18001
transform 1 0 62284 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_671
timestamp 18001
transform 1 0 62836 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_673
timestamp 1636986456
transform 1 0 63020 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_685
timestamp 1636986456
transform 1 0 64124 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_697
timestamp 1636986456
transform 1 0 65228 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_709
timestamp 1636986456
transform 1 0 66332 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_721
timestamp 18001
transform 1 0 67436 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_727
timestamp 18001
transform 1 0 67988 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_729
timestamp 1636986456
transform 1 0 68172 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_741
timestamp 1636986456
transform 1 0 69276 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_753
timestamp 1636986456
transform 1 0 70380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_765
timestamp 1636986456
transform 1 0 71484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_777
timestamp 18001
transform 1 0 72588 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_783
timestamp 18001
transform 1 0 73140 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_785
timestamp 1636986456
transform 1 0 73324 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_797
timestamp 1636986456
transform 1 0 74428 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_809
timestamp 1636986456
transform 1 0 75532 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_821
timestamp 1636986456
transform 1 0 76636 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_833
timestamp 18001
transform 1 0 77740 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_839
timestamp 18001
transform 1 0 78292 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_841
timestamp 1636986456
transform 1 0 78476 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_853
timestamp 1636986456
transform 1 0 79580 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_865
timestamp 1636986456
transform 1 0 80684 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_877
timestamp 1636986456
transform 1 0 81788 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_889
timestamp 18001
transform 1 0 82892 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_895
timestamp 18001
transform 1 0 83444 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_897
timestamp 1636986456
transform 1 0 83628 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_909
timestamp 18001
transform 1 0 84732 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_917
timestamp 18001
transform 1 0 85468 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1636986456
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1636986456
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 18001
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1636986456
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1636986456
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_53
timestamp 18001
transform 1 0 5980 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_57
timestamp 1636986456
transform 1 0 6348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_69
timestamp 1636986456
transform 1 0 7452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_81
timestamp 18001
transform 1 0 8556 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_85
timestamp 18001
transform 1 0 8924 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_95
timestamp 18001
transform 1 0 9844 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_103
timestamp 18001
transform 1 0 10580 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_107
timestamp 18001
transform 1 0 10948 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_111
timestamp 18001
transform 1 0 11316 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_113
timestamp 18001
transform 1 0 11500 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_119
timestamp 18001
transform 1 0 12052 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_127
timestamp 18001
transform 1 0 12788 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_131
timestamp 18001
transform 1 0 13156 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 18001
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1636986456
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1636986456
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_165
timestamp 18001
transform 1 0 16284 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_169
timestamp 1636986456
transform 1 0 16652 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_181
timestamp 1636986456
transform 1 0 17756 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_193
timestamp 18001
transform 1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1636986456
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1636986456
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_221
timestamp 18001
transform 1 0 21436 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_225
timestamp 1636986456
transform 1 0 21804 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_237
timestamp 1636986456
transform 1 0 22908 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_249
timestamp 18001
transform 1 0 24012 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1636986456
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1636986456
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_277
timestamp 18001
transform 1 0 26588 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_281
timestamp 1636986456
transform 1 0 26956 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_293
timestamp 1636986456
transform 1 0 28060 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_305
timestamp 18001
transform 1 0 29164 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1636986456
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1636986456
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_333
timestamp 18001
transform 1 0 31740 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_337
timestamp 1636986456
transform 1 0 32108 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_349
timestamp 1636986456
transform 1 0 33212 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_361
timestamp 18001
transform 1 0 34316 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1636986456
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1636986456
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_389
timestamp 18001
transform 1 0 36892 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_393
timestamp 1636986456
transform 1 0 37260 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_405
timestamp 1636986456
transform 1 0 38364 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_417
timestamp 18001
transform 1 0 39468 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1636986456
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1636986456
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_445
timestamp 18001
transform 1 0 42044 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_449
timestamp 1636986456
transform 1 0 42412 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_461
timestamp 1636986456
transform 1 0 43516 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_473
timestamp 18001
transform 1 0 44620 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1636986456
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1636986456
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_501
timestamp 18001
transform 1 0 47196 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_505
timestamp 1636986456
transform 1 0 47564 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_517
timestamp 18001
transform 1 0 48668 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_525
timestamp 18001
transform 1 0 49404 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_530
timestamp 18001
transform 1 0 49864 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_533
timestamp 18001
transform 1 0 50140 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_536
timestamp 18001
transform 1 0 50416 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_542
timestamp 18001
transform 1 0 50968 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_548
timestamp 18001
transform 1 0 51520 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_554
timestamp 18001
transform 1 0 52072 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_561
timestamp 18001
transform 1 0 52716 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_566
timestamp 18001
transform 1 0 53176 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_572
timestamp 1636986456
transform 1 0 53728 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_584
timestamp 18001
transform 1 0 54832 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_589
timestamp 1636986456
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_601
timestamp 1636986456
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_613
timestamp 18001
transform 1 0 57500 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_617
timestamp 1636986456
transform 1 0 57868 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_629
timestamp 1636986456
transform 1 0 58972 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_641
timestamp 18001
transform 1 0 60076 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_645
timestamp 1636986456
transform 1 0 60444 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_657
timestamp 1636986456
transform 1 0 61548 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_669
timestamp 18001
transform 1 0 62652 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_673
timestamp 1636986456
transform 1 0 63020 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_685
timestamp 1636986456
transform 1 0 64124 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_697
timestamp 18001
transform 1 0 65228 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_701
timestamp 1636986456
transform 1 0 65596 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_713
timestamp 1636986456
transform 1 0 66700 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_725
timestamp 18001
transform 1 0 67804 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_729
timestamp 1636986456
transform 1 0 68172 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_741
timestamp 1636986456
transform 1 0 69276 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_753
timestamp 18001
transform 1 0 70380 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_757
timestamp 1636986456
transform 1 0 70748 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_769
timestamp 1636986456
transform 1 0 71852 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_781
timestamp 18001
transform 1 0 72956 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_785
timestamp 1636986456
transform 1 0 73324 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_797
timestamp 1636986456
transform 1 0 74428 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_809
timestamp 18001
transform 1 0 75532 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_813
timestamp 1636986456
transform 1 0 75900 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_825
timestamp 1636986456
transform 1 0 77004 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_837
timestamp 18001
transform 1 0 78108 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_841
timestamp 1636986456
transform 1 0 78476 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_853
timestamp 1636986456
transform 1 0 79580 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_865
timestamp 18001
transform 1 0 80684 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_869
timestamp 1636986456
transform 1 0 81052 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_881
timestamp 1636986456
transform 1 0 82156 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_893
timestamp 18001
transform 1 0 83260 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_897
timestamp 1636986456
transform 1 0 83628 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1636986456
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1636986456
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1636986456
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_39
timestamp 18001
transform 1 0 4692 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_47
timestamp 18001
transform 1 0 5428 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1636986456
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1636986456
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 18001
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1636986456
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_41
timestamp 18001
transform 1 0 4876 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_49
timestamp 18001
transform 1 0 5612 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1636986456
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1636986456
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1636986456
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_39
timestamp 18001
transform 1 0 4692 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_47
timestamp 18001
transform 1 0 5428 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1636986456
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1636986456
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 18001
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1636986456
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_41
timestamp 18001
transform 1 0 4876 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_49
timestamp 18001
transform 1 0 5612 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1636986456
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1636986456
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1636986456
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_39
timestamp 18001
transform 1 0 4692 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_47
timestamp 18001
transform 1 0 5428 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1636986456
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1636986456
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 18001
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1636986456
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_41
timestamp 18001
transform 1 0 4876 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_49
timestamp 18001
transform 1 0 5612 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1636986456
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1636986456
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1636986456
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_39
timestamp 18001
transform 1 0 4692 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_47
timestamp 18001
transform 1 0 5428 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1636986456
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1636986456
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 18001
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1636986456
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_41
timestamp 18001
transform 1 0 4876 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_49
timestamp 18001
transform 1 0 5612 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1636986456
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1636986456
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1636986456
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_39
timestamp 18001
transform 1 0 4692 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_47
timestamp 18001
transform 1 0 5428 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1636986456
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1636986456
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 18001
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1636986456
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_41
timestamp 18001
transform 1 0 4876 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_49
timestamp 18001
transform 1 0 5612 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_8
timestamp 1636986456
transform 1 0 1840 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_20
timestamp 1636986456
transform 1 0 2944 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_32
timestamp 1636986456
transform 1 0 4048 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_44
timestamp 18001
transform 1 0 5152 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1636986456
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1636986456
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 18001
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1636986456
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_41
timestamp 18001
transform 1 0 4876 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_49
timestamp 18001
transform 1 0 5612 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1636986456
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1636986456
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1636986456
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_39
timestamp 18001
transform 1 0 4692 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_47
timestamp 18001
transform 1 0 5428 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_8
timestamp 1636986456
transform 1 0 1840 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_20
timestamp 18001
transform 1 0 2944 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1636986456
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_41
timestamp 18001
transform 1 0 4876 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_49
timestamp 18001
transform 1 0 5612 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1636986456
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1636986456
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1636986456
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_39
timestamp 18001
transform 1 0 4692 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_47
timestamp 18001
transform 1 0 5428 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_8
timestamp 1636986456
transform 1 0 1840 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_20
timestamp 18001
transform 1 0 2944 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1636986456
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_41
timestamp 18001
transform 1 0 4876 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_49
timestamp 18001
transform 1 0 5612 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1636986456
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1636986456
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1636986456
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_39
timestamp 18001
transform 1 0 4692 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_47
timestamp 18001
transform 1 0 5428 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1636986456
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1636986456
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 18001
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1636986456
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_41
timestamp 18001
transform 1 0 4876 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_49
timestamp 18001
transform 1 0 5612 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_8
timestamp 1636986456
transform 1 0 1840 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_20
timestamp 1636986456
transform 1 0 2944 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_32
timestamp 1636986456
transform 1 0 4048 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_44
timestamp 18001
transform 1 0 5152 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1636986456
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1636986456
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 18001
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1636986456
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_41
timestamp 18001
transform 1 0 4876 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_49
timestamp 18001
transform 1 0 5612 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_8
timestamp 1636986456
transform 1 0 1840 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_20
timestamp 1636986456
transform 1 0 2944 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_32
timestamp 1636986456
transform 1 0 4048 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_44
timestamp 18001
transform 1 0 5152 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1636986456
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1636986456
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 18001
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1636986456
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_41
timestamp 18001
transform 1 0 4876 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_49
timestamp 18001
transform 1 0 5612 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1636986456
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1636986456
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1636986456
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_39
timestamp 18001
transform 1 0 4692 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_47
timestamp 18001
transform 1 0 5428 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_8
timestamp 1636986456
transform 1 0 1840 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_20
timestamp 18001
transform 1 0 2944 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1636986456
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_41
timestamp 18001
transform 1 0 4876 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_49
timestamp 18001
transform 1 0 5612 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1636986456
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1636986456
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1636986456
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_39
timestamp 18001
transform 1 0 4692 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_47
timestamp 18001
transform 1 0 5428 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_8
timestamp 1636986456
transform 1 0 1840 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_20
timestamp 18001
transform 1 0 2944 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1636986456
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_41
timestamp 18001
transform 1 0 4876 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_49
timestamp 18001
transform 1 0 5612 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1636986456
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1636986456
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1636986456
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_39
timestamp 18001
transform 1 0 4692 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_47
timestamp 18001
transform 1 0 5428 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1636986456
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1636986456
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 18001
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1636986456
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_41
timestamp 18001
transform 1 0 4876 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_49
timestamp 18001
transform 1 0 5612 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_8
timestamp 1636986456
transform 1 0 1840 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_20
timestamp 1636986456
transform 1 0 2944 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_32
timestamp 1636986456
transform 1 0 4048 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_44
timestamp 18001
transform 1 0 5152 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1636986456
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1636986456
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 18001
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1636986456
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_41
timestamp 18001
transform 1 0 4876 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_49
timestamp 18001
transform 1 0 5612 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_8
timestamp 1636986456
transform 1 0 1840 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_20
timestamp 1636986456
transform 1 0 2944 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_32
timestamp 1636986456
transform 1 0 4048 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_44
timestamp 18001
transform 1 0 5152 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1636986456
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1636986456
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 18001
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1636986456
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_41
timestamp 18001
transform 1 0 4876 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_49
timestamp 18001
transform 1 0 5612 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1636986456
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1636986456
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1636986456
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_39
timestamp 18001
transform 1 0 4692 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_47
timestamp 18001
transform 1 0 5428 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_8
timestamp 1636986456
transform 1 0 1840 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_20
timestamp 18001
transform 1 0 2944 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1636986456
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_41
timestamp 18001
transform 1 0 4876 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_49
timestamp 18001
transform 1 0 5612 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1636986456
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1636986456
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1636986456
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_39
timestamp 18001
transform 1 0 4692 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_47
timestamp 18001
transform 1 0 5428 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_8
timestamp 1636986456
transform 1 0 1840 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_20
timestamp 18001
transform 1 0 2944 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1636986456
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_41
timestamp 18001
transform 1 0 4876 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1636986456
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1636986456
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1636986456
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_39
timestamp 18001
transform 1 0 4692 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_47
timestamp 18001
transform 1 0 5428 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1636986456
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1636986456
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 18001
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1636986456
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_41
timestamp 18001
transform 1 0 4876 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_49
timestamp 18001
transform 1 0 5612 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_8
timestamp 1636986456
transform 1 0 1840 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_20
timestamp 1636986456
transform 1 0 2944 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_32
timestamp 1636986456
transform 1 0 4048 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1636986456
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1636986456
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 18001
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1636986456
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_41
timestamp 18001
transform 1 0 4876 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_49
timestamp 18001
transform 1 0 5612 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_7
timestamp 1636986456
transform 1 0 1748 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_19
timestamp 1636986456
transform 1 0 2852 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_31
timestamp 1636986456
transform 1 0 3956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1636986456
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1636986456
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 18001
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1636986456
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_41
timestamp 18001
transform 1 0 4876 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_49
timestamp 18001
transform 1 0 5612 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1636986456
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1636986456
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1636986456
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_39
timestamp 18001
transform 1 0 4692 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_47
timestamp 18001
transform 1 0 5428 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_7
timestamp 1636986456
transform 1 0 1748 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_19
timestamp 18001
transform 1 0 2852 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 18001
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1636986456
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_41
timestamp 18001
transform 1 0 4876 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1636986456
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1636986456
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1636986456
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_39
timestamp 18001
transform 1 0 4692 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_47
timestamp 18001
transform 1 0 5428 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_7
timestamp 1636986456
transform 1 0 1748 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_19
timestamp 18001
transform 1 0 2852 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 18001
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1636986456
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_41
timestamp 18001
transform 1 0 4876 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1636986456
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1636986456
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1636986456
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_39
timestamp 18001
transform 1 0 4692 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_47
timestamp 18001
transform 1 0 5428 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1636986456
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1636986456
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 18001
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1636986456
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_41
timestamp 18001
transform 1 0 4876 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_49
timestamp 18001
transform 1 0 5612 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_7
timestamp 1636986456
transform 1 0 1748 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_19
timestamp 1636986456
transform 1 0 2852 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_31
timestamp 1636986456
transform 1 0 3956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1636986456
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1636986456
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 18001
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1636986456
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_41
timestamp 18001
transform 1 0 4876 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_49
timestamp 18001
transform 1 0 5612 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_7
timestamp 1636986456
transform 1 0 1748 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_19
timestamp 1636986456
transform 1 0 2852 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_31
timestamp 1636986456
transform 1 0 3956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1636986456
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1636986456
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 18001
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1636986456
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_41
timestamp 18001
transform 1 0 4876 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_49
timestamp 18001
transform 1 0 5612 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1636986456
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1636986456
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1636986456
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_39
timestamp 18001
transform 1 0 4692 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_47
timestamp 18001
transform 1 0 5428 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_7
timestamp 1636986456
transform 1 0 1748 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_19
timestamp 18001
transform 1 0 2852 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 18001
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1636986456
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_41
timestamp 18001
transform 1 0 4876 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1636986456
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1636986456
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1636986456
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_39
timestamp 18001
transform 1 0 4692 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_47
timestamp 18001
transform 1 0 5428 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_62_7
timestamp 1636986456
transform 1 0 1748 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_19
timestamp 18001
transform 1 0 2852 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 18001
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1636986456
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_41
timestamp 18001
transform 1 0 4876 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1636986456
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1636986456
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1636986456
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_39
timestamp 18001
transform 1 0 4692 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_47
timestamp 18001
transform 1 0 5428 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1636986456
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1636986456
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 18001
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1636986456
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_41
timestamp 18001
transform 1 0 4876 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_49
timestamp 18001
transform 1 0 5612 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_7
timestamp 1636986456
transform 1 0 1748 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_19
timestamp 1636986456
transform 1 0 2852 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_31
timestamp 18001
transform 1 0 3956 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_39
timestamp 18001
transform 1 0 4692 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1636986456
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 1636986456
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 18001
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1636986456
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_41
timestamp 18001
transform 1 0 4876 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_49
timestamp 18001
transform 1 0 5612 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_7
timestamp 1636986456
transform 1 0 1748 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_19
timestamp 1636986456
transform 1 0 2852 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_31
timestamp 1636986456
transform 1 0 3956 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1636986456
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1636986456
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 18001
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1636986456
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_41
timestamp 18001
transform 1 0 4876 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_49
timestamp 18001
transform 1 0 5612 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1636986456
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1636986456
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1636986456
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_39
timestamp 18001
transform 1 0 4692 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_69_47
timestamp 18001
transform 1 0 5428 0 -1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_70_7
timestamp 1636986456
transform 1 0 1748 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_19
timestamp 18001
transform 1 0 2852 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 18001
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1636986456
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_41
timestamp 18001
transform 1 0 4876 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1636986456
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1636986456
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 1636986456
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_39
timestamp 18001
transform 1 0 4692 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_47
timestamp 18001
transform 1 0 5428 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_72_7
timestamp 1636986456
transform 1 0 1748 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_19
timestamp 18001
transform 1 0 2852 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 18001
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1636986456
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_41
timestamp 18001
transform 1 0 4876 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1636986456
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1636986456
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1636986456
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_39
timestamp 18001
transform 1 0 4692 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_73_47
timestamp 18001
transform 1 0 5428 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1636986456
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1636986456
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 18001
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1636986456
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_41
timestamp 18001
transform 1 0 4876 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_49
timestamp 18001
transform 1 0 5612 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_7
timestamp 1636986456
transform 1 0 1748 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_19
timestamp 1636986456
transform 1 0 2852 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_31
timestamp 18001
transform 1 0 3956 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_39
timestamp 18001
transform 1 0 4692 0 -1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_76_11
timestamp 1636986456
transform 1 0 2116 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_23
timestamp 18001
transform 1 0 3220 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 18001
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1636986456
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_41
timestamp 18001
transform 1 0 4876 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_76_49
timestamp 18001
transform 1 0 5612 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_7
timestamp 1636986456
transform 1 0 1748 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_19
timestamp 1636986456
transform 1 0 2852 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_31
timestamp 18001
transform 1 0 3956 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_77_39
timestamp 18001
transform 1 0 4692 0 -1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1636986456
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1636986456
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 18001
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1636986456
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_41
timestamp 18001
transform 1 0 4876 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_78_49
timestamp 18001
transform 1 0 5612 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_6
timestamp 1636986456
transform 1 0 1656 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_18
timestamp 1636986456
transform 1 0 2760 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_30
timestamp 1636986456
transform 1 0 3864 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_42
timestamp 18001
transform 1 0 4968 0 -1 45696
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_80_7
timestamp 1636986456
transform 1 0 1748 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_19
timestamp 18001
transform 1 0 2852 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 18001
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1636986456
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_41
timestamp 18001
transform 1 0 4876 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_6
timestamp 1636986456
transform 1 0 1656 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_18
timestamp 1636986456
transform 1 0 2760 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_30
timestamp 1636986456
transform 1 0 3864 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_42
timestamp 18001
transform 1 0 4968 0 -1 46784
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_82_6
timestamp 1636986456
transform 1 0 1656 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_18
timestamp 18001
transform 1 0 2760 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_26
timestamp 18001
transform 1 0 3496 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1636986456
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_41
timestamp 18001
transform 1 0 4876 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_83_3
timestamp 1636986456
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_15
timestamp 1636986456
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_27
timestamp 1636986456
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_39
timestamp 18001
transform 1 0 4692 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_83_47
timestamp 18001
transform 1 0 5428 0 -1 47872
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_84_6
timestamp 1636986456
transform 1 0 1656 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_18
timestamp 18001
transform 1 0 2760 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_84_26
timestamp 18001
transform 1 0 3496 0 1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1636986456
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_41
timestamp 18001
transform 1 0 4876 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_84_49
timestamp 18001
transform 1 0 5612 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_8
timestamp 1636986456
transform 1 0 1840 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_20
timestamp 1636986456
transform 1 0 2944 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_32
timestamp 1636986456
transform 1 0 4048 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_44
timestamp 18001
transform 1 0 5152 0 -1 48960
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_86_6
timestamp 1636986456
transform 1 0 1656 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_18
timestamp 18001
transform 1 0 2760 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_86_26
timestamp 18001
transform 1 0 3496 0 1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_86_29
timestamp 1636986456
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_41
timestamp 18001
transform 1 0 4876 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_86_49
timestamp 18001
transform 1 0 5612 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_6
timestamp 1636986456
transform 1 0 1656 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_18
timestamp 1636986456
transform 1 0 2760 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_30
timestamp 1636986456
transform 1 0 3864 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_42
timestamp 18001
transform 1 0 4968 0 -1 50048
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_88_3
timestamp 1636986456
transform 1 0 1380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_15
timestamp 1636986456
transform 1 0 2484 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_27
timestamp 18001
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_29
timestamp 1636986456
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_41
timestamp 18001
transform 1 0 4876 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_45
timestamp 18001
transform 1 0 5244 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_6
timestamp 1636986456
transform 1 0 1656 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_18
timestamp 1636986456
transform 1 0 2760 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_30
timestamp 18001
transform 1 0 3864 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_89_38
timestamp 18001
transform 1 0 4600 0 -1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_90_6
timestamp 1636986456
transform 1 0 1656 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_90_18
timestamp 18001
transform 1 0 2760 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_90_26
timestamp 18001
transform 1 0 3496 0 1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_90_29
timestamp 1636986456
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_90_41
timestamp 18001
transform 1 0 4876 0 1 51136
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_91_6
timestamp 1636986456
transform 1 0 1656 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_18
timestamp 1636986456
transform 1 0 2760 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_30
timestamp 1636986456
transform 1 0 3864 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_42
timestamp 18001
transform 1 0 4968 0 -1 52224
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_92_6
timestamp 1636986456
transform 1 0 1656 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_18
timestamp 18001
transform 1 0 2760 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_92_26
timestamp 18001
transform 1 0 3496 0 1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_92_29
timestamp 1636986456
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_92_41
timestamp 18001
transform 1 0 4876 0 1 52224
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_93_3
timestamp 1636986456
transform 1 0 1380 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_15
timestamp 1636986456
transform 1 0 2484 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_27
timestamp 1636986456
transform 1 0 3588 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_39
timestamp 18001
transform 1 0 4692 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_93_47
timestamp 18001
transform 1 0 5428 0 -1 53312
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_94_8
timestamp 1636986456
transform 1 0 1840 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_20
timestamp 18001
transform 1 0 2944 0 1 53312
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_94_29
timestamp 1636986456
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_41
timestamp 18001
transform 1 0 4876 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_94_49
timestamp 18001
transform 1 0 5612 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_6
timestamp 1636986456
transform 1 0 1656 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_18
timestamp 1636986456
transform 1 0 2760 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_30
timestamp 1636986456
transform 1 0 3864 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_95_42
timestamp 18001
transform 1 0 4968 0 -1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_96_8
timestamp 1636986456
transform 1 0 1840 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_96_20
timestamp 18001
transform 1 0 2944 0 1 54400
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_96_29
timestamp 1636986456
transform 1 0 3772 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_96_41
timestamp 18001
transform 1 0 4876 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_96_49
timestamp 18001
transform 1 0 5612 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_6
timestamp 1636986456
transform 1 0 1656 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_18
timestamp 1636986456
transform 1 0 2760 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_30
timestamp 1636986456
transform 1 0 3864 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_97_42
timestamp 18001
transform 1 0 4968 0 -1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_98_3
timestamp 1636986456
transform 1 0 1380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_15
timestamp 1636986456
transform 1 0 2484 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_27
timestamp 18001
transform 1 0 3588 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_29
timestamp 1636986456
transform 1 0 3772 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_41
timestamp 18001
transform 1 0 4876 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_98_49
timestamp 18001
transform 1 0 5612 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_8
timestamp 1636986456
transform 1 0 1840 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_20
timestamp 1636986456
transform 1 0 2944 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_32
timestamp 1636986456
transform 1 0 4048 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_6
timestamp 1636986456
transform 1 0 1656 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_18
timestamp 18001
transform 1 0 2760 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_100_26
timestamp 18001
transform 1 0 3496 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_100_29
timestamp 18001
transform 1 0 3772 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_8
timestamp 1636986456
transform 1 0 1840 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_20
timestamp 1636986456
transform 1 0 2944 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_32
timestamp 1636986456
transform 1 0 4048 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_101_44
timestamp 18001
transform 1 0 5152 0 -1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_102_6
timestamp 1636986456
transform 1 0 1656 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_102_18
timestamp 18001
transform 1 0 2760 0 1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_102_26
timestamp 18001
transform 1 0 3496 0 1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_102_29
timestamp 1636986456
transform 1 0 3772 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_102_41
timestamp 18001
transform 1 0 4876 0 1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_103_3
timestamp 1636986456
transform 1 0 1380 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_15
timestamp 1636986456
transform 1 0 2484 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_27
timestamp 1636986456
transform 1 0 3588 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_103_39
timestamp 18001
transform 1 0 4692 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_103_47
timestamp 18001
transform 1 0 5428 0 -1 58752
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_104_8
timestamp 1636986456
transform 1 0 1840 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_104_20
timestamp 18001
transform 1 0 2944 0 1 58752
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_104_29
timestamp 1636986456
transform 1 0 3772 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_104_41
timestamp 18001
transform 1 0 4876 0 1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_104_49
timestamp 18001
transform 1 0 5612 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_6
timestamp 1636986456
transform 1 0 1656 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_18
timestamp 1636986456
transform 1 0 2760 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_30
timestamp 1636986456
transform 1 0 3864 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_105_42
timestamp 18001
transform 1 0 4968 0 -1 59840
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_106_8
timestamp 1636986456
transform 1 0 1840 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_106_20
timestamp 18001
transform 1 0 2944 0 1 59840
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_106_29
timestamp 1636986456
transform 1 0 3772 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_106_41
timestamp 18001
transform 1 0 4876 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_106_49
timestamp 18001
transform 1 0 5612 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_6
timestamp 1636986456
transform 1 0 1656 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_18
timestamp 1636986456
transform 1 0 2760 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_30
timestamp 1636986456
transform 1 0 3864 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_107_42
timestamp 18001
transform 1 0 4968 0 -1 60928
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_108_3
timestamp 1636986456
transform 1 0 1380 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_15
timestamp 1636986456
transform 1 0 2484 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_108_27
timestamp 18001
transform 1 0 3588 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_29
timestamp 1636986456
transform 1 0 3772 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_108_41
timestamp 18001
transform 1 0 4876 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_108_49
timestamp 18001
transform 1 0 5612 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_8
timestamp 1636986456
transform 1 0 1840 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_20
timestamp 1636986456
transform 1 0 2944 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_32
timestamp 1636986456
transform 1 0 4048 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_44
timestamp 18001
transform 1 0 5152 0 -1 62016
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_110_8
timestamp 1636986456
transform 1 0 1840 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_110_20
timestamp 18001
transform 1 0 2944 0 1 62016
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_110_29
timestamp 1636986456
transform 1 0 3772 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_110_41
timestamp 18001
transform 1 0 4876 0 1 62016
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_111_3
timestamp 1636986456
transform 1 0 1380 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_15
timestamp 1636986456
transform 1 0 2484 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_27
timestamp 1636986456
transform 1 0 3588 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_111_39
timestamp 18001
transform 1 0 4692 0 -1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_111_47
timestamp 18001
transform 1 0 5428 0 -1 63104
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_112_8
timestamp 1636986456
transform 1 0 1840 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_112_20
timestamp 18001
transform 1 0 2944 0 1 63104
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_112_29
timestamp 1636986456
transform 1 0 3772 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_112_41
timestamp 18001
transform 1 0 4876 0 1 63104
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_113_3
timestamp 1636986456
transform 1 0 1380 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_15
timestamp 1636986456
transform 1 0 2484 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_27
timestamp 1636986456
transform 1 0 3588 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_113_39
timestamp 18001
transform 1 0 4692 0 -1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_113_47
timestamp 18001
transform 1 0 5428 0 -1 64192
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_114_3
timestamp 1636986456
transform 1 0 1380 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_15
timestamp 1636986456
transform 1 0 2484 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_114_27
timestamp 18001
transform 1 0 3588 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_29
timestamp 1636986456
transform 1 0 3772 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_114_41
timestamp 18001
transform 1 0 4876 0 1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_114_49
timestamp 18001
transform 1 0 5612 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_8
timestamp 1636986456
transform 1 0 1840 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_20
timestamp 1636986456
transform 1 0 2944 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_32
timestamp 1636986456
transform 1 0 4048 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_3
timestamp 1636986456
transform 1 0 1380 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_15
timestamp 1636986456
transform 1 0 2484 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_116_27
timestamp 18001
transform 1 0 3588 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_29
timestamp 1636986456
transform 1 0 3772 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_116_41
timestamp 18001
transform 1 0 4876 0 1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_116_49
timestamp 18001
transform 1 0 5612 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_8
timestamp 1636986456
transform 1 0 1840 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_20
timestamp 1636986456
transform 1 0 2944 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_32
timestamp 1636986456
transform 1 0 4048 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_3
timestamp 1636986456
transform 1 0 1380 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_15
timestamp 1636986456
transform 1 0 2484 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_118_27
timestamp 18001
transform 1 0 3588 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_29
timestamp 1636986456
transform 1 0 3772 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_118_41
timestamp 18001
transform 1 0 4876 0 1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_118_49
timestamp 18001
transform 1 0 5612 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_3
timestamp 1636986456
transform 1 0 1380 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_15
timestamp 1636986456
transform 1 0 2484 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_27
timestamp 1636986456
transform 1 0 3588 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_119_39
timestamp 18001
transform 1 0 4692 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_119_47
timestamp 18001
transform 1 0 5428 0 -1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_120_8
timestamp 1636986456
transform 1 0 1840 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_120_20
timestamp 18001
transform 1 0 2944 0 1 67456
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_120_29
timestamp 1636986456
transform 1 0 3772 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_120_41
timestamp 18001
transform 1 0 4876 0 1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_121_3
timestamp 1636986456
transform 1 0 1380 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_15
timestamp 1636986456
transform 1 0 2484 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_27
timestamp 1636986456
transform 1 0 3588 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_121_39
timestamp 18001
transform 1 0 4692 0 -1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_121_47
timestamp 18001
transform 1 0 5428 0 -1 68544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_122_8
timestamp 1636986456
transform 1 0 1840 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_122_20
timestamp 18001
transform 1 0 2944 0 1 68544
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_122_29
timestamp 1636986456
transform 1 0 3772 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_122_41
timestamp 18001
transform 1 0 4876 0 1 68544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_123_3
timestamp 1636986456
transform 1 0 1380 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_15
timestamp 1636986456
transform 1 0 2484 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_27
timestamp 1636986456
transform 1 0 3588 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_123_39
timestamp 18001
transform 1 0 4692 0 -1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_123_47
timestamp 18001
transform 1 0 5428 0 -1 69632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_124_3
timestamp 1636986456
transform 1 0 1380 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_15
timestamp 1636986456
transform 1 0 2484 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_124_27
timestamp 18001
transform 1 0 3588 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_29
timestamp 1636986456
transform 1 0 3772 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_124_41
timestamp 18001
transform 1 0 4876 0 1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_124_49
timestamp 18001
transform 1 0 5612 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_7
timestamp 1636986456
transform 1 0 1748 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_19
timestamp 1636986456
transform 1 0 2852 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_31
timestamp 1636986456
transform 1 0 3956 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_3
timestamp 1636986456
transform 1 0 1380 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_15
timestamp 1636986456
transform 1 0 2484 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_126_27
timestamp 18001
transform 1 0 3588 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_29
timestamp 1636986456
transform 1 0 3772 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_126_41
timestamp 18001
transform 1 0 4876 0 1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_126_49
timestamp 18001
transform 1 0 5612 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_7
timestamp 1636986456
transform 1 0 1748 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_19
timestamp 1636986456
transform 1 0 2852 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_31
timestamp 1636986456
transform 1 0 3956 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_3
timestamp 1636986456
transform 1 0 1380 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_15
timestamp 1636986456
transform 1 0 2484 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_128_27
timestamp 18001
transform 1 0 3588 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_29
timestamp 1636986456
transform 1 0 3772 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_128_41
timestamp 18001
transform 1 0 4876 0 1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_128_49
timestamp 18001
transform 1 0 5612 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_3
timestamp 1636986456
transform 1 0 1380 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_15
timestamp 1636986456
transform 1 0 2484 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_27
timestamp 1636986456
transform 1 0 3588 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_129_39
timestamp 18001
transform 1 0 4692 0 -1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_129_47
timestamp 18001
transform 1 0 5428 0 -1 72896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_130_7
timestamp 1636986456
transform 1 0 1748 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_130_19
timestamp 18001
transform 1 0 2852 0 1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_130_27
timestamp 18001
transform 1 0 3588 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_29
timestamp 1636986456
transform 1 0 3772 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_130_41
timestamp 18001
transform 1 0 4876 0 1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_130_49
timestamp 18001
transform 1 0 5612 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_3
timestamp 1636986456
transform 1 0 1380 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_15
timestamp 1636986456
transform 1 0 2484 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_27
timestamp 1636986456
transform 1 0 3588 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_131_39
timestamp 18001
transform 1 0 4692 0 -1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_131_47
timestamp 18001
transform 1 0 5428 0 -1 73984
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_132_7
timestamp 1636986456
transform 1 0 1748 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_132_19
timestamp 18001
transform 1 0 2852 0 1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_132_27
timestamp 18001
transform 1 0 3588 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_29
timestamp 1636986456
transform 1 0 3772 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_132_41
timestamp 18001
transform 1 0 4876 0 1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_132_49
timestamp 18001
transform 1 0 5612 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_3
timestamp 1636986456
transform 1 0 1380 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_15
timestamp 1636986456
transform 1 0 2484 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_27
timestamp 1636986456
transform 1 0 3588 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_133_39
timestamp 18001
transform 1 0 4692 0 -1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_133_47
timestamp 18001
transform 1 0 5428 0 -1 75072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_134_3
timestamp 1636986456
transform 1 0 1380 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_15
timestamp 1636986456
transform 1 0 2484 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_134_27
timestamp 18001
transform 1 0 3588 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_29
timestamp 1636986456
transform 1 0 3772 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_134_41
timestamp 18001
transform 1 0 4876 0 1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_134_49
timestamp 18001
transform 1 0 5612 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_7
timestamp 1636986456
transform 1 0 1748 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_19
timestamp 1636986456
transform 1 0 2852 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_31
timestamp 1636986456
transform 1 0 3956 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_43
timestamp 18001
transform 1 0 5060 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_49
timestamp 18001
transform 1 0 5612 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_3
timestamp 1636986456
transform 1 0 1380 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_15
timestamp 1636986456
transform 1 0 2484 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_136_27
timestamp 18001
transform 1 0 3588 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_29
timestamp 1636986456
transform 1 0 3772 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_136_41
timestamp 18001
transform 1 0 4876 0 1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_136_49
timestamp 18001
transform 1 0 5612 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_7
timestamp 1636986456
transform 1 0 1748 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_19
timestamp 1636986456
transform 1 0 2852 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_31
timestamp 1636986456
transform 1 0 3956 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_43
timestamp 18001
transform 1 0 5060 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_49
timestamp 18001
transform 1 0 5612 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_138_3
timestamp 1636986456
transform 1 0 1380 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_15
timestamp 1636986456
transform 1 0 2484 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_138_27
timestamp 18001
transform 1 0 3588 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_138_29
timestamp 1636986456
transform 1 0 3772 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_138_41
timestamp 18001
transform 1 0 4876 0 1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_138_49
timestamp 18001
transform 1 0 5612 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_139_3
timestamp 1636986456
transform 1 0 1380 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_15
timestamp 1636986456
transform 1 0 2484 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_27
timestamp 1636986456
transform 1 0 3588 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_139_39
timestamp 18001
transform 1 0 4692 0 -1 78336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_139_47
timestamp 18001
transform 1 0 5428 0 -1 78336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_140_7
timestamp 1636986456
transform 1 0 1748 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_140_19
timestamp 18001
transform 1 0 2852 0 1 78336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_140_27
timestamp 18001
transform 1 0 3588 0 1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_140_29
timestamp 1636986456
transform 1 0 3772 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_140_41
timestamp 18001
transform 1 0 4876 0 1 78336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_140_49
timestamp 18001
transform 1 0 5612 0 1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_141_3
timestamp 1636986456
transform 1 0 1380 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_15
timestamp 1636986456
transform 1 0 2484 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_27
timestamp 1636986456
transform 1 0 3588 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_141_39
timestamp 18001
transform 1 0 4692 0 -1 79424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_141_47
timestamp 18001
transform 1 0 5428 0 -1 79424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_142_7
timestamp 1636986456
transform 1 0 1748 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_142_19
timestamp 18001
transform 1 0 2852 0 1 79424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_142_27
timestamp 18001
transform 1 0 3588 0 1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_142_29
timestamp 1636986456
transform 1 0 3772 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_142_41
timestamp 18001
transform 1 0 4876 0 1 79424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_142_49
timestamp 18001
transform 1 0 5612 0 1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_143_3
timestamp 1636986456
transform 1 0 1380 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_15
timestamp 1636986456
transform 1 0 2484 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_27
timestamp 1636986456
transform 1 0 3588 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_143_39
timestamp 18001
transform 1 0 4692 0 -1 80512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_143_47
timestamp 18001
transform 1 0 5428 0 -1 80512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_144_3
timestamp 1636986456
transform 1 0 1380 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_15
timestamp 1636986456
transform 1 0 2484 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_144_27
timestamp 18001
transform 1 0 3588 0 1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_144_29
timestamp 1636986456
transform 1 0 3772 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_144_41
timestamp 18001
transform 1 0 4876 0 1 80512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_144_49
timestamp 18001
transform 1 0 5612 0 1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_145_7
timestamp 1636986456
transform 1 0 1748 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_19
timestamp 1636986456
transform 1 0 2852 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_31
timestamp 1636986456
transform 1 0 3956 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_145_43
timestamp 18001
transform 1 0 5060 0 -1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_145_49
timestamp 18001
transform 1 0 5612 0 -1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_146_3
timestamp 1636986456
transform 1 0 1380 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_15
timestamp 1636986456
transform 1 0 2484 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_146_27
timestamp 18001
transform 1 0 3588 0 1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_146_29
timestamp 1636986456
transform 1 0 3772 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_146_41
timestamp 18001
transform 1 0 4876 0 1 81600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_146_49
timestamp 18001
transform 1 0 5612 0 1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_7
timestamp 1636986456
transform 1 0 1748 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_19
timestamp 1636986456
transform 1 0 2852 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_31
timestamp 1636986456
transform 1 0 3956 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_43
timestamp 18001
transform 1 0 5060 0 -1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_49
timestamp 18001
transform 1 0 5612 0 -1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_3
timestamp 1636986456
transform 1 0 1380 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_15
timestamp 1636986456
transform 1 0 2484 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_148_27
timestamp 18001
transform 1 0 3588 0 1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_29
timestamp 1636986456
transform 1 0 3772 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_148_41
timestamp 18001
transform 1 0 4876 0 1 82688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_148_49
timestamp 18001
transform 1 0 5612 0 1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_3
timestamp 1636986456
transform 1 0 1380 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_15
timestamp 1636986456
transform 1 0 2484 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_27
timestamp 1636986456
transform 1 0 3588 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_149_39
timestamp 18001
transform 1 0 4692 0 -1 83776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_149_47
timestamp 18001
transform 1 0 5428 0 -1 83776
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_150_7
timestamp 1636986456
transform 1 0 1748 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_150_19
timestamp 18001
transform 1 0 2852 0 1 83776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_150_27
timestamp 18001
transform 1 0 3588 0 1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_29
timestamp 1636986456
transform 1 0 3772 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_150_41
timestamp 18001
transform 1 0 4876 0 1 83776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_150_49
timestamp 18001
transform 1 0 5612 0 1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_151_3
timestamp 1636986456
transform 1 0 1380 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_15
timestamp 1636986456
transform 1 0 2484 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_27
timestamp 1636986456
transform 1 0 3588 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_151_39
timestamp 18001
transform 1 0 4692 0 -1 84864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_151_47
timestamp 18001
transform 1 0 5428 0 -1 84864
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_152_7
timestamp 1636986456
transform 1 0 1748 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_152_19
timestamp 18001
transform 1 0 2852 0 1 84864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_152_27
timestamp 18001
transform 1 0 3588 0 1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_152_29
timestamp 1636986456
transform 1 0 3772 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_152_41
timestamp 18001
transform 1 0 4876 0 1 84864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_152_49
timestamp 18001
transform 1 0 5612 0 1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_153_3
timestamp 1636986456
transform 1 0 1380 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_15
timestamp 1636986456
transform 1 0 2484 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_27
timestamp 1636986456
transform 1 0 3588 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_153_39
timestamp 18001
transform 1 0 4692 0 -1 85952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_153_47
timestamp 18001
transform 1 0 5428 0 -1 85952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_154_3
timestamp 1636986456
transform 1 0 1380 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_15
timestamp 1636986456
transform 1 0 2484 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_154_27
timestamp 18001
transform 1 0 3588 0 1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_154_29
timestamp 1636986456
transform 1 0 3772 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_154_41
timestamp 18001
transform 1 0 4876 0 1 85952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_154_49
timestamp 18001
transform 1 0 5612 0 1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_155_7
timestamp 1636986456
transform 1 0 1748 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_19
timestamp 1636986456
transform 1 0 2852 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_31
timestamp 1636986456
transform 1 0 3956 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_155_43
timestamp 18001
transform 1 0 5060 0 -1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_155_49
timestamp 18001
transform 1 0 5612 0 -1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_156_3
timestamp 1636986456
transform 1 0 1380 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_15
timestamp 1636986456
transform 1 0 2484 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_156_27
timestamp 18001
transform 1 0 3588 0 1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_156_29
timestamp 1636986456
transform 1 0 3772 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_156_41
timestamp 18001
transform 1 0 4876 0 1 87040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_156_49
timestamp 18001
transform 1 0 5612 0 1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_157_3
timestamp 1636986456
transform 1 0 1380 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_15
timestamp 1636986456
transform 1 0 2484 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_27
timestamp 1636986456
transform 1 0 3588 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_157_39
timestamp 18001
transform 1 0 4692 0 -1 88128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_157_47
timestamp 18001
transform 1 0 5428 0 -1 88128
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_158_3
timestamp 1636986456
transform 1 0 1380 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_15
timestamp 1636986456
transform 1 0 2484 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_158_27
timestamp 18001
transform 1 0 3588 0 1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_158_29
timestamp 1636986456
transform 1 0 3772 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_158_41
timestamp 18001
transform 1 0 4876 0 1 88128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_158_49
timestamp 18001
transform 1 0 5612 0 1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_159_3
timestamp 1636986456
transform 1 0 1380 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_15
timestamp 1636986456
transform 1 0 2484 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_27
timestamp 1636986456
transform 1 0 3588 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_159_39
timestamp 18001
transform 1 0 4692 0 -1 89216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_159_47
timestamp 18001
transform 1 0 5428 0 -1 89216
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_160_3
timestamp 1636986456
transform 1 0 1380 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_15
timestamp 1636986456
transform 1 0 2484 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_160_27
timestamp 18001
transform 1 0 3588 0 1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_160_29
timestamp 1636986456
transform 1 0 3772 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_160_41
timestamp 18001
transform 1 0 4876 0 1 89216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_160_49
timestamp 18001
transform 1 0 5612 0 1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_161_3
timestamp 1636986456
transform 1 0 1380 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_15
timestamp 1636986456
transform 1 0 2484 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_27
timestamp 1636986456
transform 1 0 3588 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_161_39
timestamp 18001
transform 1 0 4692 0 -1 90304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_161_47
timestamp 18001
transform 1 0 5428 0 -1 90304
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_162_3
timestamp 1636986456
transform 1 0 1380 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_15
timestamp 1636986456
transform 1 0 2484 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_162_27
timestamp 18001
transform 1 0 3588 0 1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_162_29
timestamp 1636986456
transform 1 0 3772 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_162_41
timestamp 18001
transform 1 0 4876 0 1 90304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_162_49
timestamp 18001
transform 1 0 5612 0 1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_163_3
timestamp 1636986456
transform 1 0 1380 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_15
timestamp 1636986456
transform 1 0 2484 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_27
timestamp 1636986456
transform 1 0 3588 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_163_39
timestamp 18001
transform 1 0 4692 0 -1 91392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_163_47
timestamp 18001
transform 1 0 5428 0 -1 91392
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_164_3
timestamp 1636986456
transform 1 0 1380 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_15
timestamp 1636986456
transform 1 0 2484 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_164_27
timestamp 18001
transform 1 0 3588 0 1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_164_29
timestamp 1636986456
transform 1 0 3772 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_41
timestamp 1636986456
transform 1 0 4876 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_164_53
timestamp 18001
transform 1 0 5980 0 1 91392
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_164_57
timestamp 1636986456
transform 1 0 6348 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_69
timestamp 1636986456
transform 1 0 7452 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_164_81
timestamp 18001
transform 1 0 8556 0 1 91392
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_164_85
timestamp 1636986456
transform 1 0 8924 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_164_97
timestamp 18001
transform 1 0 10028 0 1 91392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_164_101
timestamp 18001
transform 1 0 10396 0 1 91392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_164_109
timestamp 18001
transform 1 0 11132 0 1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_164_115
timestamp 18001
transform 1 0 11684 0 1 91392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_164_125
timestamp 18001
transform 1 0 12604 0 1 91392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_164_133
timestamp 18001
transform 1 0 13340 0 1 91392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_164_137
timestamp 18001
transform 1 0 13708 0 1 91392
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_164_141
timestamp 1636986456
transform 1 0 14076 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_153
timestamp 1636986456
transform 1 0 15180 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_164_165
timestamp 18001
transform 1 0 16284 0 1 91392
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_164_169
timestamp 1636986456
transform 1 0 16652 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_181
timestamp 1636986456
transform 1 0 17756 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_164_193
timestamp 18001
transform 1 0 18860 0 1 91392
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_164_197
timestamp 1636986456
transform 1 0 19228 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_209
timestamp 1636986456
transform 1 0 20332 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_164_221
timestamp 18001
transform 1 0 21436 0 1 91392
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_164_225
timestamp 1636986456
transform 1 0 21804 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_237
timestamp 1636986456
transform 1 0 22908 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_164_249
timestamp 18001
transform 1 0 24012 0 1 91392
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_164_253
timestamp 1636986456
transform 1 0 24380 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_265
timestamp 1636986456
transform 1 0 25484 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_164_277
timestamp 18001
transform 1 0 26588 0 1 91392
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_164_281
timestamp 1636986456
transform 1 0 26956 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_293
timestamp 1636986456
transform 1 0 28060 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_164_305
timestamp 18001
transform 1 0 29164 0 1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_164_309
timestamp 18001
transform 1 0 29532 0 1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_164_315
timestamp 18001
transform 1 0 30084 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_164_337
timestamp 18001
transform 1 0 32108 0 1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_164_342
timestamp 1636986456
transform 1 0 32568 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_164_354
timestamp 18001
transform 1 0 33672 0 1 91392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_164_362
timestamp 18001
transform 1 0 34408 0 1 91392
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_164_365
timestamp 1636986456
transform 1 0 34684 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_377
timestamp 1636986456
transform 1 0 35788 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_164_389
timestamp 18001
transform 1 0 36892 0 1 91392
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_164_393
timestamp 1636986456
transform 1 0 37260 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_405
timestamp 1636986456
transform 1 0 38364 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_164_417
timestamp 18001
transform 1 0 39468 0 1 91392
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_164_421
timestamp 1636986456
transform 1 0 39836 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_433
timestamp 1636986456
transform 1 0 40940 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_164_445
timestamp 18001
transform 1 0 42044 0 1 91392
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_164_449
timestamp 1636986456
transform 1 0 42412 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_461
timestamp 1636986456
transform 1 0 43516 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_164_473
timestamp 18001
transform 1 0 44620 0 1 91392
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_164_477
timestamp 1636986456
transform 1 0 44988 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_489
timestamp 1636986456
transform 1 0 46092 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_164_501
timestamp 18001
transform 1 0 47196 0 1 91392
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_164_505
timestamp 1636986456
transform 1 0 47564 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_164_517
timestamp 18001
transform 1 0 48668 0 1 91392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_164_525
timestamp 18001
transform 1 0 49404 0 1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_164_530
timestamp 18001
transform 1 0 49864 0 1 91392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_164_533
timestamp 18001
transform 1 0 50140 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_164_536
timestamp 18001
transform 1 0 50416 0 1 91392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_164_583
timestamp 18001
transform 1 0 54740 0 1 91392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_164_587
timestamp 18001
transform 1 0 55108 0 1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_164_589
timestamp 1636986456
transform 1 0 55292 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_601
timestamp 1636986456
transform 1 0 56396 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_164_613
timestamp 18001
transform 1 0 57500 0 1 91392
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_164_617
timestamp 1636986456
transform 1 0 57868 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_629
timestamp 1636986456
transform 1 0 58972 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_164_641
timestamp 18001
transform 1 0 60076 0 1 91392
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_164_645
timestamp 1636986456
transform 1 0 60444 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_657
timestamp 1636986456
transform 1 0 61548 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_164_669
timestamp 18001
transform 1 0 62652 0 1 91392
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_164_673
timestamp 1636986456
transform 1 0 63020 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_685
timestamp 1636986456
transform 1 0 64124 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_164_697
timestamp 18001
transform 1 0 65228 0 1 91392
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_164_701
timestamp 1636986456
transform 1 0 65596 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_713
timestamp 1636986456
transform 1 0 66700 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_164_725
timestamp 18001
transform 1 0 67804 0 1 91392
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_164_729
timestamp 1636986456
transform 1 0 68172 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_741
timestamp 1636986456
transform 1 0 69276 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_164_753
timestamp 18001
transform 1 0 70380 0 1 91392
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_164_757
timestamp 1636986456
transform 1 0 70748 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_769
timestamp 1636986456
transform 1 0 71852 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_164_781
timestamp 18001
transform 1 0 72956 0 1 91392
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_164_785
timestamp 1636986456
transform 1 0 73324 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_797
timestamp 1636986456
transform 1 0 74428 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_164_809
timestamp 18001
transform 1 0 75532 0 1 91392
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_164_813
timestamp 1636986456
transform 1 0 75900 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_825
timestamp 1636986456
transform 1 0 77004 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_164_837
timestamp 18001
transform 1 0 78108 0 1 91392
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_164_841
timestamp 1636986456
transform 1 0 78476 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_853
timestamp 1636986456
transform 1 0 79580 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_164_865
timestamp 18001
transform 1 0 80684 0 1 91392
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_164_869
timestamp 1636986456
transform 1 0 81052 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_881
timestamp 1636986456
transform 1 0 82156 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_164_893
timestamp 18001
transform 1 0 83260 0 1 91392
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_164_897
timestamp 1636986456
transform 1 0 83628 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_164_909
timestamp 18001
transform 1 0 84732 0 1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_164_925
timestamp 18001
transform 1 0 86204 0 1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_165_3
timestamp 1636986456
transform 1 0 1380 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_15
timestamp 1636986456
transform 1 0 2484 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_27
timestamp 1636986456
transform 1 0 3588 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_39
timestamp 1636986456
transform 1 0 4692 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_165_51
timestamp 18001
transform 1 0 5796 0 -1 92480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_165_55
timestamp 18001
transform 1 0 6164 0 -1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_165_57
timestamp 1636986456
transform 1 0 6348 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_69
timestamp 1636986456
transform 1 0 7452 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_81
timestamp 1636986456
transform 1 0 8556 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_93
timestamp 1636986456
transform 1 0 9660 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_165_105
timestamp 18001
transform 1 0 10764 0 -1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_165_111
timestamp 18001
transform 1 0 11316 0 -1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_165_113
timestamp 1636986456
transform 1 0 11500 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_125
timestamp 1636986456
transform 1 0 12604 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_137
timestamp 1636986456
transform 1 0 13708 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_149
timestamp 1636986456
transform 1 0 14812 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_165_161
timestamp 18001
transform 1 0 15916 0 -1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_165_167
timestamp 18001
transform 1 0 16468 0 -1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_165_169
timestamp 1636986456
transform 1 0 16652 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_181
timestamp 1636986456
transform 1 0 17756 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_193
timestamp 1636986456
transform 1 0 18860 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_205
timestamp 1636986456
transform 1 0 19964 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_165_217
timestamp 18001
transform 1 0 21068 0 -1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_165_223
timestamp 18001
transform 1 0 21620 0 -1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_165_225
timestamp 1636986456
transform 1 0 21804 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_237
timestamp 1636986456
transform 1 0 22908 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_249
timestamp 1636986456
transform 1 0 24012 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_261
timestamp 1636986456
transform 1 0 25116 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_165_273
timestamp 18001
transform 1 0 26220 0 -1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_165_279
timestamp 18001
transform 1 0 26772 0 -1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_165_281
timestamp 1636986456
transform 1 0 26956 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_293
timestamp 1636986456
transform 1 0 28060 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_165_305
timestamp 18001
transform 1 0 29164 0 -1 92480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_165_313
timestamp 18001
transform 1 0 29900 0 -1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_165_337
timestamp 18001
transform 1 0 32108 0 -1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_165_342
timestamp 1636986456
transform 1 0 32568 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_354
timestamp 1636986456
transform 1 0 33672 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_366
timestamp 1636986456
transform 1 0 34776 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_378
timestamp 1636986456
transform 1 0 35880 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_165_390
timestamp 18001
transform 1 0 36984 0 -1 92480
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_165_393
timestamp 1636986456
transform 1 0 37260 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_405
timestamp 1636986456
transform 1 0 38364 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_417
timestamp 1636986456
transform 1 0 39468 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_429
timestamp 1636986456
transform 1 0 40572 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_165_441
timestamp 18001
transform 1 0 41676 0 -1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_165_447
timestamp 18001
transform 1 0 42228 0 -1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_165_449
timestamp 1636986456
transform 1 0 42412 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_461
timestamp 1636986456
transform 1 0 43516 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_473
timestamp 1636986456
transform 1 0 44620 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_485
timestamp 1636986456
transform 1 0 45724 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_165_497
timestamp 18001
transform 1 0 46828 0 -1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_165_503
timestamp 18001
transform 1 0 47380 0 -1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_165_505
timestamp 1636986456
transform 1 0 47564 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_517
timestamp 1636986456
transform 1 0 48668 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_529
timestamp 1636986456
transform 1 0 49772 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_165_541
timestamp 18001
transform 1 0 50876 0 -1 92480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_165_549
timestamp 18001
transform 1 0 51612 0 -1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_165_554
timestamp 18001
transform 1 0 52072 0 -1 92480
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_165_567
timestamp 1636986456
transform 1 0 53268 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_579
timestamp 1636986456
transform 1 0 54372 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_591
timestamp 1636986456
transform 1 0 55476 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_603
timestamp 1636986456
transform 1 0 56580 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_165_615
timestamp 18001
transform 1 0 57684 0 -1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_165_617
timestamp 1636986456
transform 1 0 57868 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_629
timestamp 1636986456
transform 1 0 58972 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_641
timestamp 1636986456
transform 1 0 60076 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_653
timestamp 1636986456
transform 1 0 61180 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_165_665
timestamp 18001
transform 1 0 62284 0 -1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_165_671
timestamp 18001
transform 1 0 62836 0 -1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_165_673
timestamp 1636986456
transform 1 0 63020 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_685
timestamp 1636986456
transform 1 0 64124 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_697
timestamp 1636986456
transform 1 0 65228 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_709
timestamp 1636986456
transform 1 0 66332 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_165_721
timestamp 18001
transform 1 0 67436 0 -1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_165_727
timestamp 18001
transform 1 0 67988 0 -1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_165_729
timestamp 1636986456
transform 1 0 68172 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_741
timestamp 1636986456
transform 1 0 69276 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_753
timestamp 1636986456
transform 1 0 70380 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_765
timestamp 1636986456
transform 1 0 71484 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_165_777
timestamp 18001
transform 1 0 72588 0 -1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_165_783
timestamp 18001
transform 1 0 73140 0 -1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_165_785
timestamp 1636986456
transform 1 0 73324 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_797
timestamp 1636986456
transform 1 0 74428 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_809
timestamp 1636986456
transform 1 0 75532 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_821
timestamp 1636986456
transform 1 0 76636 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_165_833
timestamp 18001
transform 1 0 77740 0 -1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_165_839
timestamp 18001
transform 1 0 78292 0 -1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_165_841
timestamp 1636986456
transform 1 0 78476 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_853
timestamp 1636986456
transform 1 0 79580 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_865
timestamp 1636986456
transform 1 0 80684 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_877
timestamp 1636986456
transform 1 0 81788 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_165_889
timestamp 18001
transform 1 0 82892 0 -1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_165_895
timestamp 18001
transform 1 0 83444 0 -1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_165_897
timestamp 1636986456
transform 1 0 83628 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_165_909
timestamp 18001
transform 1 0 84732 0 -1 92480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_165_917
timestamp 18001
transform 1 0 85468 0 -1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_165_933
timestamp 18001
transform 1 0 86940 0 -1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_3
timestamp 1636986456
transform 1 0 1380 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_15
timestamp 1636986456
transform 1 0 2484 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_166_27
timestamp 18001
transform 1 0 3588 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_29
timestamp 1636986456
transform 1 0 3772 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_41
timestamp 1636986456
transform 1 0 4876 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_53
timestamp 1636986456
transform 1 0 5980 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_65
timestamp 1636986456
transform 1 0 7084 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_77
timestamp 18001
transform 1 0 8188 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_83
timestamp 18001
transform 1 0 8740 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_85
timestamp 1636986456
transform 1 0 8924 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_97
timestamp 1636986456
transform 1 0 10028 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_109
timestamp 1636986456
transform 1 0 11132 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_121
timestamp 1636986456
transform 1 0 12236 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_133
timestamp 18001
transform 1 0 13340 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_139
timestamp 18001
transform 1 0 13892 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_141
timestamp 1636986456
transform 1 0 14076 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_153
timestamp 1636986456
transform 1 0 15180 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_165
timestamp 1636986456
transform 1 0 16284 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_177
timestamp 1636986456
transform 1 0 17388 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_189
timestamp 18001
transform 1 0 18492 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_195
timestamp 18001
transform 1 0 19044 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_197
timestamp 1636986456
transform 1 0 19228 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_209
timestamp 1636986456
transform 1 0 20332 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_221
timestamp 1636986456
transform 1 0 21436 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_233
timestamp 1636986456
transform 1 0 22540 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_245
timestamp 18001
transform 1 0 23644 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_251
timestamp 18001
transform 1 0 24196 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_253
timestamp 1636986456
transform 1 0 24380 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_265
timestamp 1636986456
transform 1 0 25484 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_277
timestamp 1636986456
transform 1 0 26588 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_289
timestamp 1636986456
transform 1 0 27692 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_301
timestamp 18001
transform 1 0 28796 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_307
timestamp 18001
transform 1 0 29348 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_309
timestamp 1636986456
transform 1 0 29532 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_321
timestamp 1636986456
transform 1 0 30636 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_333
timestamp 1636986456
transform 1 0 31740 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_345
timestamp 1636986456
transform 1 0 32844 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_357
timestamp 18001
transform 1 0 33948 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_363
timestamp 18001
transform 1 0 34500 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_365
timestamp 1636986456
transform 1 0 34684 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_377
timestamp 1636986456
transform 1 0 35788 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_389
timestamp 1636986456
transform 1 0 36892 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_401
timestamp 1636986456
transform 1 0 37996 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_413
timestamp 18001
transform 1 0 39100 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_419
timestamp 18001
transform 1 0 39652 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_421
timestamp 1636986456
transform 1 0 39836 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_433
timestamp 1636986456
transform 1 0 40940 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_445
timestamp 1636986456
transform 1 0 42044 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_457
timestamp 1636986456
transform 1 0 43148 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_469
timestamp 18001
transform 1 0 44252 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_475
timestamp 18001
transform 1 0 44804 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_477
timestamp 1636986456
transform 1 0 44988 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_489
timestamp 1636986456
transform 1 0 46092 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_501
timestamp 1636986456
transform 1 0 47196 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_513
timestamp 1636986456
transform 1 0 48300 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_525
timestamp 18001
transform 1 0 49404 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_531
timestamp 18001
transform 1 0 49956 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_533
timestamp 1636986456
transform 1 0 50140 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_545
timestamp 1636986456
transform 1 0 51244 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_557
timestamp 1636986456
transform 1 0 52348 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_569
timestamp 1636986456
transform 1 0 53452 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_581
timestamp 18001
transform 1 0 54556 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_587
timestamp 18001
transform 1 0 55108 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_589
timestamp 1636986456
transform 1 0 55292 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_601
timestamp 1636986456
transform 1 0 56396 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_613
timestamp 1636986456
transform 1 0 57500 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_625
timestamp 1636986456
transform 1 0 58604 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_637
timestamp 18001
transform 1 0 59708 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_643
timestamp 18001
transform 1 0 60260 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_645
timestamp 1636986456
transform 1 0 60444 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_657
timestamp 1636986456
transform 1 0 61548 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_669
timestamp 1636986456
transform 1 0 62652 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_681
timestamp 1636986456
transform 1 0 63756 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_693
timestamp 18001
transform 1 0 64860 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_699
timestamp 18001
transform 1 0 65412 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_701
timestamp 1636986456
transform 1 0 65596 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_713
timestamp 1636986456
transform 1 0 66700 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_725
timestamp 1636986456
transform 1 0 67804 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_737
timestamp 1636986456
transform 1 0 68908 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_749
timestamp 18001
transform 1 0 70012 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_755
timestamp 18001
transform 1 0 70564 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_757
timestamp 1636986456
transform 1 0 70748 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_769
timestamp 1636986456
transform 1 0 71852 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_781
timestamp 1636986456
transform 1 0 72956 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_793
timestamp 1636986456
transform 1 0 74060 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_805
timestamp 18001
transform 1 0 75164 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_811
timestamp 18001
transform 1 0 75716 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_813
timestamp 1636986456
transform 1 0 75900 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_825
timestamp 1636986456
transform 1 0 77004 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_837
timestamp 1636986456
transform 1 0 78108 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_849
timestamp 1636986456
transform 1 0 79212 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_861
timestamp 18001
transform 1 0 80316 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_867
timestamp 18001
transform 1 0 80868 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_869
timestamp 1636986456
transform 1 0 81052 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_881
timestamp 1636986456
transform 1 0 82156 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_893
timestamp 1636986456
transform 1 0 83260 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_905
timestamp 1636986456
transform 1 0 84364 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_917
timestamp 18001
transform 1 0 85468 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_923
timestamp 18001
transform 1 0 86020 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_166_925
timestamp 18001
transform 1 0 86204 0 1 92480
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_167_3
timestamp 1636986456
transform 1 0 1380 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_15
timestamp 1636986456
transform 1 0 2484 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_27
timestamp 1636986456
transform 1 0 3588 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_39
timestamp 1636986456
transform 1 0 4692 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_167_51
timestamp 18001
transform 1 0 5796 0 -1 93568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_167_55
timestamp 18001
transform 1 0 6164 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_57
timestamp 1636986456
transform 1 0 6348 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_69
timestamp 1636986456
transform 1 0 7452 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_81
timestamp 1636986456
transform 1 0 8556 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_93
timestamp 1636986456
transform 1 0 9660 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_105
timestamp 18001
transform 1 0 10764 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_111
timestamp 18001
transform 1 0 11316 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_113
timestamp 1636986456
transform 1 0 11500 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_125
timestamp 1636986456
transform 1 0 12604 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_137
timestamp 1636986456
transform 1 0 13708 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_149
timestamp 1636986456
transform 1 0 14812 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_161
timestamp 18001
transform 1 0 15916 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_167
timestamp 18001
transform 1 0 16468 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_169
timestamp 1636986456
transform 1 0 16652 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_181
timestamp 1636986456
transform 1 0 17756 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_193
timestamp 1636986456
transform 1 0 18860 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_205
timestamp 1636986456
transform 1 0 19964 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_217
timestamp 18001
transform 1 0 21068 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_223
timestamp 18001
transform 1 0 21620 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_225
timestamp 1636986456
transform 1 0 21804 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_237
timestamp 1636986456
transform 1 0 22908 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_249
timestamp 1636986456
transform 1 0 24012 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_261
timestamp 1636986456
transform 1 0 25116 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_273
timestamp 18001
transform 1 0 26220 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_279
timestamp 18001
transform 1 0 26772 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_281
timestamp 1636986456
transform 1 0 26956 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_293
timestamp 1636986456
transform 1 0 28060 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_305
timestamp 1636986456
transform 1 0 29164 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_317
timestamp 1636986456
transform 1 0 30268 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_329
timestamp 18001
transform 1 0 31372 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_335
timestamp 18001
transform 1 0 31924 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_337
timestamp 1636986456
transform 1 0 32108 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_349
timestamp 1636986456
transform 1 0 33212 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_361
timestamp 1636986456
transform 1 0 34316 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_373
timestamp 1636986456
transform 1 0 35420 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_385
timestamp 18001
transform 1 0 36524 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_391
timestamp 18001
transform 1 0 37076 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_393
timestamp 1636986456
transform 1 0 37260 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_405
timestamp 1636986456
transform 1 0 38364 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_417
timestamp 1636986456
transform 1 0 39468 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_429
timestamp 1636986456
transform 1 0 40572 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_441
timestamp 18001
transform 1 0 41676 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_447
timestamp 18001
transform 1 0 42228 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_449
timestamp 1636986456
transform 1 0 42412 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_461
timestamp 1636986456
transform 1 0 43516 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_473
timestamp 1636986456
transform 1 0 44620 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_485
timestamp 1636986456
transform 1 0 45724 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_497
timestamp 18001
transform 1 0 46828 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_503
timestamp 18001
transform 1 0 47380 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_505
timestamp 1636986456
transform 1 0 47564 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_517
timestamp 1636986456
transform 1 0 48668 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_529
timestamp 1636986456
transform 1 0 49772 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_541
timestamp 1636986456
transform 1 0 50876 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_553
timestamp 18001
transform 1 0 51980 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_559
timestamp 18001
transform 1 0 52532 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_561
timestamp 1636986456
transform 1 0 52716 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_573
timestamp 1636986456
transform 1 0 53820 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_585
timestamp 1636986456
transform 1 0 54924 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_597
timestamp 1636986456
transform 1 0 56028 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_609
timestamp 18001
transform 1 0 57132 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_615
timestamp 18001
transform 1 0 57684 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_617
timestamp 1636986456
transform 1 0 57868 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_629
timestamp 1636986456
transform 1 0 58972 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_641
timestamp 1636986456
transform 1 0 60076 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_653
timestamp 1636986456
transform 1 0 61180 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_665
timestamp 18001
transform 1 0 62284 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_671
timestamp 18001
transform 1 0 62836 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_673
timestamp 1636986456
transform 1 0 63020 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_685
timestamp 1636986456
transform 1 0 64124 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_697
timestamp 1636986456
transform 1 0 65228 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_709
timestamp 1636986456
transform 1 0 66332 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_721
timestamp 18001
transform 1 0 67436 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_727
timestamp 18001
transform 1 0 67988 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_729
timestamp 1636986456
transform 1 0 68172 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_741
timestamp 1636986456
transform 1 0 69276 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_753
timestamp 1636986456
transform 1 0 70380 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_765
timestamp 1636986456
transform 1 0 71484 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_777
timestamp 18001
transform 1 0 72588 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_783
timestamp 18001
transform 1 0 73140 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_785
timestamp 1636986456
transform 1 0 73324 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_797
timestamp 1636986456
transform 1 0 74428 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_809
timestamp 1636986456
transform 1 0 75532 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_821
timestamp 1636986456
transform 1 0 76636 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_833
timestamp 18001
transform 1 0 77740 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_839
timestamp 18001
transform 1 0 78292 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_841
timestamp 1636986456
transform 1 0 78476 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_853
timestamp 1636986456
transform 1 0 79580 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_865
timestamp 1636986456
transform 1 0 80684 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_877
timestamp 1636986456
transform 1 0 81788 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_889
timestamp 18001
transform 1 0 82892 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_895
timestamp 18001
transform 1 0 83444 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_897
timestamp 1636986456
transform 1 0 83628 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_909
timestamp 1636986456
transform 1 0 84732 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_921
timestamp 1636986456
transform 1 0 85836 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_167_933
timestamp 18001
transform 1 0 86940 0 -1 93568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_167_939
timestamp 18001
transform 1 0 87492 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_167_942
timestamp 18001
transform 1 0 87768 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_3
timestamp 1636986456
transform 1 0 1380 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_15
timestamp 1636986456
transform 1 0 2484 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_168_27
timestamp 18001
transform 1 0 3588 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_29
timestamp 1636986456
transform 1 0 3772 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_41
timestamp 1636986456
transform 1 0 4876 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_53
timestamp 1636986456
transform 1 0 5980 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_65
timestamp 1636986456
transform 1 0 7084 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_77
timestamp 18001
transform 1 0 8188 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_83
timestamp 18001
transform 1 0 8740 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_85
timestamp 1636986456
transform 1 0 8924 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_97
timestamp 1636986456
transform 1 0 10028 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_109
timestamp 1636986456
transform 1 0 11132 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_121
timestamp 1636986456
transform 1 0 12236 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_133
timestamp 18001
transform 1 0 13340 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_139
timestamp 18001
transform 1 0 13892 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_141
timestamp 1636986456
transform 1 0 14076 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_153
timestamp 1636986456
transform 1 0 15180 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_165
timestamp 1636986456
transform 1 0 16284 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_177
timestamp 1636986456
transform 1 0 17388 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_189
timestamp 18001
transform 1 0 18492 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_195
timestamp 18001
transform 1 0 19044 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_197
timestamp 1636986456
transform 1 0 19228 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_209
timestamp 1636986456
transform 1 0 20332 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_221
timestamp 1636986456
transform 1 0 21436 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_233
timestamp 1636986456
transform 1 0 22540 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_245
timestamp 18001
transform 1 0 23644 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_251
timestamp 18001
transform 1 0 24196 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_253
timestamp 1636986456
transform 1 0 24380 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_265
timestamp 1636986456
transform 1 0 25484 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_277
timestamp 1636986456
transform 1 0 26588 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_289
timestamp 1636986456
transform 1 0 27692 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_301
timestamp 18001
transform 1 0 28796 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_307
timestamp 18001
transform 1 0 29348 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_309
timestamp 1636986456
transform 1 0 29532 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_321
timestamp 1636986456
transform 1 0 30636 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_333
timestamp 1636986456
transform 1 0 31740 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_345
timestamp 1636986456
transform 1 0 32844 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_357
timestamp 18001
transform 1 0 33948 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_363
timestamp 18001
transform 1 0 34500 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_365
timestamp 1636986456
transform 1 0 34684 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_377
timestamp 1636986456
transform 1 0 35788 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_389
timestamp 1636986456
transform 1 0 36892 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_401
timestamp 1636986456
transform 1 0 37996 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_413
timestamp 18001
transform 1 0 39100 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_419
timestamp 18001
transform 1 0 39652 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_421
timestamp 1636986456
transform 1 0 39836 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_433
timestamp 1636986456
transform 1 0 40940 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_445
timestamp 1636986456
transform 1 0 42044 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_457
timestamp 1636986456
transform 1 0 43148 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_469
timestamp 18001
transform 1 0 44252 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_475
timestamp 18001
transform 1 0 44804 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_477
timestamp 1636986456
transform 1 0 44988 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_489
timestamp 1636986456
transform 1 0 46092 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_501
timestamp 1636986456
transform 1 0 47196 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_513
timestamp 1636986456
transform 1 0 48300 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_525
timestamp 18001
transform 1 0 49404 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_531
timestamp 18001
transform 1 0 49956 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_533
timestamp 1636986456
transform 1 0 50140 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_545
timestamp 1636986456
transform 1 0 51244 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_557
timestamp 1636986456
transform 1 0 52348 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_569
timestamp 1636986456
transform 1 0 53452 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_581
timestamp 18001
transform 1 0 54556 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_587
timestamp 18001
transform 1 0 55108 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_589
timestamp 1636986456
transform 1 0 55292 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_601
timestamp 1636986456
transform 1 0 56396 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_613
timestamp 1636986456
transform 1 0 57500 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_625
timestamp 1636986456
transform 1 0 58604 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_637
timestamp 18001
transform 1 0 59708 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_643
timestamp 18001
transform 1 0 60260 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_645
timestamp 1636986456
transform 1 0 60444 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_657
timestamp 1636986456
transform 1 0 61548 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_669
timestamp 1636986456
transform 1 0 62652 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_681
timestamp 1636986456
transform 1 0 63756 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_693
timestamp 18001
transform 1 0 64860 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_699
timestamp 18001
transform 1 0 65412 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_701
timestamp 1636986456
transform 1 0 65596 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_713
timestamp 1636986456
transform 1 0 66700 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_725
timestamp 1636986456
transform 1 0 67804 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_737
timestamp 1636986456
transform 1 0 68908 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_749
timestamp 18001
transform 1 0 70012 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_755
timestamp 18001
transform 1 0 70564 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_757
timestamp 1636986456
transform 1 0 70748 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_769
timestamp 1636986456
transform 1 0 71852 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_781
timestamp 1636986456
transform 1 0 72956 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_793
timestamp 1636986456
transform 1 0 74060 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_805
timestamp 18001
transform 1 0 75164 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_811
timestamp 18001
transform 1 0 75716 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_813
timestamp 1636986456
transform 1 0 75900 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_825
timestamp 1636986456
transform 1 0 77004 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_837
timestamp 1636986456
transform 1 0 78108 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_849
timestamp 1636986456
transform 1 0 79212 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_861
timestamp 18001
transform 1 0 80316 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_867
timestamp 18001
transform 1 0 80868 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_869
timestamp 1636986456
transform 1 0 81052 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_881
timestamp 1636986456
transform 1 0 82156 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_893
timestamp 1636986456
transform 1 0 83260 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_905
timestamp 1636986456
transform 1 0 84364 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_917
timestamp 18001
transform 1 0 85468 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_923
timestamp 18001
transform 1 0 86020 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_925
timestamp 1636986456
transform 1 0 86204 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_168_937
timestamp 18001
transform 1 0 87308 0 1 93568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_168_941
timestamp 18001
transform 1 0 87676 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_168_946
timestamp 18001
transform 1 0 88136 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_3
timestamp 1636986456
transform 1 0 1380 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_15
timestamp 1636986456
transform 1 0 2484 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_27
timestamp 1636986456
transform 1 0 3588 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_39
timestamp 1636986456
transform 1 0 4692 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_169_51
timestamp 18001
transform 1 0 5796 0 -1 94656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_169_55
timestamp 18001
transform 1 0 6164 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_57
timestamp 1636986456
transform 1 0 6348 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_69
timestamp 1636986456
transform 1 0 7452 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_81
timestamp 1636986456
transform 1 0 8556 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_93
timestamp 1636986456
transform 1 0 9660 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_105
timestamp 18001
transform 1 0 10764 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_111
timestamp 18001
transform 1 0 11316 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_113
timestamp 1636986456
transform 1 0 11500 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_125
timestamp 1636986456
transform 1 0 12604 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_137
timestamp 1636986456
transform 1 0 13708 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_149
timestamp 1636986456
transform 1 0 14812 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_161
timestamp 18001
transform 1 0 15916 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_167
timestamp 18001
transform 1 0 16468 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_169
timestamp 1636986456
transform 1 0 16652 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_181
timestamp 1636986456
transform 1 0 17756 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_193
timestamp 1636986456
transform 1 0 18860 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_205
timestamp 1636986456
transform 1 0 19964 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_217
timestamp 18001
transform 1 0 21068 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_223
timestamp 18001
transform 1 0 21620 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_225
timestamp 1636986456
transform 1 0 21804 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_237
timestamp 1636986456
transform 1 0 22908 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_249
timestamp 1636986456
transform 1 0 24012 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_261
timestamp 1636986456
transform 1 0 25116 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_273
timestamp 18001
transform 1 0 26220 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_279
timestamp 18001
transform 1 0 26772 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_281
timestamp 1636986456
transform 1 0 26956 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_293
timestamp 1636986456
transform 1 0 28060 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_305
timestamp 1636986456
transform 1 0 29164 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_317
timestamp 1636986456
transform 1 0 30268 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_329
timestamp 18001
transform 1 0 31372 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_335
timestamp 18001
transform 1 0 31924 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_337
timestamp 1636986456
transform 1 0 32108 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_349
timestamp 1636986456
transform 1 0 33212 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_361
timestamp 1636986456
transform 1 0 34316 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_373
timestamp 1636986456
transform 1 0 35420 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_385
timestamp 18001
transform 1 0 36524 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_391
timestamp 18001
transform 1 0 37076 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_393
timestamp 1636986456
transform 1 0 37260 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_405
timestamp 1636986456
transform 1 0 38364 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_417
timestamp 1636986456
transform 1 0 39468 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_429
timestamp 1636986456
transform 1 0 40572 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_441
timestamp 18001
transform 1 0 41676 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_447
timestamp 18001
transform 1 0 42228 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_449
timestamp 1636986456
transform 1 0 42412 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_461
timestamp 1636986456
transform 1 0 43516 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_473
timestamp 1636986456
transform 1 0 44620 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_485
timestamp 1636986456
transform 1 0 45724 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_497
timestamp 18001
transform 1 0 46828 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_503
timestamp 18001
transform 1 0 47380 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_505
timestamp 1636986456
transform 1 0 47564 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_517
timestamp 1636986456
transform 1 0 48668 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_529
timestamp 1636986456
transform 1 0 49772 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_541
timestamp 1636986456
transform 1 0 50876 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_553
timestamp 18001
transform 1 0 51980 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_559
timestamp 18001
transform 1 0 52532 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_561
timestamp 1636986456
transform 1 0 52716 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_573
timestamp 1636986456
transform 1 0 53820 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_585
timestamp 1636986456
transform 1 0 54924 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_597
timestamp 1636986456
transform 1 0 56028 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_609
timestamp 18001
transform 1 0 57132 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_615
timestamp 18001
transform 1 0 57684 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_617
timestamp 1636986456
transform 1 0 57868 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_629
timestamp 1636986456
transform 1 0 58972 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_641
timestamp 1636986456
transform 1 0 60076 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_653
timestamp 1636986456
transform 1 0 61180 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_665
timestamp 18001
transform 1 0 62284 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_671
timestamp 18001
transform 1 0 62836 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_673
timestamp 1636986456
transform 1 0 63020 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_685
timestamp 1636986456
transform 1 0 64124 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_697
timestamp 1636986456
transform 1 0 65228 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_709
timestamp 1636986456
transform 1 0 66332 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_721
timestamp 18001
transform 1 0 67436 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_727
timestamp 18001
transform 1 0 67988 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_729
timestamp 1636986456
transform 1 0 68172 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_741
timestamp 1636986456
transform 1 0 69276 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_753
timestamp 1636986456
transform 1 0 70380 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_765
timestamp 1636986456
transform 1 0 71484 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_777
timestamp 18001
transform 1 0 72588 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_783
timestamp 18001
transform 1 0 73140 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_785
timestamp 1636986456
transform 1 0 73324 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_797
timestamp 1636986456
transform 1 0 74428 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_809
timestamp 1636986456
transform 1 0 75532 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_821
timestamp 1636986456
transform 1 0 76636 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_833
timestamp 18001
transform 1 0 77740 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_839
timestamp 18001
transform 1 0 78292 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_841
timestamp 1636986456
transform 1 0 78476 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_853
timestamp 1636986456
transform 1 0 79580 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_865
timestamp 1636986456
transform 1 0 80684 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_877
timestamp 1636986456
transform 1 0 81788 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_889
timestamp 18001
transform 1 0 82892 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_895
timestamp 18001
transform 1 0 83444 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_897
timestamp 1636986456
transform 1 0 83628 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_909
timestamp 1636986456
transform 1 0 84732 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_921
timestamp 1636986456
transform 1 0 85836 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_933
timestamp 1636986456
transform 1 0 86940 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_169_945
timestamp 18001
transform 1 0 88044 0 -1 94656
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_170_3
timestamp 1636986456
transform 1 0 1380 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_15
timestamp 1636986456
transform 1 0 2484 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_170_27
timestamp 18001
transform 1 0 3588 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_29
timestamp 1636986456
transform 1 0 3772 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_41
timestamp 1636986456
transform 1 0 4876 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_53
timestamp 1636986456
transform 1 0 5980 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_65
timestamp 1636986456
transform 1 0 7084 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_77
timestamp 18001
transform 1 0 8188 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_83
timestamp 18001
transform 1 0 8740 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_85
timestamp 1636986456
transform 1 0 8924 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_97
timestamp 1636986456
transform 1 0 10028 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_109
timestamp 1636986456
transform 1 0 11132 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_121
timestamp 1636986456
transform 1 0 12236 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_133
timestamp 18001
transform 1 0 13340 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_139
timestamp 18001
transform 1 0 13892 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_141
timestamp 1636986456
transform 1 0 14076 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_153
timestamp 1636986456
transform 1 0 15180 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_165
timestamp 1636986456
transform 1 0 16284 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_177
timestamp 1636986456
transform 1 0 17388 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_189
timestamp 18001
transform 1 0 18492 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_195
timestamp 18001
transform 1 0 19044 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_197
timestamp 1636986456
transform 1 0 19228 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_209
timestamp 1636986456
transform 1 0 20332 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_221
timestamp 1636986456
transform 1 0 21436 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_233
timestamp 1636986456
transform 1 0 22540 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_245
timestamp 18001
transform 1 0 23644 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_251
timestamp 18001
transform 1 0 24196 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_253
timestamp 1636986456
transform 1 0 24380 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_265
timestamp 1636986456
transform 1 0 25484 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_277
timestamp 1636986456
transform 1 0 26588 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_289
timestamp 1636986456
transform 1 0 27692 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_301
timestamp 18001
transform 1 0 28796 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_307
timestamp 18001
transform 1 0 29348 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_309
timestamp 1636986456
transform 1 0 29532 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_321
timestamp 1636986456
transform 1 0 30636 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_333
timestamp 1636986456
transform 1 0 31740 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_345
timestamp 1636986456
transform 1 0 32844 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_357
timestamp 18001
transform 1 0 33948 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_363
timestamp 18001
transform 1 0 34500 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_365
timestamp 1636986456
transform 1 0 34684 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_377
timestamp 1636986456
transform 1 0 35788 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_389
timestamp 1636986456
transform 1 0 36892 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_401
timestamp 1636986456
transform 1 0 37996 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_413
timestamp 18001
transform 1 0 39100 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_419
timestamp 18001
transform 1 0 39652 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_421
timestamp 1636986456
transform 1 0 39836 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_433
timestamp 1636986456
transform 1 0 40940 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_445
timestamp 1636986456
transform 1 0 42044 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_457
timestamp 1636986456
transform 1 0 43148 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_469
timestamp 18001
transform 1 0 44252 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_475
timestamp 18001
transform 1 0 44804 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_477
timestamp 1636986456
transform 1 0 44988 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_489
timestamp 1636986456
transform 1 0 46092 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_501
timestamp 1636986456
transform 1 0 47196 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_513
timestamp 1636986456
transform 1 0 48300 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_525
timestamp 18001
transform 1 0 49404 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_531
timestamp 18001
transform 1 0 49956 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_533
timestamp 1636986456
transform 1 0 50140 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_545
timestamp 1636986456
transform 1 0 51244 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_170_557
timestamp 18001
transform 1 0 52348 0 1 94656
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_170_561
timestamp 1636986456
transform 1 0 52716 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_573
timestamp 1636986456
transform 1 0 53820 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_170_585
timestamp 18001
transform 1 0 54924 0 1 94656
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_170_589
timestamp 1636986456
transform 1 0 55292 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_601
timestamp 1636986456
transform 1 0 56396 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_613
timestamp 1636986456
transform 1 0 57500 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_625
timestamp 1636986456
transform 1 0 58604 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_637
timestamp 18001
transform 1 0 59708 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_643
timestamp 18001
transform 1 0 60260 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_645
timestamp 1636986456
transform 1 0 60444 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_657
timestamp 1636986456
transform 1 0 61548 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_669
timestamp 1636986456
transform 1 0 62652 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_681
timestamp 1636986456
transform 1 0 63756 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_693
timestamp 18001
transform 1 0 64860 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_699
timestamp 18001
transform 1 0 65412 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_701
timestamp 1636986456
transform 1 0 65596 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_713
timestamp 1636986456
transform 1 0 66700 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_725
timestamp 1636986456
transform 1 0 67804 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_737
timestamp 1636986456
transform 1 0 68908 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_749
timestamp 18001
transform 1 0 70012 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_755
timestamp 18001
transform 1 0 70564 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_757
timestamp 1636986456
transform 1 0 70748 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_769
timestamp 1636986456
transform 1 0 71852 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_781
timestamp 1636986456
transform 1 0 72956 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_793
timestamp 1636986456
transform 1 0 74060 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_805
timestamp 18001
transform 1 0 75164 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_811
timestamp 18001
transform 1 0 75716 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_813
timestamp 1636986456
transform 1 0 75900 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_825
timestamp 1636986456
transform 1 0 77004 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_837
timestamp 1636986456
transform 1 0 78108 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_849
timestamp 1636986456
transform 1 0 79212 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_861
timestamp 18001
transform 1 0 80316 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_867
timestamp 18001
transform 1 0 80868 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_869
timestamp 1636986456
transform 1 0 81052 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_881
timestamp 1636986456
transform 1 0 82156 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_893
timestamp 1636986456
transform 1 0 83260 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_905
timestamp 1636986456
transform 1 0 84364 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_917
timestamp 18001
transform 1 0 85468 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_923
timestamp 18001
transform 1 0 86020 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_925
timestamp 1636986456
transform 1 0 86204 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_937
timestamp 1636986456
transform 1 0 87308 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_170_949
timestamp 18001
transform 1 0 88412 0 1 94656
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_171_3
timestamp 1636986456
transform 1 0 1380 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_15
timestamp 1636986456
transform 1 0 2484 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_171_27
timestamp 18001
transform 1 0 3588 0 -1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_171_29
timestamp 1636986456
transform 1 0 3772 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_41
timestamp 1636986456
transform 1 0 4876 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_171_53
timestamp 18001
transform 1 0 5980 0 -1 95744
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_171_57
timestamp 1636986456
transform 1 0 6348 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_171_69
timestamp 18001
transform 1 0 7452 0 -1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_171_77
timestamp 18001
transform 1 0 8188 0 -1 95744
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_171_85
timestamp 1636986456
transform 1 0 8924 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_97
timestamp 1636986456
transform 1 0 10028 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_171_109
timestamp 18001
transform 1 0 11132 0 -1 95744
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_171_113
timestamp 1636986456
transform 1 0 11500 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_125
timestamp 1636986456
transform 1 0 12604 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_171_137
timestamp 18001
transform 1 0 13708 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_171_141
timestamp 18001
transform 1 0 14076 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_147
timestamp 18001
transform 1 0 14628 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_171_156
timestamp 18001
transform 1 0 15456 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_171_163
timestamp 18001
transform 1 0 16100 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_171_167
timestamp 18001
transform 1 0 16468 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_171_175
timestamp 18001
transform 1 0 17204 0 -1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_171_189
timestamp 18001
transform 1 0 18492 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_195
timestamp 18001
transform 1 0 19044 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_171_205
timestamp 18001
transform 1 0 19964 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_171_212
timestamp 18001
transform 1 0 20608 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_171_225
timestamp 18001
transform 1 0 21804 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_231
timestamp 18001
transform 1 0 22356 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_171_238
timestamp 18001
transform 1 0 23000 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_171_251
timestamp 18001
transform 1 0 24196 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_171_259
timestamp 18001
transform 1 0 24932 0 -1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_171_273
timestamp 18001
transform 1 0 26220 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_279
timestamp 18001
transform 1 0 26772 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_171_287
timestamp 18001
transform 1 0 27508 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_171_293
timestamp 18001
transform 1 0 28060 0 -1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_171_301
timestamp 18001
transform 1 0 28796 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_171_307
timestamp 18001
transform 1 0 29348 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_171_309
timestamp 18001
transform 1 0 29532 0 -1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_171_317
timestamp 18001
transform 1 0 30268 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_171_322
timestamp 18001
transform 1 0 30728 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_171_329
timestamp 18001
transform 1 0 31372 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_335
timestamp 18001
transform 1 0 31924 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_171_337
timestamp 18001
transform 1 0 32108 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_171_343
timestamp 18001
transform 1 0 32660 0 -1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_171_351
timestamp 18001
transform 1 0 33396 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_171_357
timestamp 18001
transform 1 0 33948 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_363
timestamp 18001
transform 1 0 34500 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_171_365
timestamp 18001
transform 1 0 34684 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_171_371
timestamp 18001
transform 1 0 35236 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_171_378
timestamp 18001
transform 1 0 35880 0 -1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_171_386
timestamp 18001
transform 1 0 36616 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_171_393
timestamp 18001
transform 1 0 37260 0 -1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_171_401
timestamp 18001
transform 1 0 37996 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_171_406
timestamp 18001
transform 1 0 38456 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_171_413
timestamp 18001
transform 1 0 39100 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_419
timestamp 18001
transform 1 0 39652 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_171_421
timestamp 18001
transform 1 0 39836 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_171_427
timestamp 18001
transform 1 0 40388 0 -1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_171_435
timestamp 18001
transform 1 0 41124 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_171_441
timestamp 18001
transform 1 0 41676 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_447
timestamp 18001
transform 1 0 42228 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_171_449
timestamp 18001
transform 1 0 42412 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_171_455
timestamp 18001
transform 1 0 42964 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_171_462
timestamp 18001
transform 1 0 43608 0 -1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_171_470
timestamp 18001
transform 1 0 44344 0 -1 95744
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_171_477
timestamp 1636986456
transform 1 0 44988 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_489
timestamp 1636986456
transform 1 0 46092 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_171_501
timestamp 18001
transform 1 0 47196 0 -1 95744
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_171_505
timestamp 1636986456
transform 1 0 47564 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_517
timestamp 1636986456
transform 1 0 48668 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_171_529
timestamp 18001
transform 1 0 49772 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_171_533
timestamp 18001
transform 1 0 50140 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_539
timestamp 18001
transform 1 0 50692 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_171_579
timestamp 18001
transform 1 0 54372 0 -1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_171_587
timestamp 18001
transform 1 0 55108 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_171_597
timestamp 18001
transform 1 0 56028 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_171_604
timestamp 18001
transform 1 0 56672 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_171_611
timestamp 18001
transform 1 0 57316 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_171_615
timestamp 18001
transform 1 0 57684 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_171_623
timestamp 18001
transform 1 0 58420 0 -1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_171_639
timestamp 18001
transform 1 0 59892 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_171_647
timestamp 18001
transform 1 0 60628 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_171_651
timestamp 18001
transform 1 0 60996 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_171_658
timestamp 18001
transform 1 0 61640 0 -1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_171_673
timestamp 18001
transform 1 0 63020 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_679
timestamp 18001
transform 1 0 63572 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_171_698
timestamp 18001
transform 1 0 65320 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_171_707
timestamp 18001
transform 1 0 66148 0 -1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_171_721
timestamp 18001
transform 1 0 67436 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_171_727
timestamp 18001
transform 1 0 67988 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_171_729
timestamp 18001
transform 1 0 68172 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_735
timestamp 18001
transform 1 0 68724 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_171_741
timestamp 18001
transform 1 0 69276 0 -1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_171_749
timestamp 18001
transform 1 0 70012 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_171_757
timestamp 18001
transform 1 0 70748 0 -1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_171_765
timestamp 18001
transform 1 0 71484 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_171_770
timestamp 18001
transform 1 0 71944 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_171_777
timestamp 18001
transform 1 0 72588 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_783
timestamp 18001
transform 1 0 73140 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_171_785
timestamp 18001
transform 1 0 73324 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_171_791
timestamp 18001
transform 1 0 73876 0 -1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_171_799
timestamp 18001
transform 1 0 74612 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_171_805
timestamp 18001
transform 1 0 75164 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_171_813
timestamp 18001
transform 1 0 75900 0 -1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_171_821
timestamp 18001
transform 1 0 76636 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_171_826
timestamp 18001
transform 1 0 77096 0 -1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_171_834
timestamp 18001
transform 1 0 77832 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_171_841
timestamp 18001
transform 1 0 78476 0 -1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_171_849
timestamp 18001
transform 1 0 79212 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_171_854
timestamp 18001
transform 1 0 79672 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_171_861
timestamp 18001
transform 1 0 80316 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_867
timestamp 18001
transform 1 0 80868 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_171_869
timestamp 18001
transform 1 0 81052 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_171_875
timestamp 18001
transform 1 0 81604 0 -1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_171_883
timestamp 18001
transform 1 0 82340 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_171_889
timestamp 18001
transform 1 0 82892 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_895
timestamp 18001
transform 1 0 83444 0 -1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_171_897
timestamp 1636986456
transform 1 0 83628 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_909
timestamp 1636986456
transform 1 0 84732 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_171_921
timestamp 18001
transform 1 0 85836 0 -1 95744
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_171_925
timestamp 1636986456
transform 1 0 86204 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_937
timestamp 1636986456
transform 1 0 87308 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_171_949
timestamp 18001
transform 1 0 88412 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  fpga_234
timestamp 18001
transform -1 0 1656 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_235
timestamp 18001
transform -1 0 1656 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_236
timestamp 18001
transform -1 0 1656 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_237
timestamp 18001
transform -1 0 1656 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_238
timestamp 18001
transform -1 0 1656 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_239
timestamp 18001
transform -1 0 1656 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_240
timestamp 18001
transform -1 0 1656 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_241
timestamp 18001
transform -1 0 1656 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_242
timestamp 18001
transform -1 0 1656 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_243
timestamp 18001
transform -1 0 1656 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_244
timestamp 18001
transform -1 0 1656 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_245
timestamp 18001
transform -1 0 1656 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_246
timestamp 18001
transform -1 0 1656 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_247
timestamp 18001
transform -1 0 1656 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_248
timestamp 18001
transform -1 0 1656 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_249
timestamp 18001
transform -1 0 1656 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input1
timestamp 18001
transform 1 0 1380 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__buf_12  input2
timestamp 18001
transform 1 0 52716 0 -1 95744
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 18001
transform -1 0 5704 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 18001
transform 1 0 5336 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 18001
transform -1 0 5704 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input6
timestamp 18001
transform -1 0 5704 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 18001
transform 1 0 5336 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 18001
transform -1 0 5704 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 18001
transform -1 0 5704 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 18001
transform 1 0 87584 0 -1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input11
timestamp 18001
transform 1 0 87952 0 1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 18001
transform 1 0 5428 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 18001
transform -1 0 87584 0 -1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 18001
transform -1 0 87952 0 1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 18001
transform -1 0 87308 0 -1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 18001
transform -1 0 88596 0 1 91392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 18001
transform -1 0 86756 0 1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp 18001
transform -1 0 88228 0 1 91392
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 18001
transform -1 0 88596 0 -1 92480
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 18001
transform -1 0 87860 0 1 91392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input21
timestamp 18001
transform -1 0 88228 0 -1 92480
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input22
timestamp 18001
transform -1 0 87492 0 1 91392
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 18001
transform 1 0 5428 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input24
timestamp 18001
transform -1 0 5704 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input25
timestamp 18001
transform -1 0 5704 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input26
timestamp 18001
transform 1 0 5428 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input27
timestamp 18001
transform 1 0 5428 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input28
timestamp 18001
transform -1 0 5704 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input29
timestamp 18001
transform -1 0 5704 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input30
timestamp 18001
transform 1 0 5336 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input31
timestamp 18001
transform 1 0 14904 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 18001
transform -1 0 26220 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input33
timestamp 18001
transform -1 0 27508 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input34
timestamp 18001
transform 1 0 27784 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input35
timestamp 18001
transform -1 0 29348 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input36
timestamp 18001
transform -1 0 55844 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input37
timestamp 18001
transform -1 0 56488 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input38
timestamp 18001
transform -1 0 57132 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input39
timestamp 18001
transform 1 0 58052 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input40
timestamp 18001
transform 1 0 15548 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input41
timestamp 18001
transform 1 0 59340 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input42
timestamp 18001
transform 1 0 59984 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input43
timestamp 18001
transform 1 0 61272 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp 18001
transform -1 0 62928 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input45
timestamp 18001
transform 1 0 63848 0 -1 95744
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input46
timestamp 18001
transform -1 0 65136 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input47
timestamp 18001
transform -1 0 66148 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input48
timestamp 18001
transform -1 0 67436 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input49
timestamp 18001
transform 1 0 67712 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input50
timestamp 18001
transform -1 0 69276 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input51
timestamp 18001
transform 1 0 16836 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input52
timestamp 18001
transform 1 0 18124 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input53
timestamp 18001
transform 1 0 19412 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input54
timestamp 18001
transform -1 0 20424 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input55
timestamp 18001
transform 1 0 21344 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input56
timestamp 18001
transform -1 0 23000 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input57
timestamp 18001
transform 1 0 23276 0 -1 95744
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input58
timestamp 18001
transform 1 0 24564 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 18001
transform 1 0 31004 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input60
timestamp 18001
transform -1 0 42320 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input61
timestamp 18001
transform 1 0 42596 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input62
timestamp 18001
transform -1 0 44252 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input63
timestamp 18001
transform -1 0 45448 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 18001
transform 1 0 70932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 18001
transform -1 0 71852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input66
timestamp 18001
transform -1 0 73140 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input67
timestamp 18001
transform -1 0 74428 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 18001
transform -1 0 31924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input69
timestamp 18001
transform -1 0 75716 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input70
timestamp 18001
transform 1 0 76084 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input71
timestamp 18001
transform -1 0 77648 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input72
timestamp 18001
transform 1 0 78660 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input73
timestamp 18001
transform -1 0 79948 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input74
timestamp 18001
transform -1 0 80960 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input75
timestamp 18001
transform -1 0 82248 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input76
timestamp 18001
transform -1 0 83536 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input77
timestamp 18001
transform -1 0 87124 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input78
timestamp 18001
transform -1 0 86112 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input79
timestamp 18001
transform -1 0 33212 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input80
timestamp 18001
transform -1 0 34500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input81
timestamp 18001
transform 1 0 34868 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input82
timestamp 18001
transform -1 0 36432 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input83
timestamp 18001
transform -1 0 37720 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input84
timestamp 18001
transform 1 0 38732 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input85
timestamp 18001
transform -1 0 40204 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input86
timestamp 18001
transform -1 0 41032 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input87
timestamp 18001
transform 1 0 7820 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input88
timestamp 18001
transform 1 0 1380 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input89
timestamp 18001
transform 1 0 1380 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input90
timestamp 18001
transform 1 0 1380 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input91
timestamp 18001
transform 1 0 1380 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input92
timestamp 18001
transform 1 0 1380 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input93
timestamp 18001
transform 1 0 1380 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input94
timestamp 18001
transform 1 0 1380 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input95
timestamp 18001
transform 1 0 1380 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input96
timestamp 18001
transform -1 0 8740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input97
timestamp 18001
transform 1 0 1380 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input98
timestamp 18001
transform 1 0 1380 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input99
timestamp 18001
transform 1 0 1380 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input100
timestamp 18001
transform 1 0 1380 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input101
timestamp 18001
transform 1 0 1380 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input102
timestamp 18001
transform 1 0 1380 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input103
timestamp 18001
transform 1 0 1380 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input104
timestamp 18001
transform 1 0 1380 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input105
timestamp 18001
transform 1 0 1380 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input106
timestamp 18001
transform 1 0 1380 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input107
timestamp 18001
transform 1 0 1380 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input108
timestamp 18001
transform 1 0 1380 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input109
timestamp 18001
transform 1 0 1380 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input110
timestamp 18001
transform 1 0 1380 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input111
timestamp 18001
transform 1 0 1380 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input112
timestamp 18001
transform 1 0 1380 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input113
timestamp 18001
transform 1 0 1380 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input114
timestamp 18001
transform 1 0 1380 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  input115
timestamp 18001
transform -1 0 11408 0 1 2176
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  input116
timestamp 18001
transform 1 0 12328 0 1 2176
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  input117
timestamp 18001
transform 1 0 14076 0 1 2176
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_12  input118
timestamp 18001
transform 1 0 50968 0 -1 95744
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  max_cap232
timestamp 18001
transform 1 0 52716 0 1 91392
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  max_cap233
timestamp 18001
transform 1 0 51152 0 1 91392
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  output119
timestamp 18001
transform 1 0 5336 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output120
timestamp 18001
transform 1 0 86388 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output121
timestamp 18001
transform 1 0 87860 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output122
timestamp 18001
transform 1 0 88228 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp 18001
transform 1 0 5336 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output124
timestamp 18001
transform 1 0 5336 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output125
timestamp 18001
transform 1 0 5336 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output126
timestamp 18001
transform 1 0 5336 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output127
timestamp 18001
transform 1 0 5336 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output128
timestamp 18001
transform 1 0 5336 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output129
timestamp 18001
transform 1 0 87124 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output130
timestamp 18001
transform 1 0 5336 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output131
timestamp 18001
transform 1 0 5336 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output132
timestamp 18001
transform 1 0 5336 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output133
timestamp 18001
transform 1 0 5336 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output134
timestamp 18001
transform 1 0 5336 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output135
timestamp 18001
transform 1 0 5336 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output136
timestamp 18001
transform 1 0 5336 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output137
timestamp 18001
transform 1 0 5336 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output138
timestamp 18001
transform 1 0 5336 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp 18001
transform 1 0 5336 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output140
timestamp 18001
transform 1 0 87860 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output141
timestamp 18001
transform 1 0 87492 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output142
timestamp 18001
transform 1 0 88228 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output143
timestamp 18001
transform 1 0 86756 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output144
timestamp 18001
transform 1 0 87124 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output145
timestamp 18001
transform 1 0 87860 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output146
timestamp 18001
transform 1 0 87492 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output147
timestamp 18001
transform 1 0 88228 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output148
timestamp 18001
transform 1 0 30360 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output149
timestamp 18001
transform 1 0 41308 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output150
timestamp 18001
transform 1 0 42596 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output151
timestamp 18001
transform -1 0 43608 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output152
timestamp 18001
transform 1 0 44528 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output153
timestamp 18001
transform 1 0 70288 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output154
timestamp 18001
transform 1 0 71576 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output155
timestamp 18001
transform 1 0 72220 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output156
timestamp 18001
transform 1 0 73508 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output157
timestamp 18001
transform -1 0 31372 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output158
timestamp 18001
transform 1 0 74796 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output159
timestamp 18001
transform -1 0 75808 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output160
timestamp 18001
transform 1 0 76728 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output161
timestamp 18001
transform 1 0 78016 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output162
timestamp 18001
transform 1 0 79304 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output163
timestamp 18001
transform 1 0 79948 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output164
timestamp 18001
transform 1 0 81236 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output165
timestamp 18001
transform 1 0 82524 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output166
timestamp 18001
transform 1 0 88228 0 1 92480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output167
timestamp 18001
transform 1 0 86756 0 1 91392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output168
timestamp 18001
transform 1 0 32292 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output169
timestamp 18001
transform 1 0 33580 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output170
timestamp 18001
transform 1 0 34868 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output171
timestamp 18001
transform -1 0 35880 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output172
timestamp 18001
transform 1 0 36800 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output173
timestamp 18001
transform 1 0 38088 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output174
timestamp 18001
transform -1 0 39100 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output175
timestamp 18001
transform 1 0 40020 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output176
timestamp 18001
transform 1 0 15548 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output177
timestamp 18001
transform 1 0 26496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output178
timestamp 18001
transform -1 0 27508 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output179
timestamp 18001
transform 1 0 28428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output180
timestamp 18001
transform 1 0 29716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output181
timestamp 18001
transform 1 0 55476 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output182
timestamp 18001
transform -1 0 56488 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output183
timestamp 18001
transform 1 0 57408 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output184
timestamp 18001
transform 1 0 58696 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output185
timestamp 18001
transform -1 0 16560 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output186
timestamp 18001
transform 1 0 59984 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output187
timestamp 18001
transform 1 0 60628 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output188
timestamp 18001
transform 1 0 61916 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output189
timestamp 18001
transform 1 0 63204 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output190
timestamp 18001
transform -1 0 64216 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output191
timestamp 18001
transform 1 0 65136 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output192
timestamp 18001
transform 1 0 66424 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output193
timestamp 18001
transform 1 0 67712 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output194
timestamp 18001
transform 1 0 68356 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output195
timestamp 18001
transform 1 0 69644 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output196
timestamp 18001
transform 1 0 17480 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output197
timestamp 18001
transform 1 0 18768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output198
timestamp 18001
transform -1 0 19780 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output199
timestamp 18001
transform 1 0 20700 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output200
timestamp 18001
transform 1 0 21988 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output201
timestamp 18001
transform 1 0 23276 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output202
timestamp 18001
transform -1 0 24288 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output203
timestamp 18001
transform 1 0 25208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output204
timestamp 18001
transform -1 0 1748 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output205
timestamp 18001
transform -1 0 1748 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output206
timestamp 18001
transform -1 0 1748 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output207
timestamp 18001
transform -1 0 1748 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output208
timestamp 18001
transform -1 0 1748 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output209
timestamp 18001
transform -1 0 1748 0 -1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output210
timestamp 18001
transform -1 0 1748 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output211
timestamp 18001
transform -1 0 1748 0 1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output212
timestamp 18001
transform -1 0 1748 0 1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output213
timestamp 18001
transform -1 0 1748 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output214
timestamp 18001
transform -1 0 1748 0 -1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output215
timestamp 18001
transform -1 0 1748 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output216
timestamp 18001
transform -1 0 1748 0 1 78336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output217
timestamp 18001
transform -1 0 1748 0 1 79424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output218
timestamp 18001
transform -1 0 1748 0 -1 81600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output219
timestamp 18001
transform -1 0 1748 0 -1 82688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output220
timestamp 18001
transform -1 0 1748 0 1 83776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output221
timestamp 18001
transform -1 0 1748 0 1 84864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output222
timestamp 18001
transform -1 0 1748 0 -1 87040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output223
timestamp 18001
transform 1 0 8464 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output224
timestamp 18001
transform -1 0 1748 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output225
timestamp 18001
transform -1 0 1748 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output226
timestamp 18001
transform -1 0 1748 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output227
timestamp 18001
transform -1 0 1748 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output228
timestamp 18001
transform -1 0 1748 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output229
timestamp 18001
transform -1 0 1748 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output230
timestamp 18001
transform -1 0 1748 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output231
timestamp 18001
transform -1 0 1748 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_172
timestamp 18001
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 18001
transform -1 0 88872 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_173
timestamp 18001
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 18001
transform -1 0 88872 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_174
timestamp 18001
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 18001
transform -1 0 88872 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_175
timestamp 18001
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 18001
transform -1 0 88872 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_176
timestamp 18001
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 18001
transform -1 0 88872 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_177
timestamp 18001
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 18001
transform -1 0 88872 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_178
timestamp 18001
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 18001
transform -1 0 88872 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_1_Left_343
timestamp 18001
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_1_Right_163
timestamp 18001
transform -1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_1_Left_179
timestamp 18001
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_1_Right_7
timestamp 18001
transform -1 0 5980 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_1_Left_180
timestamp 18001
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_1_Right_8
timestamp 18001
transform -1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_1_Left_181
timestamp 18001
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_1_Right_9
timestamp 18001
transform -1 0 5980 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_1_Left_182
timestamp 18001
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_1_Right_10
timestamp 18001
transform -1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_1_Left_183
timestamp 18001
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_1_Right_11
timestamp 18001
transform -1 0 5980 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_1_Left_184
timestamp 18001
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_1_Right_12
timestamp 18001
transform -1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_1_Left_185
timestamp 18001
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_1_Right_13
timestamp 18001
transform -1 0 5980 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_1_Left_186
timestamp 18001
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_1_Right_14
timestamp 18001
transform -1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_1_Left_187
timestamp 18001
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_1_Right_15
timestamp 18001
transform -1 0 5980 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_1_Left_188
timestamp 18001
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_1_Right_16
timestamp 18001
transform -1 0 5980 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_1_Left_189
timestamp 18001
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_1_Right_17
timestamp 18001
transform -1 0 5980 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_1_Left_190
timestamp 18001
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_1_Right_18
timestamp 18001
transform -1 0 5980 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_1_Left_191
timestamp 18001
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_1_Right_19
timestamp 18001
transform -1 0 5980 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_1_Left_192
timestamp 18001
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_1_Right_20
timestamp 18001
transform -1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_1_Left_193
timestamp 18001
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_1_Right_21
timestamp 18001
transform -1 0 5980 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_1_Left_194
timestamp 18001
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_1_Right_22
timestamp 18001
transform -1 0 5980 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_1_Left_195
timestamp 18001
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_1_Right_23
timestamp 18001
transform -1 0 5980 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_1_Left_196
timestamp 18001
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_1_Right_24
timestamp 18001
transform -1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_1_Left_197
timestamp 18001
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_1_Right_25
timestamp 18001
transform -1 0 5980 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_1_Left_198
timestamp 18001
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_1_Right_26
timestamp 18001
transform -1 0 5980 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_1_Left_199
timestamp 18001
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_1_Right_27
timestamp 18001
transform -1 0 5980 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_1_Left_200
timestamp 18001
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_1_Right_28
timestamp 18001
transform -1 0 5980 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_1_Left_201
timestamp 18001
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_1_Right_29
timestamp 18001
transform -1 0 5980 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_1_Left_202
timestamp 18001
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_1_Right_30
timestamp 18001
transform -1 0 5980 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_1_Left_203
timestamp 18001
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_1_Right_31
timestamp 18001
transform -1 0 5980 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_1_Left_204
timestamp 18001
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_1_Right_32
timestamp 18001
transform -1 0 5980 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_1_Left_205
timestamp 18001
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_1_Right_33
timestamp 18001
transform -1 0 5980 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_1_Left_206
timestamp 18001
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_1_Right_34
timestamp 18001
transform -1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_1_Left_207
timestamp 18001
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_1_Right_35
timestamp 18001
transform -1 0 5980 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_1_Left_208
timestamp 18001
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_1_Right_36
timestamp 18001
transform -1 0 5980 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_1_Left_209
timestamp 18001
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_1_Right_37
timestamp 18001
transform -1 0 5980 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_1_Left_210
timestamp 18001
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_1_Right_38
timestamp 18001
transform -1 0 5980 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_1_Left_211
timestamp 18001
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_1_Right_39
timestamp 18001
transform -1 0 5980 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_1_Left_212
timestamp 18001
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_1_Right_40
timestamp 18001
transform -1 0 5980 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_1_Left_213
timestamp 18001
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_1_Right_41
timestamp 18001
transform -1 0 5980 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_1_Left_214
timestamp 18001
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_1_Right_42
timestamp 18001
transform -1 0 5980 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_1_Left_215
timestamp 18001
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_1_Right_43
timestamp 18001
transform -1 0 5980 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_1_Left_216
timestamp 18001
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_1_Right_44
timestamp 18001
transform -1 0 5980 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_1_Left_217
timestamp 18001
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_1_Right_45
timestamp 18001
transform -1 0 5980 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_1_Left_218
timestamp 18001
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_1_Right_46
timestamp 18001
transform -1 0 5980 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_1_Left_219
timestamp 18001
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_1_Right_47
timestamp 18001
transform -1 0 5980 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_1_Left_220
timestamp 18001
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_1_Right_48
timestamp 18001
transform -1 0 5980 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_1_Left_221
timestamp 18001
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_1_Right_49
timestamp 18001
transform -1 0 5980 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_1_Left_222
timestamp 18001
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_1_Right_50
timestamp 18001
transform -1 0 5980 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_1_Left_223
timestamp 18001
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_1_Right_51
timestamp 18001
transform -1 0 5980 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_1_Left_224
timestamp 18001
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_1_Right_52
timestamp 18001
transform -1 0 5980 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_1_Left_225
timestamp 18001
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_1_Right_53
timestamp 18001
transform -1 0 5980 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_1_Left_226
timestamp 18001
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_1_Right_54
timestamp 18001
transform -1 0 5980 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_1_Left_227
timestamp 18001
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_1_Right_55
timestamp 18001
transform -1 0 5980 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_1_Left_228
timestamp 18001
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_1_Right_56
timestamp 18001
transform -1 0 5980 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_1_Left_229
timestamp 18001
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_1_Right_57
timestamp 18001
transform -1 0 5980 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_1_Left_230
timestamp 18001
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_1_Right_58
timestamp 18001
transform -1 0 5980 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_1_Left_231
timestamp 18001
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_1_Right_59
timestamp 18001
transform -1 0 5980 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_1_Left_232
timestamp 18001
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_1_Right_60
timestamp 18001
transform -1 0 5980 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_1_Left_233
timestamp 18001
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_1_Right_61
timestamp 18001
transform -1 0 5980 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_1_Left_234
timestamp 18001
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_1_Right_62
timestamp 18001
transform -1 0 5980 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_1_Left_235
timestamp 18001
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_1_Right_63
timestamp 18001
transform -1 0 5980 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_1_Left_236
timestamp 18001
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_1_Right_64
timestamp 18001
transform -1 0 5980 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_1_Left_237
timestamp 18001
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_1_Right_65
timestamp 18001
transform -1 0 5980 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_1_Left_238
timestamp 18001
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_1_Right_66
timestamp 18001
transform -1 0 5980 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_1_Left_239
timestamp 18001
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_1_Right_67
timestamp 18001
transform -1 0 5980 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_1_Left_240
timestamp 18001
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_1_Right_68
timestamp 18001
transform -1 0 5980 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_1_Left_241
timestamp 18001
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_1_Right_69
timestamp 18001
transform -1 0 5980 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_1_Left_242
timestamp 18001
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_1_Right_70
timestamp 18001
transform -1 0 5980 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_1_Left_243
timestamp 18001
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_1_Right_71
timestamp 18001
transform -1 0 5980 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_1_Left_244
timestamp 18001
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_1_Right_72
timestamp 18001
transform -1 0 5980 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_1_Left_245
timestamp 18001
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_1_Right_73
timestamp 18001
transform -1 0 5980 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_1_Left_246
timestamp 18001
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_1_Right_74
timestamp 18001
transform -1 0 5980 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_1_Left_247
timestamp 18001
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_1_Right_75
timestamp 18001
transform -1 0 5980 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_1_Left_248
timestamp 18001
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_1_Right_76
timestamp 18001
transform -1 0 5980 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_1_Left_249
timestamp 18001
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_1_Right_77
timestamp 18001
transform -1 0 5980 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_1_Left_250
timestamp 18001
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_1_Right_78
timestamp 18001
transform -1 0 5980 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_1_Left_251
timestamp 18001
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_1_Right_79
timestamp 18001
transform -1 0 5980 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_1_Left_252
timestamp 18001
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_1_Right_80
timestamp 18001
transform -1 0 5980 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_1_Left_253
timestamp 18001
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_1_Right_81
timestamp 18001
transform -1 0 5980 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_1_Left_254
timestamp 18001
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_1_Right_82
timestamp 18001
transform -1 0 5980 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_1_Left_255
timestamp 18001
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_1_Right_83
timestamp 18001
transform -1 0 5980 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_1_Left_256
timestamp 18001
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_1_Right_84
timestamp 18001
transform -1 0 5980 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_1_Left_257
timestamp 18001
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_1_Right_85
timestamp 18001
transform -1 0 5980 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_1_Left_258
timestamp 18001
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_1_Right_86
timestamp 18001
transform -1 0 5980 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_1_Left_259
timestamp 18001
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_1_Right_87
timestamp 18001
transform -1 0 5980 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_1_Left_260
timestamp 18001
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_1_Right_88
timestamp 18001
transform -1 0 5980 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_1_Left_261
timestamp 18001
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_1_Right_89
timestamp 18001
transform -1 0 5980 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_1_Left_262
timestamp 18001
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_1_Right_90
timestamp 18001
transform -1 0 5980 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_1_Left_263
timestamp 18001
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_1_Right_91
timestamp 18001
transform -1 0 5980 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_1_Left_264
timestamp 18001
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_1_Right_92
timestamp 18001
transform -1 0 5980 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_1_Left_265
timestamp 18001
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_1_Right_93
timestamp 18001
transform -1 0 5980 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_1_Left_266
timestamp 18001
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_1_Right_94
timestamp 18001
transform -1 0 5980 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_1_Left_267
timestamp 18001
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_1_Right_95
timestamp 18001
transform -1 0 5980 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_1_Left_268
timestamp 18001
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_1_Right_96
timestamp 18001
transform -1 0 5980 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_1_Left_269
timestamp 18001
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_1_Right_97
timestamp 18001
transform -1 0 5980 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_1_Left_270
timestamp 18001
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_1_Right_98
timestamp 18001
transform -1 0 5980 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_1_Left_271
timestamp 18001
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_1_Right_99
timestamp 18001
transform -1 0 5980 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_1_Left_272
timestamp 18001
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_1_Right_100
timestamp 18001
transform -1 0 5980 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_1_Left_273
timestamp 18001
transform 1 0 1104 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_1_Right_101
timestamp 18001
transform -1 0 5980 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_1_Left_274
timestamp 18001
transform 1 0 1104 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_1_Right_102
timestamp 18001
transform -1 0 5980 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_1_Left_275
timestamp 18001
transform 1 0 1104 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_1_Right_103
timestamp 18001
transform -1 0 5980 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_1_Left_276
timestamp 18001
transform 1 0 1104 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_1_Right_104
timestamp 18001
transform -1 0 5980 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_1_Left_277
timestamp 18001
transform 1 0 1104 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_1_Right_105
timestamp 18001
transform -1 0 5980 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_1_Left_278
timestamp 18001
transform 1 0 1104 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_1_Right_106
timestamp 18001
transform -1 0 5980 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_1_Left_279
timestamp 18001
transform 1 0 1104 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_1_Right_107
timestamp 18001
transform -1 0 5980 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_1_Left_280
timestamp 18001
transform 1 0 1104 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_1_Right_108
timestamp 18001
transform -1 0 5980 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_1_Left_281
timestamp 18001
transform 1 0 1104 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_1_Right_109
timestamp 18001
transform -1 0 5980 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_1_Left_282
timestamp 18001
transform 1 0 1104 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_1_Right_110
timestamp 18001
transform -1 0 5980 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_1_Left_283
timestamp 18001
transform 1 0 1104 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_1_Right_111
timestamp 18001
transform -1 0 5980 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_1_Left_284
timestamp 18001
transform 1 0 1104 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_1_Right_112
timestamp 18001
transform -1 0 5980 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_1_Left_285
timestamp 18001
transform 1 0 1104 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_1_Right_113
timestamp 18001
transform -1 0 5980 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_1_Left_286
timestamp 18001
transform 1 0 1104 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_1_Right_114
timestamp 18001
transform -1 0 5980 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_1_Left_287
timestamp 18001
transform 1 0 1104 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_1_Right_115
timestamp 18001
transform -1 0 5980 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_117_1_Left_288
timestamp 18001
transform 1 0 1104 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_117_1_Right_116
timestamp 18001
transform -1 0 5980 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_118_1_Left_289
timestamp 18001
transform 1 0 1104 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_118_1_Right_117
timestamp 18001
transform -1 0 5980 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_119_1_Left_290
timestamp 18001
transform 1 0 1104 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_119_1_Right_118
timestamp 18001
transform -1 0 5980 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_120_1_Left_291
timestamp 18001
transform 1 0 1104 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_120_1_Right_119
timestamp 18001
transform -1 0 5980 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_121_1_Left_292
timestamp 18001
transform 1 0 1104 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_121_1_Right_120
timestamp 18001
transform -1 0 5980 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_122_1_Left_293
timestamp 18001
transform 1 0 1104 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_122_1_Right_121
timestamp 18001
transform -1 0 5980 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_123_1_Left_294
timestamp 18001
transform 1 0 1104 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_123_1_Right_122
timestamp 18001
transform -1 0 5980 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_124_1_Left_295
timestamp 18001
transform 1 0 1104 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_124_1_Right_123
timestamp 18001
transform -1 0 5980 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_125_1_Left_296
timestamp 18001
transform 1 0 1104 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_125_1_Right_124
timestamp 18001
transform -1 0 5980 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_126_1_Left_297
timestamp 18001
transform 1 0 1104 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_126_1_Right_125
timestamp 18001
transform -1 0 5980 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_127_1_Left_298
timestamp 18001
transform 1 0 1104 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_127_1_Right_126
timestamp 18001
transform -1 0 5980 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_128_1_Left_299
timestamp 18001
transform 1 0 1104 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_128_1_Right_127
timestamp 18001
transform -1 0 5980 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_129_1_Left_300
timestamp 18001
transform 1 0 1104 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_129_1_Right_128
timestamp 18001
transform -1 0 5980 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_130_1_Left_301
timestamp 18001
transform 1 0 1104 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_130_1_Right_129
timestamp 18001
transform -1 0 5980 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_131_1_Left_302
timestamp 18001
transform 1 0 1104 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_131_1_Right_130
timestamp 18001
transform -1 0 5980 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_132_1_Left_303
timestamp 18001
transform 1 0 1104 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_132_1_Right_131
timestamp 18001
transform -1 0 5980 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_133_1_Left_304
timestamp 18001
transform 1 0 1104 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_133_1_Right_132
timestamp 18001
transform -1 0 5980 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_134_1_Left_305
timestamp 18001
transform 1 0 1104 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_134_1_Right_133
timestamp 18001
transform -1 0 5980 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_135_1_Left_306
timestamp 18001
transform 1 0 1104 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_135_1_Right_134
timestamp 18001
transform -1 0 5980 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_136_1_Left_307
timestamp 18001
transform 1 0 1104 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_136_1_Right_135
timestamp 18001
transform -1 0 5980 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_137_1_Left_308
timestamp 18001
transform 1 0 1104 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_137_1_Right_136
timestamp 18001
transform -1 0 5980 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_138_1_Left_309
timestamp 18001
transform 1 0 1104 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_138_1_Right_137
timestamp 18001
transform -1 0 5980 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_139_1_Left_310
timestamp 18001
transform 1 0 1104 0 -1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_139_1_Right_138
timestamp 18001
transform -1 0 5980 0 -1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_140_1_Left_311
timestamp 18001
transform 1 0 1104 0 1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_140_1_Right_139
timestamp 18001
transform -1 0 5980 0 1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_141_1_Left_312
timestamp 18001
transform 1 0 1104 0 -1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_141_1_Right_140
timestamp 18001
transform -1 0 5980 0 -1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_142_1_Left_313
timestamp 18001
transform 1 0 1104 0 1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_142_1_Right_141
timestamp 18001
transform -1 0 5980 0 1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_143_1_Left_314
timestamp 18001
transform 1 0 1104 0 -1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_143_1_Right_142
timestamp 18001
transform -1 0 5980 0 -1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_144_1_Left_315
timestamp 18001
transform 1 0 1104 0 1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_144_1_Right_143
timestamp 18001
transform -1 0 5980 0 1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_145_1_Left_316
timestamp 18001
transform 1 0 1104 0 -1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_145_1_Right_144
timestamp 18001
transform -1 0 5980 0 -1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_146_1_Left_317
timestamp 18001
transform 1 0 1104 0 1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_146_1_Right_145
timestamp 18001
transform -1 0 5980 0 1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_147_1_Left_318
timestamp 18001
transform 1 0 1104 0 -1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_147_1_Right_146
timestamp 18001
transform -1 0 5980 0 -1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_148_1_Left_319
timestamp 18001
transform 1 0 1104 0 1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_148_1_Right_147
timestamp 18001
transform -1 0 5980 0 1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_149_1_Left_320
timestamp 18001
transform 1 0 1104 0 -1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_149_1_Right_148
timestamp 18001
transform -1 0 5980 0 -1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_150_1_Left_321
timestamp 18001
transform 1 0 1104 0 1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_150_1_Right_149
timestamp 18001
transform -1 0 5980 0 1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_151_1_Left_322
timestamp 18001
transform 1 0 1104 0 -1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_151_1_Right_150
timestamp 18001
transform -1 0 5980 0 -1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_152_1_Left_323
timestamp 18001
transform 1 0 1104 0 1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_152_1_Right_151
timestamp 18001
transform -1 0 5980 0 1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_153_1_Left_324
timestamp 18001
transform 1 0 1104 0 -1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_153_1_Right_152
timestamp 18001
transform -1 0 5980 0 -1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_154_1_Left_325
timestamp 18001
transform 1 0 1104 0 1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_154_1_Right_153
timestamp 18001
transform -1 0 5980 0 1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_155_1_Left_326
timestamp 18001
transform 1 0 1104 0 -1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_155_1_Right_154
timestamp 18001
transform -1 0 5980 0 -1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_156_1_Left_327
timestamp 18001
transform 1 0 1104 0 1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_156_1_Right_155
timestamp 18001
transform -1 0 5980 0 1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_157_1_Left_328
timestamp 18001
transform 1 0 1104 0 -1 88128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_157_1_Right_156
timestamp 18001
transform -1 0 5980 0 -1 88128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_158_1_Left_329
timestamp 18001
transform 1 0 1104 0 1 88128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_158_1_Right_157
timestamp 18001
transform -1 0 5980 0 1 88128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_159_1_Left_330
timestamp 18001
transform 1 0 1104 0 -1 89216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_159_1_Right_158
timestamp 18001
transform -1 0 5980 0 -1 89216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_160_1_Left_331
timestamp 18001
transform 1 0 1104 0 1 89216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_160_1_Right_159
timestamp 18001
transform -1 0 5980 0 1 89216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_161_1_Left_332
timestamp 18001
transform 1 0 1104 0 -1 90304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_161_1_Right_160
timestamp 18001
transform -1 0 5980 0 -1 90304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_162_1_Left_333
timestamp 18001
transform 1 0 1104 0 1 90304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_162_1_Right_161
timestamp 18001
transform -1 0 5980 0 1 90304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_163_1_Left_334
timestamp 18001
transform 1 0 1104 0 -1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_163_1_Right_162
timestamp 18001
transform -1 0 5980 0 -1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_164_Left_335
timestamp 18001
transform 1 0 1104 0 1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_164_Right_164
timestamp 18001
transform -1 0 88872 0 1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_165_Left_336
timestamp 18001
transform 1 0 1104 0 -1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_165_Right_165
timestamp 18001
transform -1 0 88872 0 -1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_166_Left_337
timestamp 18001
transform 1 0 1104 0 1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_166_Right_166
timestamp 18001
transform -1 0 88872 0 1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_167_Left_338
timestamp 18001
transform 1 0 1104 0 -1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_167_Right_167
timestamp 18001
transform -1 0 88872 0 -1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_168_Left_339
timestamp 18001
transform 1 0 1104 0 1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_168_Right_168
timestamp 18001
transform -1 0 88872 0 1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_169_Left_340
timestamp 18001
transform 1 0 1104 0 -1 94656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_169_Right_169
timestamp 18001
transform -1 0 88872 0 -1 94656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_170_Left_341
timestamp 18001
transform 1 0 1104 0 1 94656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_170_Right_170
timestamp 18001
transform -1 0 88872 0 1 94656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_171_Left_342
timestamp 18001
transform 1 0 1104 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_171_Right_171
timestamp 18001
transform -1 0 88872 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_344
timestamp 18001
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_345
timestamp 18001
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_346
timestamp 18001
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_347
timestamp 18001
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_348
timestamp 18001
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_349
timestamp 18001
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_350
timestamp 18001
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_351
timestamp 18001
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_352
timestamp 18001
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_353
timestamp 18001
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_354
timestamp 18001
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_355
timestamp 18001
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_356
timestamp 18001
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_357
timestamp 18001
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_358
timestamp 18001
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_359
timestamp 18001
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_360
timestamp 18001
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_361
timestamp 18001
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_362
timestamp 18001
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_363
timestamp 18001
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_364
timestamp 18001
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_365
timestamp 18001
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_366
timestamp 18001
transform 1 0 60352 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_367
timestamp 18001
transform 1 0 62928 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_368
timestamp 18001
transform 1 0 65504 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_369
timestamp 18001
transform 1 0 68080 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_370
timestamp 18001
transform 1 0 70656 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_371
timestamp 18001
transform 1 0 73232 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_372
timestamp 18001
transform 1 0 75808 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_373
timestamp 18001
transform 1 0 78384 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_374
timestamp 18001
transform 1 0 80960 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_375
timestamp 18001
transform 1 0 83536 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_376
timestamp 18001
transform 1 0 86112 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_377
timestamp 18001
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_378
timestamp 18001
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_379
timestamp 18001
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_380
timestamp 18001
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_381
timestamp 18001
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_382
timestamp 18001
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_383
timestamp 18001
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_384
timestamp 18001
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_385
timestamp 18001
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_386
timestamp 18001
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_387
timestamp 18001
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_388
timestamp 18001
transform 1 0 62928 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_389
timestamp 18001
transform 1 0 68080 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_390
timestamp 18001
transform 1 0 73232 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_391
timestamp 18001
transform 1 0 78384 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_392
timestamp 18001
transform 1 0 83536 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_393
timestamp 18001
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_394
timestamp 18001
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_395
timestamp 18001
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_396
timestamp 18001
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_397
timestamp 18001
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_398
timestamp 18001
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_399
timestamp 18001
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_400
timestamp 18001
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_401
timestamp 18001
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_402
timestamp 18001
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_403
timestamp 18001
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_404
timestamp 18001
transform 1 0 60352 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_405
timestamp 18001
transform 1 0 65504 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_406
timestamp 18001
transform 1 0 70656 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_407
timestamp 18001
transform 1 0 75808 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_408
timestamp 18001
transform 1 0 80960 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_409
timestamp 18001
transform 1 0 86112 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_410
timestamp 18001
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_411
timestamp 18001
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_412
timestamp 18001
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_413
timestamp 18001
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_414
timestamp 18001
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_415
timestamp 18001
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_416
timestamp 18001
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_417
timestamp 18001
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_418
timestamp 18001
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_419
timestamp 18001
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_420
timestamp 18001
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_421
timestamp 18001
transform 1 0 62928 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_422
timestamp 18001
transform 1 0 68080 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_423
timestamp 18001
transform 1 0 73232 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_424
timestamp 18001
transform 1 0 78384 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_425
timestamp 18001
transform 1 0 83536 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_426
timestamp 18001
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_427
timestamp 18001
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_428
timestamp 18001
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_429
timestamp 18001
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_430
timestamp 18001
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_431
timestamp 18001
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_432
timestamp 18001
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_433
timestamp 18001
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_434
timestamp 18001
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_435
timestamp 18001
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_436
timestamp 18001
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_437
timestamp 18001
transform 1 0 60352 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_438
timestamp 18001
transform 1 0 65504 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_439
timestamp 18001
transform 1 0 70656 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_440
timestamp 18001
transform 1 0 75808 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_441
timestamp 18001
transform 1 0 80960 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_442
timestamp 18001
transform 1 0 86112 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_443
timestamp 18001
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_444
timestamp 18001
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_445
timestamp 18001
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_446
timestamp 18001
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_447
timestamp 18001
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_448
timestamp 18001
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_449
timestamp 18001
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_450
timestamp 18001
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_451
timestamp 18001
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_452
timestamp 18001
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_453
timestamp 18001
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_454
timestamp 18001
transform 1 0 62928 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_455
timestamp 18001
transform 1 0 68080 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_456
timestamp 18001
transform 1 0 73232 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_457
timestamp 18001
transform 1 0 78384 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_458
timestamp 18001
transform 1 0 83536 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_459
timestamp 18001
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_460
timestamp 18001
transform 1 0 6256 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_461
timestamp 18001
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_462
timestamp 18001
transform 1 0 11408 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_463
timestamp 18001
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_464
timestamp 18001
transform 1 0 16560 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_465
timestamp 18001
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_466
timestamp 18001
transform 1 0 21712 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_467
timestamp 18001
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_468
timestamp 18001
transform 1 0 26864 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_469
timestamp 18001
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_470
timestamp 18001
transform 1 0 32016 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_471
timestamp 18001
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_472
timestamp 18001
transform 1 0 37168 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_473
timestamp 18001
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_474
timestamp 18001
transform 1 0 42320 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_475
timestamp 18001
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_476
timestamp 18001
transform 1 0 47472 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_477
timestamp 18001
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_478
timestamp 18001
transform 1 0 52624 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_479
timestamp 18001
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_480
timestamp 18001
transform 1 0 57776 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_481
timestamp 18001
transform 1 0 60352 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_482
timestamp 18001
transform 1 0 62928 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_483
timestamp 18001
transform 1 0 65504 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_484
timestamp 18001
transform 1 0 68080 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_485
timestamp 18001
transform 1 0 70656 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_486
timestamp 18001
transform 1 0 73232 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_487
timestamp 18001
transform 1 0 75808 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_488
timestamp 18001
transform 1 0 78384 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_489
timestamp 18001
transform 1 0 80960 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_490
timestamp 18001
transform 1 0 83536 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_491
timestamp 18001
transform 1 0 86112 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1_492
timestamp 18001
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_1_493
timestamp 18001
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_1_494
timestamp 18001
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_1_495
timestamp 18001
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_1_496
timestamp 18001
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_1_497
timestamp 18001
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_1_498
timestamp 18001
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_1_499
timestamp 18001
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_1_500
timestamp 18001
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_1_501
timestamp 18001
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_1_502
timestamp 18001
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_1_503
timestamp 18001
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_1_504
timestamp 18001
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_1_505
timestamp 18001
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_1_506
timestamp 18001
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_1_507
timestamp 18001
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_1_508
timestamp 18001
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_1_509
timestamp 18001
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_1_510
timestamp 18001
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_1_511
timestamp 18001
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_1_512
timestamp 18001
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_1_513
timestamp 18001
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_1_514
timestamp 18001
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_1_515
timestamp 18001
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_1_516
timestamp 18001
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_1_517
timestamp 18001
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1_518
timestamp 18001
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1_519
timestamp 18001
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1_520
timestamp 18001
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_1_521
timestamp 18001
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_1_522
timestamp 18001
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_1_523
timestamp 18001
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1_524
timestamp 18001
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1_525
timestamp 18001
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1_526
timestamp 18001
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1_527
timestamp 18001
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1_528
timestamp 18001
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1_529
timestamp 18001
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1_530
timestamp 18001
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1_531
timestamp 18001
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1_532
timestamp 18001
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1_533
timestamp 18001
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1_534
timestamp 18001
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1_535
timestamp 18001
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1_536
timestamp 18001
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1_537
timestamp 18001
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1_538
timestamp 18001
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_1_539
timestamp 18001
transform 1 0 3680 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_1_540
timestamp 18001
transform 1 0 3680 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_1_541
timestamp 18001
transform 1 0 3680 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_1_542
timestamp 18001
transform 1 0 3680 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_1_543
timestamp 18001
transform 1 0 3680 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_1_544
timestamp 18001
transform 1 0 3680 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_1_545
timestamp 18001
transform 1 0 3680 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_1_546
timestamp 18001
transform 1 0 3680 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1_547
timestamp 18001
transform 1 0 3680 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1_548
timestamp 18001
transform 1 0 3680 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1_549
timestamp 18001
transform 1 0 3680 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1_550
timestamp 18001
transform 1 0 3680 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1_551
timestamp 18001
transform 1 0 3680 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1_552
timestamp 18001
transform 1 0 3680 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1_553
timestamp 18001
transform 1 0 3680 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1_554
timestamp 18001
transform 1 0 3680 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1_555
timestamp 18001
transform 1 0 3680 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1_556
timestamp 18001
transform 1 0 3680 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1_557
timestamp 18001
transform 1 0 3680 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_140_1_558
timestamp 18001
transform 1 0 3680 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_142_1_559
timestamp 18001
transform 1 0 3680 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_144_1_560
timestamp 18001
transform 1 0 3680 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_1_561
timestamp 18001
transform 1 0 3680 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_1_562
timestamp 18001
transform 1 0 3680 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_1_563
timestamp 18001
transform 1 0 3680 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_1_564
timestamp 18001
transform 1 0 3680 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_1_565
timestamp 18001
transform 1 0 3680 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_156_1_566
timestamp 18001
transform 1 0 3680 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_158_1_567
timestamp 18001
transform 1 0 3680 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_160_1_568
timestamp 18001
transform 1 0 3680 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_162_1_569
timestamp 18001
transform 1 0 3680 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_570
timestamp 18001
transform 1 0 3680 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_571
timestamp 18001
transform 1 0 6256 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_572
timestamp 18001
transform 1 0 8832 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_573
timestamp 18001
transform 1 0 11408 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_574
timestamp 18001
transform 1 0 13984 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_575
timestamp 18001
transform 1 0 16560 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_576
timestamp 18001
transform 1 0 19136 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_577
timestamp 18001
transform 1 0 21712 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_578
timestamp 18001
transform 1 0 24288 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_579
timestamp 18001
transform 1 0 26864 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_580
timestamp 18001
transform 1 0 29440 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_581
timestamp 18001
transform 1 0 32016 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_582
timestamp 18001
transform 1 0 34592 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_583
timestamp 18001
transform 1 0 37168 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_584
timestamp 18001
transform 1 0 39744 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_585
timestamp 18001
transform 1 0 42320 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_586
timestamp 18001
transform 1 0 44896 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_587
timestamp 18001
transform 1 0 47472 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_588
timestamp 18001
transform 1 0 50048 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_589
timestamp 18001
transform 1 0 52624 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_590
timestamp 18001
transform 1 0 55200 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_591
timestamp 18001
transform 1 0 57776 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_592
timestamp 18001
transform 1 0 60352 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_593
timestamp 18001
transform 1 0 62928 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_594
timestamp 18001
transform 1 0 65504 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_595
timestamp 18001
transform 1 0 68080 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_596
timestamp 18001
transform 1 0 70656 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_597
timestamp 18001
transform 1 0 73232 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_598
timestamp 18001
transform 1 0 75808 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_599
timestamp 18001
transform 1 0 78384 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_600
timestamp 18001
transform 1 0 80960 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_601
timestamp 18001
transform 1 0 83536 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_602
timestamp 18001
transform 1 0 86112 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_603
timestamp 18001
transform 1 0 6256 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_604
timestamp 18001
transform 1 0 11408 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_605
timestamp 18001
transform 1 0 16560 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_606
timestamp 18001
transform 1 0 21712 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_607
timestamp 18001
transform 1 0 26864 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_608
timestamp 18001
transform 1 0 32016 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_609
timestamp 18001
transform 1 0 37168 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_610
timestamp 18001
transform 1 0 42320 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_611
timestamp 18001
transform 1 0 47472 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_612
timestamp 18001
transform 1 0 52624 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_613
timestamp 18001
transform 1 0 57776 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_614
timestamp 18001
transform 1 0 62928 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_615
timestamp 18001
transform 1 0 68080 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_616
timestamp 18001
transform 1 0 73232 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_617
timestamp 18001
transform 1 0 78384 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_618
timestamp 18001
transform 1 0 83536 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_619
timestamp 18001
transform 1 0 3680 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_620
timestamp 18001
transform 1 0 8832 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_621
timestamp 18001
transform 1 0 13984 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_622
timestamp 18001
transform 1 0 19136 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_623
timestamp 18001
transform 1 0 24288 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_624
timestamp 18001
transform 1 0 29440 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_625
timestamp 18001
transform 1 0 34592 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_626
timestamp 18001
transform 1 0 39744 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_627
timestamp 18001
transform 1 0 44896 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_628
timestamp 18001
transform 1 0 50048 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_629
timestamp 18001
transform 1 0 55200 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_630
timestamp 18001
transform 1 0 60352 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_631
timestamp 18001
transform 1 0 65504 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_632
timestamp 18001
transform 1 0 70656 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_633
timestamp 18001
transform 1 0 75808 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_634
timestamp 18001
transform 1 0 80960 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_635
timestamp 18001
transform 1 0 86112 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_636
timestamp 18001
transform 1 0 6256 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_637
timestamp 18001
transform 1 0 11408 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_638
timestamp 18001
transform 1 0 16560 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_639
timestamp 18001
transform 1 0 21712 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_640
timestamp 18001
transform 1 0 26864 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_641
timestamp 18001
transform 1 0 32016 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_642
timestamp 18001
transform 1 0 37168 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_643
timestamp 18001
transform 1 0 42320 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_644
timestamp 18001
transform 1 0 47472 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_645
timestamp 18001
transform 1 0 52624 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_646
timestamp 18001
transform 1 0 57776 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_647
timestamp 18001
transform 1 0 62928 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_648
timestamp 18001
transform 1 0 68080 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_649
timestamp 18001
transform 1 0 73232 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_650
timestamp 18001
transform 1 0 78384 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_651
timestamp 18001
transform 1 0 83536 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_652
timestamp 18001
transform 1 0 3680 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_653
timestamp 18001
transform 1 0 8832 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_654
timestamp 18001
transform 1 0 13984 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_655
timestamp 18001
transform 1 0 19136 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_656
timestamp 18001
transform 1 0 24288 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_657
timestamp 18001
transform 1 0 29440 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_658
timestamp 18001
transform 1 0 34592 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_659
timestamp 18001
transform 1 0 39744 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_660
timestamp 18001
transform 1 0 44896 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_661
timestamp 18001
transform 1 0 50048 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_662
timestamp 18001
transform 1 0 55200 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_663
timestamp 18001
transform 1 0 60352 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_664
timestamp 18001
transform 1 0 65504 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_665
timestamp 18001
transform 1 0 70656 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_666
timestamp 18001
transform 1 0 75808 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_667
timestamp 18001
transform 1 0 80960 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_668
timestamp 18001
transform 1 0 86112 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_669
timestamp 18001
transform 1 0 6256 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_670
timestamp 18001
transform 1 0 11408 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_671
timestamp 18001
transform 1 0 16560 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_672
timestamp 18001
transform 1 0 21712 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_673
timestamp 18001
transform 1 0 26864 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_674
timestamp 18001
transform 1 0 32016 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_675
timestamp 18001
transform 1 0 37168 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_676
timestamp 18001
transform 1 0 42320 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_677
timestamp 18001
transform 1 0 47472 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_678
timestamp 18001
transform 1 0 52624 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_679
timestamp 18001
transform 1 0 57776 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_680
timestamp 18001
transform 1 0 62928 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_681
timestamp 18001
transform 1 0 68080 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_682
timestamp 18001
transform 1 0 73232 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_683
timestamp 18001
transform 1 0 78384 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_684
timestamp 18001
transform 1 0 83536 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_685
timestamp 18001
transform 1 0 3680 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_686
timestamp 18001
transform 1 0 8832 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_687
timestamp 18001
transform 1 0 13984 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_688
timestamp 18001
transform 1 0 19136 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_689
timestamp 18001
transform 1 0 24288 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_690
timestamp 18001
transform 1 0 29440 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_691
timestamp 18001
transform 1 0 34592 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_692
timestamp 18001
transform 1 0 39744 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_693
timestamp 18001
transform 1 0 44896 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_694
timestamp 18001
transform 1 0 50048 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_695
timestamp 18001
transform 1 0 55200 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_696
timestamp 18001
transform 1 0 60352 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_697
timestamp 18001
transform 1 0 65504 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_698
timestamp 18001
transform 1 0 70656 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_699
timestamp 18001
transform 1 0 75808 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_700
timestamp 18001
transform 1 0 80960 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_701
timestamp 18001
transform 1 0 86112 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_702
timestamp 18001
transform 1 0 3680 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_703
timestamp 18001
transform 1 0 6256 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_704
timestamp 18001
transform 1 0 8832 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_705
timestamp 18001
transform 1 0 11408 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_706
timestamp 18001
transform 1 0 13984 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_707
timestamp 18001
transform 1 0 16560 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_708
timestamp 18001
transform 1 0 19136 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_709
timestamp 18001
transform 1 0 21712 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_710
timestamp 18001
transform 1 0 24288 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_711
timestamp 18001
transform 1 0 26864 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_712
timestamp 18001
transform 1 0 29440 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_713
timestamp 18001
transform 1 0 32016 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_714
timestamp 18001
transform 1 0 34592 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_715
timestamp 18001
transform 1 0 37168 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_716
timestamp 18001
transform 1 0 39744 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_717
timestamp 18001
transform 1 0 42320 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_718
timestamp 18001
transform 1 0 44896 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_719
timestamp 18001
transform 1 0 47472 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_720
timestamp 18001
transform 1 0 50048 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_721
timestamp 18001
transform 1 0 52624 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_722
timestamp 18001
transform 1 0 55200 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_723
timestamp 18001
transform 1 0 57776 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_724
timestamp 18001
transform 1 0 60352 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_725
timestamp 18001
transform 1 0 62928 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_726
timestamp 18001
transform 1 0 65504 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_727
timestamp 18001
transform 1 0 68080 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_728
timestamp 18001
transform 1 0 70656 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_729
timestamp 18001
transform 1 0 73232 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_730
timestamp 18001
transform 1 0 75808 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_731
timestamp 18001
transform 1 0 78384 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_732
timestamp 18001
transform 1 0 80960 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_733
timestamp 18001
transform 1 0 83536 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_734
timestamp 18001
transform 1 0 86112 0 -1 95744
box -38 -48 130 592
<< labels >>
flabel metal2 s 49606 97200 49662 98000 0 FreeSans 224 90 0 0 clk
port 0 nsew signal input
flabel metal3 s 0 43528 800 43648 0 FreeSans 480 0 0 0 config_data_in
port 1 nsew signal input
flabel metal3 s 89200 50328 90000 50448 0 FreeSans 480 0 0 0 config_data_out
port 2 nsew signal output
flabel metal2 s 52182 97200 52238 98000 0 FreeSans 224 90 0 0 config_en
port 3 nsew signal input
flabel metal3 s 89200 27888 90000 28008 0 FreeSans 480 0 0 0 io_east_in[0]
port 4 nsew signal input
flabel metal3 s 89200 41488 90000 41608 0 FreeSans 480 0 0 0 io_east_in[10]
port 5 nsew signal input
flabel metal3 s 89200 42848 90000 42968 0 FreeSans 480 0 0 0 io_east_in[11]
port 6 nsew signal input
flabel metal3 s 89200 44208 90000 44328 0 FreeSans 480 0 0 0 io_east_in[12]
port 7 nsew signal input
flabel metal3 s 89200 45568 90000 45688 0 FreeSans 480 0 0 0 io_east_in[13]
port 8 nsew signal input
flabel metal2 s 662 0 718 800 0 FreeSans 224 90 0 0 io_east_in[14]
port 9 nsew signal input
flabel metal2 s 1306 0 1362 800 0 FreeSans 224 90 0 0 io_east_in[15]
port 10 nsew signal input
flabel metal3 s 89200 70048 90000 70168 0 FreeSans 480 0 0 0 io_east_in[16]
port 11 nsew signal input
flabel metal3 s 89200 71408 90000 71528 0 FreeSans 480 0 0 0 io_east_in[17]
port 12 nsew signal input
flabel metal3 s 89200 72768 90000 72888 0 FreeSans 480 0 0 0 io_east_in[18]
port 13 nsew signal input
flabel metal3 s 89200 74128 90000 74248 0 FreeSans 480 0 0 0 io_east_in[19]
port 14 nsew signal input
flabel metal3 s 89200 29248 90000 29368 0 FreeSans 480 0 0 0 io_east_in[1]
port 15 nsew signal input
flabel metal3 s 89200 75488 90000 75608 0 FreeSans 480 0 0 0 io_east_in[20]
port 16 nsew signal input
flabel metal3 s 89200 76848 90000 76968 0 FreeSans 480 0 0 0 io_east_in[21]
port 17 nsew signal input
flabel metal3 s 89200 78208 90000 78328 0 FreeSans 480 0 0 0 io_east_in[22]
port 18 nsew signal input
flabel metal3 s 89200 79568 90000 79688 0 FreeSans 480 0 0 0 io_east_in[23]
port 19 nsew signal input
flabel metal3 s 89200 80928 90000 81048 0 FreeSans 480 0 0 0 io_east_in[24]
port 20 nsew signal input
flabel metal3 s 89200 82288 90000 82408 0 FreeSans 480 0 0 0 io_east_in[25]
port 21 nsew signal input
flabel metal3 s 89200 83648 90000 83768 0 FreeSans 480 0 0 0 io_east_in[26]
port 22 nsew signal input
flabel metal3 s 89200 85008 90000 85128 0 FreeSans 480 0 0 0 io_east_in[27]
port 23 nsew signal input
flabel metal3 s 89200 86368 90000 86488 0 FreeSans 480 0 0 0 io_east_in[28]
port 24 nsew signal input
flabel metal3 s 89200 87728 90000 87848 0 FreeSans 480 0 0 0 io_east_in[29]
port 25 nsew signal input
flabel metal3 s 89200 30608 90000 30728 0 FreeSans 480 0 0 0 io_east_in[2]
port 26 nsew signal input
flabel metal2 s 1950 0 2006 800 0 FreeSans 224 90 0 0 io_east_in[30]
port 27 nsew signal input
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 io_east_in[31]
port 28 nsew signal input
flabel metal3 s 89200 31968 90000 32088 0 FreeSans 480 0 0 0 io_east_in[3]
port 29 nsew signal input
flabel metal3 s 89200 33328 90000 33448 0 FreeSans 480 0 0 0 io_east_in[4]
port 30 nsew signal input
flabel metal3 s 89200 34688 90000 34808 0 FreeSans 480 0 0 0 io_east_in[5]
port 31 nsew signal input
flabel metal3 s 89200 36048 90000 36168 0 FreeSans 480 0 0 0 io_east_in[6]
port 32 nsew signal input
flabel metal3 s 89200 37408 90000 37528 0 FreeSans 480 0 0 0 io_east_in[7]
port 33 nsew signal input
flabel metal3 s 89200 38768 90000 38888 0 FreeSans 480 0 0 0 io_east_in[8]
port 34 nsew signal input
flabel metal3 s 89200 40128 90000 40248 0 FreeSans 480 0 0 0 io_east_in[9]
port 35 nsew signal input
flabel metal3 s 89200 9528 90000 9648 0 FreeSans 480 0 0 0 io_east_out[0]
port 36 nsew signal output
flabel metal3 s 89200 22448 90000 22568 0 FreeSans 480 0 0 0 io_east_out[10]
port 37 nsew signal output
flabel metal3 s 89200 23808 90000 23928 0 FreeSans 480 0 0 0 io_east_out[11]
port 38 nsew signal output
flabel metal3 s 89200 25168 90000 25288 0 FreeSans 480 0 0 0 io_east_out[12]
port 39 nsew signal output
flabel metal3 s 89200 26528 90000 26648 0 FreeSans 480 0 0 0 io_east_out[13]
port 40 nsew signal output
flabel metal3 s 0 52368 800 52488 0 FreeSans 480 0 0 0 io_east_out[14]
port 41 nsew signal output
flabel metal3 s 0 60528 800 60648 0 FreeSans 480 0 0 0 io_east_out[15]
port 42 nsew signal output
flabel metal3 s 89200 51008 90000 51128 0 FreeSans 480 0 0 0 io_east_out[16]
port 43 nsew signal output
flabel metal3 s 89200 52368 90000 52488 0 FreeSans 480 0 0 0 io_east_out[17]
port 44 nsew signal output
flabel metal3 s 89200 53728 90000 53848 0 FreeSans 480 0 0 0 io_east_out[18]
port 45 nsew signal output
flabel metal3 s 89200 55088 90000 55208 0 FreeSans 480 0 0 0 io_east_out[19]
port 46 nsew signal output
flabel metal3 s 89200 10208 90000 10328 0 FreeSans 480 0 0 0 io_east_out[1]
port 47 nsew signal output
flabel metal3 s 89200 56448 90000 56568 0 FreeSans 480 0 0 0 io_east_out[20]
port 48 nsew signal output
flabel metal3 s 89200 57808 90000 57928 0 FreeSans 480 0 0 0 io_east_out[21]
port 49 nsew signal output
flabel metal3 s 89200 59168 90000 59288 0 FreeSans 480 0 0 0 io_east_out[22]
port 50 nsew signal output
flabel metal3 s 89200 60528 90000 60648 0 FreeSans 480 0 0 0 io_east_out[23]
port 51 nsew signal output
flabel metal3 s 89200 61888 90000 62008 0 FreeSans 480 0 0 0 io_east_out[24]
port 52 nsew signal output
flabel metal3 s 89200 63248 90000 63368 0 FreeSans 480 0 0 0 io_east_out[25]
port 53 nsew signal output
flabel metal3 s 89200 64608 90000 64728 0 FreeSans 480 0 0 0 io_east_out[26]
port 54 nsew signal output
flabel metal3 s 89200 65968 90000 66088 0 FreeSans 480 0 0 0 io_east_out[27]
port 55 nsew signal output
flabel metal3 s 89200 67328 90000 67448 0 FreeSans 480 0 0 0 io_east_out[28]
port 56 nsew signal output
flabel metal3 s 89200 68688 90000 68808 0 FreeSans 480 0 0 0 io_east_out[29]
port 57 nsew signal output
flabel metal3 s 89200 11568 90000 11688 0 FreeSans 480 0 0 0 io_east_out[2]
port 58 nsew signal output
flabel metal3 s 0 50328 800 50448 0 FreeSans 480 0 0 0 io_east_out[30]
port 59 nsew signal output
flabel metal3 s 0 48968 800 49088 0 FreeSans 480 0 0 0 io_east_out[31]
port 60 nsew signal output
flabel metal3 s 89200 12928 90000 13048 0 FreeSans 480 0 0 0 io_east_out[3]
port 61 nsew signal output
flabel metal3 s 89200 14288 90000 14408 0 FreeSans 480 0 0 0 io_east_out[4]
port 62 nsew signal output
flabel metal3 s 89200 15648 90000 15768 0 FreeSans 480 0 0 0 io_east_out[5]
port 63 nsew signal output
flabel metal3 s 89200 17008 90000 17128 0 FreeSans 480 0 0 0 io_east_out[6]
port 64 nsew signal output
flabel metal3 s 89200 18368 90000 18488 0 FreeSans 480 0 0 0 io_east_out[7]
port 65 nsew signal output
flabel metal3 s 89200 19728 90000 19848 0 FreeSans 480 0 0 0 io_east_out[8]
port 66 nsew signal output
flabel metal3 s 89200 21088 90000 21208 0 FreeSans 480 0 0 0 io_east_out[9]
port 67 nsew signal output
flabel metal2 s 14830 97200 14886 98000 0 FreeSans 224 90 0 0 io_north_in[0]
port 68 nsew signal input
flabel metal2 s 25778 97200 25834 98000 0 FreeSans 224 90 0 0 io_north_in[10]
port 69 nsew signal input
flabel metal2 s 27066 97200 27122 98000 0 FreeSans 224 90 0 0 io_north_in[11]
port 70 nsew signal input
flabel metal2 s 27710 97200 27766 98000 0 FreeSans 224 90 0 0 io_north_in[12]
port 71 nsew signal input
flabel metal2 s 28998 97200 29054 98000 0 FreeSans 224 90 0 0 io_north_in[13]
port 72 nsew signal input
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 io_north_in[14]
port 73 nsew signal input
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 io_north_in[15]
port 74 nsew signal input
flabel metal2 s 54758 97200 54814 98000 0 FreeSans 224 90 0 0 io_north_in[16]
port 75 nsew signal input
flabel metal2 s 56046 97200 56102 98000 0 FreeSans 224 90 0 0 io_north_in[17]
port 76 nsew signal input
flabel metal2 s 56690 97200 56746 98000 0 FreeSans 224 90 0 0 io_north_in[18]
port 77 nsew signal input
flabel metal2 s 57978 97200 58034 98000 0 FreeSans 224 90 0 0 io_north_in[19]
port 78 nsew signal input
flabel metal2 s 15474 97200 15530 98000 0 FreeSans 224 90 0 0 io_north_in[1]
port 79 nsew signal input
flabel metal2 s 59266 97200 59322 98000 0 FreeSans 224 90 0 0 io_north_in[20]
port 80 nsew signal input
flabel metal2 s 59910 97200 59966 98000 0 FreeSans 224 90 0 0 io_north_in[21]
port 81 nsew signal input
flabel metal2 s 61198 97200 61254 98000 0 FreeSans 224 90 0 0 io_north_in[22]
port 82 nsew signal input
flabel metal2 s 62486 97200 62542 98000 0 FreeSans 224 90 0 0 io_north_in[23]
port 83 nsew signal input
flabel metal2 s 63774 97200 63830 98000 0 FreeSans 224 90 0 0 io_north_in[24]
port 84 nsew signal input
flabel metal2 s 64418 97200 64474 98000 0 FreeSans 224 90 0 0 io_north_in[25]
port 85 nsew signal input
flabel metal2 s 65706 97200 65762 98000 0 FreeSans 224 90 0 0 io_north_in[26]
port 86 nsew signal input
flabel metal2 s 66994 97200 67050 98000 0 FreeSans 224 90 0 0 io_north_in[27]
port 87 nsew signal input
flabel metal2 s 67638 97200 67694 98000 0 FreeSans 224 90 0 0 io_north_in[28]
port 88 nsew signal input
flabel metal2 s 68926 97200 68982 98000 0 FreeSans 224 90 0 0 io_north_in[29]
port 89 nsew signal input
flabel metal2 s 16762 97200 16818 98000 0 FreeSans 224 90 0 0 io_north_in[2]
port 90 nsew signal input
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 io_north_in[30]
port 91 nsew signal input
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 io_north_in[31]
port 92 nsew signal input
flabel metal2 s 18050 97200 18106 98000 0 FreeSans 224 90 0 0 io_north_in[3]
port 93 nsew signal input
flabel metal2 s 19338 97200 19394 98000 0 FreeSans 224 90 0 0 io_north_in[4]
port 94 nsew signal input
flabel metal2 s 19982 97200 20038 98000 0 FreeSans 224 90 0 0 io_north_in[5]
port 95 nsew signal input
flabel metal2 s 21270 97200 21326 98000 0 FreeSans 224 90 0 0 io_north_in[6]
port 96 nsew signal input
flabel metal2 s 22558 97200 22614 98000 0 FreeSans 224 90 0 0 io_north_in[7]
port 97 nsew signal input
flabel metal2 s 23202 97200 23258 98000 0 FreeSans 224 90 0 0 io_north_in[8]
port 98 nsew signal input
flabel metal2 s 24490 97200 24546 98000 0 FreeSans 224 90 0 0 io_north_in[9]
port 99 nsew signal input
flabel metal2 s 30286 97200 30342 98000 0 FreeSans 224 90 0 0 io_north_out[0]
port 100 nsew signal output
flabel metal2 s 41234 97200 41290 98000 0 FreeSans 224 90 0 0 io_north_out[10]
port 101 nsew signal output
flabel metal2 s 42522 97200 42578 98000 0 FreeSans 224 90 0 0 io_north_out[11]
port 102 nsew signal output
flabel metal2 s 43166 97200 43222 98000 0 FreeSans 224 90 0 0 io_north_out[12]
port 103 nsew signal output
flabel metal2 s 44454 97200 44510 98000 0 FreeSans 224 90 0 0 io_north_out[13]
port 104 nsew signal output
flabel metal3 s 0 57808 800 57928 0 FreeSans 480 0 0 0 io_north_out[14]
port 105 nsew signal output
flabel metal3 s 0 51688 800 51808 0 FreeSans 480 0 0 0 io_north_out[15]
port 106 nsew signal output
flabel metal2 s 70214 97200 70270 98000 0 FreeSans 224 90 0 0 io_north_out[16]
port 107 nsew signal output
flabel metal2 s 71502 97200 71558 98000 0 FreeSans 224 90 0 0 io_north_out[17]
port 108 nsew signal output
flabel metal2 s 72146 97200 72202 98000 0 FreeSans 224 90 0 0 io_north_out[18]
port 109 nsew signal output
flabel metal2 s 73434 97200 73490 98000 0 FreeSans 224 90 0 0 io_north_out[19]
port 110 nsew signal output
flabel metal2 s 30930 97200 30986 98000 0 FreeSans 224 90 0 0 io_north_out[1]
port 111 nsew signal output
flabel metal2 s 74722 97200 74778 98000 0 FreeSans 224 90 0 0 io_north_out[20]
port 112 nsew signal output
flabel metal2 s 75366 97200 75422 98000 0 FreeSans 224 90 0 0 io_north_out[21]
port 113 nsew signal output
flabel metal2 s 76654 97200 76710 98000 0 FreeSans 224 90 0 0 io_north_out[22]
port 114 nsew signal output
flabel metal2 s 77942 97200 77998 98000 0 FreeSans 224 90 0 0 io_north_out[23]
port 115 nsew signal output
flabel metal2 s 79230 97200 79286 98000 0 FreeSans 224 90 0 0 io_north_out[24]
port 116 nsew signal output
flabel metal2 s 79874 97200 79930 98000 0 FreeSans 224 90 0 0 io_north_out[25]
port 117 nsew signal output
flabel metal2 s 81162 97200 81218 98000 0 FreeSans 224 90 0 0 io_north_out[26]
port 118 nsew signal output
flabel metal2 s 82450 97200 82506 98000 0 FreeSans 224 90 0 0 io_north_out[27]
port 119 nsew signal output
flabel metal3 s 89200 89088 90000 89208 0 FreeSans 480 0 0 0 io_north_out[28]
port 120 nsew signal output
flabel metal3 s 89200 88408 90000 88528 0 FreeSans 480 0 0 0 io_north_out[29]
port 121 nsew signal output
flabel metal2 s 32218 97200 32274 98000 0 FreeSans 224 90 0 0 io_north_out[2]
port 122 nsew signal output
flabel metal3 s 0 46928 800 47048 0 FreeSans 480 0 0 0 io_north_out[30]
port 123 nsew signal output
flabel metal3 s 0 55088 800 55208 0 FreeSans 480 0 0 0 io_north_out[31]
port 124 nsew signal output
flabel metal2 s 33506 97200 33562 98000 0 FreeSans 224 90 0 0 io_north_out[3]
port 125 nsew signal output
flabel metal2 s 34794 97200 34850 98000 0 FreeSans 224 90 0 0 io_north_out[4]
port 126 nsew signal output
flabel metal2 s 35438 97200 35494 98000 0 FreeSans 224 90 0 0 io_north_out[5]
port 127 nsew signal output
flabel metal2 s 36726 97200 36782 98000 0 FreeSans 224 90 0 0 io_north_out[6]
port 128 nsew signal output
flabel metal2 s 38014 97200 38070 98000 0 FreeSans 224 90 0 0 io_north_out[7]
port 129 nsew signal output
flabel metal2 s 38658 97200 38714 98000 0 FreeSans 224 90 0 0 io_north_out[8]
port 130 nsew signal output
flabel metal2 s 39946 97200 40002 98000 0 FreeSans 224 90 0 0 io_north_out[9]
port 131 nsew signal output
flabel metal2 s 30930 0 30986 800 0 FreeSans 224 90 0 0 io_south_in[0]
port 132 nsew signal input
flabel metal2 s 41878 0 41934 800 0 FreeSans 224 90 0 0 io_south_in[10]
port 133 nsew signal input
flabel metal2 s 42522 0 42578 800 0 FreeSans 224 90 0 0 io_south_in[11]
port 134 nsew signal input
flabel metal2 s 43810 0 43866 800 0 FreeSans 224 90 0 0 io_south_in[12]
port 135 nsew signal input
flabel metal2 s 45098 0 45154 800 0 FreeSans 224 90 0 0 io_south_in[13]
port 136 nsew signal input
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 io_south_in[14]
port 137 nsew signal input
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 io_south_in[15]
port 138 nsew signal input
flabel metal2 s 70858 0 70914 800 0 FreeSans 224 90 0 0 io_south_in[16]
port 139 nsew signal input
flabel metal2 s 71502 0 71558 800 0 FreeSans 224 90 0 0 io_south_in[17]
port 140 nsew signal input
flabel metal2 s 72790 0 72846 800 0 FreeSans 224 90 0 0 io_south_in[18]
port 141 nsew signal input
flabel metal2 s 74078 0 74134 800 0 FreeSans 224 90 0 0 io_south_in[19]
port 142 nsew signal input
flabel metal2 s 31574 0 31630 800 0 FreeSans 224 90 0 0 io_south_in[1]
port 143 nsew signal input
flabel metal2 s 75366 0 75422 800 0 FreeSans 224 90 0 0 io_south_in[20]
port 144 nsew signal input
flabel metal2 s 76010 0 76066 800 0 FreeSans 224 90 0 0 io_south_in[21]
port 145 nsew signal input
flabel metal2 s 77298 0 77354 800 0 FreeSans 224 90 0 0 io_south_in[22]
port 146 nsew signal input
flabel metal2 s 78586 0 78642 800 0 FreeSans 224 90 0 0 io_south_in[23]
port 147 nsew signal input
flabel metal2 s 79230 0 79286 800 0 FreeSans 224 90 0 0 io_south_in[24]
port 148 nsew signal input
flabel metal2 s 80518 0 80574 800 0 FreeSans 224 90 0 0 io_south_in[25]
port 149 nsew signal input
flabel metal2 s 81806 0 81862 800 0 FreeSans 224 90 0 0 io_south_in[26]
port 150 nsew signal input
flabel metal2 s 83094 0 83150 800 0 FreeSans 224 90 0 0 io_south_in[27]
port 151 nsew signal input
flabel metal3 s 89200 8848 90000 8968 0 FreeSans 480 0 0 0 io_south_in[28]
port 152 nsew signal input
flabel metal3 s 89200 8168 90000 8288 0 FreeSans 480 0 0 0 io_south_in[29]
port 153 nsew signal input
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 io_south_in[2]
port 154 nsew signal input
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 io_south_in[30]
port 155 nsew signal input
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 io_south_in[31]
port 156 nsew signal input
flabel metal2 s 34150 0 34206 800 0 FreeSans 224 90 0 0 io_south_in[3]
port 157 nsew signal input
flabel metal2 s 34794 0 34850 800 0 FreeSans 224 90 0 0 io_south_in[4]
port 158 nsew signal input
flabel metal2 s 36082 0 36138 800 0 FreeSans 224 90 0 0 io_south_in[5]
port 159 nsew signal input
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 io_south_in[6]
port 160 nsew signal input
flabel metal2 s 38658 0 38714 800 0 FreeSans 224 90 0 0 io_south_in[7]
port 161 nsew signal input
flabel metal2 s 39302 0 39358 800 0 FreeSans 224 90 0 0 io_south_in[8]
port 162 nsew signal input
flabel metal2 s 40590 0 40646 800 0 FreeSans 224 90 0 0 io_south_in[9]
port 163 nsew signal input
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 io_south_out[0]
port 164 nsew signal output
flabel metal2 s 26422 0 26478 800 0 FreeSans 224 90 0 0 io_south_out[10]
port 165 nsew signal output
flabel metal2 s 27066 0 27122 800 0 FreeSans 224 90 0 0 io_south_out[11]
port 166 nsew signal output
flabel metal2 s 28354 0 28410 800 0 FreeSans 224 90 0 0 io_south_out[12]
port 167 nsew signal output
flabel metal2 s 29642 0 29698 800 0 FreeSans 224 90 0 0 io_south_out[13]
port 168 nsew signal output
flabel metal3 s 0 53728 800 53848 0 FreeSans 480 0 0 0 io_south_out[14]
port 169 nsew signal output
flabel metal3 s 0 59168 800 59288 0 FreeSans 480 0 0 0 io_south_out[15]
port 170 nsew signal output
flabel metal2 s 55402 0 55458 800 0 FreeSans 224 90 0 0 io_south_out[16]
port 171 nsew signal output
flabel metal2 s 56046 0 56102 800 0 FreeSans 224 90 0 0 io_south_out[17]
port 172 nsew signal output
flabel metal2 s 57334 0 57390 800 0 FreeSans 224 90 0 0 io_south_out[18]
port 173 nsew signal output
flabel metal2 s 58622 0 58678 800 0 FreeSans 224 90 0 0 io_south_out[19]
port 174 nsew signal output
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 io_south_out[1]
port 175 nsew signal output
flabel metal2 s 59910 0 59966 800 0 FreeSans 224 90 0 0 io_south_out[20]
port 176 nsew signal output
flabel metal2 s 60554 0 60610 800 0 FreeSans 224 90 0 0 io_south_out[21]
port 177 nsew signal output
flabel metal2 s 61842 0 61898 800 0 FreeSans 224 90 0 0 io_south_out[22]
port 178 nsew signal output
flabel metal2 s 63130 0 63186 800 0 FreeSans 224 90 0 0 io_south_out[23]
port 179 nsew signal output
flabel metal2 s 63774 0 63830 800 0 FreeSans 224 90 0 0 io_south_out[24]
port 180 nsew signal output
flabel metal2 s 65062 0 65118 800 0 FreeSans 224 90 0 0 io_south_out[25]
port 181 nsew signal output
flabel metal2 s 66350 0 66406 800 0 FreeSans 224 90 0 0 io_south_out[26]
port 182 nsew signal output
flabel metal2 s 67638 0 67694 800 0 FreeSans 224 90 0 0 io_south_out[27]
port 183 nsew signal output
flabel metal2 s 68282 0 68338 800 0 FreeSans 224 90 0 0 io_south_out[28]
port 184 nsew signal output
flabel metal2 s 69570 0 69626 800 0 FreeSans 224 90 0 0 io_south_out[29]
port 185 nsew signal output
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 io_south_out[2]
port 186 nsew signal output
flabel metal3 s 0 47608 800 47728 0 FreeSans 480 0 0 0 io_south_out[30]
port 187 nsew signal output
flabel metal3 s 0 51008 800 51128 0 FreeSans 480 0 0 0 io_south_out[31]
port 188 nsew signal output
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 io_south_out[3]
port 189 nsew signal output
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 io_south_out[4]
port 190 nsew signal output
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 io_south_out[5]
port 191 nsew signal output
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 io_south_out[6]
port 192 nsew signal output
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 io_south_out[7]
port 193 nsew signal output
flabel metal2 s 23846 0 23902 800 0 FreeSans 224 90 0 0 io_south_out[8]
port 194 nsew signal output
flabel metal2 s 25134 0 25190 800 0 FreeSans 224 90 0 0 io_south_out[9]
port 195 nsew signal output
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 io_west_in[0]
port 196 nsew signal input
flabel metal3 s 0 22448 800 22568 0 FreeSans 480 0 0 0 io_west_in[10]
port 197 nsew signal input
flabel metal3 s 0 23808 800 23928 0 FreeSans 480 0 0 0 io_west_in[11]
port 198 nsew signal input
flabel metal3 s 0 25168 800 25288 0 FreeSans 480 0 0 0 io_west_in[12]
port 199 nsew signal input
flabel metal3 s 0 26528 800 26648 0 FreeSans 480 0 0 0 io_west_in[13]
port 200 nsew signal input
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 io_west_in[14]
port 201 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 io_west_in[15]
port 202 nsew signal input
flabel metal3 s 0 48288 800 48408 0 FreeSans 480 0 0 0 io_west_in[16]
port 203 nsew signal input
flabel metal3 s 0 53048 800 53168 0 FreeSans 480 0 0 0 io_west_in[17]
port 204 nsew signal input
flabel metal3 s 0 54408 800 54528 0 FreeSans 480 0 0 0 io_west_in[18]
port 205 nsew signal input
flabel metal3 s 0 55768 800 55888 0 FreeSans 480 0 0 0 io_west_in[19]
port 206 nsew signal input
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 io_west_in[1]
port 207 nsew signal input
flabel metal3 s 0 57128 800 57248 0 FreeSans 480 0 0 0 io_west_in[20]
port 208 nsew signal input
flabel metal3 s 0 58488 800 58608 0 FreeSans 480 0 0 0 io_west_in[21]
port 209 nsew signal input
flabel metal3 s 0 59848 800 59968 0 FreeSans 480 0 0 0 io_west_in[22]
port 210 nsew signal input
flabel metal3 s 0 61208 800 61328 0 FreeSans 480 0 0 0 io_west_in[23]
port 211 nsew signal input
flabel metal3 s 0 61888 800 62008 0 FreeSans 480 0 0 0 io_west_in[24]
port 212 nsew signal input
flabel metal3 s 0 63248 800 63368 0 FreeSans 480 0 0 0 io_west_in[25]
port 213 nsew signal input
flabel metal3 s 0 64608 800 64728 0 FreeSans 480 0 0 0 io_west_in[26]
port 214 nsew signal input
flabel metal3 s 0 65968 800 66088 0 FreeSans 480 0 0 0 io_west_in[27]
port 215 nsew signal input
flabel metal3 s 0 67328 800 67448 0 FreeSans 480 0 0 0 io_west_in[28]
port 216 nsew signal input
flabel metal3 s 0 68688 800 68808 0 FreeSans 480 0 0 0 io_west_in[29]
port 217 nsew signal input
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 io_west_in[2]
port 218 nsew signal input
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 io_west_in[30]
port 219 nsew signal input
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 io_west_in[31]
port 220 nsew signal input
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 io_west_in[3]
port 221 nsew signal input
flabel metal3 s 0 14288 800 14408 0 FreeSans 480 0 0 0 io_west_in[4]
port 222 nsew signal input
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 io_west_in[5]
port 223 nsew signal input
flabel metal3 s 0 17008 800 17128 0 FreeSans 480 0 0 0 io_west_in[6]
port 224 nsew signal input
flabel metal3 s 0 18368 800 18488 0 FreeSans 480 0 0 0 io_west_in[7]
port 225 nsew signal input
flabel metal3 s 0 19728 800 19848 0 FreeSans 480 0 0 0 io_west_in[8]
port 226 nsew signal input
flabel metal3 s 0 21088 800 21208 0 FreeSans 480 0 0 0 io_west_in[9]
port 227 nsew signal input
flabel metal3 s 0 27888 800 28008 0 FreeSans 480 0 0 0 io_west_out[0]
port 228 nsew signal output
flabel metal3 s 0 41488 800 41608 0 FreeSans 480 0 0 0 io_west_out[10]
port 229 nsew signal output
flabel metal3 s 0 42848 800 42968 0 FreeSans 480 0 0 0 io_west_out[11]
port 230 nsew signal output
flabel metal3 s 0 44208 800 44328 0 FreeSans 480 0 0 0 io_west_out[12]
port 231 nsew signal output
flabel metal3 s 0 45568 800 45688 0 FreeSans 480 0 0 0 io_west_out[13]
port 232 nsew signal output
flabel metal3 s 0 56448 800 56568 0 FreeSans 480 0 0 0 io_west_out[14]
port 233 nsew signal output
flabel metal3 s 0 46248 800 46368 0 FreeSans 480 0 0 0 io_west_out[15]
port 234 nsew signal output
flabel metal3 s 0 70048 800 70168 0 FreeSans 480 0 0 0 io_west_out[16]
port 235 nsew signal output
flabel metal3 s 0 71408 800 71528 0 FreeSans 480 0 0 0 io_west_out[17]
port 236 nsew signal output
flabel metal3 s 0 72768 800 72888 0 FreeSans 480 0 0 0 io_west_out[18]
port 237 nsew signal output
flabel metal3 s 0 74128 800 74248 0 FreeSans 480 0 0 0 io_west_out[19]
port 238 nsew signal output
flabel metal3 s 0 29248 800 29368 0 FreeSans 480 0 0 0 io_west_out[1]
port 239 nsew signal output
flabel metal3 s 0 75488 800 75608 0 FreeSans 480 0 0 0 io_west_out[20]
port 240 nsew signal output
flabel metal3 s 0 76848 800 76968 0 FreeSans 480 0 0 0 io_west_out[21]
port 241 nsew signal output
flabel metal3 s 0 78208 800 78328 0 FreeSans 480 0 0 0 io_west_out[22]
port 242 nsew signal output
flabel metal3 s 0 79568 800 79688 0 FreeSans 480 0 0 0 io_west_out[23]
port 243 nsew signal output
flabel metal3 s 0 80928 800 81048 0 FreeSans 480 0 0 0 io_west_out[24]
port 244 nsew signal output
flabel metal3 s 0 82288 800 82408 0 FreeSans 480 0 0 0 io_west_out[25]
port 245 nsew signal output
flabel metal3 s 0 83648 800 83768 0 FreeSans 480 0 0 0 io_west_out[26]
port 246 nsew signal output
flabel metal3 s 0 85008 800 85128 0 FreeSans 480 0 0 0 io_west_out[27]
port 247 nsew signal output
flabel metal3 s 0 86368 800 86488 0 FreeSans 480 0 0 0 io_west_out[28]
port 248 nsew signal output
flabel metal2 s 8390 97200 8446 98000 0 FreeSans 224 90 0 0 io_west_out[29]
port 249 nsew signal output
flabel metal3 s 0 30608 800 30728 0 FreeSans 480 0 0 0 io_west_out[2]
port 250 nsew signal output
flabel metal3 s 0 49648 800 49768 0 FreeSans 480 0 0 0 io_west_out[30]
port 251 nsew signal output
flabel metal3 s 0 44888 800 45008 0 FreeSans 480 0 0 0 io_west_out[31]
port 252 nsew signal output
flabel metal3 s 0 31968 800 32088 0 FreeSans 480 0 0 0 io_west_out[3]
port 253 nsew signal output
flabel metal3 s 0 33328 800 33448 0 FreeSans 480 0 0 0 io_west_out[4]
port 254 nsew signal output
flabel metal3 s 0 34688 800 34808 0 FreeSans 480 0 0 0 io_west_out[5]
port 255 nsew signal output
flabel metal3 s 0 36048 800 36168 0 FreeSans 480 0 0 0 io_west_out[6]
port 256 nsew signal output
flabel metal3 s 0 37408 800 37528 0 FreeSans 480 0 0 0 io_west_out[7]
port 257 nsew signal output
flabel metal3 s 0 38768 800 38888 0 FreeSans 480 0 0 0 io_west_out[8]
port 258 nsew signal output
flabel metal3 s 0 40128 800 40248 0 FreeSans 480 0 0 0 io_west_out[9]
port 259 nsew signal output
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 le_clk
port 260 nsew signal input
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 le_en
port 261 nsew signal input
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 le_nrst
port 262 nsew signal input
flabel metal2 s 50894 97200 50950 98000 0 FreeSans 224 90 0 0 nrst
port 263 nsew signal input
flabel metal4 s -416 656 -96 97264 0 FreeSans 1920 90 0 0 vccd1
port 264 nsew power bidirectional
flabel metal5 s -416 656 90392 976 0 FreeSans 2560 0 0 0 vccd1
port 264 nsew power bidirectional
flabel metal5 s -416 96944 90392 97264 0 FreeSans 2560 0 0 0 vccd1
port 264 nsew power bidirectional
flabel metal4 s 90072 656 90392 97264 0 FreeSans 1920 90 0 0 vccd1
port 264 nsew power bidirectional
flabel metal4 s 36944 -4 37264 8559 0 FreeSans 1920 90 0 0 vccd1
port 264 nsew power bidirectional
flabel metal4 s 36944 90377 37264 97924 0 FreeSans 1920 90 0 0 vccd1
port 264 nsew power bidirectional
flabel metal4 s 72944 -4 73264 8559 0 FreeSans 1920 90 0 0 vccd1
port 264 nsew power bidirectional
flabel metal4 s 72944 90377 73264 97924 0 FreeSans 1920 90 0 0 vccd1
port 264 nsew power bidirectional
flabel metal5 s -1076 35416 91052 35736 0 FreeSans 2560 0 0 0 vccd1
port 264 nsew power bidirectional
flabel metal5 s -1076 68816 91052 69136 0 FreeSans 2560 0 0 0 vccd1
port 264 nsew power bidirectional
flabel metal4 s 3060 5392 3380 91984 0 FreeSans 1920 90 0 0 vccd1
port 264 nsew power bidirectional
flabel metal4 s -1076 -4 -756 97924 0 FreeSans 1920 90 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal5 s -1076 -4 91052 316 0 FreeSans 2560 0 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal5 s -1076 97604 91052 97924 0 FreeSans 2560 0 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal4 s 90732 -4 91052 97924 0 FreeSans 1920 90 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal4 s 37604 -4 37924 8559 0 FreeSans 1920 90 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal4 s 37604 90377 37924 97924 0 FreeSans 1920 90 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal4 s 73604 -4 73924 8559 0 FreeSans 1920 90 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal4 s 73604 90377 73924 97924 0 FreeSans 1920 90 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal5 s -1076 36076 91052 36396 0 FreeSans 2560 0 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal5 s -1076 69476 91052 69796 0 FreeSans 2560 0 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal4 s 3796 5392 4116 91984 0 FreeSans 1920 90 0 0 vssd1
port 265 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 90000 98000
<< end >>
