magic
tech sky130A
magscale 1 2
timestamp 1752462437
<< viali >>
rect 14105 95625 14139 95659
rect 15393 95625 15427 95659
rect 16681 95625 16715 95659
rect 17325 95625 17359 95659
rect 18613 95625 18647 95659
rect 19901 95625 19935 95659
rect 21189 95625 21223 95659
rect 21833 95625 21867 95659
rect 23121 95625 23155 95659
rect 25053 95625 25087 95659
rect 26341 95625 26375 95659
rect 27629 95625 27663 95659
rect 29009 95625 29043 95659
rect 29561 95625 29595 95659
rect 30849 95625 30883 95659
rect 32505 95625 32539 95659
rect 33057 95625 33091 95659
rect 34437 95625 34471 95659
rect 35725 95625 35759 95659
rect 37013 95625 37047 95659
rect 37565 95625 37599 95659
rect 38945 95625 38979 95659
rect 40233 95625 40267 95659
rect 40785 95625 40819 95659
rect 42165 95625 42199 95659
rect 43453 95625 43487 95659
rect 44741 95625 44775 95659
rect 45293 95625 45327 95659
rect 46673 95625 46707 95659
rect 47961 95625 47995 95659
rect 48513 95625 48547 95659
rect 50905 95625 50939 95659
rect 55045 95625 55079 95659
rect 57161 95625 57195 95659
rect 58541 95625 58575 95659
rect 59829 95625 59863 95659
rect 60473 95625 60507 95659
rect 61761 95625 61795 95659
rect 63049 95625 63083 95659
rect 63693 95625 63727 95659
rect 64981 95625 65015 95659
rect 66361 95625 66395 95659
rect 67925 95625 67959 95659
rect 69397 95625 69431 95659
rect 69949 95625 69983 95659
rect 70777 95625 70811 95659
rect 71421 95625 71455 95659
rect 72709 95625 72743 95659
rect 74365 95625 74399 95659
rect 75653 95625 75687 95659
rect 76205 95625 76239 95659
rect 77585 95625 77619 95659
rect 78873 95625 78907 95659
rect 79425 95625 79459 95659
rect 80805 95625 80839 95659
rect 82093 95625 82127 95659
rect 83381 95625 83415 95659
rect 83933 95625 83967 95659
rect 85313 95625 85347 95659
rect 86601 95625 86635 95659
rect 87153 95625 87187 95659
rect 88533 95625 88567 95659
rect 89821 95625 89855 95659
rect 91109 95625 91143 95659
rect 17601 95557 17635 95591
rect 18981 95557 19015 95591
rect 20269 95557 20303 95591
rect 21557 95557 21591 95591
rect 23489 95557 23523 95591
rect 60197 95557 60231 95591
rect 60749 95557 60783 95591
rect 62129 95557 62163 95591
rect 63417 95557 63451 95591
rect 65349 95557 65383 95591
rect 14289 95489 14323 95523
rect 15577 95489 15611 95523
rect 16865 95489 16899 95523
rect 22017 95489 22051 95523
rect 25237 95489 25271 95523
rect 26709 95489 26743 95523
rect 27997 95489 28031 95523
rect 29285 95489 29319 95523
rect 29745 95489 29779 95523
rect 31217 95489 31251 95523
rect 32321 95489 32355 95523
rect 33241 95489 33275 95523
rect 34253 95489 34287 95523
rect 35541 95489 35575 95523
rect 36829 95489 36863 95523
rect 37749 95489 37783 95523
rect 38761 95489 38795 95523
rect 40049 95489 40083 95523
rect 40969 95489 41003 95523
rect 41981 95489 42015 95523
rect 43269 95489 43303 95523
rect 44557 95489 44591 95523
rect 45477 95489 45511 95523
rect 46489 95489 46523 95523
rect 47777 95489 47811 95523
rect 48697 95489 48731 95523
rect 51089 95489 51123 95523
rect 52469 95489 52503 95523
rect 52745 95489 52779 95523
rect 52929 95489 52963 95523
rect 55321 95489 55355 95523
rect 57069 95489 57103 95523
rect 57713 95489 57747 95523
rect 57897 95489 57931 95523
rect 58725 95489 58759 95523
rect 63877 95489 63911 95523
rect 66453 95489 66487 95523
rect 68201 95489 68235 95523
rect 69305 95489 69339 95523
rect 69857 95489 69891 95523
rect 71145 95489 71179 95523
rect 71605 95489 71639 95523
rect 72893 95489 72927 95523
rect 74181 95489 74215 95523
rect 75469 95489 75503 95523
rect 76389 95489 76423 95523
rect 77401 95489 77435 95523
rect 78689 95489 78723 95523
rect 79609 95489 79643 95523
rect 80621 95489 80655 95523
rect 81909 95489 81943 95523
rect 83197 95489 83231 95523
rect 84117 95489 84151 95523
rect 85129 95489 85163 95523
rect 86417 95489 86451 95523
rect 87337 95489 87371 95523
rect 88349 95489 88383 95523
rect 89637 95489 89671 95523
rect 90925 95489 90959 95523
rect 25513 95421 25547 95455
rect 52101 95421 52135 95455
rect 54125 95421 54159 95455
rect 54401 95421 54435 95455
rect 56517 95421 56551 95455
rect 66729 95421 66763 95455
rect 68477 95421 68511 95455
rect 18797 95353 18831 95387
rect 20085 95353 20119 95387
rect 21373 95353 21407 95387
rect 23305 95353 23339 95387
rect 29101 95353 29135 95387
rect 60013 95353 60047 95387
rect 61945 95353 61979 95387
rect 63233 95353 63267 95387
rect 14473 95285 14507 95319
rect 15761 95285 15795 95319
rect 17049 95285 17083 95319
rect 17693 95285 17727 95319
rect 22201 95285 22235 95319
rect 26525 95285 26559 95319
rect 27813 95285 27847 95319
rect 29929 95285 29963 95319
rect 31033 95285 31067 95319
rect 56885 95285 56919 95319
rect 57529 95285 57563 95319
rect 58909 95285 58943 95319
rect 60841 95285 60875 95319
rect 64061 95285 64095 95319
rect 65257 95285 65291 95319
rect 69121 95285 69155 95319
rect 69673 95285 69707 95319
rect 70961 95285 70995 95319
rect 71789 95285 71823 95319
rect 73077 95285 73111 95319
rect 24409 95081 24443 95115
rect 52837 95081 52871 95115
rect 56793 95081 56827 95115
rect 24593 94945 24627 94979
rect 52929 94945 52963 94979
rect 24869 94877 24903 94911
rect 51181 94741 51215 94775
rect 54585 93993 54619 94027
rect 54769 93925 54803 93959
rect 54309 93857 54343 93891
rect 53113 93789 53147 93823
rect 56793 93449 56827 93483
rect 31677 93313 31711 93347
rect 40509 93313 40543 93347
rect 52745 93313 52779 93347
rect 56701 93313 56735 93347
rect 32137 93245 32171 93279
rect 40325 93245 40359 93279
rect 42257 93245 42291 93279
rect 42441 93245 42475 93279
rect 50905 93245 50939 93279
rect 53941 93245 53975 93279
rect 54401 93245 54435 93279
rect 56241 93245 56275 93279
rect 52469 93177 52503 93211
rect 8953 93109 8987 93143
rect 10057 93109 10091 93143
rect 11161 93109 11195 93143
rect 12265 93109 12299 93143
rect 13277 93109 13311 93143
rect 30389 93109 30423 93143
rect 31861 93109 31895 93143
rect 51089 93109 51123 93143
rect 52009 93109 52043 93143
rect 52377 93109 52411 93143
rect 54217 93109 54251 93143
rect 55137 93109 55171 93143
rect 57069 93109 57103 93143
rect 97365 87397 97399 87431
rect 1685 87261 1719 87295
rect 97273 87261 97307 87295
rect 97549 87261 97583 87295
rect 1501 87125 1535 87159
rect 1685 86785 1719 86819
rect 97273 86785 97307 86819
rect 97549 86785 97583 86819
rect 1501 86581 1535 86615
rect 97365 86581 97399 86615
rect 97365 85221 97399 85255
rect 1685 85085 1719 85119
rect 97273 85085 97307 85119
rect 97549 85085 97583 85119
rect 1501 84949 1535 84983
rect 1685 84609 1719 84643
rect 97273 84609 97307 84643
rect 97549 84609 97583 84643
rect 1501 84473 1535 84507
rect 97365 84405 97399 84439
rect 1685 83521 1719 83555
rect 97273 83521 97307 83555
rect 97549 83521 97583 83555
rect 1501 83317 1535 83351
rect 97365 83317 97399 83351
rect 97365 81957 97399 81991
rect 1685 81821 1719 81855
rect 97273 81821 97307 81855
rect 97549 81821 97583 81855
rect 1501 81685 1535 81719
rect 1685 81345 1719 81379
rect 97273 81345 97307 81379
rect 97549 81345 97583 81379
rect 1501 81141 1535 81175
rect 97365 81141 97399 81175
rect 97365 79781 97399 79815
rect 1685 79645 1719 79679
rect 97273 79645 97307 79679
rect 97549 79645 97583 79679
rect 1501 79509 1535 79543
rect 1685 79169 1719 79203
rect 97181 79169 97215 79203
rect 97457 79169 97491 79203
rect 1501 79033 1535 79067
rect 97273 79033 97307 79067
rect 1685 78081 1719 78115
rect 97273 78081 97307 78115
rect 97549 78081 97583 78115
rect 1501 77877 1535 77911
rect 97365 77877 97399 77911
rect 97365 76517 97399 76551
rect 1685 76381 1719 76415
rect 97273 76381 97307 76415
rect 97549 76381 97583 76415
rect 1501 76245 1535 76279
rect 1501 76041 1535 76075
rect 1685 75905 1719 75939
rect 97273 75905 97307 75939
rect 97549 75905 97583 75939
rect 97365 75701 97399 75735
rect 97273 74341 97307 74375
rect 1685 74205 1719 74239
rect 97181 74137 97215 74171
rect 97457 74137 97491 74171
rect 1501 74069 1535 74103
rect 1685 73729 1719 73763
rect 97273 73729 97307 73763
rect 97549 73729 97583 73763
rect 1501 73593 1535 73627
rect 97365 73525 97399 73559
rect 1685 72641 1719 72675
rect 97273 72573 97307 72607
rect 97549 72573 97583 72607
rect 1501 72437 1535 72471
rect 97549 72165 97583 72199
rect 97365 71077 97399 71111
rect 1685 70941 1719 70975
rect 97273 70941 97307 70975
rect 97549 70941 97583 70975
rect 1501 70805 1535 70839
rect 5549 70601 5583 70635
rect 97457 70601 97491 70635
rect 1409 70465 1443 70499
rect 1685 70465 1719 70499
rect 97273 70465 97307 70499
rect 1593 70261 1627 70295
rect 5641 69853 5675 69887
rect 4353 69717 4387 69751
rect 5641 69513 5675 69547
rect 97273 68765 97307 68799
rect 1501 68697 1535 68731
rect 1685 68697 1719 68731
rect 1777 68629 1811 68663
rect 97457 68629 97491 68663
rect 1501 68289 1535 68323
rect 1777 68289 1811 68323
rect 97273 68289 97307 68323
rect 1685 68153 1719 68187
rect 97457 68085 97491 68119
rect 1501 67201 1535 67235
rect 1777 67201 1811 67235
rect 97273 67201 97307 67235
rect 1685 67065 1719 67099
rect 97457 66997 97491 67031
rect 1685 65637 1719 65671
rect 97273 65501 97307 65535
rect 1501 65433 1535 65467
rect 1777 65433 1811 65467
rect 97457 65365 97491 65399
rect 1501 65025 1535 65059
rect 1777 65025 1811 65059
rect 97273 65025 97307 65059
rect 1685 64889 1719 64923
rect 97457 64889 97491 64923
rect 97273 63325 97307 63359
rect 1501 63257 1535 63291
rect 1685 63257 1719 63291
rect 1777 63189 1811 63223
rect 97457 63189 97491 63223
rect 1501 62849 1535 62883
rect 1961 62849 1995 62883
rect 97273 62849 97307 62883
rect 1777 62713 1811 62747
rect 97457 62645 97491 62679
rect 1501 61761 1535 61795
rect 1777 61761 1811 61795
rect 97273 61761 97307 61795
rect 1685 61625 1719 61659
rect 97457 61557 97491 61591
rect 1777 60265 1811 60299
rect 97273 60061 97307 60095
rect 1501 59993 1535 60027
rect 1961 59993 1995 60027
rect 97457 59925 97491 59959
rect 1409 59585 1443 59619
rect 1777 59585 1811 59619
rect 97273 59585 97307 59619
rect 1593 59381 1627 59415
rect 97457 59381 97491 59415
rect 1409 57885 1443 57919
rect 1777 57885 1811 57919
rect 97273 57885 97307 57919
rect 1593 57749 1627 57783
rect 97457 57749 97491 57783
rect 1501 57409 1535 57443
rect 1961 57409 1995 57443
rect 97273 57409 97307 57443
rect 1777 57273 1811 57307
rect 97457 57205 97491 57239
rect 1501 56321 1535 56355
rect 1961 56321 1995 56355
rect 97273 56321 97307 56355
rect 1777 56185 1811 56219
rect 97457 56117 97491 56151
rect 1593 54825 1627 54859
rect 1409 54621 1443 54655
rect 1777 54621 1811 54655
rect 97273 54621 97307 54655
rect 97457 54485 97491 54519
rect 1409 54145 1443 54179
rect 1777 54145 1811 54179
rect 97273 54145 97307 54179
rect 1593 53941 1627 53975
rect 97457 53941 97491 53975
rect 5641 51017 5675 51051
rect 5273 50813 5307 50847
rect 94697 50813 94731 50847
rect 5457 50745 5491 50779
rect 94513 50745 94547 50779
rect 94329 50677 94363 50711
rect 5641 50133 5675 50167
rect 1593 48841 1627 48875
rect 5549 48841 5583 48875
rect 94697 48773 94731 48807
rect 1409 48705 1443 48739
rect 1777 48705 1811 48739
rect 94329 48705 94363 48739
rect 5273 48637 5307 48671
rect 94513 48637 94547 48671
rect 5457 48569 5491 48603
rect 94881 48501 94915 48535
rect 5641 48229 5675 48263
rect 1685 45917 1719 45951
rect 97273 45917 97307 45951
rect 97549 45917 97583 45951
rect 1501 45781 1535 45815
rect 97365 45781 97399 45815
rect 1501 44489 1535 44523
rect 1685 44353 1719 44387
rect 97273 44353 97307 44387
rect 97549 44353 97583 44387
rect 97365 44217 97399 44251
rect 1685 43265 1719 43299
rect 97273 43265 97307 43299
rect 97549 43265 97583 43299
rect 97365 43129 97399 43163
rect 1501 43061 1535 43095
rect 1685 42653 1719 42687
rect 97273 42653 97307 42687
rect 97549 42653 97583 42687
rect 1501 42517 1535 42551
rect 97365 42517 97399 42551
rect 97365 41225 97399 41259
rect 1685 41089 1719 41123
rect 97273 41089 97307 41123
rect 97549 41089 97583 41123
rect 1501 40953 1535 40987
rect 1685 40477 1719 40511
rect 97273 40477 97307 40511
rect 97549 40477 97583 40511
rect 1501 40341 1535 40375
rect 97365 40341 97399 40375
rect 97365 39049 97399 39083
rect 1685 38913 1719 38947
rect 97273 38913 97307 38947
rect 97549 38913 97583 38947
rect 1501 38709 1535 38743
rect 97365 37961 97399 37995
rect 1685 37825 1719 37859
rect 97273 37825 97307 37859
rect 97549 37825 97583 37859
rect 1501 37621 1535 37655
rect 97273 37281 97307 37315
rect 1685 37213 1719 37247
rect 97181 37145 97215 37179
rect 97457 37145 97491 37179
rect 1501 37077 1535 37111
rect 97365 35785 97399 35819
rect 1685 35649 1719 35683
rect 97273 35649 97307 35683
rect 97549 35649 97583 35683
rect 1501 35513 1535 35547
rect 1685 35037 1719 35071
rect 97273 35037 97307 35071
rect 97549 35037 97583 35071
rect 1501 34901 1535 34935
rect 97365 34901 97399 34935
rect 97365 33609 97399 33643
rect 1685 33473 1719 33507
rect 97273 33473 97307 33507
rect 97549 33473 97583 33507
rect 1501 33269 1535 33303
rect 97273 32453 97307 32487
rect 1685 32385 1719 32419
rect 97181 32385 97215 32419
rect 97457 32385 97491 32419
rect 1501 32181 1535 32215
rect 1501 31909 1535 31943
rect 97365 31909 97399 31943
rect 1685 31773 1719 31807
rect 97273 31773 97307 31807
rect 97549 31773 97583 31807
rect 97549 30549 97583 30583
rect 1685 30209 1719 30243
rect 97273 30209 97307 30243
rect 97549 30141 97583 30175
rect 1501 30073 1535 30107
rect 1685 29597 1719 29631
rect 97273 29597 97307 29631
rect 97549 29597 97583 29631
rect 1501 29461 1535 29495
rect 97365 29461 97399 29495
rect 1593 28169 1627 28203
rect 1409 28033 1443 28067
rect 1685 28033 1719 28067
rect 97273 28033 97307 28067
rect 97457 27897 97491 27931
rect 1501 26945 1535 26979
rect 1685 26945 1719 26979
rect 97273 26945 97307 26979
rect 1777 26877 1811 26911
rect 97457 26741 97491 26775
rect 97457 26469 97491 26503
rect 1501 26333 1535 26367
rect 1777 26333 1811 26367
rect 97273 26333 97307 26367
rect 1685 26265 1719 26299
rect 1501 24769 1535 24803
rect 1685 24769 1719 24803
rect 97273 24769 97307 24803
rect 1777 24701 1811 24735
rect 97457 24565 97491 24599
rect 97273 24157 97307 24191
rect 1501 24089 1535 24123
rect 1685 24089 1719 24123
rect 1777 24021 1811 24055
rect 97457 24021 97491 24055
rect 1501 22593 1535 22627
rect 1685 22593 1719 22627
rect 97273 22593 97307 22627
rect 1777 22525 1811 22559
rect 97457 22457 97491 22491
rect 1501 21505 1535 21539
rect 1685 21505 1719 21539
rect 97273 21505 97307 21539
rect 1777 21437 1811 21471
rect 97457 21301 97491 21335
rect 97273 20893 97307 20927
rect 1501 20825 1535 20859
rect 1869 20825 1903 20859
rect 1961 20757 1995 20791
rect 97457 20757 97491 20791
rect 97457 19465 97491 19499
rect 1501 19329 1535 19363
rect 1777 19329 1811 19363
rect 97273 19329 97307 19363
rect 1685 19193 1719 19227
rect 97273 18717 97307 18751
rect 1501 18649 1535 18683
rect 1869 18649 1903 18683
rect 1961 18581 1995 18615
rect 97457 18581 97491 18615
rect 1593 17289 1627 17323
rect 1409 17153 1443 17187
rect 1777 17153 1811 17187
rect 97273 17153 97307 17187
rect 97457 17017 97491 17051
rect 1593 16201 1627 16235
rect 1409 16065 1443 16099
rect 1777 16065 1811 16099
rect 97273 16065 97307 16099
rect 97457 15861 97491 15895
rect 97273 15453 97307 15487
rect 1501 15385 1535 15419
rect 1869 15385 1903 15419
rect 1961 15317 1995 15351
rect 97457 15317 97491 15351
rect 97457 14025 97491 14059
rect 1501 13889 1535 13923
rect 1869 13889 1903 13923
rect 97273 13889 97307 13923
rect 1961 13821 1995 13855
rect 1593 13413 1627 13447
rect 1409 13277 1443 13311
rect 1777 13277 1811 13311
rect 97273 13277 97307 13311
rect 97457 13141 97491 13175
rect 1593 11849 1627 11883
rect 1409 11713 1443 11747
rect 1777 11713 1811 11747
rect 97273 11713 97307 11747
rect 97457 11577 97491 11611
rect 97181 8449 97215 8483
rect 97549 8449 97583 8483
rect 97365 8313 97399 8347
rect 8953 5865 8987 5899
rect 12173 5865 12207 5899
rect 50905 5865 50939 5899
rect 51089 5865 51123 5899
rect 10057 5729 10091 5763
rect 52009 5729 52043 5763
rect 11161 5661 11195 5695
rect 53113 5661 53147 5695
rect 54217 5593 54251 5627
rect 13185 3145 13219 3179
rect 12909 3077 12943 3111
rect 11713 3009 11747 3043
rect 11621 2805 11655 2839
rect 89545 2805 89579 2839
rect 11621 2601 11655 2635
rect 32321 2601 32355 2635
rect 33149 2601 33183 2635
rect 34253 2601 34287 2635
rect 35541 2601 35575 2635
rect 36829 2601 36863 2635
rect 37657 2601 37691 2635
rect 38761 2601 38795 2635
rect 40049 2601 40083 2635
rect 40877 2601 40911 2635
rect 41981 2601 42015 2635
rect 43269 2601 43303 2635
rect 48789 2601 48823 2635
rect 74181 2601 74215 2635
rect 75469 2601 75503 2635
rect 76297 2601 76331 2635
rect 77401 2601 77435 2635
rect 78689 2601 78723 2635
rect 79517 2601 79551 2635
rect 80805 2601 80839 2635
rect 81909 2601 81943 2635
rect 83197 2601 83231 2635
rect 84025 2601 84059 2635
rect 85129 2601 85163 2635
rect 44557 2533 44591 2567
rect 86417 2533 86451 2567
rect 10885 2465 10919 2499
rect 12817 2465 12851 2499
rect 13829 2465 13863 2499
rect 45477 2465 45511 2499
rect 46765 2465 46799 2499
rect 48053 2465 48087 2499
rect 87337 2465 87371 2499
rect 89085 2465 89119 2499
rect 90005 2465 90039 2499
rect 11161 2397 11195 2431
rect 11805 2397 11839 2431
rect 12357 2397 12391 2431
rect 14565 2397 14599 2431
rect 15577 2397 15611 2431
rect 16865 2397 16899 2431
rect 17785 2397 17819 2431
rect 18797 2397 18831 2431
rect 20085 2397 20119 2431
rect 21373 2397 21407 2431
rect 22293 2397 22327 2431
rect 23305 2397 23339 2431
rect 24593 2397 24627 2431
rect 25513 2397 25547 2431
rect 26525 2397 26559 2431
rect 27813 2397 27847 2431
rect 29101 2397 29135 2431
rect 30021 2397 30055 2431
rect 31033 2397 31067 2431
rect 32505 2397 32539 2431
rect 32965 2397 32999 2431
rect 34437 2397 34471 2431
rect 35725 2397 35759 2431
rect 37013 2397 37047 2431
rect 37473 2397 37507 2431
rect 38945 2397 38979 2431
rect 40233 2397 40267 2431
rect 40693 2397 40727 2431
rect 42165 2397 42199 2431
rect 43453 2397 43487 2431
rect 45201 2397 45235 2431
rect 46489 2397 46523 2431
rect 47777 2397 47811 2431
rect 48973 2397 49007 2431
rect 56425 2397 56459 2431
rect 57437 2397 57471 2431
rect 58725 2397 58759 2431
rect 60013 2397 60047 2431
rect 60933 2397 60967 2431
rect 61945 2397 61979 2431
rect 63233 2397 63267 2431
rect 64153 2397 64187 2431
rect 65165 2397 65199 2431
rect 66453 2397 66487 2431
rect 67741 2397 67775 2431
rect 68661 2397 68695 2431
rect 69673 2397 69707 2431
rect 70961 2397 70995 2431
rect 71881 2397 71915 2431
rect 72893 2397 72927 2431
rect 74365 2397 74399 2431
rect 75653 2397 75687 2431
rect 76113 2397 76147 2431
rect 77585 2397 77619 2431
rect 78873 2397 78907 2431
rect 79333 2397 79367 2431
rect 80621 2397 80655 2431
rect 82093 2397 82127 2431
rect 83381 2397 83415 2431
rect 83841 2397 83875 2431
rect 85313 2397 85347 2431
rect 87061 2397 87095 2431
rect 88809 2397 88843 2431
rect 89729 2397 89763 2431
rect 44741 2329 44775 2363
rect 86601 2329 86635 2363
rect 12265 2261 12299 2295
rect 14381 2261 14415 2295
rect 15761 2261 15795 2295
rect 17049 2261 17083 2295
rect 17601 2261 17635 2295
rect 18981 2261 19015 2295
rect 20269 2261 20303 2295
rect 21557 2261 21591 2295
rect 22109 2261 22143 2295
rect 23489 2261 23523 2295
rect 24777 2261 24811 2295
rect 25329 2261 25363 2295
rect 26709 2261 26743 2295
rect 27997 2261 28031 2295
rect 29285 2261 29319 2295
rect 29837 2261 29871 2295
rect 31217 2261 31251 2295
rect 32229 2261 32263 2295
rect 32873 2261 32907 2295
rect 34161 2261 34195 2295
rect 35449 2261 35483 2295
rect 36737 2261 36771 2295
rect 37381 2261 37415 2295
rect 38669 2261 38703 2295
rect 39957 2261 39991 2295
rect 40601 2261 40635 2295
rect 41889 2261 41923 2295
rect 43177 2261 43211 2295
rect 44465 2261 44499 2295
rect 45109 2261 45143 2295
rect 46397 2261 46431 2295
rect 47685 2261 47719 2295
rect 49065 2261 49099 2295
rect 56241 2261 56275 2295
rect 57621 2261 57655 2295
rect 58909 2261 58943 2295
rect 60197 2261 60231 2295
rect 60749 2261 60783 2295
rect 62129 2261 62163 2295
rect 63417 2261 63451 2295
rect 63969 2261 64003 2295
rect 65349 2261 65383 2295
rect 66637 2261 66671 2295
rect 67925 2261 67959 2295
rect 68477 2261 68511 2295
rect 69857 2261 69891 2295
rect 71145 2261 71179 2295
rect 71697 2261 71731 2295
rect 73077 2261 73111 2295
rect 74089 2261 74123 2295
rect 75377 2261 75411 2295
rect 76021 2261 76055 2295
rect 77309 2261 77343 2295
rect 78597 2261 78631 2295
rect 79241 2261 79275 2295
rect 80529 2261 80563 2295
rect 81817 2261 81851 2295
rect 83105 2261 83139 2295
rect 83749 2261 83783 2295
rect 85037 2261 85071 2295
rect 86325 2261 86359 2295
rect 86969 2261 87003 2295
rect 88533 2261 88567 2295
<< metal1 >>
rect 1104 95770 97888 95792
rect 1104 95718 4874 95770
rect 4926 95718 4938 95770
rect 4990 95718 5002 95770
rect 5054 95718 5066 95770
rect 5118 95718 5130 95770
rect 5182 95718 35594 95770
rect 35646 95718 35658 95770
rect 35710 95718 35722 95770
rect 35774 95718 35786 95770
rect 35838 95718 35850 95770
rect 35902 95718 66314 95770
rect 66366 95718 66378 95770
rect 66430 95718 66442 95770
rect 66494 95718 66506 95770
rect 66558 95718 66570 95770
rect 66622 95718 97034 95770
rect 97086 95718 97098 95770
rect 97150 95718 97162 95770
rect 97214 95718 97226 95770
rect 97278 95718 97290 95770
rect 97342 95718 97888 95770
rect 1104 95696 97888 95718
rect 14090 95616 14096 95668
rect 14148 95616 14154 95668
rect 15378 95616 15384 95668
rect 15436 95616 15442 95668
rect 16666 95616 16672 95668
rect 16724 95616 16730 95668
rect 17310 95616 17316 95668
rect 17368 95656 17374 95668
rect 17368 95628 17632 95656
rect 17368 95616 17374 95628
rect 14108 95520 14136 95616
rect 14277 95523 14335 95529
rect 14277 95520 14289 95523
rect 14108 95492 14289 95520
rect 14277 95489 14289 95492
rect 14323 95489 14335 95523
rect 15396 95520 15424 95616
rect 15565 95523 15623 95529
rect 15565 95520 15577 95523
rect 15396 95492 15577 95520
rect 14277 95483 14335 95489
rect 15565 95489 15577 95492
rect 15611 95489 15623 95523
rect 16684 95520 16712 95616
rect 17604 95597 17632 95628
rect 18598 95616 18604 95668
rect 18656 95656 18662 95668
rect 18656 95628 19012 95656
rect 18656 95616 18662 95628
rect 18984 95597 19012 95628
rect 19886 95616 19892 95668
rect 19944 95656 19950 95668
rect 19944 95628 20300 95656
rect 19944 95616 19950 95628
rect 20272 95597 20300 95628
rect 21174 95616 21180 95668
rect 21232 95656 21238 95668
rect 21232 95628 21588 95656
rect 21232 95616 21238 95628
rect 21560 95597 21588 95628
rect 21818 95616 21824 95668
rect 21876 95616 21882 95668
rect 23106 95616 23112 95668
rect 23164 95656 23170 95668
rect 23164 95628 23520 95656
rect 23164 95616 23170 95628
rect 17589 95591 17647 95597
rect 17589 95557 17601 95591
rect 17635 95557 17647 95591
rect 17589 95551 17647 95557
rect 18969 95591 19027 95597
rect 18969 95557 18981 95591
rect 19015 95557 19027 95591
rect 18969 95551 19027 95557
rect 20257 95591 20315 95597
rect 20257 95557 20269 95591
rect 20303 95557 20315 95591
rect 20257 95551 20315 95557
rect 21545 95591 21603 95597
rect 21545 95557 21557 95591
rect 21591 95557 21603 95591
rect 21545 95551 21603 95557
rect 16853 95523 16911 95529
rect 16853 95520 16865 95523
rect 16684 95492 16865 95520
rect 15565 95483 15623 95489
rect 16853 95489 16865 95492
rect 16899 95489 16911 95523
rect 21836 95520 21864 95616
rect 23492 95597 23520 95628
rect 25038 95616 25044 95668
rect 25096 95616 25102 95668
rect 26326 95616 26332 95668
rect 26384 95616 26390 95668
rect 27614 95616 27620 95668
rect 27672 95616 27678 95668
rect 28997 95659 29055 95665
rect 28997 95625 29009 95659
rect 29043 95656 29055 95659
rect 29086 95656 29092 95668
rect 29043 95628 29092 95656
rect 29043 95625 29055 95628
rect 28997 95619 29055 95625
rect 29086 95616 29092 95628
rect 29144 95616 29150 95668
rect 29546 95616 29552 95668
rect 29604 95616 29610 95668
rect 30834 95616 30840 95668
rect 30892 95616 30898 95668
rect 32490 95616 32496 95668
rect 32548 95616 32554 95668
rect 33042 95616 33048 95668
rect 33100 95616 33106 95668
rect 34422 95616 34428 95668
rect 34480 95616 34486 95668
rect 35342 95616 35348 95668
rect 35400 95656 35406 95668
rect 35713 95659 35771 95665
rect 35713 95656 35725 95659
rect 35400 95628 35725 95656
rect 35400 95616 35406 95628
rect 35713 95625 35725 95628
rect 35759 95625 35771 95659
rect 35713 95619 35771 95625
rect 36998 95616 37004 95668
rect 37056 95616 37062 95668
rect 37550 95616 37556 95668
rect 37608 95616 37614 95668
rect 38930 95616 38936 95668
rect 38988 95616 38994 95668
rect 39850 95616 39856 95668
rect 39908 95656 39914 95668
rect 40221 95659 40279 95665
rect 40221 95656 40233 95659
rect 39908 95628 40233 95656
rect 39908 95616 39914 95628
rect 40221 95625 40233 95628
rect 40267 95625 40279 95659
rect 40221 95619 40279 95625
rect 40770 95616 40776 95668
rect 40828 95616 40834 95668
rect 42150 95616 42156 95668
rect 42208 95616 42214 95668
rect 43438 95616 43444 95668
rect 43496 95616 43502 95668
rect 44726 95616 44732 95668
rect 44784 95616 44790 95668
rect 45278 95616 45284 95668
rect 45336 95616 45342 95668
rect 46658 95616 46664 95668
rect 46716 95616 46722 95668
rect 47946 95616 47952 95668
rect 48004 95616 48010 95668
rect 48498 95616 48504 95668
rect 48556 95616 48562 95668
rect 50893 95659 50951 95665
rect 50893 95625 50905 95659
rect 50939 95656 50951 95659
rect 50982 95656 50988 95668
rect 50939 95628 50988 95656
rect 50939 95625 50951 95628
rect 50893 95619 50951 95625
rect 50982 95616 50988 95628
rect 51040 95616 51046 95668
rect 54386 95616 54392 95668
rect 54444 95656 54450 95668
rect 55033 95659 55091 95665
rect 55033 95656 55045 95659
rect 54444 95628 55045 95656
rect 54444 95616 54450 95628
rect 55033 95625 55045 95628
rect 55079 95656 55091 95659
rect 55079 95628 55214 95656
rect 55079 95625 55091 95628
rect 55033 95619 55091 95625
rect 23477 95591 23535 95597
rect 23477 95557 23489 95591
rect 23523 95557 23535 95591
rect 23477 95551 23535 95557
rect 22005 95523 22063 95529
rect 22005 95520 22017 95523
rect 21836 95492 22017 95520
rect 16853 95483 16911 95489
rect 22005 95489 22017 95492
rect 22051 95489 22063 95523
rect 25056 95520 25084 95616
rect 25225 95523 25283 95529
rect 25225 95520 25237 95523
rect 25056 95492 25237 95520
rect 22005 95483 22063 95489
rect 25225 95489 25237 95492
rect 25271 95489 25283 95523
rect 26344 95520 26372 95616
rect 26697 95523 26755 95529
rect 26697 95520 26709 95523
rect 26344 95492 26709 95520
rect 25225 95483 25283 95489
rect 26697 95489 26709 95492
rect 26743 95489 26755 95523
rect 27632 95520 27660 95616
rect 27985 95523 28043 95529
rect 27985 95520 27997 95523
rect 27632 95492 27997 95520
rect 26697 95483 26755 95489
rect 27985 95489 27997 95492
rect 28031 95489 28043 95523
rect 29104 95520 29132 95616
rect 29273 95523 29331 95529
rect 29273 95520 29285 95523
rect 29104 95492 29285 95520
rect 27985 95483 28043 95489
rect 29273 95489 29285 95492
rect 29319 95489 29331 95523
rect 29564 95520 29592 95616
rect 29733 95523 29791 95529
rect 29733 95520 29745 95523
rect 29564 95492 29745 95520
rect 29273 95483 29331 95489
rect 29733 95489 29745 95492
rect 29779 95489 29791 95523
rect 30852 95520 30880 95616
rect 31205 95523 31263 95529
rect 31205 95520 31217 95523
rect 30852 95492 31217 95520
rect 29733 95483 29791 95489
rect 31205 95489 31217 95492
rect 31251 95489 31263 95523
rect 31205 95483 31263 95489
rect 32306 95480 32312 95532
rect 32364 95480 32370 95532
rect 33226 95480 33232 95532
rect 33284 95480 33290 95532
rect 34238 95480 34244 95532
rect 34296 95480 34302 95532
rect 35342 95480 35348 95532
rect 35400 95520 35406 95532
rect 35529 95523 35587 95529
rect 35529 95520 35541 95523
rect 35400 95492 35541 95520
rect 35400 95480 35406 95492
rect 35529 95489 35541 95492
rect 35575 95489 35587 95523
rect 35529 95483 35587 95489
rect 36446 95480 36452 95532
rect 36504 95520 36510 95532
rect 36817 95523 36875 95529
rect 36817 95520 36829 95523
rect 36504 95492 36829 95520
rect 36504 95480 36510 95492
rect 36817 95489 36829 95492
rect 36863 95489 36875 95523
rect 36817 95483 36875 95489
rect 37734 95480 37740 95532
rect 37792 95480 37798 95532
rect 38746 95480 38752 95532
rect 38804 95480 38810 95532
rect 39758 95480 39764 95532
rect 39816 95520 39822 95532
rect 40037 95523 40095 95529
rect 40037 95520 40049 95523
rect 39816 95492 40049 95520
rect 39816 95480 39822 95492
rect 40037 95489 40049 95492
rect 40083 95489 40095 95523
rect 40037 95483 40095 95489
rect 40954 95480 40960 95532
rect 41012 95480 41018 95532
rect 41966 95480 41972 95532
rect 42024 95480 42030 95532
rect 43254 95480 43260 95532
rect 43312 95480 43318 95532
rect 44174 95480 44180 95532
rect 44232 95520 44238 95532
rect 44545 95523 44603 95529
rect 44545 95520 44557 95523
rect 44232 95492 44557 95520
rect 44232 95480 44238 95492
rect 44545 95489 44557 95492
rect 44591 95489 44603 95523
rect 44545 95483 44603 95489
rect 45462 95480 45468 95532
rect 45520 95480 45526 95532
rect 46474 95480 46480 95532
rect 46532 95480 46538 95532
rect 47762 95480 47768 95532
rect 47820 95480 47826 95532
rect 48682 95480 48688 95532
rect 48740 95480 48746 95532
rect 51074 95480 51080 95532
rect 51132 95480 51138 95532
rect 51810 95480 51816 95532
rect 51868 95520 51874 95532
rect 52457 95523 52515 95529
rect 52457 95520 52469 95523
rect 51868 95492 52469 95520
rect 51868 95480 51874 95492
rect 52457 95489 52469 95492
rect 52503 95520 52515 95523
rect 52733 95523 52791 95529
rect 52733 95520 52745 95523
rect 52503 95492 52745 95520
rect 52503 95489 52515 95492
rect 52457 95483 52515 95489
rect 52733 95489 52745 95492
rect 52779 95489 52791 95523
rect 52733 95483 52791 95489
rect 52914 95480 52920 95532
rect 52972 95480 52978 95532
rect 55186 95520 55214 95628
rect 56410 95616 56416 95668
rect 56468 95656 56474 95668
rect 57149 95659 57207 95665
rect 57149 95656 57161 95659
rect 56468 95628 57161 95656
rect 56468 95616 56474 95628
rect 57072 95529 57100 95628
rect 57149 95625 57161 95628
rect 57195 95625 57207 95659
rect 57149 95619 57207 95625
rect 58526 95616 58532 95668
rect 58584 95616 58590 95668
rect 59814 95616 59820 95668
rect 59872 95656 59878 95668
rect 59872 95628 60228 95656
rect 59872 95616 59878 95628
rect 55309 95523 55367 95529
rect 55309 95520 55321 95523
rect 55186 95492 55321 95520
rect 55309 95489 55321 95492
rect 55355 95489 55367 95523
rect 55309 95483 55367 95489
rect 57057 95523 57115 95529
rect 57057 95489 57069 95523
rect 57103 95489 57115 95523
rect 57057 95483 57115 95489
rect 57698 95480 57704 95532
rect 57756 95520 57762 95532
rect 57885 95523 57943 95529
rect 57885 95520 57897 95523
rect 57756 95492 57897 95520
rect 57756 95480 57762 95492
rect 57885 95489 57897 95492
rect 57931 95489 57943 95523
rect 58544 95520 58572 95616
rect 60200 95597 60228 95628
rect 60458 95616 60464 95668
rect 60516 95656 60522 95668
rect 60516 95628 60780 95656
rect 60516 95616 60522 95628
rect 60752 95597 60780 95628
rect 61746 95616 61752 95668
rect 61804 95656 61810 95668
rect 61804 95628 62160 95656
rect 61804 95616 61810 95628
rect 62132 95597 62160 95628
rect 63034 95616 63040 95668
rect 63092 95656 63098 95668
rect 63092 95628 63448 95656
rect 63092 95616 63098 95628
rect 63420 95597 63448 95628
rect 63678 95616 63684 95668
rect 63736 95616 63742 95668
rect 64966 95616 64972 95668
rect 65024 95656 65030 95668
rect 66349 95659 66407 95665
rect 65024 95628 65380 95656
rect 65024 95616 65030 95628
rect 60185 95591 60243 95597
rect 60185 95557 60197 95591
rect 60231 95557 60243 95591
rect 60185 95551 60243 95557
rect 60737 95591 60795 95597
rect 60737 95557 60749 95591
rect 60783 95557 60795 95591
rect 60737 95551 60795 95557
rect 62117 95591 62175 95597
rect 62117 95557 62129 95591
rect 62163 95557 62175 95591
rect 62117 95551 62175 95557
rect 63405 95591 63463 95597
rect 63405 95557 63417 95591
rect 63451 95557 63463 95591
rect 63405 95551 63463 95557
rect 58713 95523 58771 95529
rect 58713 95520 58725 95523
rect 58544 95492 58725 95520
rect 57885 95483 57943 95489
rect 58713 95489 58725 95492
rect 58759 95489 58771 95523
rect 63696 95520 63724 95616
rect 65352 95597 65380 95628
rect 66349 95625 66361 95659
rect 66395 95656 66407 95659
rect 66714 95656 66720 95668
rect 66395 95628 66720 95656
rect 66395 95625 66407 95628
rect 66349 95619 66407 95625
rect 65337 95591 65395 95597
rect 65337 95557 65349 95591
rect 65383 95557 65395 95591
rect 65337 95551 65395 95557
rect 66456 95529 66484 95628
rect 66714 95616 66720 95628
rect 66772 95616 66778 95668
rect 67910 95616 67916 95668
rect 67968 95616 67974 95668
rect 68554 95616 68560 95668
rect 68612 95656 68618 95668
rect 69385 95659 69443 95665
rect 69385 95656 69397 95659
rect 68612 95628 69397 95656
rect 68612 95616 68618 95628
rect 63865 95523 63923 95529
rect 63865 95520 63877 95523
rect 63696 95492 63877 95520
rect 58713 95483 58771 95489
rect 63865 95489 63877 95492
rect 63911 95489 63923 95523
rect 63865 95483 63923 95489
rect 66441 95523 66499 95529
rect 66441 95489 66453 95523
rect 66487 95489 66499 95523
rect 67928 95520 67956 95616
rect 69308 95529 69336 95628
rect 69385 95625 69397 95628
rect 69431 95625 69443 95659
rect 69385 95619 69443 95625
rect 69842 95616 69848 95668
rect 69900 95656 69906 95668
rect 69937 95659 69995 95665
rect 69937 95656 69949 95659
rect 69900 95628 69949 95656
rect 69900 95616 69906 95628
rect 69937 95625 69949 95628
rect 69983 95625 69995 95659
rect 69937 95619 69995 95625
rect 70762 95616 70768 95668
rect 70820 95616 70826 95668
rect 71406 95616 71412 95668
rect 71464 95616 71470 95668
rect 72694 95616 72700 95668
rect 72752 95616 72758 95668
rect 74350 95616 74356 95668
rect 74408 95616 74414 95668
rect 75638 95616 75644 95668
rect 75696 95616 75702 95668
rect 76190 95616 76196 95668
rect 76248 95616 76254 95668
rect 77570 95616 77576 95668
rect 77628 95616 77634 95668
rect 78490 95616 78496 95668
rect 78548 95656 78554 95668
rect 78861 95659 78919 95665
rect 78861 95656 78873 95659
rect 78548 95628 78873 95656
rect 78548 95616 78554 95628
rect 78861 95625 78873 95628
rect 78907 95625 78919 95659
rect 78861 95619 78919 95625
rect 79410 95616 79416 95668
rect 79468 95616 79474 95668
rect 80790 95616 80796 95668
rect 80848 95616 80854 95668
rect 82078 95616 82084 95668
rect 82136 95616 82142 95668
rect 83366 95616 83372 95668
rect 83424 95616 83430 95668
rect 83918 95616 83924 95668
rect 83976 95616 83982 95668
rect 85298 95616 85304 95668
rect 85356 95616 85362 95668
rect 86586 95616 86592 95668
rect 86644 95616 86650 95668
rect 87138 95616 87144 95668
rect 87196 95616 87202 95668
rect 88150 95616 88156 95668
rect 88208 95656 88214 95668
rect 88521 95659 88579 95665
rect 88521 95656 88533 95659
rect 88208 95628 88533 95656
rect 88208 95616 88214 95628
rect 88521 95625 88533 95628
rect 88567 95625 88579 95659
rect 88521 95619 88579 95625
rect 89622 95616 89628 95668
rect 89680 95656 89686 95668
rect 89809 95659 89867 95665
rect 89809 95656 89821 95659
rect 89680 95628 89821 95656
rect 89680 95616 89686 95628
rect 89809 95625 89821 95628
rect 89855 95625 89867 95659
rect 89809 95619 89867 95625
rect 91002 95616 91008 95668
rect 91060 95656 91066 95668
rect 91097 95659 91155 95665
rect 91097 95656 91109 95659
rect 91060 95628 91109 95656
rect 91060 95616 91066 95628
rect 91097 95625 91109 95628
rect 91143 95625 91155 95659
rect 91097 95619 91155 95625
rect 69860 95529 69888 95616
rect 68189 95523 68247 95529
rect 68189 95520 68201 95523
rect 67928 95492 68201 95520
rect 66441 95483 66499 95489
rect 68189 95489 68201 95492
rect 68235 95489 68247 95523
rect 68189 95483 68247 95489
rect 69293 95523 69351 95529
rect 69293 95489 69305 95523
rect 69339 95489 69351 95523
rect 69293 95483 69351 95489
rect 69845 95523 69903 95529
rect 69845 95489 69857 95523
rect 69891 95489 69903 95523
rect 70780 95520 70808 95616
rect 71133 95523 71191 95529
rect 71133 95520 71145 95523
rect 70780 95492 71145 95520
rect 69845 95483 69903 95489
rect 71133 95489 71145 95492
rect 71179 95489 71191 95523
rect 71424 95520 71452 95616
rect 71593 95523 71651 95529
rect 71593 95520 71605 95523
rect 71424 95492 71605 95520
rect 71133 95483 71191 95489
rect 71593 95489 71605 95492
rect 71639 95489 71651 95523
rect 72712 95520 72740 95616
rect 72881 95523 72939 95529
rect 72881 95520 72893 95523
rect 72712 95492 72893 95520
rect 71593 95483 71651 95489
rect 72881 95489 72893 95492
rect 72927 95489 72939 95523
rect 72881 95483 72939 95489
rect 74166 95480 74172 95532
rect 74224 95480 74230 95532
rect 75454 95480 75460 95532
rect 75512 95480 75518 95532
rect 76374 95480 76380 95532
rect 76432 95480 76438 95532
rect 77386 95480 77392 95532
rect 77444 95480 77450 95532
rect 78582 95480 78588 95532
rect 78640 95520 78646 95532
rect 78677 95523 78735 95529
rect 78677 95520 78689 95523
rect 78640 95492 78689 95520
rect 78640 95480 78646 95492
rect 78677 95489 78689 95492
rect 78723 95489 78735 95523
rect 78677 95483 78735 95489
rect 79594 95480 79600 95532
rect 79652 95480 79658 95532
rect 80606 95480 80612 95532
rect 80664 95480 80670 95532
rect 81894 95480 81900 95532
rect 81952 95480 81958 95532
rect 83182 95480 83188 95532
rect 83240 95480 83246 95532
rect 84102 95480 84108 95532
rect 84160 95480 84166 95532
rect 85114 95480 85120 95532
rect 85172 95480 85178 95532
rect 86402 95480 86408 95532
rect 86460 95480 86466 95532
rect 87322 95480 87328 95532
rect 87380 95480 87386 95532
rect 88334 95480 88340 95532
rect 88392 95480 88398 95532
rect 89622 95480 89628 95532
rect 89680 95480 89686 95532
rect 90910 95480 90916 95532
rect 90968 95480 90974 95532
rect 25498 95412 25504 95464
rect 25556 95412 25562 95464
rect 52089 95455 52147 95461
rect 52089 95421 52101 95455
rect 52135 95452 52147 95455
rect 52362 95452 52368 95464
rect 52135 95424 52368 95452
rect 52135 95421 52147 95424
rect 52089 95415 52147 95421
rect 52362 95412 52368 95424
rect 52420 95412 52426 95464
rect 54110 95412 54116 95464
rect 54168 95452 54174 95464
rect 54389 95455 54447 95461
rect 54389 95452 54401 95455
rect 54168 95424 54401 95452
rect 54168 95412 54174 95424
rect 54389 95421 54401 95424
rect 54435 95421 54447 95455
rect 54389 95415 54447 95421
rect 56505 95455 56563 95461
rect 56505 95421 56517 95455
rect 56551 95452 56563 95455
rect 56778 95452 56784 95464
rect 56551 95424 56784 95452
rect 56551 95421 56563 95424
rect 56505 95415 56563 95421
rect 56778 95412 56784 95424
rect 56836 95412 56842 95464
rect 66714 95412 66720 95464
rect 66772 95412 66778 95464
rect 67450 95412 67456 95464
rect 67508 95452 67514 95464
rect 68465 95455 68523 95461
rect 68465 95452 68477 95455
rect 67508 95424 68477 95452
rect 67508 95412 67514 95424
rect 68465 95421 68477 95424
rect 68511 95421 68523 95455
rect 68465 95415 68523 95421
rect 18782 95344 18788 95396
rect 18840 95344 18846 95396
rect 20070 95344 20076 95396
rect 20128 95344 20134 95396
rect 20990 95344 20996 95396
rect 21048 95384 21054 95396
rect 21361 95387 21419 95393
rect 21361 95384 21373 95387
rect 21048 95356 21373 95384
rect 21048 95344 21054 95356
rect 21361 95353 21373 95356
rect 21407 95353 21419 95387
rect 21361 95347 21419 95353
rect 23290 95344 23296 95396
rect 23348 95344 23354 95396
rect 28718 95344 28724 95396
rect 28776 95384 28782 95396
rect 29089 95387 29147 95393
rect 29089 95384 29101 95387
rect 28776 95356 29101 95384
rect 28776 95344 28782 95356
rect 29089 95353 29101 95356
rect 29135 95353 29147 95387
rect 29089 95347 29147 95353
rect 59998 95344 60004 95396
rect 60056 95344 60062 95396
rect 61930 95344 61936 95396
rect 61988 95344 61994 95396
rect 63218 95344 63224 95396
rect 63276 95344 63282 95396
rect 14458 95276 14464 95328
rect 14516 95276 14522 95328
rect 15746 95276 15752 95328
rect 15804 95276 15810 95328
rect 16574 95276 16580 95328
rect 16632 95316 16638 95328
rect 17037 95319 17095 95325
rect 17037 95316 17049 95319
rect 16632 95288 17049 95316
rect 16632 95276 16638 95288
rect 17037 95285 17049 95288
rect 17083 95285 17095 95319
rect 17037 95279 17095 95285
rect 17678 95276 17684 95328
rect 17736 95276 17742 95328
rect 22186 95276 22192 95328
rect 22244 95276 22250 95328
rect 26510 95276 26516 95328
rect 26568 95276 26574 95328
rect 27798 95276 27804 95328
rect 27856 95276 27862 95328
rect 29914 95276 29920 95328
rect 29972 95276 29978 95328
rect 31018 95276 31024 95328
rect 31076 95276 31082 95328
rect 56502 95276 56508 95328
rect 56560 95316 56566 95328
rect 56873 95319 56931 95325
rect 56873 95316 56885 95319
rect 56560 95288 56885 95316
rect 56560 95276 56566 95288
rect 56873 95285 56885 95288
rect 56919 95285 56931 95319
rect 56873 95279 56931 95285
rect 57514 95276 57520 95328
rect 57572 95276 57578 95328
rect 58894 95276 58900 95328
rect 58952 95276 58958 95328
rect 60826 95276 60832 95328
rect 60884 95276 60890 95328
rect 64046 95276 64052 95328
rect 64104 95276 64110 95328
rect 65242 95276 65248 95328
rect 65300 95276 65306 95328
rect 68830 95276 68836 95328
rect 68888 95316 68894 95328
rect 69109 95319 69167 95325
rect 69109 95316 69121 95319
rect 68888 95288 69121 95316
rect 68888 95276 68894 95288
rect 69109 95285 69121 95288
rect 69155 95285 69167 95319
rect 69109 95279 69167 95285
rect 69658 95276 69664 95328
rect 69716 95276 69722 95328
rect 70946 95276 70952 95328
rect 71004 95276 71010 95328
rect 71774 95276 71780 95328
rect 71832 95276 71838 95328
rect 73062 95276 73068 95328
rect 73120 95276 73126 95328
rect 1104 95226 97888 95248
rect 1104 95174 4214 95226
rect 4266 95174 4278 95226
rect 4330 95174 4342 95226
rect 4394 95174 4406 95226
rect 4458 95174 4470 95226
rect 4522 95174 34934 95226
rect 34986 95174 34998 95226
rect 35050 95174 35062 95226
rect 35114 95174 35126 95226
rect 35178 95174 35190 95226
rect 35242 95174 65654 95226
rect 65706 95174 65718 95226
rect 65770 95174 65782 95226
rect 65834 95174 65846 95226
rect 65898 95174 65910 95226
rect 65962 95174 96374 95226
rect 96426 95174 96438 95226
rect 96490 95174 96502 95226
rect 96554 95174 96566 95226
rect 96618 95174 96630 95226
rect 96682 95174 97888 95226
rect 1104 95152 97888 95174
rect 24394 95072 24400 95124
rect 24452 95072 24458 95124
rect 52825 95115 52883 95121
rect 52825 95081 52837 95115
rect 52871 95112 52883 95115
rect 52914 95112 52920 95124
rect 52871 95084 52920 95112
rect 52871 95081 52883 95084
rect 52825 95075 52883 95081
rect 52914 95072 52920 95084
rect 52972 95072 52978 95124
rect 56778 95072 56784 95124
rect 56836 95072 56842 95124
rect 24412 94976 24440 95072
rect 24581 94979 24639 94985
rect 24581 94976 24593 94979
rect 24412 94948 24593 94976
rect 24581 94945 24593 94948
rect 24627 94945 24639 94979
rect 24581 94939 24639 94945
rect 52454 94936 52460 94988
rect 52512 94976 52518 94988
rect 52914 94976 52920 94988
rect 52512 94948 52920 94976
rect 52512 94936 52518 94948
rect 52914 94936 52920 94948
rect 52972 94936 52978 94988
rect 24302 94868 24308 94920
rect 24360 94908 24366 94920
rect 24857 94911 24915 94917
rect 24857 94908 24869 94911
rect 24360 94880 24869 94908
rect 24360 94868 24366 94880
rect 24857 94877 24869 94880
rect 24903 94877 24915 94911
rect 24857 94871 24915 94877
rect 51074 94732 51080 94784
rect 51132 94772 51138 94784
rect 51169 94775 51227 94781
rect 51169 94772 51181 94775
rect 51132 94744 51181 94772
rect 51132 94732 51138 94744
rect 51169 94741 51181 94744
rect 51215 94741 51227 94775
rect 51169 94735 51227 94741
rect 1104 94682 97888 94704
rect 1104 94630 4874 94682
rect 4926 94630 4938 94682
rect 4990 94630 5002 94682
rect 5054 94630 5066 94682
rect 5118 94630 5130 94682
rect 5182 94630 35594 94682
rect 35646 94630 35658 94682
rect 35710 94630 35722 94682
rect 35774 94630 35786 94682
rect 35838 94630 35850 94682
rect 35902 94630 66314 94682
rect 66366 94630 66378 94682
rect 66430 94630 66442 94682
rect 66494 94630 66506 94682
rect 66558 94630 66570 94682
rect 66622 94630 97034 94682
rect 97086 94630 97098 94682
rect 97150 94630 97162 94682
rect 97214 94630 97226 94682
rect 97278 94630 97290 94682
rect 97342 94630 97888 94682
rect 1104 94608 97888 94630
rect 1104 94138 97888 94160
rect 1104 94086 4214 94138
rect 4266 94086 4278 94138
rect 4330 94086 4342 94138
rect 4394 94086 4406 94138
rect 4458 94086 4470 94138
rect 4522 94086 34934 94138
rect 34986 94086 34998 94138
rect 35050 94086 35062 94138
rect 35114 94086 35126 94138
rect 35178 94086 35190 94138
rect 35242 94086 65654 94138
rect 65706 94086 65718 94138
rect 65770 94086 65782 94138
rect 65834 94086 65846 94138
rect 65898 94086 65910 94138
rect 65962 94086 96374 94138
rect 96426 94086 96438 94138
rect 96490 94086 96502 94138
rect 96554 94086 96566 94138
rect 96618 94086 96630 94138
rect 96682 94086 97888 94138
rect 1104 94064 97888 94086
rect 54110 93984 54116 94036
rect 54168 94024 54174 94036
rect 54573 94027 54631 94033
rect 54573 94024 54585 94027
rect 54168 93996 54585 94024
rect 54168 93984 54174 93996
rect 54573 93993 54585 93996
rect 54619 93993 54631 94027
rect 54573 93987 54631 93993
rect 54757 93959 54815 93965
rect 54757 93956 54769 93959
rect 54312 93928 54769 93956
rect 54110 93888 54116 93900
rect 53852 93860 54116 93888
rect 52546 93780 52552 93832
rect 52604 93820 52610 93832
rect 53101 93823 53159 93829
rect 53101 93820 53113 93823
rect 52604 93792 53113 93820
rect 52604 93780 52610 93792
rect 53101 93789 53113 93792
rect 53147 93820 53159 93823
rect 53852 93820 53880 93860
rect 54110 93848 54116 93860
rect 54168 93848 54174 93900
rect 54312 93897 54340 93928
rect 54757 93925 54769 93928
rect 54803 93956 54815 93959
rect 54803 93928 55214 93956
rect 54803 93925 54815 93928
rect 54757 93919 54815 93925
rect 54297 93891 54355 93897
rect 54297 93857 54309 93891
rect 54343 93857 54355 93891
rect 55186 93888 55214 93928
rect 91646 93888 91652 93900
rect 55186 93860 91652 93888
rect 54297 93851 54355 93857
rect 91646 93848 91652 93860
rect 91704 93848 91710 93900
rect 53147 93792 53880 93820
rect 53147 93789 53159 93792
rect 53101 93783 53159 93789
rect 1104 93594 97888 93616
rect 1104 93542 4874 93594
rect 4926 93542 4938 93594
rect 4990 93542 5002 93594
rect 5054 93542 5066 93594
rect 5118 93542 5130 93594
rect 5182 93542 35594 93594
rect 35646 93542 35658 93594
rect 35710 93542 35722 93594
rect 35774 93542 35786 93594
rect 35838 93542 35850 93594
rect 35902 93542 66314 93594
rect 66366 93542 66378 93594
rect 66430 93542 66442 93594
rect 66494 93542 66506 93594
rect 66558 93542 66570 93594
rect 66622 93542 97034 93594
rect 97086 93542 97098 93594
rect 97150 93542 97162 93594
rect 97214 93542 97226 93594
rect 97278 93542 97290 93594
rect 97342 93542 97888 93594
rect 1104 93520 97888 93542
rect 56778 93480 56784 93492
rect 56704 93452 56784 93480
rect 31665 93347 31723 93353
rect 31665 93313 31677 93347
rect 31711 93344 31723 93347
rect 31846 93344 31852 93356
rect 31711 93316 31852 93344
rect 31711 93313 31723 93316
rect 31665 93307 31723 93313
rect 31846 93304 31852 93316
rect 31904 93304 31910 93356
rect 40497 93347 40555 93353
rect 40497 93344 40509 93347
rect 40328 93316 40509 93344
rect 40328 93285 40356 93316
rect 40497 93313 40509 93316
rect 40543 93313 40555 93347
rect 52733 93347 52791 93353
rect 52733 93344 52745 93347
rect 40497 93307 40555 93313
rect 52472 93316 52745 93344
rect 32125 93279 32183 93285
rect 32125 93276 32137 93279
rect 31726 93248 32137 93276
rect 5534 93168 5540 93220
rect 5592 93208 5598 93220
rect 5592 93180 16574 93208
rect 5592 93168 5598 93180
rect 8938 93100 8944 93152
rect 8996 93100 9002 93152
rect 10042 93100 10048 93152
rect 10100 93100 10106 93152
rect 11146 93100 11152 93152
rect 11204 93100 11210 93152
rect 12250 93100 12256 93152
rect 12308 93100 12314 93152
rect 13262 93100 13268 93152
rect 13320 93100 13326 93152
rect 16546 93140 16574 93180
rect 30377 93143 30435 93149
rect 30377 93140 30389 93143
rect 16546 93112 30389 93140
rect 30377 93109 30389 93112
rect 30423 93140 30435 93143
rect 31726 93140 31754 93248
rect 32125 93245 32137 93248
rect 32171 93276 32183 93279
rect 40313 93279 40371 93285
rect 40313 93276 40325 93279
rect 32171 93248 40325 93276
rect 32171 93245 32183 93248
rect 32125 93239 32183 93245
rect 40313 93245 40325 93248
rect 40359 93245 40371 93279
rect 40313 93239 40371 93245
rect 42245 93279 42303 93285
rect 42245 93245 42257 93279
rect 42291 93276 42303 93279
rect 42429 93279 42487 93285
rect 42429 93276 42441 93279
rect 42291 93248 42441 93276
rect 42291 93245 42303 93248
rect 42245 93239 42303 93245
rect 42429 93245 42441 93248
rect 42475 93276 42487 93279
rect 50706 93276 50712 93288
rect 42475 93248 50712 93276
rect 42475 93245 42487 93248
rect 42429 93239 42487 93245
rect 50706 93236 50712 93248
rect 50764 93276 50770 93288
rect 50893 93279 50951 93285
rect 50893 93276 50905 93279
rect 50764 93248 50905 93276
rect 50764 93236 50770 93248
rect 50893 93245 50905 93248
rect 50939 93245 50951 93279
rect 50893 93239 50951 93245
rect 52472 93217 52500 93316
rect 52733 93313 52745 93316
rect 52779 93344 52791 93347
rect 52914 93344 52920 93356
rect 52779 93316 52920 93344
rect 52779 93313 52791 93316
rect 52733 93307 52791 93313
rect 52914 93304 52920 93316
rect 52972 93304 52978 93356
rect 54202 93304 54208 93356
rect 54260 93344 54266 93356
rect 56704 93353 56732 93452
rect 56778 93440 56784 93452
rect 56836 93440 56842 93492
rect 56689 93347 56747 93353
rect 56689 93344 56701 93347
rect 54260 93316 56701 93344
rect 54260 93304 54266 93316
rect 56689 93313 56701 93316
rect 56735 93313 56747 93347
rect 56689 93307 56747 93313
rect 53929 93279 53987 93285
rect 53929 93245 53941 93279
rect 53975 93276 53987 93279
rect 54389 93279 54447 93285
rect 54389 93276 54401 93279
rect 53975 93248 54401 93276
rect 53975 93245 53987 93248
rect 53929 93239 53987 93245
rect 54389 93245 54401 93248
rect 54435 93276 54447 93279
rect 56229 93279 56287 93285
rect 54435 93248 55214 93276
rect 54435 93245 54447 93248
rect 54389 93239 54447 93245
rect 52457 93211 52515 93217
rect 52457 93208 52469 93211
rect 52012 93180 52469 93208
rect 52012 93152 52040 93180
rect 52457 93177 52469 93180
rect 52503 93177 52515 93211
rect 55186 93208 55214 93248
rect 56229 93245 56241 93279
rect 56275 93276 56287 93279
rect 57054 93276 57060 93288
rect 56275 93248 57060 93276
rect 56275 93245 56287 93248
rect 56229 93239 56287 93245
rect 57054 93236 57060 93248
rect 57112 93236 57118 93288
rect 55186 93180 64874 93208
rect 52457 93171 52515 93177
rect 30423 93112 31754 93140
rect 30423 93109 30435 93112
rect 30377 93103 30435 93109
rect 31846 93100 31852 93152
rect 31904 93140 31910 93152
rect 49878 93140 49884 93152
rect 31904 93112 49884 93140
rect 31904 93100 31910 93112
rect 49878 93100 49884 93112
rect 49936 93100 49942 93152
rect 51074 93100 51080 93152
rect 51132 93100 51138 93152
rect 51994 93100 52000 93152
rect 52052 93100 52058 93152
rect 52365 93143 52423 93149
rect 52365 93109 52377 93143
rect 52411 93140 52423 93143
rect 52546 93140 52552 93152
rect 52411 93112 52552 93140
rect 52411 93109 52423 93112
rect 52365 93103 52423 93109
rect 52546 93100 52552 93112
rect 52604 93100 52610 93152
rect 54202 93100 54208 93152
rect 54260 93100 54266 93152
rect 55122 93100 55128 93152
rect 55180 93100 55186 93152
rect 57054 93100 57060 93152
rect 57112 93100 57118 93152
rect 64846 93140 64874 93180
rect 91738 93140 91744 93152
rect 64846 93112 91744 93140
rect 91738 93100 91744 93112
rect 91796 93100 91802 93152
rect 1104 93050 97888 93072
rect 1104 92998 4214 93050
rect 4266 92998 4278 93050
rect 4330 92998 4342 93050
rect 4394 92998 4406 93050
rect 4458 92998 4470 93050
rect 4522 92998 34934 93050
rect 34986 92998 34998 93050
rect 35050 92998 35062 93050
rect 35114 92998 35126 93050
rect 35178 92998 35190 93050
rect 35242 92998 65654 93050
rect 65706 92998 65718 93050
rect 65770 92998 65782 93050
rect 65834 92998 65846 93050
rect 65898 92998 65910 93050
rect 65962 92998 96374 93050
rect 96426 92998 96438 93050
rect 96490 92998 96502 93050
rect 96554 92998 96566 93050
rect 96618 92998 96630 93050
rect 96682 92998 97888 93050
rect 1104 92976 97888 92998
rect 57054 92896 57060 92948
rect 57112 92936 57118 92948
rect 91830 92936 91836 92948
rect 57112 92908 91836 92936
rect 57112 92896 57118 92908
rect 91830 92896 91836 92908
rect 91888 92896 91894 92948
rect 10042 92828 10048 92880
rect 10100 92868 10106 92880
rect 51994 92868 52000 92880
rect 10100 92840 52000 92868
rect 10100 92828 10106 92840
rect 51994 92828 52000 92840
rect 52052 92828 52058 92880
rect 12250 92760 12256 92812
rect 12308 92800 12314 92812
rect 54202 92800 54208 92812
rect 12308 92772 54208 92800
rect 12308 92760 12314 92772
rect 54202 92760 54208 92772
rect 54260 92760 54266 92812
rect 11146 92692 11152 92744
rect 11204 92732 11210 92744
rect 52546 92732 52552 92744
rect 11204 92704 52552 92732
rect 11204 92692 11210 92704
rect 52546 92692 52552 92704
rect 52604 92692 52610 92744
rect 1104 92506 5980 92528
rect 1104 92454 4874 92506
rect 4926 92454 4938 92506
rect 4990 92454 5002 92506
rect 5054 92454 5066 92506
rect 5118 92454 5130 92506
rect 5182 92454 5980 92506
rect 94024 92506 97888 92528
rect 1104 92432 5980 92454
rect 50522 92420 50528 92472
rect 50580 92460 50586 92472
rect 51074 92460 51080 92472
rect 50580 92432 51080 92460
rect 50580 92420 50586 92432
rect 51074 92420 51080 92432
rect 51132 92420 51138 92472
rect 94024 92454 97034 92506
rect 97086 92454 97098 92506
rect 97150 92454 97162 92506
rect 97214 92454 97226 92506
rect 97278 92454 97290 92506
rect 97342 92454 97888 92506
rect 94024 92432 97888 92454
rect 1104 91962 5980 91984
rect 1104 91910 4214 91962
rect 4266 91910 4278 91962
rect 4330 91910 4342 91962
rect 4394 91910 4406 91962
rect 4458 91910 4470 91962
rect 4522 91910 5980 91962
rect 1104 91888 5980 91910
rect 94024 91962 97888 91984
rect 94024 91910 96374 91962
rect 96426 91910 96438 91962
rect 96490 91910 96502 91962
rect 96554 91910 96566 91962
rect 96618 91910 96630 91962
rect 96682 91910 97888 91962
rect 94024 91888 97888 91910
rect 1104 91418 5980 91440
rect 1104 91366 4874 91418
rect 4926 91366 4938 91418
rect 4990 91366 5002 91418
rect 5054 91366 5066 91418
rect 5118 91366 5130 91418
rect 5182 91366 5980 91418
rect 1104 91344 5980 91366
rect 94024 91418 97888 91440
rect 94024 91366 97034 91418
rect 97086 91366 97098 91418
rect 97150 91366 97162 91418
rect 97214 91366 97226 91418
rect 97278 91366 97290 91418
rect 97342 91366 97888 91418
rect 94024 91344 97888 91366
rect 1104 90874 5980 90896
rect 1104 90822 4214 90874
rect 4266 90822 4278 90874
rect 4330 90822 4342 90874
rect 4394 90822 4406 90874
rect 4458 90822 4470 90874
rect 4522 90822 5980 90874
rect 1104 90800 5980 90822
rect 94024 90874 97888 90896
rect 94024 90822 96374 90874
rect 96426 90822 96438 90874
rect 96490 90822 96502 90874
rect 96554 90822 96566 90874
rect 96618 90822 96630 90874
rect 96682 90822 97888 90874
rect 94024 90800 97888 90822
rect 5718 90448 5724 90500
rect 5776 90488 5782 90500
rect 55122 90488 55128 90500
rect 5776 90460 55128 90488
rect 5776 90448 5782 90460
rect 55122 90448 55128 90460
rect 55180 90448 55186 90500
rect 1104 90330 5980 90352
rect 1104 90278 4874 90330
rect 4926 90278 4938 90330
rect 4990 90278 5002 90330
rect 5054 90278 5066 90330
rect 5118 90278 5130 90330
rect 5182 90278 5980 90330
rect 1104 90256 5980 90278
rect 94024 90330 97888 90352
rect 94024 90278 97034 90330
rect 97086 90278 97098 90330
rect 97150 90278 97162 90330
rect 97214 90278 97226 90330
rect 97278 90278 97290 90330
rect 97342 90278 97888 90330
rect 94024 90256 97888 90278
rect 5626 90108 5632 90160
rect 5684 90148 5690 90160
rect 8478 90148 8484 90160
rect 5684 90120 8484 90148
rect 5684 90108 5690 90120
rect 8478 90108 8484 90120
rect 8536 90108 8542 90160
rect 1104 89786 5980 89808
rect 1104 89734 4214 89786
rect 4266 89734 4278 89786
rect 4330 89734 4342 89786
rect 4394 89734 4406 89786
rect 4458 89734 4470 89786
rect 4522 89734 5980 89786
rect 1104 89712 5980 89734
rect 94024 89786 97888 89808
rect 94024 89734 96374 89786
rect 96426 89734 96438 89786
rect 96490 89734 96502 89786
rect 96554 89734 96566 89786
rect 96618 89734 96630 89786
rect 96682 89734 97888 89786
rect 94024 89712 97888 89734
rect 1104 89242 5980 89264
rect 1104 89190 4874 89242
rect 4926 89190 4938 89242
rect 4990 89190 5002 89242
rect 5054 89190 5066 89242
rect 5118 89190 5130 89242
rect 5182 89190 5980 89242
rect 1104 89168 5980 89190
rect 94024 89242 97888 89264
rect 94024 89190 97034 89242
rect 97086 89190 97098 89242
rect 97150 89190 97162 89242
rect 97214 89190 97226 89242
rect 97278 89190 97290 89242
rect 97342 89190 97888 89242
rect 94024 89168 97888 89190
rect 1104 88698 5980 88720
rect 1104 88646 4214 88698
rect 4266 88646 4278 88698
rect 4330 88646 4342 88698
rect 4394 88646 4406 88698
rect 4458 88646 4470 88698
rect 4522 88646 5980 88698
rect 1104 88624 5980 88646
rect 94024 88698 97888 88720
rect 94024 88646 96374 88698
rect 96426 88646 96438 88698
rect 96490 88646 96502 88698
rect 96554 88646 96566 88698
rect 96618 88646 96630 88698
rect 96682 88646 97888 88698
rect 94024 88624 97888 88646
rect 1104 88154 5980 88176
rect 1104 88102 4874 88154
rect 4926 88102 4938 88154
rect 4990 88102 5002 88154
rect 5054 88102 5066 88154
rect 5118 88102 5130 88154
rect 5182 88102 5980 88154
rect 1104 88080 5980 88102
rect 94024 88154 97888 88176
rect 94024 88102 97034 88154
rect 97086 88102 97098 88154
rect 97150 88102 97162 88154
rect 97214 88102 97226 88154
rect 97278 88102 97290 88154
rect 97342 88102 97888 88154
rect 94024 88080 97888 88102
rect 1104 87610 5980 87632
rect 1104 87558 4214 87610
rect 4266 87558 4278 87610
rect 4330 87558 4342 87610
rect 4394 87558 4406 87610
rect 4458 87558 4470 87610
rect 4522 87558 5980 87610
rect 1104 87536 5980 87558
rect 94024 87610 97888 87632
rect 94024 87558 96374 87610
rect 96426 87558 96438 87610
rect 96490 87558 96502 87610
rect 96554 87558 96566 87610
rect 96618 87558 96630 87610
rect 96682 87558 97888 87610
rect 94024 87536 97888 87558
rect 97350 87388 97356 87440
rect 97408 87388 97414 87440
rect 1673 87295 1731 87301
rect 1673 87261 1685 87295
rect 1719 87292 1731 87295
rect 8294 87292 8300 87304
rect 1719 87264 8300 87292
rect 1719 87261 1731 87264
rect 1673 87255 1731 87261
rect 8294 87252 8300 87264
rect 8352 87252 8358 87304
rect 97261 87295 97319 87301
rect 97261 87261 97273 87295
rect 97307 87292 97319 87295
rect 97534 87292 97540 87304
rect 97307 87264 97540 87292
rect 97307 87261 97319 87264
rect 97261 87255 97319 87261
rect 97534 87252 97540 87264
rect 97592 87252 97598 87304
rect 842 87116 848 87168
rect 900 87156 906 87168
rect 1489 87159 1547 87165
rect 1489 87156 1501 87159
rect 900 87128 1501 87156
rect 900 87116 906 87128
rect 1489 87125 1501 87128
rect 1535 87125 1547 87159
rect 1489 87119 1547 87125
rect 1104 87066 5980 87088
rect 1104 87014 4874 87066
rect 4926 87014 4938 87066
rect 4990 87014 5002 87066
rect 5054 87014 5066 87066
rect 5118 87014 5130 87066
rect 5182 87014 5980 87066
rect 1104 86992 5980 87014
rect 94024 87066 97888 87088
rect 94024 87014 97034 87066
rect 97086 87014 97098 87066
rect 97150 87014 97162 87066
rect 97214 87014 97226 87066
rect 97278 87014 97290 87066
rect 97342 87014 97888 87066
rect 94024 86992 97888 87014
rect 1673 86819 1731 86825
rect 1673 86785 1685 86819
rect 1719 86816 1731 86819
rect 8294 86816 8300 86828
rect 1719 86788 8300 86816
rect 1719 86785 1731 86788
rect 1673 86779 1731 86785
rect 8294 86776 8300 86788
rect 8352 86776 8358 86828
rect 97261 86819 97319 86825
rect 97261 86785 97273 86819
rect 97307 86816 97319 86819
rect 97534 86816 97540 86828
rect 97307 86788 97540 86816
rect 97307 86785 97319 86788
rect 97261 86779 97319 86785
rect 97534 86776 97540 86788
rect 97592 86776 97598 86828
rect 842 86572 848 86624
rect 900 86612 906 86624
rect 1489 86615 1547 86621
rect 1489 86612 1501 86615
rect 900 86584 1501 86612
rect 900 86572 906 86584
rect 1489 86581 1501 86584
rect 1535 86581 1547 86615
rect 1489 86575 1547 86581
rect 97350 86572 97356 86624
rect 97408 86572 97414 86624
rect 1104 86522 5980 86544
rect 1104 86470 4214 86522
rect 4266 86470 4278 86522
rect 4330 86470 4342 86522
rect 4394 86470 4406 86522
rect 4458 86470 4470 86522
rect 4522 86470 5980 86522
rect 1104 86448 5980 86470
rect 94024 86522 97888 86544
rect 94024 86470 96374 86522
rect 96426 86470 96438 86522
rect 96490 86470 96502 86522
rect 96554 86470 96566 86522
rect 96618 86470 96630 86522
rect 96682 86470 97888 86522
rect 94024 86448 97888 86470
rect 1104 85978 5980 86000
rect 1104 85926 4874 85978
rect 4926 85926 4938 85978
rect 4990 85926 5002 85978
rect 5054 85926 5066 85978
rect 5118 85926 5130 85978
rect 5182 85926 5980 85978
rect 1104 85904 5980 85926
rect 94024 85978 97888 86000
rect 94024 85926 97034 85978
rect 97086 85926 97098 85978
rect 97150 85926 97162 85978
rect 97214 85926 97226 85978
rect 97278 85926 97290 85978
rect 97342 85926 97888 85978
rect 94024 85904 97888 85926
rect 1104 85434 5980 85456
rect 1104 85382 4214 85434
rect 4266 85382 4278 85434
rect 4330 85382 4342 85434
rect 4394 85382 4406 85434
rect 4458 85382 4470 85434
rect 4522 85382 5980 85434
rect 1104 85360 5980 85382
rect 94024 85434 97888 85456
rect 94024 85382 96374 85434
rect 96426 85382 96438 85434
rect 96490 85382 96502 85434
rect 96554 85382 96566 85434
rect 96618 85382 96630 85434
rect 96682 85382 97888 85434
rect 94024 85360 97888 85382
rect 97350 85212 97356 85264
rect 97408 85212 97414 85264
rect 1673 85119 1731 85125
rect 1673 85085 1685 85119
rect 1719 85116 1731 85119
rect 8294 85116 8300 85128
rect 1719 85088 8300 85116
rect 1719 85085 1731 85088
rect 1673 85079 1731 85085
rect 8294 85076 8300 85088
rect 8352 85076 8358 85128
rect 97261 85119 97319 85125
rect 97261 85085 97273 85119
rect 97307 85116 97319 85119
rect 97534 85116 97540 85128
rect 97307 85088 97540 85116
rect 97307 85085 97319 85088
rect 97261 85079 97319 85085
rect 97534 85076 97540 85088
rect 97592 85076 97598 85128
rect 842 84940 848 84992
rect 900 84980 906 84992
rect 1489 84983 1547 84989
rect 1489 84980 1501 84983
rect 900 84952 1501 84980
rect 900 84940 906 84952
rect 1489 84949 1501 84952
rect 1535 84949 1547 84983
rect 1489 84943 1547 84949
rect 1104 84890 5980 84912
rect 1104 84838 4874 84890
rect 4926 84838 4938 84890
rect 4990 84838 5002 84890
rect 5054 84838 5066 84890
rect 5118 84838 5130 84890
rect 5182 84838 5980 84890
rect 1104 84816 5980 84838
rect 94024 84890 97888 84912
rect 94024 84838 97034 84890
rect 97086 84838 97098 84890
rect 97150 84838 97162 84890
rect 97214 84838 97226 84890
rect 97278 84838 97290 84890
rect 97342 84838 97888 84890
rect 94024 84816 97888 84838
rect 1670 84600 1676 84652
rect 1728 84600 1734 84652
rect 97261 84643 97319 84649
rect 97261 84609 97273 84643
rect 97307 84640 97319 84643
rect 97534 84640 97540 84652
rect 97307 84612 97540 84640
rect 97307 84609 97319 84612
rect 97261 84603 97319 84609
rect 97534 84600 97540 84612
rect 97592 84600 97598 84652
rect 842 84464 848 84516
rect 900 84504 906 84516
rect 1489 84507 1547 84513
rect 1489 84504 1501 84507
rect 900 84476 1501 84504
rect 900 84464 906 84476
rect 1489 84473 1501 84476
rect 1535 84473 1547 84507
rect 1489 84467 1547 84473
rect 97350 84396 97356 84448
rect 97408 84396 97414 84448
rect 1104 84346 5980 84368
rect 1104 84294 4214 84346
rect 4266 84294 4278 84346
rect 4330 84294 4342 84346
rect 4394 84294 4406 84346
rect 4458 84294 4470 84346
rect 4522 84294 5980 84346
rect 1104 84272 5980 84294
rect 94024 84346 97888 84368
rect 94024 84294 96374 84346
rect 96426 84294 96438 84346
rect 96490 84294 96502 84346
rect 96554 84294 96566 84346
rect 96618 84294 96630 84346
rect 96682 84294 97888 84346
rect 94024 84272 97888 84294
rect 1104 83802 5980 83824
rect 1104 83750 4874 83802
rect 4926 83750 4938 83802
rect 4990 83750 5002 83802
rect 5054 83750 5066 83802
rect 5118 83750 5130 83802
rect 5182 83750 5980 83802
rect 1104 83728 5980 83750
rect 94024 83802 97888 83824
rect 94024 83750 97034 83802
rect 97086 83750 97098 83802
rect 97150 83750 97162 83802
rect 97214 83750 97226 83802
rect 97278 83750 97290 83802
rect 97342 83750 97888 83802
rect 94024 83728 97888 83750
rect 1673 83555 1731 83561
rect 1673 83521 1685 83555
rect 1719 83552 1731 83555
rect 8294 83552 8300 83564
rect 1719 83524 8300 83552
rect 1719 83521 1731 83524
rect 1673 83515 1731 83521
rect 8294 83512 8300 83524
rect 8352 83512 8358 83564
rect 97261 83555 97319 83561
rect 97261 83521 97273 83555
rect 97307 83552 97319 83555
rect 97534 83552 97540 83564
rect 97307 83524 97540 83552
rect 97307 83521 97319 83524
rect 97261 83515 97319 83521
rect 97534 83512 97540 83524
rect 97592 83512 97598 83564
rect 842 83308 848 83360
rect 900 83348 906 83360
rect 1489 83351 1547 83357
rect 1489 83348 1501 83351
rect 900 83320 1501 83348
rect 900 83308 906 83320
rect 1489 83317 1501 83320
rect 1535 83317 1547 83351
rect 1489 83311 1547 83317
rect 97350 83308 97356 83360
rect 97408 83308 97414 83360
rect 1104 83258 5980 83280
rect 1104 83206 4214 83258
rect 4266 83206 4278 83258
rect 4330 83206 4342 83258
rect 4394 83206 4406 83258
rect 4458 83206 4470 83258
rect 4522 83206 5980 83258
rect 1104 83184 5980 83206
rect 94024 83258 97888 83280
rect 94024 83206 96374 83258
rect 96426 83206 96438 83258
rect 96490 83206 96502 83258
rect 96554 83206 96566 83258
rect 96618 83206 96630 83258
rect 96682 83206 97888 83258
rect 94024 83184 97888 83206
rect 1104 82714 5980 82736
rect 1104 82662 4874 82714
rect 4926 82662 4938 82714
rect 4990 82662 5002 82714
rect 5054 82662 5066 82714
rect 5118 82662 5130 82714
rect 5182 82662 5980 82714
rect 1104 82640 5980 82662
rect 94024 82714 97888 82736
rect 94024 82662 97034 82714
rect 97086 82662 97098 82714
rect 97150 82662 97162 82714
rect 97214 82662 97226 82714
rect 97278 82662 97290 82714
rect 97342 82662 97888 82714
rect 94024 82640 97888 82662
rect 1104 82170 5980 82192
rect 1104 82118 4214 82170
rect 4266 82118 4278 82170
rect 4330 82118 4342 82170
rect 4394 82118 4406 82170
rect 4458 82118 4470 82170
rect 4522 82118 5980 82170
rect 1104 82096 5980 82118
rect 94024 82170 97888 82192
rect 94024 82118 96374 82170
rect 96426 82118 96438 82170
rect 96490 82118 96502 82170
rect 96554 82118 96566 82170
rect 96618 82118 96630 82170
rect 96682 82118 97888 82170
rect 94024 82096 97888 82118
rect 97350 81948 97356 82000
rect 97408 81948 97414 82000
rect 1673 81855 1731 81861
rect 1673 81821 1685 81855
rect 1719 81852 1731 81855
rect 8294 81852 8300 81864
rect 1719 81824 8300 81852
rect 1719 81821 1731 81824
rect 1673 81815 1731 81821
rect 8294 81812 8300 81824
rect 8352 81812 8358 81864
rect 97261 81855 97319 81861
rect 97261 81821 97273 81855
rect 97307 81852 97319 81855
rect 97534 81852 97540 81864
rect 97307 81824 97540 81852
rect 97307 81821 97319 81824
rect 97261 81815 97319 81821
rect 97534 81812 97540 81824
rect 97592 81812 97598 81864
rect 842 81676 848 81728
rect 900 81716 906 81728
rect 1489 81719 1547 81725
rect 1489 81716 1501 81719
rect 900 81688 1501 81716
rect 900 81676 906 81688
rect 1489 81685 1501 81688
rect 1535 81685 1547 81719
rect 1489 81679 1547 81685
rect 1104 81626 5980 81648
rect 1104 81574 4874 81626
rect 4926 81574 4938 81626
rect 4990 81574 5002 81626
rect 5054 81574 5066 81626
rect 5118 81574 5130 81626
rect 5182 81574 5980 81626
rect 1104 81552 5980 81574
rect 94024 81626 97888 81648
rect 94024 81574 97034 81626
rect 97086 81574 97098 81626
rect 97150 81574 97162 81626
rect 97214 81574 97226 81626
rect 97278 81574 97290 81626
rect 97342 81574 97888 81626
rect 94024 81552 97888 81574
rect 1673 81379 1731 81385
rect 1673 81345 1685 81379
rect 1719 81376 1731 81379
rect 8294 81376 8300 81388
rect 1719 81348 8300 81376
rect 1719 81345 1731 81348
rect 1673 81339 1731 81345
rect 8294 81336 8300 81348
rect 8352 81336 8358 81388
rect 97261 81379 97319 81385
rect 97261 81345 97273 81379
rect 97307 81376 97319 81379
rect 97534 81376 97540 81388
rect 97307 81348 97540 81376
rect 97307 81345 97319 81348
rect 97261 81339 97319 81345
rect 97534 81336 97540 81348
rect 97592 81336 97598 81388
rect 842 81132 848 81184
rect 900 81172 906 81184
rect 1489 81175 1547 81181
rect 1489 81172 1501 81175
rect 900 81144 1501 81172
rect 900 81132 906 81144
rect 1489 81141 1501 81144
rect 1535 81141 1547 81175
rect 1489 81135 1547 81141
rect 97350 81132 97356 81184
rect 97408 81132 97414 81184
rect 1104 81082 5980 81104
rect 1104 81030 4214 81082
rect 4266 81030 4278 81082
rect 4330 81030 4342 81082
rect 4394 81030 4406 81082
rect 4458 81030 4470 81082
rect 4522 81030 5980 81082
rect 1104 81008 5980 81030
rect 94024 81082 97888 81104
rect 94024 81030 96374 81082
rect 96426 81030 96438 81082
rect 96490 81030 96502 81082
rect 96554 81030 96566 81082
rect 96618 81030 96630 81082
rect 96682 81030 97888 81082
rect 94024 81008 97888 81030
rect 1104 80538 5980 80560
rect 1104 80486 4874 80538
rect 4926 80486 4938 80538
rect 4990 80486 5002 80538
rect 5054 80486 5066 80538
rect 5118 80486 5130 80538
rect 5182 80486 5980 80538
rect 1104 80464 5980 80486
rect 94024 80538 97888 80560
rect 94024 80486 97034 80538
rect 97086 80486 97098 80538
rect 97150 80486 97162 80538
rect 97214 80486 97226 80538
rect 97278 80486 97290 80538
rect 97342 80486 97888 80538
rect 94024 80464 97888 80486
rect 1104 79994 5980 80016
rect 1104 79942 4214 79994
rect 4266 79942 4278 79994
rect 4330 79942 4342 79994
rect 4394 79942 4406 79994
rect 4458 79942 4470 79994
rect 4522 79942 5980 79994
rect 1104 79920 5980 79942
rect 94024 79994 97888 80016
rect 94024 79942 96374 79994
rect 96426 79942 96438 79994
rect 96490 79942 96502 79994
rect 96554 79942 96566 79994
rect 96618 79942 96630 79994
rect 96682 79942 97888 79994
rect 94024 79920 97888 79942
rect 97350 79772 97356 79824
rect 97408 79772 97414 79824
rect 1673 79679 1731 79685
rect 1673 79645 1685 79679
rect 1719 79676 1731 79679
rect 8294 79676 8300 79688
rect 1719 79648 8300 79676
rect 1719 79645 1731 79648
rect 1673 79639 1731 79645
rect 8294 79636 8300 79648
rect 8352 79636 8358 79688
rect 97261 79679 97319 79685
rect 97261 79645 97273 79679
rect 97307 79676 97319 79679
rect 97534 79676 97540 79688
rect 97307 79648 97540 79676
rect 97307 79645 97319 79648
rect 97261 79639 97319 79645
rect 97534 79636 97540 79648
rect 97592 79636 97598 79688
rect 842 79500 848 79552
rect 900 79540 906 79552
rect 1489 79543 1547 79549
rect 1489 79540 1501 79543
rect 900 79512 1501 79540
rect 900 79500 906 79512
rect 1489 79509 1501 79512
rect 1535 79509 1547 79543
rect 1489 79503 1547 79509
rect 1104 79450 5980 79472
rect 1104 79398 4874 79450
rect 4926 79398 4938 79450
rect 4990 79398 5002 79450
rect 5054 79398 5066 79450
rect 5118 79398 5130 79450
rect 5182 79398 5980 79450
rect 1104 79376 5980 79398
rect 94024 79450 97888 79472
rect 94024 79398 97034 79450
rect 97086 79398 97098 79450
rect 97150 79398 97162 79450
rect 97214 79398 97226 79450
rect 97278 79398 97290 79450
rect 97342 79398 97888 79450
rect 94024 79376 97888 79398
rect 1673 79203 1731 79209
rect 1673 79169 1685 79203
rect 1719 79200 1731 79203
rect 8294 79200 8300 79212
rect 1719 79172 8300 79200
rect 1719 79169 1731 79172
rect 1673 79163 1731 79169
rect 8294 79160 8300 79172
rect 8352 79160 8358 79212
rect 97169 79203 97227 79209
rect 97169 79169 97181 79203
rect 97215 79200 97227 79203
rect 97442 79200 97448 79212
rect 97215 79172 97448 79200
rect 97215 79169 97227 79172
rect 97169 79163 97227 79169
rect 97442 79160 97448 79172
rect 97500 79160 97506 79212
rect 842 79024 848 79076
rect 900 79064 906 79076
rect 1489 79067 1547 79073
rect 1489 79064 1501 79067
rect 900 79036 1501 79064
rect 900 79024 906 79036
rect 1489 79033 1501 79036
rect 1535 79033 1547 79067
rect 1489 79027 1547 79033
rect 97258 79024 97264 79076
rect 97316 79024 97322 79076
rect 1104 78906 5980 78928
rect 1104 78854 4214 78906
rect 4266 78854 4278 78906
rect 4330 78854 4342 78906
rect 4394 78854 4406 78906
rect 4458 78854 4470 78906
rect 4522 78854 5980 78906
rect 1104 78832 5980 78854
rect 94024 78906 97888 78928
rect 94024 78854 96374 78906
rect 96426 78854 96438 78906
rect 96490 78854 96502 78906
rect 96554 78854 96566 78906
rect 96618 78854 96630 78906
rect 96682 78854 97888 78906
rect 94024 78832 97888 78854
rect 1104 78362 5980 78384
rect 1104 78310 4874 78362
rect 4926 78310 4938 78362
rect 4990 78310 5002 78362
rect 5054 78310 5066 78362
rect 5118 78310 5130 78362
rect 5182 78310 5980 78362
rect 1104 78288 5980 78310
rect 94024 78362 97888 78384
rect 94024 78310 97034 78362
rect 97086 78310 97098 78362
rect 97150 78310 97162 78362
rect 97214 78310 97226 78362
rect 97278 78310 97290 78362
rect 97342 78310 97888 78362
rect 94024 78288 97888 78310
rect 1673 78115 1731 78121
rect 1673 78081 1685 78115
rect 1719 78112 1731 78115
rect 8294 78112 8300 78124
rect 1719 78084 8300 78112
rect 1719 78081 1731 78084
rect 1673 78075 1731 78081
rect 8294 78072 8300 78084
rect 8352 78072 8358 78124
rect 97261 78115 97319 78121
rect 97261 78081 97273 78115
rect 97307 78112 97319 78115
rect 97534 78112 97540 78124
rect 97307 78084 97540 78112
rect 97307 78081 97319 78084
rect 97261 78075 97319 78081
rect 97534 78072 97540 78084
rect 97592 78072 97598 78124
rect 842 77868 848 77920
rect 900 77908 906 77920
rect 1489 77911 1547 77917
rect 1489 77908 1501 77911
rect 900 77880 1501 77908
rect 900 77868 906 77880
rect 1489 77877 1501 77880
rect 1535 77877 1547 77911
rect 1489 77871 1547 77877
rect 97350 77868 97356 77920
rect 97408 77868 97414 77920
rect 1104 77818 5980 77840
rect 1104 77766 4214 77818
rect 4266 77766 4278 77818
rect 4330 77766 4342 77818
rect 4394 77766 4406 77818
rect 4458 77766 4470 77818
rect 4522 77766 5980 77818
rect 1104 77744 5980 77766
rect 94024 77818 97888 77840
rect 94024 77766 96374 77818
rect 96426 77766 96438 77818
rect 96490 77766 96502 77818
rect 96554 77766 96566 77818
rect 96618 77766 96630 77818
rect 96682 77766 97888 77818
rect 94024 77744 97888 77766
rect 1104 77274 5980 77296
rect 1104 77222 4874 77274
rect 4926 77222 4938 77274
rect 4990 77222 5002 77274
rect 5054 77222 5066 77274
rect 5118 77222 5130 77274
rect 5182 77222 5980 77274
rect 1104 77200 5980 77222
rect 94024 77274 97888 77296
rect 94024 77222 97034 77274
rect 97086 77222 97098 77274
rect 97150 77222 97162 77274
rect 97214 77222 97226 77274
rect 97278 77222 97290 77274
rect 97342 77222 97888 77274
rect 94024 77200 97888 77222
rect 1104 76730 5980 76752
rect 1104 76678 4214 76730
rect 4266 76678 4278 76730
rect 4330 76678 4342 76730
rect 4394 76678 4406 76730
rect 4458 76678 4470 76730
rect 4522 76678 5980 76730
rect 1104 76656 5980 76678
rect 94024 76730 97888 76752
rect 94024 76678 96374 76730
rect 96426 76678 96438 76730
rect 96490 76678 96502 76730
rect 96554 76678 96566 76730
rect 96618 76678 96630 76730
rect 96682 76678 97888 76730
rect 94024 76656 97888 76678
rect 97350 76508 97356 76560
rect 97408 76508 97414 76560
rect 1673 76415 1731 76421
rect 1673 76381 1685 76415
rect 1719 76412 1731 76415
rect 8294 76412 8300 76424
rect 1719 76384 8300 76412
rect 1719 76381 1731 76384
rect 1673 76375 1731 76381
rect 8294 76372 8300 76384
rect 8352 76372 8358 76424
rect 97261 76415 97319 76421
rect 97261 76381 97273 76415
rect 97307 76412 97319 76415
rect 97534 76412 97540 76424
rect 97307 76384 97540 76412
rect 97307 76381 97319 76384
rect 97261 76375 97319 76381
rect 97534 76372 97540 76384
rect 97592 76372 97598 76424
rect 842 76236 848 76288
rect 900 76276 906 76288
rect 1489 76279 1547 76285
rect 1489 76276 1501 76279
rect 900 76248 1501 76276
rect 900 76236 906 76248
rect 1489 76245 1501 76248
rect 1535 76245 1547 76279
rect 1489 76239 1547 76245
rect 1104 76186 5980 76208
rect 1104 76134 4874 76186
rect 4926 76134 4938 76186
rect 4990 76134 5002 76186
rect 5054 76134 5066 76186
rect 5118 76134 5130 76186
rect 5182 76134 5980 76186
rect 1104 76112 5980 76134
rect 94024 76186 97888 76208
rect 94024 76134 97034 76186
rect 97086 76134 97098 76186
rect 97150 76134 97162 76186
rect 97214 76134 97226 76186
rect 97278 76134 97290 76186
rect 97342 76134 97888 76186
rect 94024 76112 97888 76134
rect 842 76032 848 76084
rect 900 76072 906 76084
rect 1489 76075 1547 76081
rect 1489 76072 1501 76075
rect 900 76044 1501 76072
rect 900 76032 906 76044
rect 1489 76041 1501 76044
rect 1535 76041 1547 76075
rect 1489 76035 1547 76041
rect 1670 75896 1676 75948
rect 1728 75896 1734 75948
rect 97261 75939 97319 75945
rect 97261 75905 97273 75939
rect 97307 75936 97319 75939
rect 97534 75936 97540 75948
rect 97307 75908 97540 75936
rect 97307 75905 97319 75908
rect 97261 75899 97319 75905
rect 97534 75896 97540 75908
rect 97592 75896 97598 75948
rect 97350 75692 97356 75744
rect 97408 75692 97414 75744
rect 1104 75642 5980 75664
rect 1104 75590 4214 75642
rect 4266 75590 4278 75642
rect 4330 75590 4342 75642
rect 4394 75590 4406 75642
rect 4458 75590 4470 75642
rect 4522 75590 5980 75642
rect 1104 75568 5980 75590
rect 94024 75642 97888 75664
rect 94024 75590 96374 75642
rect 96426 75590 96438 75642
rect 96490 75590 96502 75642
rect 96554 75590 96566 75642
rect 96618 75590 96630 75642
rect 96682 75590 97888 75642
rect 94024 75568 97888 75590
rect 1104 75098 5980 75120
rect 1104 75046 4874 75098
rect 4926 75046 4938 75098
rect 4990 75046 5002 75098
rect 5054 75046 5066 75098
rect 5118 75046 5130 75098
rect 5182 75046 5980 75098
rect 1104 75024 5980 75046
rect 94024 75098 97888 75120
rect 94024 75046 97034 75098
rect 97086 75046 97098 75098
rect 97150 75046 97162 75098
rect 97214 75046 97226 75098
rect 97278 75046 97290 75098
rect 97342 75046 97888 75098
rect 94024 75024 97888 75046
rect 1104 74554 5980 74576
rect 1104 74502 4214 74554
rect 4266 74502 4278 74554
rect 4330 74502 4342 74554
rect 4394 74502 4406 74554
rect 4458 74502 4470 74554
rect 4522 74502 5980 74554
rect 1104 74480 5980 74502
rect 94024 74554 97888 74576
rect 94024 74502 96374 74554
rect 96426 74502 96438 74554
rect 96490 74502 96502 74554
rect 96554 74502 96566 74554
rect 96618 74502 96630 74554
rect 96682 74502 97888 74554
rect 94024 74480 97888 74502
rect 97258 74332 97264 74384
rect 97316 74332 97322 74384
rect 1673 74239 1731 74245
rect 1673 74205 1685 74239
rect 1719 74236 1731 74239
rect 8294 74236 8300 74248
rect 1719 74208 8300 74236
rect 1719 74205 1731 74208
rect 1673 74199 1731 74205
rect 8294 74196 8300 74208
rect 8352 74196 8358 74248
rect 97169 74171 97227 74177
rect 97169 74137 97181 74171
rect 97215 74168 97227 74171
rect 97442 74168 97448 74180
rect 97215 74140 97448 74168
rect 97215 74137 97227 74140
rect 97169 74131 97227 74137
rect 97442 74128 97448 74140
rect 97500 74128 97506 74180
rect 842 74060 848 74112
rect 900 74100 906 74112
rect 1489 74103 1547 74109
rect 1489 74100 1501 74103
rect 900 74072 1501 74100
rect 900 74060 906 74072
rect 1489 74069 1501 74072
rect 1535 74069 1547 74103
rect 1489 74063 1547 74069
rect 1104 74010 5980 74032
rect 1104 73958 4874 74010
rect 4926 73958 4938 74010
rect 4990 73958 5002 74010
rect 5054 73958 5066 74010
rect 5118 73958 5130 74010
rect 5182 73958 5980 74010
rect 1104 73936 5980 73958
rect 94024 74010 97888 74032
rect 94024 73958 97034 74010
rect 97086 73958 97098 74010
rect 97150 73958 97162 74010
rect 97214 73958 97226 74010
rect 97278 73958 97290 74010
rect 97342 73958 97888 74010
rect 94024 73936 97888 73958
rect 1673 73763 1731 73769
rect 1673 73729 1685 73763
rect 1719 73760 1731 73763
rect 8294 73760 8300 73772
rect 1719 73732 8300 73760
rect 1719 73729 1731 73732
rect 1673 73723 1731 73729
rect 8294 73720 8300 73732
rect 8352 73720 8358 73772
rect 97261 73763 97319 73769
rect 97261 73729 97273 73763
rect 97307 73760 97319 73763
rect 97534 73760 97540 73772
rect 97307 73732 97540 73760
rect 97307 73729 97319 73732
rect 97261 73723 97319 73729
rect 97534 73720 97540 73732
rect 97592 73720 97598 73772
rect 842 73584 848 73636
rect 900 73624 906 73636
rect 1489 73627 1547 73633
rect 1489 73624 1501 73627
rect 900 73596 1501 73624
rect 900 73584 906 73596
rect 1489 73593 1501 73596
rect 1535 73593 1547 73627
rect 1489 73587 1547 73593
rect 97350 73516 97356 73568
rect 97408 73516 97414 73568
rect 1104 73466 5980 73488
rect 1104 73414 4214 73466
rect 4266 73414 4278 73466
rect 4330 73414 4342 73466
rect 4394 73414 4406 73466
rect 4458 73414 4470 73466
rect 4522 73414 5980 73466
rect 1104 73392 5980 73414
rect 94024 73466 97888 73488
rect 94024 73414 96374 73466
rect 96426 73414 96438 73466
rect 96490 73414 96502 73466
rect 96554 73414 96566 73466
rect 96618 73414 96630 73466
rect 96682 73414 97888 73466
rect 94024 73392 97888 73414
rect 1104 72922 5980 72944
rect 1104 72870 4874 72922
rect 4926 72870 4938 72922
rect 4990 72870 5002 72922
rect 5054 72870 5066 72922
rect 5118 72870 5130 72922
rect 5182 72870 5980 72922
rect 1104 72848 5980 72870
rect 94024 72922 97888 72944
rect 94024 72870 97034 72922
rect 97086 72870 97098 72922
rect 97150 72870 97162 72922
rect 97214 72870 97226 72922
rect 97278 72870 97290 72922
rect 97342 72870 97888 72922
rect 94024 72848 97888 72870
rect 1673 72675 1731 72681
rect 1673 72641 1685 72675
rect 1719 72672 1731 72675
rect 8294 72672 8300 72684
rect 1719 72644 8300 72672
rect 1719 72641 1731 72644
rect 1673 72635 1731 72641
rect 8294 72632 8300 72644
rect 8352 72632 8358 72684
rect 97258 72564 97264 72616
rect 97316 72564 97322 72616
rect 97534 72564 97540 72616
rect 97592 72564 97598 72616
rect 842 72428 848 72480
rect 900 72468 906 72480
rect 1489 72471 1547 72477
rect 1489 72468 1501 72471
rect 900 72440 1501 72468
rect 900 72428 906 72440
rect 1489 72437 1501 72440
rect 1535 72437 1547 72471
rect 1489 72431 1547 72437
rect 1104 72378 5980 72400
rect 1104 72326 4214 72378
rect 4266 72326 4278 72378
rect 4330 72326 4342 72378
rect 4394 72326 4406 72378
rect 4458 72326 4470 72378
rect 4522 72326 5980 72378
rect 1104 72304 5980 72326
rect 94024 72378 97888 72400
rect 94024 72326 96374 72378
rect 96426 72326 96438 72378
rect 96490 72326 96502 72378
rect 96554 72326 96566 72378
rect 96618 72326 96630 72378
rect 96682 72326 97888 72378
rect 94024 72304 97888 72326
rect 97534 72156 97540 72208
rect 97592 72156 97598 72208
rect 1104 71834 5980 71856
rect 1104 71782 4874 71834
rect 4926 71782 4938 71834
rect 4990 71782 5002 71834
rect 5054 71782 5066 71834
rect 5118 71782 5130 71834
rect 5182 71782 5980 71834
rect 1104 71760 5980 71782
rect 94024 71834 97888 71856
rect 94024 71782 97034 71834
rect 97086 71782 97098 71834
rect 97150 71782 97162 71834
rect 97214 71782 97226 71834
rect 97278 71782 97290 71834
rect 97342 71782 97888 71834
rect 94024 71760 97888 71782
rect 1104 71290 5980 71312
rect 1104 71238 4214 71290
rect 4266 71238 4278 71290
rect 4330 71238 4342 71290
rect 4394 71238 4406 71290
rect 4458 71238 4470 71290
rect 4522 71238 5980 71290
rect 1104 71216 5980 71238
rect 94024 71290 97888 71312
rect 94024 71238 96374 71290
rect 96426 71238 96438 71290
rect 96490 71238 96502 71290
rect 96554 71238 96566 71290
rect 96618 71238 96630 71290
rect 96682 71238 97888 71290
rect 94024 71216 97888 71238
rect 97350 71068 97356 71120
rect 97408 71068 97414 71120
rect 1673 70975 1731 70981
rect 1673 70941 1685 70975
rect 1719 70972 1731 70975
rect 8294 70972 8300 70984
rect 1719 70944 8300 70972
rect 1719 70941 1731 70944
rect 1673 70935 1731 70941
rect 8294 70932 8300 70944
rect 8352 70932 8358 70984
rect 97261 70975 97319 70981
rect 97261 70941 97273 70975
rect 97307 70972 97319 70975
rect 97534 70972 97540 70984
rect 97307 70944 97540 70972
rect 97307 70941 97319 70944
rect 97261 70935 97319 70941
rect 97534 70932 97540 70944
rect 97592 70932 97598 70984
rect 842 70796 848 70848
rect 900 70836 906 70848
rect 1489 70839 1547 70845
rect 1489 70836 1501 70839
rect 900 70808 1501 70836
rect 900 70796 906 70808
rect 1489 70805 1501 70808
rect 1535 70805 1547 70839
rect 1489 70799 1547 70805
rect 1104 70746 5980 70768
rect 1104 70694 4874 70746
rect 4926 70694 4938 70746
rect 4990 70694 5002 70746
rect 5054 70694 5066 70746
rect 5118 70694 5130 70746
rect 5182 70694 5980 70746
rect 1104 70672 5980 70694
rect 94024 70746 97888 70768
rect 94024 70694 97034 70746
rect 97086 70694 97098 70746
rect 97150 70694 97162 70746
rect 97214 70694 97226 70746
rect 97278 70694 97290 70746
rect 97342 70694 97888 70746
rect 94024 70672 97888 70694
rect 5534 70592 5540 70644
rect 5592 70592 5598 70644
rect 97442 70592 97448 70644
rect 97500 70592 97506 70644
rect 1302 70456 1308 70508
rect 1360 70496 1366 70508
rect 1397 70499 1455 70505
rect 1397 70496 1409 70499
rect 1360 70468 1409 70496
rect 1360 70456 1366 70468
rect 1397 70465 1409 70468
rect 1443 70496 1455 70499
rect 1673 70499 1731 70505
rect 1673 70496 1685 70499
rect 1443 70468 1685 70496
rect 1443 70465 1455 70468
rect 1397 70459 1455 70465
rect 1673 70465 1685 70468
rect 1719 70465 1731 70499
rect 1673 70459 1731 70465
rect 97258 70456 97264 70508
rect 97316 70456 97322 70508
rect 1578 70252 1584 70304
rect 1636 70252 1642 70304
rect 1104 70202 5980 70224
rect 1104 70150 4214 70202
rect 4266 70150 4278 70202
rect 4330 70150 4342 70202
rect 4394 70150 4406 70202
rect 4458 70150 4470 70202
rect 4522 70150 5980 70202
rect 1104 70128 5980 70150
rect 94024 70202 97888 70224
rect 94024 70150 96374 70202
rect 96426 70150 96438 70202
rect 96490 70150 96502 70202
rect 96554 70150 96566 70202
rect 96618 70150 96630 70202
rect 96682 70150 97888 70202
rect 94024 70128 97888 70150
rect 5534 69844 5540 69896
rect 5592 69884 5598 69896
rect 5629 69887 5687 69893
rect 5629 69884 5641 69887
rect 5592 69856 5641 69884
rect 5592 69844 5598 69856
rect 5629 69853 5641 69856
rect 5675 69853 5687 69887
rect 5629 69847 5687 69853
rect 4341 69751 4399 69757
rect 4341 69717 4353 69751
rect 4387 69748 4399 69751
rect 5626 69748 5632 69760
rect 4387 69720 5632 69748
rect 4387 69717 4399 69720
rect 4341 69711 4399 69717
rect 5626 69708 5632 69720
rect 5684 69708 5690 69760
rect 1104 69658 5980 69680
rect 1104 69606 4874 69658
rect 4926 69606 4938 69658
rect 4990 69606 5002 69658
rect 5054 69606 5066 69658
rect 5118 69606 5130 69658
rect 5182 69606 5980 69658
rect 1104 69584 5980 69606
rect 94024 69658 97888 69680
rect 94024 69606 97034 69658
rect 97086 69606 97098 69658
rect 97150 69606 97162 69658
rect 97214 69606 97226 69658
rect 97278 69606 97290 69658
rect 97342 69606 97888 69658
rect 94024 69584 97888 69606
rect 5626 69504 5632 69556
rect 5684 69504 5690 69556
rect 1104 69114 5980 69136
rect 1104 69062 4214 69114
rect 4266 69062 4278 69114
rect 4330 69062 4342 69114
rect 4394 69062 4406 69114
rect 4458 69062 4470 69114
rect 4522 69062 5980 69114
rect 1104 69040 5980 69062
rect 94024 69114 97888 69136
rect 94024 69062 96374 69114
rect 96426 69062 96438 69114
rect 96490 69062 96502 69114
rect 96554 69062 96566 69114
rect 96618 69062 96630 69114
rect 96682 69062 97888 69114
rect 94024 69040 97888 69062
rect 97258 68756 97264 68808
rect 97316 68756 97322 68808
rect 1118 68688 1124 68740
rect 1176 68728 1182 68740
rect 1489 68731 1547 68737
rect 1489 68728 1501 68731
rect 1176 68700 1501 68728
rect 1176 68688 1182 68700
rect 1489 68697 1501 68700
rect 1535 68697 1547 68731
rect 1489 68691 1547 68697
rect 1673 68731 1731 68737
rect 1673 68697 1685 68731
rect 1719 68728 1731 68731
rect 8294 68728 8300 68740
rect 1719 68700 8300 68728
rect 1719 68697 1731 68700
rect 1673 68691 1731 68697
rect 1504 68660 1532 68691
rect 8294 68688 8300 68700
rect 8352 68688 8358 68740
rect 1765 68663 1823 68669
rect 1765 68660 1777 68663
rect 1504 68632 1777 68660
rect 1765 68629 1777 68632
rect 1811 68629 1823 68663
rect 1765 68623 1823 68629
rect 97442 68620 97448 68672
rect 97500 68620 97506 68672
rect 1104 68570 5980 68592
rect 1104 68518 4874 68570
rect 4926 68518 4938 68570
rect 4990 68518 5002 68570
rect 5054 68518 5066 68570
rect 5118 68518 5130 68570
rect 5182 68518 5980 68570
rect 1104 68496 5980 68518
rect 94024 68570 97888 68592
rect 94024 68518 97034 68570
rect 97086 68518 97098 68570
rect 97150 68518 97162 68570
rect 97214 68518 97226 68570
rect 97278 68518 97290 68570
rect 97342 68518 97888 68570
rect 94024 68496 97888 68518
rect 1302 68280 1308 68332
rect 1360 68320 1366 68332
rect 1489 68323 1547 68329
rect 1489 68320 1501 68323
rect 1360 68292 1501 68320
rect 1360 68280 1366 68292
rect 1489 68289 1501 68292
rect 1535 68320 1547 68323
rect 1765 68323 1823 68329
rect 1765 68320 1777 68323
rect 1535 68292 1777 68320
rect 1535 68289 1547 68292
rect 1489 68283 1547 68289
rect 1765 68289 1777 68292
rect 1811 68289 1823 68323
rect 1765 68283 1823 68289
rect 97258 68280 97264 68332
rect 97316 68280 97322 68332
rect 1673 68187 1731 68193
rect 1673 68153 1685 68187
rect 1719 68184 1731 68187
rect 8294 68184 8300 68196
rect 1719 68156 8300 68184
rect 1719 68153 1731 68156
rect 1673 68147 1731 68153
rect 8294 68144 8300 68156
rect 8352 68144 8358 68196
rect 97442 68076 97448 68128
rect 97500 68076 97506 68128
rect 1104 68026 5980 68048
rect 1104 67974 4214 68026
rect 4266 67974 4278 68026
rect 4330 67974 4342 68026
rect 4394 67974 4406 68026
rect 4458 67974 4470 68026
rect 4522 67974 5980 68026
rect 1104 67952 5980 67974
rect 94024 68026 97888 68048
rect 94024 67974 96374 68026
rect 96426 67974 96438 68026
rect 96490 67974 96502 68026
rect 96554 67974 96566 68026
rect 96618 67974 96630 68026
rect 96682 67974 97888 68026
rect 94024 67952 97888 67974
rect 1104 67482 5980 67504
rect 1104 67430 4874 67482
rect 4926 67430 4938 67482
rect 4990 67430 5002 67482
rect 5054 67430 5066 67482
rect 5118 67430 5130 67482
rect 5182 67430 5980 67482
rect 1104 67408 5980 67430
rect 94024 67482 97888 67504
rect 94024 67430 97034 67482
rect 97086 67430 97098 67482
rect 97150 67430 97162 67482
rect 97214 67430 97226 67482
rect 97278 67430 97290 67482
rect 97342 67430 97888 67482
rect 94024 67408 97888 67430
rect 1302 67192 1308 67244
rect 1360 67232 1366 67244
rect 1489 67235 1547 67241
rect 1489 67232 1501 67235
rect 1360 67204 1501 67232
rect 1360 67192 1366 67204
rect 1489 67201 1501 67204
rect 1535 67232 1547 67235
rect 1765 67235 1823 67241
rect 1765 67232 1777 67235
rect 1535 67204 1777 67232
rect 1535 67201 1547 67204
rect 1489 67195 1547 67201
rect 1765 67201 1777 67204
rect 1811 67201 1823 67235
rect 1765 67195 1823 67201
rect 97258 67192 97264 67244
rect 97316 67192 97322 67244
rect 1673 67099 1731 67105
rect 1673 67065 1685 67099
rect 1719 67096 1731 67099
rect 8294 67096 8300 67108
rect 1719 67068 8300 67096
rect 1719 67065 1731 67068
rect 1673 67059 1731 67065
rect 8294 67056 8300 67068
rect 8352 67056 8358 67108
rect 97442 66988 97448 67040
rect 97500 66988 97506 67040
rect 1104 66938 5980 66960
rect 1104 66886 4214 66938
rect 4266 66886 4278 66938
rect 4330 66886 4342 66938
rect 4394 66886 4406 66938
rect 4458 66886 4470 66938
rect 4522 66886 5980 66938
rect 1104 66864 5980 66886
rect 94024 66938 97888 66960
rect 94024 66886 96374 66938
rect 96426 66886 96438 66938
rect 96490 66886 96502 66938
rect 96554 66886 96566 66938
rect 96618 66886 96630 66938
rect 96682 66886 97888 66938
rect 94024 66864 97888 66886
rect 1104 66394 5980 66416
rect 1104 66342 4874 66394
rect 4926 66342 4938 66394
rect 4990 66342 5002 66394
rect 5054 66342 5066 66394
rect 5118 66342 5130 66394
rect 5182 66342 5980 66394
rect 1104 66320 5980 66342
rect 94024 66394 97888 66416
rect 94024 66342 97034 66394
rect 97086 66342 97098 66394
rect 97150 66342 97162 66394
rect 97214 66342 97226 66394
rect 97278 66342 97290 66394
rect 97342 66342 97888 66394
rect 94024 66320 97888 66342
rect 1104 65850 5980 65872
rect 1104 65798 4214 65850
rect 4266 65798 4278 65850
rect 4330 65798 4342 65850
rect 4394 65798 4406 65850
rect 4458 65798 4470 65850
rect 4522 65798 5980 65850
rect 1104 65776 5980 65798
rect 94024 65850 97888 65872
rect 94024 65798 96374 65850
rect 96426 65798 96438 65850
rect 96490 65798 96502 65850
rect 96554 65798 96566 65850
rect 96618 65798 96630 65850
rect 96682 65798 97888 65850
rect 94024 65776 97888 65798
rect 1673 65671 1731 65677
rect 1673 65637 1685 65671
rect 1719 65668 1731 65671
rect 8294 65668 8300 65680
rect 1719 65640 8300 65668
rect 1719 65637 1731 65640
rect 1673 65631 1731 65637
rect 8294 65628 8300 65640
rect 8352 65628 8358 65680
rect 97258 65492 97264 65544
rect 97316 65492 97322 65544
rect 1118 65424 1124 65476
rect 1176 65464 1182 65476
rect 1489 65467 1547 65473
rect 1489 65464 1501 65467
rect 1176 65436 1501 65464
rect 1176 65424 1182 65436
rect 1489 65433 1501 65436
rect 1535 65464 1547 65467
rect 1765 65467 1823 65473
rect 1765 65464 1777 65467
rect 1535 65436 1777 65464
rect 1535 65433 1547 65436
rect 1489 65427 1547 65433
rect 1765 65433 1777 65436
rect 1811 65433 1823 65467
rect 1765 65427 1823 65433
rect 97442 65356 97448 65408
rect 97500 65356 97506 65408
rect 1104 65306 5980 65328
rect 1104 65254 4874 65306
rect 4926 65254 4938 65306
rect 4990 65254 5002 65306
rect 5054 65254 5066 65306
rect 5118 65254 5130 65306
rect 5182 65254 5980 65306
rect 1104 65232 5980 65254
rect 94024 65306 97888 65328
rect 94024 65254 97034 65306
rect 97086 65254 97098 65306
rect 97150 65254 97162 65306
rect 97214 65254 97226 65306
rect 97278 65254 97290 65306
rect 97342 65254 97888 65306
rect 94024 65232 97888 65254
rect 1302 65016 1308 65068
rect 1360 65056 1366 65068
rect 1489 65059 1547 65065
rect 1489 65056 1501 65059
rect 1360 65028 1501 65056
rect 1360 65016 1366 65028
rect 1489 65025 1501 65028
rect 1535 65056 1547 65059
rect 1765 65059 1823 65065
rect 1765 65056 1777 65059
rect 1535 65028 1777 65056
rect 1535 65025 1547 65028
rect 1489 65019 1547 65025
rect 1765 65025 1777 65028
rect 1811 65025 1823 65059
rect 1765 65019 1823 65025
rect 97258 65016 97264 65068
rect 97316 65016 97322 65068
rect 1670 64880 1676 64932
rect 1728 64880 1734 64932
rect 97442 64880 97448 64932
rect 97500 64880 97506 64932
rect 1104 64762 5980 64784
rect 1104 64710 4214 64762
rect 4266 64710 4278 64762
rect 4330 64710 4342 64762
rect 4394 64710 4406 64762
rect 4458 64710 4470 64762
rect 4522 64710 5980 64762
rect 1104 64688 5980 64710
rect 94024 64762 97888 64784
rect 94024 64710 96374 64762
rect 96426 64710 96438 64762
rect 96490 64710 96502 64762
rect 96554 64710 96566 64762
rect 96618 64710 96630 64762
rect 96682 64710 97888 64762
rect 94024 64688 97888 64710
rect 1104 64218 5980 64240
rect 1104 64166 4874 64218
rect 4926 64166 4938 64218
rect 4990 64166 5002 64218
rect 5054 64166 5066 64218
rect 5118 64166 5130 64218
rect 5182 64166 5980 64218
rect 1104 64144 5980 64166
rect 94024 64218 97888 64240
rect 94024 64166 97034 64218
rect 97086 64166 97098 64218
rect 97150 64166 97162 64218
rect 97214 64166 97226 64218
rect 97278 64166 97290 64218
rect 97342 64166 97888 64218
rect 94024 64144 97888 64166
rect 1104 63674 5980 63696
rect 1104 63622 4214 63674
rect 4266 63622 4278 63674
rect 4330 63622 4342 63674
rect 4394 63622 4406 63674
rect 4458 63622 4470 63674
rect 4522 63622 5980 63674
rect 1104 63600 5980 63622
rect 94024 63674 97888 63696
rect 94024 63622 96374 63674
rect 96426 63622 96438 63674
rect 96490 63622 96502 63674
rect 96554 63622 96566 63674
rect 96618 63622 96630 63674
rect 96682 63622 97888 63674
rect 94024 63600 97888 63622
rect 97258 63316 97264 63368
rect 97316 63316 97322 63368
rect 1118 63248 1124 63300
rect 1176 63288 1182 63300
rect 1489 63291 1547 63297
rect 1489 63288 1501 63291
rect 1176 63260 1501 63288
rect 1176 63248 1182 63260
rect 1489 63257 1501 63260
rect 1535 63257 1547 63291
rect 1489 63251 1547 63257
rect 1673 63291 1731 63297
rect 1673 63257 1685 63291
rect 1719 63288 1731 63291
rect 8294 63288 8300 63300
rect 1719 63260 8300 63288
rect 1719 63257 1731 63260
rect 1673 63251 1731 63257
rect 1504 63220 1532 63251
rect 8294 63248 8300 63260
rect 8352 63248 8358 63300
rect 1765 63223 1823 63229
rect 1765 63220 1777 63223
rect 1504 63192 1777 63220
rect 1765 63189 1777 63192
rect 1811 63189 1823 63223
rect 1765 63183 1823 63189
rect 97442 63180 97448 63232
rect 97500 63180 97506 63232
rect 1104 63130 5980 63152
rect 1104 63078 4874 63130
rect 4926 63078 4938 63130
rect 4990 63078 5002 63130
rect 5054 63078 5066 63130
rect 5118 63078 5130 63130
rect 5182 63078 5980 63130
rect 1104 63056 5980 63078
rect 94024 63130 97888 63152
rect 94024 63078 97034 63130
rect 97086 63078 97098 63130
rect 97150 63078 97162 63130
rect 97214 63078 97226 63130
rect 97278 63078 97290 63130
rect 97342 63078 97888 63130
rect 94024 63056 97888 63078
rect 1302 62840 1308 62892
rect 1360 62880 1366 62892
rect 1489 62883 1547 62889
rect 1489 62880 1501 62883
rect 1360 62852 1501 62880
rect 1360 62840 1366 62852
rect 1489 62849 1501 62852
rect 1535 62880 1547 62883
rect 1949 62883 2007 62889
rect 1949 62880 1961 62883
rect 1535 62852 1961 62880
rect 1535 62849 1547 62852
rect 1489 62843 1547 62849
rect 1949 62849 1961 62852
rect 1995 62849 2007 62883
rect 1949 62843 2007 62849
rect 97258 62840 97264 62892
rect 97316 62840 97322 62892
rect 1765 62747 1823 62753
rect 1765 62713 1777 62747
rect 1811 62744 1823 62747
rect 8294 62744 8300 62756
rect 1811 62716 8300 62744
rect 1811 62713 1823 62716
rect 1765 62707 1823 62713
rect 8294 62704 8300 62716
rect 8352 62704 8358 62756
rect 97442 62636 97448 62688
rect 97500 62636 97506 62688
rect 1104 62586 5980 62608
rect 1104 62534 4214 62586
rect 4266 62534 4278 62586
rect 4330 62534 4342 62586
rect 4394 62534 4406 62586
rect 4458 62534 4470 62586
rect 4522 62534 5980 62586
rect 1104 62512 5980 62534
rect 94024 62586 97888 62608
rect 94024 62534 96374 62586
rect 96426 62534 96438 62586
rect 96490 62534 96502 62586
rect 96554 62534 96566 62586
rect 96618 62534 96630 62586
rect 96682 62534 97888 62586
rect 94024 62512 97888 62534
rect 1104 62042 5980 62064
rect 1104 61990 4874 62042
rect 4926 61990 4938 62042
rect 4990 61990 5002 62042
rect 5054 61990 5066 62042
rect 5118 61990 5130 62042
rect 5182 61990 5980 62042
rect 1104 61968 5980 61990
rect 94024 62042 97888 62064
rect 94024 61990 97034 62042
rect 97086 61990 97098 62042
rect 97150 61990 97162 62042
rect 97214 61990 97226 62042
rect 97278 61990 97290 62042
rect 97342 61990 97888 62042
rect 94024 61968 97888 61990
rect 1302 61752 1308 61804
rect 1360 61792 1366 61804
rect 1489 61795 1547 61801
rect 1489 61792 1501 61795
rect 1360 61764 1501 61792
rect 1360 61752 1366 61764
rect 1489 61761 1501 61764
rect 1535 61792 1547 61795
rect 1765 61795 1823 61801
rect 1765 61792 1777 61795
rect 1535 61764 1777 61792
rect 1535 61761 1547 61764
rect 1489 61755 1547 61761
rect 1765 61761 1777 61764
rect 1811 61761 1823 61795
rect 1765 61755 1823 61761
rect 97258 61752 97264 61804
rect 97316 61752 97322 61804
rect 1673 61659 1731 61665
rect 1673 61625 1685 61659
rect 1719 61656 1731 61659
rect 8294 61656 8300 61668
rect 1719 61628 8300 61656
rect 1719 61625 1731 61628
rect 1673 61619 1731 61625
rect 8294 61616 8300 61628
rect 8352 61616 8358 61668
rect 97442 61548 97448 61600
rect 97500 61548 97506 61600
rect 1104 61498 5980 61520
rect 1104 61446 4214 61498
rect 4266 61446 4278 61498
rect 4330 61446 4342 61498
rect 4394 61446 4406 61498
rect 4458 61446 4470 61498
rect 4522 61446 5980 61498
rect 1104 61424 5980 61446
rect 94024 61498 97888 61520
rect 94024 61446 96374 61498
rect 96426 61446 96438 61498
rect 96490 61446 96502 61498
rect 96554 61446 96566 61498
rect 96618 61446 96630 61498
rect 96682 61446 97888 61498
rect 94024 61424 97888 61446
rect 1104 60954 5980 60976
rect 1104 60902 4874 60954
rect 4926 60902 4938 60954
rect 4990 60902 5002 60954
rect 5054 60902 5066 60954
rect 5118 60902 5130 60954
rect 5182 60902 5980 60954
rect 1104 60880 5980 60902
rect 94024 60954 97888 60976
rect 94024 60902 97034 60954
rect 97086 60902 97098 60954
rect 97150 60902 97162 60954
rect 97214 60902 97226 60954
rect 97278 60902 97290 60954
rect 97342 60902 97888 60954
rect 94024 60880 97888 60902
rect 1104 60410 5980 60432
rect 1104 60358 4214 60410
rect 4266 60358 4278 60410
rect 4330 60358 4342 60410
rect 4394 60358 4406 60410
rect 4458 60358 4470 60410
rect 4522 60358 5980 60410
rect 1104 60336 5980 60358
rect 94024 60410 97888 60432
rect 94024 60358 96374 60410
rect 96426 60358 96438 60410
rect 96490 60358 96502 60410
rect 96554 60358 96566 60410
rect 96618 60358 96630 60410
rect 96682 60358 97888 60410
rect 94024 60336 97888 60358
rect 1765 60299 1823 60305
rect 1765 60265 1777 60299
rect 1811 60296 1823 60299
rect 8294 60296 8300 60308
rect 1811 60268 8300 60296
rect 1811 60265 1823 60268
rect 1765 60259 1823 60265
rect 8294 60256 8300 60268
rect 8352 60256 8358 60308
rect 97258 60052 97264 60104
rect 97316 60052 97322 60104
rect 1210 59984 1216 60036
rect 1268 60024 1274 60036
rect 1489 60027 1547 60033
rect 1489 60024 1501 60027
rect 1268 59996 1501 60024
rect 1268 59984 1274 59996
rect 1489 59993 1501 59996
rect 1535 60024 1547 60027
rect 1949 60027 2007 60033
rect 1949 60024 1961 60027
rect 1535 59996 1961 60024
rect 1535 59993 1547 59996
rect 1489 59987 1547 59993
rect 1949 59993 1961 59996
rect 1995 59993 2007 60027
rect 1949 59987 2007 59993
rect 50430 59984 50436 60036
rect 50488 60024 50494 60036
rect 50614 60024 50620 60036
rect 50488 59996 50620 60024
rect 50488 59984 50494 59996
rect 50614 59984 50620 59996
rect 50672 59984 50678 60036
rect 97442 59916 97448 59968
rect 97500 59916 97506 59968
rect 1104 59866 5980 59888
rect 1104 59814 4874 59866
rect 4926 59814 4938 59866
rect 4990 59814 5002 59866
rect 5054 59814 5066 59866
rect 5118 59814 5130 59866
rect 5182 59814 5980 59866
rect 1104 59792 5980 59814
rect 94024 59866 97888 59888
rect 94024 59814 97034 59866
rect 97086 59814 97098 59866
rect 97150 59814 97162 59866
rect 97214 59814 97226 59866
rect 97278 59814 97290 59866
rect 97342 59814 97888 59866
rect 94024 59792 97888 59814
rect 1210 59576 1216 59628
rect 1268 59616 1274 59628
rect 1397 59619 1455 59625
rect 1397 59616 1409 59619
rect 1268 59588 1409 59616
rect 1268 59576 1274 59588
rect 1397 59585 1409 59588
rect 1443 59616 1455 59619
rect 1765 59619 1823 59625
rect 1765 59616 1777 59619
rect 1443 59588 1777 59616
rect 1443 59585 1455 59588
rect 1397 59579 1455 59585
rect 1765 59585 1777 59588
rect 1811 59585 1823 59619
rect 1765 59579 1823 59585
rect 97258 59576 97264 59628
rect 97316 59576 97322 59628
rect 1578 59372 1584 59424
rect 1636 59372 1642 59424
rect 97442 59372 97448 59424
rect 97500 59372 97506 59424
rect 1104 59322 5980 59344
rect 1104 59270 4214 59322
rect 4266 59270 4278 59322
rect 4330 59270 4342 59322
rect 4394 59270 4406 59322
rect 4458 59270 4470 59322
rect 4522 59270 5980 59322
rect 1104 59248 5980 59270
rect 94024 59322 97888 59344
rect 94024 59270 96374 59322
rect 96426 59270 96438 59322
rect 96490 59270 96502 59322
rect 96554 59270 96566 59322
rect 96618 59270 96630 59322
rect 96682 59270 97888 59322
rect 94024 59248 97888 59270
rect 1104 58778 5980 58800
rect 1104 58726 4874 58778
rect 4926 58726 4938 58778
rect 4990 58726 5002 58778
rect 5054 58726 5066 58778
rect 5118 58726 5130 58778
rect 5182 58726 5980 58778
rect 1104 58704 5980 58726
rect 94024 58778 97888 58800
rect 94024 58726 97034 58778
rect 97086 58726 97098 58778
rect 97150 58726 97162 58778
rect 97214 58726 97226 58778
rect 97278 58726 97290 58778
rect 97342 58726 97888 58778
rect 94024 58704 97888 58726
rect 1104 58234 5980 58256
rect 1104 58182 4214 58234
rect 4266 58182 4278 58234
rect 4330 58182 4342 58234
rect 4394 58182 4406 58234
rect 4458 58182 4470 58234
rect 4522 58182 5980 58234
rect 1104 58160 5980 58182
rect 94024 58234 97888 58256
rect 94024 58182 96374 58234
rect 96426 58182 96438 58234
rect 96490 58182 96502 58234
rect 96554 58182 96566 58234
rect 96618 58182 96630 58234
rect 96682 58182 97888 58234
rect 94024 58160 97888 58182
rect 1302 57876 1308 57928
rect 1360 57916 1366 57928
rect 1397 57919 1455 57925
rect 1397 57916 1409 57919
rect 1360 57888 1409 57916
rect 1360 57876 1366 57888
rect 1397 57885 1409 57888
rect 1443 57916 1455 57919
rect 1765 57919 1823 57925
rect 1765 57916 1777 57919
rect 1443 57888 1777 57916
rect 1443 57885 1455 57888
rect 1397 57879 1455 57885
rect 1765 57885 1777 57888
rect 1811 57885 1823 57919
rect 1765 57879 1823 57885
rect 97258 57876 97264 57928
rect 97316 57876 97322 57928
rect 1578 57740 1584 57792
rect 1636 57740 1642 57792
rect 97442 57740 97448 57792
rect 97500 57740 97506 57792
rect 1104 57690 5980 57712
rect 1104 57638 4874 57690
rect 4926 57638 4938 57690
rect 4990 57638 5002 57690
rect 5054 57638 5066 57690
rect 5118 57638 5130 57690
rect 5182 57638 5980 57690
rect 1104 57616 5980 57638
rect 94024 57690 97888 57712
rect 94024 57638 97034 57690
rect 97086 57638 97098 57690
rect 97150 57638 97162 57690
rect 97214 57638 97226 57690
rect 97278 57638 97290 57690
rect 97342 57638 97888 57690
rect 94024 57616 97888 57638
rect 1302 57400 1308 57452
rect 1360 57440 1366 57452
rect 1489 57443 1547 57449
rect 1489 57440 1501 57443
rect 1360 57412 1501 57440
rect 1360 57400 1366 57412
rect 1489 57409 1501 57412
rect 1535 57440 1547 57443
rect 1949 57443 2007 57449
rect 1949 57440 1961 57443
rect 1535 57412 1961 57440
rect 1535 57409 1547 57412
rect 1489 57403 1547 57409
rect 1949 57409 1961 57412
rect 1995 57409 2007 57443
rect 1949 57403 2007 57409
rect 97258 57400 97264 57452
rect 97316 57400 97322 57452
rect 1765 57307 1823 57313
rect 1765 57273 1777 57307
rect 1811 57304 1823 57307
rect 8294 57304 8300 57316
rect 1811 57276 8300 57304
rect 1811 57273 1823 57276
rect 1765 57267 1823 57273
rect 8294 57264 8300 57276
rect 8352 57264 8358 57316
rect 97442 57196 97448 57248
rect 97500 57196 97506 57248
rect 1104 57146 5980 57168
rect 1104 57094 4214 57146
rect 4266 57094 4278 57146
rect 4330 57094 4342 57146
rect 4394 57094 4406 57146
rect 4458 57094 4470 57146
rect 4522 57094 5980 57146
rect 1104 57072 5980 57094
rect 94024 57146 97888 57168
rect 94024 57094 96374 57146
rect 96426 57094 96438 57146
rect 96490 57094 96502 57146
rect 96554 57094 96566 57146
rect 96618 57094 96630 57146
rect 96682 57094 97888 57146
rect 94024 57072 97888 57094
rect 1104 56602 5980 56624
rect 1104 56550 4874 56602
rect 4926 56550 4938 56602
rect 4990 56550 5002 56602
rect 5054 56550 5066 56602
rect 5118 56550 5130 56602
rect 5182 56550 5980 56602
rect 1104 56528 5980 56550
rect 94024 56602 97888 56624
rect 94024 56550 97034 56602
rect 97086 56550 97098 56602
rect 97150 56550 97162 56602
rect 97214 56550 97226 56602
rect 97278 56550 97290 56602
rect 97342 56550 97888 56602
rect 94024 56528 97888 56550
rect 1302 56312 1308 56364
rect 1360 56352 1366 56364
rect 1489 56355 1547 56361
rect 1489 56352 1501 56355
rect 1360 56324 1501 56352
rect 1360 56312 1366 56324
rect 1489 56321 1501 56324
rect 1535 56352 1547 56355
rect 1949 56355 2007 56361
rect 1949 56352 1961 56355
rect 1535 56324 1961 56352
rect 1535 56321 1547 56324
rect 1489 56315 1547 56321
rect 1949 56321 1961 56324
rect 1995 56321 2007 56355
rect 1949 56315 2007 56321
rect 97258 56312 97264 56364
rect 97316 56312 97322 56364
rect 1765 56219 1823 56225
rect 1765 56185 1777 56219
rect 1811 56216 1823 56219
rect 8294 56216 8300 56228
rect 1811 56188 8300 56216
rect 1811 56185 1823 56188
rect 1765 56179 1823 56185
rect 8294 56176 8300 56188
rect 8352 56176 8358 56228
rect 97442 56108 97448 56160
rect 97500 56108 97506 56160
rect 1104 56058 5980 56080
rect 1104 56006 4214 56058
rect 4266 56006 4278 56058
rect 4330 56006 4342 56058
rect 4394 56006 4406 56058
rect 4458 56006 4470 56058
rect 4522 56006 5980 56058
rect 1104 55984 5980 56006
rect 94024 56058 97888 56080
rect 94024 56006 96374 56058
rect 96426 56006 96438 56058
rect 96490 56006 96502 56058
rect 96554 56006 96566 56058
rect 96618 56006 96630 56058
rect 96682 56006 97888 56058
rect 94024 55984 97888 56006
rect 1104 55514 5980 55536
rect 1104 55462 4874 55514
rect 4926 55462 4938 55514
rect 4990 55462 5002 55514
rect 5054 55462 5066 55514
rect 5118 55462 5130 55514
rect 5182 55462 5980 55514
rect 1104 55440 5980 55462
rect 94024 55514 97888 55536
rect 94024 55462 97034 55514
rect 97086 55462 97098 55514
rect 97150 55462 97162 55514
rect 97214 55462 97226 55514
rect 97278 55462 97290 55514
rect 97342 55462 97888 55514
rect 94024 55440 97888 55462
rect 1104 54970 5980 54992
rect 1104 54918 4214 54970
rect 4266 54918 4278 54970
rect 4330 54918 4342 54970
rect 4394 54918 4406 54970
rect 4458 54918 4470 54970
rect 4522 54918 5980 54970
rect 1104 54896 5980 54918
rect 94024 54970 97888 54992
rect 94024 54918 96374 54970
rect 96426 54918 96438 54970
rect 96490 54918 96502 54970
rect 96554 54918 96566 54970
rect 96618 54918 96630 54970
rect 96682 54918 97888 54970
rect 94024 54896 97888 54918
rect 1581 54859 1639 54865
rect 1581 54825 1593 54859
rect 1627 54856 1639 54859
rect 8294 54856 8300 54868
rect 1627 54828 8300 54856
rect 1627 54825 1639 54828
rect 1581 54819 1639 54825
rect 8294 54816 8300 54828
rect 8352 54816 8358 54868
rect 1302 54612 1308 54664
rect 1360 54652 1366 54664
rect 1397 54655 1455 54661
rect 1397 54652 1409 54655
rect 1360 54624 1409 54652
rect 1360 54612 1366 54624
rect 1397 54621 1409 54624
rect 1443 54652 1455 54655
rect 1765 54655 1823 54661
rect 1765 54652 1777 54655
rect 1443 54624 1777 54652
rect 1443 54621 1455 54624
rect 1397 54615 1455 54621
rect 1765 54621 1777 54624
rect 1811 54621 1823 54655
rect 1765 54615 1823 54621
rect 97258 54612 97264 54664
rect 97316 54612 97322 54664
rect 97442 54476 97448 54528
rect 97500 54476 97506 54528
rect 1104 54426 5980 54448
rect 1104 54374 4874 54426
rect 4926 54374 4938 54426
rect 4990 54374 5002 54426
rect 5054 54374 5066 54426
rect 5118 54374 5130 54426
rect 5182 54374 5980 54426
rect 1104 54352 5980 54374
rect 94024 54426 97888 54448
rect 94024 54374 97034 54426
rect 97086 54374 97098 54426
rect 97150 54374 97162 54426
rect 97214 54374 97226 54426
rect 97278 54374 97290 54426
rect 97342 54374 97888 54426
rect 94024 54352 97888 54374
rect 1210 54136 1216 54188
rect 1268 54176 1274 54188
rect 1397 54179 1455 54185
rect 1397 54176 1409 54179
rect 1268 54148 1409 54176
rect 1268 54136 1274 54148
rect 1397 54145 1409 54148
rect 1443 54176 1455 54179
rect 1765 54179 1823 54185
rect 1765 54176 1777 54179
rect 1443 54148 1777 54176
rect 1443 54145 1455 54148
rect 1397 54139 1455 54145
rect 1765 54145 1777 54148
rect 1811 54145 1823 54179
rect 1765 54139 1823 54145
rect 97258 54136 97264 54188
rect 97316 54136 97322 54188
rect 1578 53932 1584 53984
rect 1636 53932 1642 53984
rect 97442 53932 97448 53984
rect 97500 53932 97506 53984
rect 1104 53882 5980 53904
rect 1104 53830 4214 53882
rect 4266 53830 4278 53882
rect 4330 53830 4342 53882
rect 4394 53830 4406 53882
rect 4458 53830 4470 53882
rect 4522 53830 5980 53882
rect 1104 53808 5980 53830
rect 94024 53882 97888 53904
rect 94024 53830 96374 53882
rect 96426 53830 96438 53882
rect 96490 53830 96502 53882
rect 96554 53830 96566 53882
rect 96618 53830 96630 53882
rect 96682 53830 97888 53882
rect 94024 53808 97888 53830
rect 1104 53338 5980 53360
rect 1104 53286 4874 53338
rect 4926 53286 4938 53338
rect 4990 53286 5002 53338
rect 5054 53286 5066 53338
rect 5118 53286 5130 53338
rect 5182 53286 5980 53338
rect 1104 53264 5980 53286
rect 94024 53338 97888 53360
rect 94024 53286 97034 53338
rect 97086 53286 97098 53338
rect 97150 53286 97162 53338
rect 97214 53286 97226 53338
rect 97278 53286 97290 53338
rect 97342 53286 97888 53338
rect 94024 53264 97888 53286
rect 1104 52794 5980 52816
rect 1104 52742 4214 52794
rect 4266 52742 4278 52794
rect 4330 52742 4342 52794
rect 4394 52742 4406 52794
rect 4458 52742 4470 52794
rect 4522 52742 5980 52794
rect 1104 52720 5980 52742
rect 94024 52794 97888 52816
rect 94024 52742 96374 52794
rect 96426 52742 96438 52794
rect 96490 52742 96502 52794
rect 96554 52742 96566 52794
rect 96618 52742 96630 52794
rect 96682 52742 97888 52794
rect 94024 52720 97888 52742
rect 1104 52250 5980 52272
rect 1104 52198 4874 52250
rect 4926 52198 4938 52250
rect 4990 52198 5002 52250
rect 5054 52198 5066 52250
rect 5118 52198 5130 52250
rect 5182 52198 5980 52250
rect 1104 52176 5980 52198
rect 94024 52250 97888 52272
rect 94024 52198 97034 52250
rect 97086 52198 97098 52250
rect 97150 52198 97162 52250
rect 97214 52198 97226 52250
rect 97278 52198 97290 52250
rect 97342 52198 97888 52250
rect 94024 52176 97888 52198
rect 1104 51706 5980 51728
rect 1104 51654 4214 51706
rect 4266 51654 4278 51706
rect 4330 51654 4342 51706
rect 4394 51654 4406 51706
rect 4458 51654 4470 51706
rect 4522 51654 5980 51706
rect 1104 51632 5980 51654
rect 94024 51706 97888 51728
rect 94024 51654 96374 51706
rect 96426 51654 96438 51706
rect 96490 51654 96502 51706
rect 96554 51654 96566 51706
rect 96618 51654 96630 51706
rect 96682 51654 97888 51706
rect 94024 51632 97888 51654
rect 1104 51162 5980 51184
rect 1104 51110 4874 51162
rect 4926 51110 4938 51162
rect 4990 51110 5002 51162
rect 5054 51110 5066 51162
rect 5118 51110 5130 51162
rect 5182 51110 5980 51162
rect 1104 51088 5980 51110
rect 94024 51162 97888 51184
rect 94024 51110 97034 51162
rect 97086 51110 97098 51162
rect 97150 51110 97162 51162
rect 97214 51110 97226 51162
rect 97278 51110 97290 51162
rect 97342 51110 97888 51162
rect 94024 51088 97888 51110
rect 5629 51051 5687 51057
rect 5629 51017 5641 51051
rect 5675 51048 5687 51051
rect 5718 51048 5724 51060
rect 5675 51020 5724 51048
rect 5675 51017 5687 51020
rect 5629 51011 5687 51017
rect 5718 51008 5724 51020
rect 5776 51048 5782 51060
rect 8478 51048 8484 51060
rect 5776 51020 8484 51048
rect 5776 51008 5782 51020
rect 8478 51008 8484 51020
rect 8536 51008 8542 51060
rect 5261 50847 5319 50853
rect 5261 50813 5273 50847
rect 5307 50844 5319 50847
rect 7466 50844 7472 50856
rect 5307 50816 7472 50844
rect 5307 50813 5319 50816
rect 5261 50807 5319 50813
rect 7466 50804 7472 50816
rect 7524 50804 7530 50856
rect 92106 50804 92112 50856
rect 92164 50844 92170 50856
rect 94685 50847 94743 50853
rect 94685 50844 94697 50847
rect 92164 50816 94697 50844
rect 92164 50804 92170 50816
rect 94685 50813 94697 50816
rect 94731 50813 94743 50847
rect 94685 50807 94743 50813
rect 5445 50779 5503 50785
rect 5445 50745 5457 50779
rect 5491 50776 5503 50779
rect 94501 50779 94559 50785
rect 94501 50776 94513 50779
rect 5491 50748 6500 50776
rect 5491 50745 5503 50748
rect 5445 50739 5503 50745
rect 6472 50708 6500 50748
rect 80026 50748 94513 50776
rect 6472 50680 6914 50708
rect 6886 50640 6914 50680
rect 8202 50640 8208 50652
rect 1104 50618 5980 50640
rect 1104 50566 4214 50618
rect 4266 50566 4278 50618
rect 4330 50566 4342 50618
rect 4394 50566 4406 50618
rect 4458 50566 4470 50618
rect 4522 50566 5980 50618
rect 6886 50612 8208 50640
rect 8202 50600 8208 50612
rect 8260 50640 8266 50652
rect 9858 50640 9864 50652
rect 8260 50612 9864 50640
rect 8260 50600 8266 50612
rect 9858 50600 9864 50612
rect 9916 50600 9922 50652
rect 1104 50544 5980 50566
rect 10226 50192 10232 50244
rect 10284 50232 10290 50244
rect 10284 50204 16574 50232
rect 10284 50192 10290 50204
rect 5629 50167 5687 50173
rect 5629 50133 5641 50167
rect 5675 50164 5687 50167
rect 8018 50164 8024 50176
rect 5675 50136 8024 50164
rect 5675 50133 5687 50136
rect 5629 50127 5687 50133
rect 8018 50124 8024 50136
rect 8076 50164 8082 50176
rect 11790 50164 11796 50176
rect 8076 50136 11796 50164
rect 8076 50124 8082 50136
rect 11790 50124 11796 50136
rect 11848 50124 11854 50176
rect 16546 50164 16574 50204
rect 53374 50192 53380 50244
rect 53432 50232 53438 50244
rect 80026 50232 80054 50748
rect 94501 50745 94513 50748
rect 94547 50745 94559 50779
rect 94501 50739 94559 50745
rect 94317 50711 94375 50717
rect 94317 50708 94329 50711
rect 53432 50204 80054 50232
rect 89686 50680 94329 50708
rect 53432 50192 53438 50204
rect 52270 50164 52276 50176
rect 16546 50136 52276 50164
rect 52270 50124 52276 50136
rect 52328 50164 52334 50176
rect 89686 50164 89714 50680
rect 94317 50677 94329 50680
rect 94363 50677 94375 50711
rect 94317 50671 94375 50677
rect 94024 50618 97888 50640
rect 94024 50566 96374 50618
rect 96426 50566 96438 50618
rect 96490 50566 96502 50618
rect 96554 50566 96566 50618
rect 96618 50566 96630 50618
rect 96682 50566 97888 50618
rect 94024 50544 97888 50566
rect 52328 50136 89714 50164
rect 52328 50124 52334 50136
rect 1104 50074 5980 50096
rect 1104 50022 4874 50074
rect 4926 50022 4938 50074
rect 4990 50022 5002 50074
rect 5054 50022 5066 50074
rect 5118 50022 5130 50074
rect 5182 50022 5980 50074
rect 7466 50056 7472 50108
rect 7524 50096 7530 50108
rect 8110 50096 8116 50108
rect 7524 50068 8116 50096
rect 7524 50056 7530 50068
rect 8110 50056 8116 50068
rect 8168 50096 8174 50108
rect 11146 50096 11152 50108
rect 8168 50068 11152 50096
rect 8168 50056 8174 50068
rect 11146 50056 11152 50068
rect 11204 50096 11210 50108
rect 52914 50096 52920 50108
rect 11204 50068 52920 50096
rect 11204 50056 11210 50068
rect 52914 50056 52920 50068
rect 52972 50056 52978 50108
rect 94024 50074 97888 50096
rect 1104 50000 5980 50022
rect 54478 49988 54484 50040
rect 54536 50028 54542 50040
rect 91922 50028 91928 50040
rect 54536 50000 91928 50028
rect 54536 49988 54542 50000
rect 91922 49988 91928 50000
rect 91980 50028 91986 50040
rect 92106 50028 92112 50040
rect 91980 50000 92112 50028
rect 91980 49988 91986 50000
rect 92106 49988 92112 50000
rect 92164 49988 92170 50040
rect 94024 50022 97034 50074
rect 97086 50022 97098 50074
rect 97150 50022 97162 50074
rect 97214 50022 97226 50074
rect 97278 50022 97290 50074
rect 97342 50022 97888 50074
rect 94024 50000 97888 50022
rect 1104 49530 5980 49552
rect 1104 49478 4214 49530
rect 4266 49478 4278 49530
rect 4330 49478 4342 49530
rect 4394 49478 4406 49530
rect 4458 49478 4470 49530
rect 4522 49478 5980 49530
rect 1104 49456 5980 49478
rect 94024 49530 97888 49552
rect 94024 49478 96374 49530
rect 96426 49478 96438 49530
rect 96490 49478 96502 49530
rect 96554 49478 96566 49530
rect 96618 49478 96630 49530
rect 96682 49478 97888 49530
rect 94024 49456 97888 49478
rect 1104 48986 5980 49008
rect 1104 48934 4874 48986
rect 4926 48934 4938 48986
rect 4990 48934 5002 48986
rect 5054 48934 5066 48986
rect 5118 48934 5130 48986
rect 5182 48934 5980 48986
rect 1104 48912 5980 48934
rect 94024 48986 97888 49008
rect 94024 48934 97034 48986
rect 97086 48934 97098 48986
rect 97150 48934 97162 48986
rect 97214 48934 97226 48986
rect 97278 48934 97290 48986
rect 97342 48934 97888 48986
rect 94024 48912 97888 48934
rect 1581 48875 1639 48881
rect 1581 48841 1593 48875
rect 1627 48841 1639 48875
rect 1581 48835 1639 48841
rect 1596 48804 1624 48835
rect 5534 48832 5540 48884
rect 5592 48872 5598 48884
rect 8478 48872 8484 48884
rect 5592 48844 8484 48872
rect 5592 48832 5598 48844
rect 8478 48832 8484 48844
rect 8536 48832 8542 48884
rect 12894 48804 12900 48816
rect 1596 48776 12900 48804
rect 12894 48764 12900 48776
rect 12952 48764 12958 48816
rect 52270 48764 52276 48816
rect 52328 48804 52334 48816
rect 91738 48804 91744 48816
rect 52328 48776 91744 48804
rect 52328 48764 52334 48776
rect 91738 48764 91744 48776
rect 91796 48804 91802 48816
rect 94685 48807 94743 48813
rect 94685 48804 94697 48807
rect 91796 48776 94697 48804
rect 91796 48764 91802 48776
rect 94685 48773 94697 48776
rect 94731 48773 94743 48807
rect 94685 48767 94743 48773
rect 1210 48696 1216 48748
rect 1268 48736 1274 48748
rect 1397 48739 1455 48745
rect 1397 48736 1409 48739
rect 1268 48708 1409 48736
rect 1268 48696 1274 48708
rect 1397 48705 1409 48708
rect 1443 48736 1455 48739
rect 1765 48739 1823 48745
rect 1765 48736 1777 48739
rect 1443 48708 1777 48736
rect 1443 48705 1455 48708
rect 1397 48699 1455 48705
rect 1765 48705 1777 48708
rect 1811 48705 1823 48739
rect 1765 48699 1823 48705
rect 5626 48696 5632 48748
rect 5684 48736 5690 48748
rect 11146 48736 11152 48748
rect 5684 48708 11152 48736
rect 5684 48696 5690 48708
rect 11146 48696 11152 48708
rect 11204 48696 11210 48748
rect 55582 48696 55588 48748
rect 55640 48736 55646 48748
rect 94317 48739 94375 48745
rect 94317 48736 94329 48739
rect 55640 48708 94329 48736
rect 55640 48696 55646 48708
rect 94317 48705 94329 48708
rect 94363 48705 94375 48739
rect 94317 48699 94375 48705
rect 5261 48671 5319 48677
rect 5261 48637 5273 48671
rect 5307 48668 5319 48671
rect 10226 48668 10232 48680
rect 5307 48640 10232 48668
rect 5307 48637 5319 48640
rect 5261 48631 5319 48637
rect 10226 48628 10232 48640
rect 10284 48668 10290 48680
rect 51810 48668 51816 48680
rect 10284 48640 51816 48668
rect 10284 48628 10290 48640
rect 51810 48628 51816 48640
rect 51868 48628 51874 48680
rect 54478 48628 54484 48680
rect 54536 48668 54542 48680
rect 91830 48668 91836 48680
rect 54536 48640 91836 48668
rect 54536 48628 54542 48640
rect 91830 48628 91836 48640
rect 91888 48668 91894 48680
rect 94501 48671 94559 48677
rect 94501 48668 94513 48671
rect 91888 48640 94513 48668
rect 91888 48628 91894 48640
rect 94501 48637 94513 48640
rect 94547 48637 94559 48671
rect 94501 48631 94559 48637
rect 5445 48603 5503 48609
rect 5445 48569 5457 48603
rect 5491 48600 5503 48603
rect 11882 48600 11888 48612
rect 5491 48572 11888 48600
rect 5491 48569 5503 48572
rect 5445 48563 5503 48569
rect 11882 48560 11888 48572
rect 11940 48600 11946 48612
rect 54018 48600 54024 48612
rect 11940 48572 54024 48600
rect 11940 48560 11946 48572
rect 54018 48560 54024 48572
rect 54076 48560 54082 48612
rect 50338 48492 50344 48544
rect 50396 48532 50402 48544
rect 55398 48532 55404 48544
rect 50396 48504 55404 48532
rect 50396 48492 50402 48504
rect 55398 48492 55404 48504
rect 55456 48492 55462 48544
rect 91646 48532 91652 48544
rect 80026 48504 91652 48532
rect 1104 48442 5980 48464
rect 1104 48390 4214 48442
rect 4266 48390 4278 48442
rect 4330 48390 4342 48442
rect 4394 48390 4406 48442
rect 4458 48390 4470 48442
rect 4522 48390 5980 48442
rect 11330 48424 11336 48476
rect 11388 48464 11394 48476
rect 53374 48464 53380 48476
rect 11388 48436 53380 48464
rect 11388 48424 11394 48436
rect 53374 48424 53380 48436
rect 53432 48464 53438 48476
rect 80026 48464 80054 48504
rect 91646 48492 91652 48504
rect 91704 48532 91710 48544
rect 94869 48535 94927 48541
rect 94869 48532 94881 48535
rect 91704 48504 94881 48532
rect 91704 48492 91710 48504
rect 94869 48501 94881 48504
rect 94915 48501 94927 48535
rect 94869 48495 94927 48501
rect 53432 48436 80054 48464
rect 94024 48442 97888 48464
rect 53432 48424 53438 48436
rect 1104 48368 5980 48390
rect 94024 48390 96374 48442
rect 96426 48390 96438 48442
rect 96490 48390 96502 48442
rect 96554 48390 96566 48442
rect 96618 48390 96630 48442
rect 96682 48390 97888 48442
rect 94024 48368 97888 48390
rect 5626 48220 5632 48272
rect 5684 48220 5690 48272
rect 1104 47898 5980 47920
rect 1104 47846 4874 47898
rect 4926 47846 4938 47898
rect 4990 47846 5002 47898
rect 5054 47846 5066 47898
rect 5118 47846 5130 47898
rect 5182 47846 5980 47898
rect 1104 47824 5980 47846
rect 94024 47898 97888 47920
rect 94024 47846 97034 47898
rect 97086 47846 97098 47898
rect 97150 47846 97162 47898
rect 97214 47846 97226 47898
rect 97278 47846 97290 47898
rect 97342 47846 97888 47898
rect 94024 47824 97888 47846
rect 1104 47354 5980 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 5980 47354
rect 1104 47280 5980 47302
rect 94024 47354 97888 47376
rect 94024 47302 96374 47354
rect 96426 47302 96438 47354
rect 96490 47302 96502 47354
rect 96554 47302 96566 47354
rect 96618 47302 96630 47354
rect 96682 47302 97888 47354
rect 94024 47280 97888 47302
rect 1104 46810 5980 46832
rect 1104 46758 4874 46810
rect 4926 46758 4938 46810
rect 4990 46758 5002 46810
rect 5054 46758 5066 46810
rect 5118 46758 5130 46810
rect 5182 46758 5980 46810
rect 1104 46736 5980 46758
rect 94024 46810 97888 46832
rect 94024 46758 97034 46810
rect 97086 46758 97098 46810
rect 97150 46758 97162 46810
rect 97214 46758 97226 46810
rect 97278 46758 97290 46810
rect 97342 46758 97888 46810
rect 94024 46736 97888 46758
rect 1104 46266 5980 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 5980 46266
rect 1104 46192 5980 46214
rect 94024 46266 97888 46288
rect 94024 46214 96374 46266
rect 96426 46214 96438 46266
rect 96490 46214 96502 46266
rect 96554 46214 96566 46266
rect 96618 46214 96630 46266
rect 96682 46214 97888 46266
rect 94024 46192 97888 46214
rect 1670 45908 1676 45960
rect 1728 45908 1734 45960
rect 97261 45951 97319 45957
rect 97261 45917 97273 45951
rect 97307 45948 97319 45951
rect 97534 45948 97540 45960
rect 97307 45920 97540 45948
rect 97307 45917 97319 45920
rect 97261 45911 97319 45917
rect 97534 45908 97540 45920
rect 97592 45908 97598 45960
rect 842 45772 848 45824
rect 900 45812 906 45824
rect 1489 45815 1547 45821
rect 1489 45812 1501 45815
rect 900 45784 1501 45812
rect 900 45772 906 45784
rect 1489 45781 1501 45784
rect 1535 45781 1547 45815
rect 1489 45775 1547 45781
rect 97353 45815 97411 45821
rect 97353 45781 97365 45815
rect 97399 45812 97411 45815
rect 97442 45812 97448 45824
rect 97399 45784 97448 45812
rect 97399 45781 97411 45784
rect 97353 45775 97411 45781
rect 97442 45772 97448 45784
rect 97500 45772 97506 45824
rect 1104 45722 5980 45744
rect 1104 45670 4874 45722
rect 4926 45670 4938 45722
rect 4990 45670 5002 45722
rect 5054 45670 5066 45722
rect 5118 45670 5130 45722
rect 5182 45670 5980 45722
rect 1104 45648 5980 45670
rect 94024 45722 97888 45744
rect 94024 45670 97034 45722
rect 97086 45670 97098 45722
rect 97150 45670 97162 45722
rect 97214 45670 97226 45722
rect 97278 45670 97290 45722
rect 97342 45670 97888 45722
rect 94024 45648 97888 45670
rect 1104 45178 5980 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 5980 45178
rect 1104 45104 5980 45126
rect 94024 45178 97888 45200
rect 94024 45126 96374 45178
rect 96426 45126 96438 45178
rect 96490 45126 96502 45178
rect 96554 45126 96566 45178
rect 96618 45126 96630 45178
rect 96682 45126 97888 45178
rect 94024 45104 97888 45126
rect 1104 44634 5980 44656
rect 1104 44582 4874 44634
rect 4926 44582 4938 44634
rect 4990 44582 5002 44634
rect 5054 44582 5066 44634
rect 5118 44582 5130 44634
rect 5182 44582 5980 44634
rect 1104 44560 5980 44582
rect 94024 44634 97888 44656
rect 94024 44582 97034 44634
rect 97086 44582 97098 44634
rect 97150 44582 97162 44634
rect 97214 44582 97226 44634
rect 97278 44582 97290 44634
rect 97342 44582 97888 44634
rect 94024 44560 97888 44582
rect 842 44480 848 44532
rect 900 44520 906 44532
rect 1489 44523 1547 44529
rect 1489 44520 1501 44523
rect 900 44492 1501 44520
rect 900 44480 906 44492
rect 1489 44489 1501 44492
rect 1535 44489 1547 44523
rect 1489 44483 1547 44489
rect 1673 44387 1731 44393
rect 1673 44353 1685 44387
rect 1719 44384 1731 44387
rect 8294 44384 8300 44396
rect 1719 44356 8300 44384
rect 1719 44353 1731 44356
rect 1673 44347 1731 44353
rect 8294 44344 8300 44356
rect 8352 44344 8358 44396
rect 97261 44387 97319 44393
rect 97261 44353 97273 44387
rect 97307 44384 97319 44387
rect 97534 44384 97540 44396
rect 97307 44356 97540 44384
rect 97307 44353 97319 44356
rect 97261 44347 97319 44353
rect 97534 44344 97540 44356
rect 97592 44344 97598 44396
rect 97350 44208 97356 44260
rect 97408 44208 97414 44260
rect 1104 44090 5980 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 5980 44090
rect 1104 44016 5980 44038
rect 94024 44090 97888 44112
rect 94024 44038 96374 44090
rect 96426 44038 96438 44090
rect 96490 44038 96502 44090
rect 96554 44038 96566 44090
rect 96618 44038 96630 44090
rect 96682 44038 97888 44090
rect 94024 44016 97888 44038
rect 1104 43546 5980 43568
rect 1104 43494 4874 43546
rect 4926 43494 4938 43546
rect 4990 43494 5002 43546
rect 5054 43494 5066 43546
rect 5118 43494 5130 43546
rect 5182 43494 5980 43546
rect 1104 43472 5980 43494
rect 94024 43546 97888 43568
rect 94024 43494 97034 43546
rect 97086 43494 97098 43546
rect 97150 43494 97162 43546
rect 97214 43494 97226 43546
rect 97278 43494 97290 43546
rect 97342 43494 97888 43546
rect 94024 43472 97888 43494
rect 1673 43299 1731 43305
rect 1673 43265 1685 43299
rect 1719 43296 1731 43299
rect 8294 43296 8300 43308
rect 1719 43268 8300 43296
rect 1719 43265 1731 43268
rect 1673 43259 1731 43265
rect 8294 43256 8300 43268
rect 8352 43256 8358 43308
rect 97261 43299 97319 43305
rect 97261 43265 97273 43299
rect 97307 43296 97319 43299
rect 97534 43296 97540 43308
rect 97307 43268 97540 43296
rect 97307 43265 97319 43268
rect 97261 43259 97319 43265
rect 97534 43256 97540 43268
rect 97592 43256 97598 43308
rect 97350 43120 97356 43172
rect 97408 43120 97414 43172
rect 842 43052 848 43104
rect 900 43092 906 43104
rect 1489 43095 1547 43101
rect 1489 43092 1501 43095
rect 900 43064 1501 43092
rect 900 43052 906 43064
rect 1489 43061 1501 43064
rect 1535 43061 1547 43095
rect 1489 43055 1547 43061
rect 1104 43002 5980 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 5980 43002
rect 1104 42928 5980 42950
rect 94024 43002 97888 43024
rect 94024 42950 96374 43002
rect 96426 42950 96438 43002
rect 96490 42950 96502 43002
rect 96554 42950 96566 43002
rect 96618 42950 96630 43002
rect 96682 42950 97888 43002
rect 94024 42928 97888 42950
rect 1673 42687 1731 42693
rect 1673 42653 1685 42687
rect 1719 42684 1731 42687
rect 8294 42684 8300 42696
rect 1719 42656 8300 42684
rect 1719 42653 1731 42656
rect 1673 42647 1731 42653
rect 8294 42644 8300 42656
rect 8352 42644 8358 42696
rect 97261 42687 97319 42693
rect 97261 42653 97273 42687
rect 97307 42684 97319 42687
rect 97534 42684 97540 42696
rect 97307 42656 97540 42684
rect 97307 42653 97319 42656
rect 97261 42647 97319 42653
rect 97534 42644 97540 42656
rect 97592 42644 97598 42696
rect 842 42508 848 42560
rect 900 42548 906 42560
rect 1489 42551 1547 42557
rect 1489 42548 1501 42551
rect 900 42520 1501 42548
rect 900 42508 906 42520
rect 1489 42517 1501 42520
rect 1535 42517 1547 42551
rect 1489 42511 1547 42517
rect 97353 42551 97411 42557
rect 97353 42517 97365 42551
rect 97399 42548 97411 42551
rect 97442 42548 97448 42560
rect 97399 42520 97448 42548
rect 97399 42517 97411 42520
rect 97353 42511 97411 42517
rect 97442 42508 97448 42520
rect 97500 42508 97506 42560
rect 1104 42458 5980 42480
rect 1104 42406 4874 42458
rect 4926 42406 4938 42458
rect 4990 42406 5002 42458
rect 5054 42406 5066 42458
rect 5118 42406 5130 42458
rect 5182 42406 5980 42458
rect 1104 42384 5980 42406
rect 94024 42458 97888 42480
rect 94024 42406 97034 42458
rect 97086 42406 97098 42458
rect 97150 42406 97162 42458
rect 97214 42406 97226 42458
rect 97278 42406 97290 42458
rect 97342 42406 97888 42458
rect 94024 42384 97888 42406
rect 1104 41914 5980 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 5980 41914
rect 1104 41840 5980 41862
rect 94024 41914 97888 41936
rect 94024 41862 96374 41914
rect 96426 41862 96438 41914
rect 96490 41862 96502 41914
rect 96554 41862 96566 41914
rect 96618 41862 96630 41914
rect 96682 41862 97888 41914
rect 94024 41840 97888 41862
rect 1104 41370 5980 41392
rect 1104 41318 4874 41370
rect 4926 41318 4938 41370
rect 4990 41318 5002 41370
rect 5054 41318 5066 41370
rect 5118 41318 5130 41370
rect 5182 41318 5980 41370
rect 1104 41296 5980 41318
rect 94024 41370 97888 41392
rect 94024 41318 97034 41370
rect 97086 41318 97098 41370
rect 97150 41318 97162 41370
rect 97214 41318 97226 41370
rect 97278 41318 97290 41370
rect 97342 41318 97888 41370
rect 94024 41296 97888 41318
rect 97350 41216 97356 41268
rect 97408 41216 97414 41268
rect 1673 41123 1731 41129
rect 1673 41089 1685 41123
rect 1719 41120 1731 41123
rect 8294 41120 8300 41132
rect 1719 41092 8300 41120
rect 1719 41089 1731 41092
rect 1673 41083 1731 41089
rect 8294 41080 8300 41092
rect 8352 41080 8358 41132
rect 97261 41123 97319 41129
rect 97261 41089 97273 41123
rect 97307 41120 97319 41123
rect 97534 41120 97540 41132
rect 97307 41092 97540 41120
rect 97307 41089 97319 41092
rect 97261 41083 97319 41089
rect 97534 41080 97540 41092
rect 97592 41080 97598 41132
rect 842 40944 848 40996
rect 900 40984 906 40996
rect 1489 40987 1547 40993
rect 1489 40984 1501 40987
rect 900 40956 1501 40984
rect 900 40944 906 40956
rect 1489 40953 1501 40956
rect 1535 40953 1547 40987
rect 1489 40947 1547 40953
rect 1104 40826 5980 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 5980 40826
rect 1104 40752 5980 40774
rect 94024 40826 97888 40848
rect 94024 40774 96374 40826
rect 96426 40774 96438 40826
rect 96490 40774 96502 40826
rect 96554 40774 96566 40826
rect 96618 40774 96630 40826
rect 96682 40774 97888 40826
rect 94024 40752 97888 40774
rect 1670 40468 1676 40520
rect 1728 40468 1734 40520
rect 97261 40511 97319 40517
rect 97261 40477 97273 40511
rect 97307 40508 97319 40511
rect 97534 40508 97540 40520
rect 97307 40480 97540 40508
rect 97307 40477 97319 40480
rect 97261 40471 97319 40477
rect 97534 40468 97540 40480
rect 97592 40468 97598 40520
rect 842 40332 848 40384
rect 900 40372 906 40384
rect 1489 40375 1547 40381
rect 1489 40372 1501 40375
rect 900 40344 1501 40372
rect 900 40332 906 40344
rect 1489 40341 1501 40344
rect 1535 40341 1547 40375
rect 1489 40335 1547 40341
rect 97353 40375 97411 40381
rect 97353 40341 97365 40375
rect 97399 40372 97411 40375
rect 97442 40372 97448 40384
rect 97399 40344 97448 40372
rect 97399 40341 97411 40344
rect 97353 40335 97411 40341
rect 97442 40332 97448 40344
rect 97500 40332 97506 40384
rect 1104 40282 5980 40304
rect 1104 40230 4874 40282
rect 4926 40230 4938 40282
rect 4990 40230 5002 40282
rect 5054 40230 5066 40282
rect 5118 40230 5130 40282
rect 5182 40230 5980 40282
rect 1104 40208 5980 40230
rect 94024 40282 97888 40304
rect 94024 40230 97034 40282
rect 97086 40230 97098 40282
rect 97150 40230 97162 40282
rect 97214 40230 97226 40282
rect 97278 40230 97290 40282
rect 97342 40230 97888 40282
rect 94024 40208 97888 40230
rect 1104 39738 5980 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 5980 39738
rect 1104 39664 5980 39686
rect 94024 39738 97888 39760
rect 94024 39686 96374 39738
rect 96426 39686 96438 39738
rect 96490 39686 96502 39738
rect 96554 39686 96566 39738
rect 96618 39686 96630 39738
rect 96682 39686 97888 39738
rect 94024 39664 97888 39686
rect 1104 39194 5980 39216
rect 1104 39142 4874 39194
rect 4926 39142 4938 39194
rect 4990 39142 5002 39194
rect 5054 39142 5066 39194
rect 5118 39142 5130 39194
rect 5182 39142 5980 39194
rect 1104 39120 5980 39142
rect 94024 39194 97888 39216
rect 94024 39142 97034 39194
rect 97086 39142 97098 39194
rect 97150 39142 97162 39194
rect 97214 39142 97226 39194
rect 97278 39142 97290 39194
rect 97342 39142 97888 39194
rect 94024 39120 97888 39142
rect 97350 39040 97356 39092
rect 97408 39040 97414 39092
rect 1673 38947 1731 38953
rect 1673 38913 1685 38947
rect 1719 38944 1731 38947
rect 8294 38944 8300 38956
rect 1719 38916 8300 38944
rect 1719 38913 1731 38916
rect 1673 38907 1731 38913
rect 8294 38904 8300 38916
rect 8352 38904 8358 38956
rect 97261 38947 97319 38953
rect 97261 38913 97273 38947
rect 97307 38944 97319 38947
rect 97534 38944 97540 38956
rect 97307 38916 97540 38944
rect 97307 38913 97319 38916
rect 97261 38907 97319 38913
rect 97534 38904 97540 38916
rect 97592 38904 97598 38956
rect 842 38700 848 38752
rect 900 38740 906 38752
rect 1489 38743 1547 38749
rect 1489 38740 1501 38743
rect 900 38712 1501 38740
rect 900 38700 906 38712
rect 1489 38709 1501 38712
rect 1535 38709 1547 38743
rect 1489 38703 1547 38709
rect 1104 38650 5980 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 5980 38650
rect 1104 38576 5980 38598
rect 94024 38650 97888 38672
rect 94024 38598 96374 38650
rect 96426 38598 96438 38650
rect 96490 38598 96502 38650
rect 96554 38598 96566 38650
rect 96618 38598 96630 38650
rect 96682 38598 97888 38650
rect 94024 38576 97888 38598
rect 1104 38106 5980 38128
rect 1104 38054 4874 38106
rect 4926 38054 4938 38106
rect 4990 38054 5002 38106
rect 5054 38054 5066 38106
rect 5118 38054 5130 38106
rect 5182 38054 5980 38106
rect 1104 38032 5980 38054
rect 94024 38106 97888 38128
rect 94024 38054 97034 38106
rect 97086 38054 97098 38106
rect 97150 38054 97162 38106
rect 97214 38054 97226 38106
rect 97278 38054 97290 38106
rect 97342 38054 97888 38106
rect 94024 38032 97888 38054
rect 97350 37952 97356 38004
rect 97408 37952 97414 38004
rect 1673 37859 1731 37865
rect 1673 37825 1685 37859
rect 1719 37856 1731 37859
rect 8294 37856 8300 37868
rect 1719 37828 8300 37856
rect 1719 37825 1731 37828
rect 1673 37819 1731 37825
rect 8294 37816 8300 37828
rect 8352 37816 8358 37868
rect 97261 37859 97319 37865
rect 97261 37825 97273 37859
rect 97307 37856 97319 37859
rect 97534 37856 97540 37868
rect 97307 37828 97540 37856
rect 97307 37825 97319 37828
rect 97261 37819 97319 37825
rect 97534 37816 97540 37828
rect 97592 37816 97598 37868
rect 842 37612 848 37664
rect 900 37652 906 37664
rect 1489 37655 1547 37661
rect 1489 37652 1501 37655
rect 900 37624 1501 37652
rect 900 37612 906 37624
rect 1489 37621 1501 37624
rect 1535 37621 1547 37655
rect 1489 37615 1547 37621
rect 1104 37562 5980 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 5980 37562
rect 1104 37488 5980 37510
rect 94024 37562 97888 37584
rect 94024 37510 96374 37562
rect 96426 37510 96438 37562
rect 96490 37510 96502 37562
rect 96554 37510 96566 37562
rect 96618 37510 96630 37562
rect 96682 37510 97888 37562
rect 94024 37488 97888 37510
rect 96614 37272 96620 37324
rect 96672 37312 96678 37324
rect 97261 37315 97319 37321
rect 97261 37312 97273 37315
rect 96672 37284 97273 37312
rect 96672 37272 96678 37284
rect 97261 37281 97273 37284
rect 97307 37281 97319 37315
rect 97261 37275 97319 37281
rect 1673 37247 1731 37253
rect 1673 37213 1685 37247
rect 1719 37244 1731 37247
rect 8294 37244 8300 37256
rect 1719 37216 8300 37244
rect 1719 37213 1731 37216
rect 1673 37207 1731 37213
rect 8294 37204 8300 37216
rect 8352 37204 8358 37256
rect 97169 37179 97227 37185
rect 97169 37145 97181 37179
rect 97215 37176 97227 37179
rect 97442 37176 97448 37188
rect 97215 37148 97448 37176
rect 97215 37145 97227 37148
rect 97169 37139 97227 37145
rect 97442 37136 97448 37148
rect 97500 37136 97506 37188
rect 842 37068 848 37120
rect 900 37108 906 37120
rect 1489 37111 1547 37117
rect 1489 37108 1501 37111
rect 900 37080 1501 37108
rect 900 37068 906 37080
rect 1489 37077 1501 37080
rect 1535 37077 1547 37111
rect 1489 37071 1547 37077
rect 1104 37018 5980 37040
rect 1104 36966 4874 37018
rect 4926 36966 4938 37018
rect 4990 36966 5002 37018
rect 5054 36966 5066 37018
rect 5118 36966 5130 37018
rect 5182 36966 5980 37018
rect 1104 36944 5980 36966
rect 94024 37018 97888 37040
rect 94024 36966 97034 37018
rect 97086 36966 97098 37018
rect 97150 36966 97162 37018
rect 97214 36966 97226 37018
rect 97278 36966 97290 37018
rect 97342 36966 97888 37018
rect 94024 36944 97888 36966
rect 1104 36474 5980 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 5980 36474
rect 1104 36400 5980 36422
rect 94024 36474 97888 36496
rect 94024 36422 96374 36474
rect 96426 36422 96438 36474
rect 96490 36422 96502 36474
rect 96554 36422 96566 36474
rect 96618 36422 96630 36474
rect 96682 36422 97888 36474
rect 94024 36400 97888 36422
rect 1104 35930 5980 35952
rect 1104 35878 4874 35930
rect 4926 35878 4938 35930
rect 4990 35878 5002 35930
rect 5054 35878 5066 35930
rect 5118 35878 5130 35930
rect 5182 35878 5980 35930
rect 1104 35856 5980 35878
rect 94024 35930 97888 35952
rect 94024 35878 97034 35930
rect 97086 35878 97098 35930
rect 97150 35878 97162 35930
rect 97214 35878 97226 35930
rect 97278 35878 97290 35930
rect 97342 35878 97888 35930
rect 94024 35856 97888 35878
rect 97350 35776 97356 35828
rect 97408 35776 97414 35828
rect 1673 35683 1731 35689
rect 1673 35649 1685 35683
rect 1719 35680 1731 35683
rect 8294 35680 8300 35692
rect 1719 35652 8300 35680
rect 1719 35649 1731 35652
rect 1673 35643 1731 35649
rect 8294 35640 8300 35652
rect 8352 35640 8358 35692
rect 97261 35683 97319 35689
rect 97261 35649 97273 35683
rect 97307 35680 97319 35683
rect 97534 35680 97540 35692
rect 97307 35652 97540 35680
rect 97307 35649 97319 35652
rect 97261 35643 97319 35649
rect 97534 35640 97540 35652
rect 97592 35640 97598 35692
rect 842 35504 848 35556
rect 900 35544 906 35556
rect 1489 35547 1547 35553
rect 1489 35544 1501 35547
rect 900 35516 1501 35544
rect 900 35504 906 35516
rect 1489 35513 1501 35516
rect 1535 35513 1547 35547
rect 1489 35507 1547 35513
rect 1104 35386 5980 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 5980 35386
rect 1104 35312 5980 35334
rect 94024 35386 97888 35408
rect 94024 35334 96374 35386
rect 96426 35334 96438 35386
rect 96490 35334 96502 35386
rect 96554 35334 96566 35386
rect 96618 35334 96630 35386
rect 96682 35334 97888 35386
rect 94024 35312 97888 35334
rect 1670 35028 1676 35080
rect 1728 35028 1734 35080
rect 97261 35071 97319 35077
rect 97261 35037 97273 35071
rect 97307 35068 97319 35071
rect 97534 35068 97540 35080
rect 97307 35040 97540 35068
rect 97307 35037 97319 35040
rect 97261 35031 97319 35037
rect 97534 35028 97540 35040
rect 97592 35028 97598 35080
rect 842 34892 848 34944
rect 900 34932 906 34944
rect 1489 34935 1547 34941
rect 1489 34932 1501 34935
rect 900 34904 1501 34932
rect 900 34892 906 34904
rect 1489 34901 1501 34904
rect 1535 34901 1547 34935
rect 1489 34895 1547 34901
rect 97353 34935 97411 34941
rect 97353 34901 97365 34935
rect 97399 34932 97411 34935
rect 97442 34932 97448 34944
rect 97399 34904 97448 34932
rect 97399 34901 97411 34904
rect 97353 34895 97411 34901
rect 97442 34892 97448 34904
rect 97500 34892 97506 34944
rect 1104 34842 5980 34864
rect 1104 34790 4874 34842
rect 4926 34790 4938 34842
rect 4990 34790 5002 34842
rect 5054 34790 5066 34842
rect 5118 34790 5130 34842
rect 5182 34790 5980 34842
rect 1104 34768 5980 34790
rect 94024 34842 97888 34864
rect 94024 34790 97034 34842
rect 97086 34790 97098 34842
rect 97150 34790 97162 34842
rect 97214 34790 97226 34842
rect 97278 34790 97290 34842
rect 97342 34790 97888 34842
rect 94024 34768 97888 34790
rect 1104 34298 5980 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 5980 34298
rect 1104 34224 5980 34246
rect 94024 34298 97888 34320
rect 94024 34246 96374 34298
rect 96426 34246 96438 34298
rect 96490 34246 96502 34298
rect 96554 34246 96566 34298
rect 96618 34246 96630 34298
rect 96682 34246 97888 34298
rect 94024 34224 97888 34246
rect 1104 33754 5980 33776
rect 1104 33702 4874 33754
rect 4926 33702 4938 33754
rect 4990 33702 5002 33754
rect 5054 33702 5066 33754
rect 5118 33702 5130 33754
rect 5182 33702 5980 33754
rect 1104 33680 5980 33702
rect 94024 33754 97888 33776
rect 94024 33702 97034 33754
rect 97086 33702 97098 33754
rect 97150 33702 97162 33754
rect 97214 33702 97226 33754
rect 97278 33702 97290 33754
rect 97342 33702 97888 33754
rect 94024 33680 97888 33702
rect 97350 33600 97356 33652
rect 97408 33600 97414 33652
rect 1673 33507 1731 33513
rect 1673 33473 1685 33507
rect 1719 33504 1731 33507
rect 8294 33504 8300 33516
rect 1719 33476 8300 33504
rect 1719 33473 1731 33476
rect 1673 33467 1731 33473
rect 8294 33464 8300 33476
rect 8352 33464 8358 33516
rect 97261 33507 97319 33513
rect 97261 33473 97273 33507
rect 97307 33504 97319 33507
rect 97534 33504 97540 33516
rect 97307 33476 97540 33504
rect 97307 33473 97319 33476
rect 97261 33467 97319 33473
rect 97534 33464 97540 33476
rect 97592 33464 97598 33516
rect 842 33260 848 33312
rect 900 33300 906 33312
rect 1489 33303 1547 33309
rect 1489 33300 1501 33303
rect 900 33272 1501 33300
rect 900 33260 906 33272
rect 1489 33269 1501 33272
rect 1535 33269 1547 33303
rect 1489 33263 1547 33269
rect 1104 33210 5980 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 5980 33210
rect 1104 33136 5980 33158
rect 94024 33210 97888 33232
rect 94024 33158 96374 33210
rect 96426 33158 96438 33210
rect 96490 33158 96502 33210
rect 96554 33158 96566 33210
rect 96618 33158 96630 33210
rect 96682 33158 97888 33210
rect 94024 33136 97888 33158
rect 1104 32666 5980 32688
rect 1104 32614 4874 32666
rect 4926 32614 4938 32666
rect 4990 32614 5002 32666
rect 5054 32614 5066 32666
rect 5118 32614 5130 32666
rect 5182 32614 5980 32666
rect 1104 32592 5980 32614
rect 94024 32666 97888 32688
rect 94024 32614 97034 32666
rect 97086 32614 97098 32666
rect 97150 32614 97162 32666
rect 97214 32614 97226 32666
rect 97278 32614 97290 32666
rect 97342 32614 97888 32666
rect 94024 32592 97888 32614
rect 97258 32444 97264 32496
rect 97316 32444 97322 32496
rect 1673 32419 1731 32425
rect 1673 32385 1685 32419
rect 1719 32416 1731 32419
rect 8294 32416 8300 32428
rect 1719 32388 8300 32416
rect 1719 32385 1731 32388
rect 1673 32379 1731 32385
rect 8294 32376 8300 32388
rect 8352 32376 8358 32428
rect 97169 32419 97227 32425
rect 97169 32385 97181 32419
rect 97215 32416 97227 32419
rect 97442 32416 97448 32428
rect 97215 32388 97448 32416
rect 97215 32385 97227 32388
rect 97169 32379 97227 32385
rect 97442 32376 97448 32388
rect 97500 32376 97506 32428
rect 842 32172 848 32224
rect 900 32212 906 32224
rect 1489 32215 1547 32221
rect 1489 32212 1501 32215
rect 900 32184 1501 32212
rect 900 32172 906 32184
rect 1489 32181 1501 32184
rect 1535 32181 1547 32215
rect 1489 32175 1547 32181
rect 1104 32122 5980 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 5980 32122
rect 1104 32048 5980 32070
rect 94024 32122 97888 32144
rect 94024 32070 96374 32122
rect 96426 32070 96438 32122
rect 96490 32070 96502 32122
rect 96554 32070 96566 32122
rect 96618 32070 96630 32122
rect 96682 32070 97888 32122
rect 94024 32048 97888 32070
rect 842 31900 848 31952
rect 900 31940 906 31952
rect 1489 31943 1547 31949
rect 1489 31940 1501 31943
rect 900 31912 1501 31940
rect 900 31900 906 31912
rect 1489 31909 1501 31912
rect 1535 31909 1547 31943
rect 1489 31903 1547 31909
rect 96614 31900 96620 31952
rect 96672 31940 96678 31952
rect 97353 31943 97411 31949
rect 97353 31940 97365 31943
rect 96672 31912 97365 31940
rect 96672 31900 96678 31912
rect 97353 31909 97365 31912
rect 97399 31909 97411 31943
rect 97353 31903 97411 31909
rect 1670 31764 1676 31816
rect 1728 31764 1734 31816
rect 97261 31807 97319 31813
rect 97261 31773 97273 31807
rect 97307 31804 97319 31807
rect 97534 31804 97540 31816
rect 97307 31776 97540 31804
rect 97307 31773 97319 31776
rect 97261 31767 97319 31773
rect 97534 31764 97540 31776
rect 97592 31764 97598 31816
rect 1104 31578 5980 31600
rect 1104 31526 4874 31578
rect 4926 31526 4938 31578
rect 4990 31526 5002 31578
rect 5054 31526 5066 31578
rect 5118 31526 5130 31578
rect 5182 31526 5980 31578
rect 1104 31504 5980 31526
rect 94024 31578 97888 31600
rect 94024 31526 97034 31578
rect 97086 31526 97098 31578
rect 97150 31526 97162 31578
rect 97214 31526 97226 31578
rect 97278 31526 97290 31578
rect 97342 31526 97888 31578
rect 94024 31504 97888 31526
rect 1104 31034 5980 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 5980 31034
rect 1104 30960 5980 30982
rect 94024 31034 97888 31056
rect 94024 30982 96374 31034
rect 96426 30982 96438 31034
rect 96490 30982 96502 31034
rect 96554 30982 96566 31034
rect 96618 30982 96630 31034
rect 96682 30982 97888 31034
rect 94024 30960 97888 30982
rect 97534 30540 97540 30592
rect 97592 30540 97598 30592
rect 1104 30490 5980 30512
rect 1104 30438 4874 30490
rect 4926 30438 4938 30490
rect 4990 30438 5002 30490
rect 5054 30438 5066 30490
rect 5118 30438 5130 30490
rect 5182 30438 5980 30490
rect 1104 30416 5980 30438
rect 94024 30490 97888 30512
rect 94024 30438 97034 30490
rect 97086 30438 97098 30490
rect 97150 30438 97162 30490
rect 97214 30438 97226 30490
rect 97278 30438 97290 30490
rect 97342 30438 97888 30490
rect 94024 30416 97888 30438
rect 1673 30243 1731 30249
rect 1673 30209 1685 30243
rect 1719 30240 1731 30243
rect 8294 30240 8300 30252
rect 1719 30212 8300 30240
rect 1719 30209 1731 30212
rect 1673 30203 1731 30209
rect 8294 30200 8300 30212
rect 8352 30200 8358 30252
rect 97258 30200 97264 30252
rect 97316 30200 97322 30252
rect 97534 30132 97540 30184
rect 97592 30132 97598 30184
rect 842 30064 848 30116
rect 900 30104 906 30116
rect 1489 30107 1547 30113
rect 1489 30104 1501 30107
rect 900 30076 1501 30104
rect 900 30064 906 30076
rect 1489 30073 1501 30076
rect 1535 30073 1547 30107
rect 1489 30067 1547 30073
rect 1104 29946 5980 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 5980 29946
rect 1104 29872 5980 29894
rect 94024 29946 97888 29968
rect 94024 29894 96374 29946
rect 96426 29894 96438 29946
rect 96490 29894 96502 29946
rect 96554 29894 96566 29946
rect 96618 29894 96630 29946
rect 96682 29894 97888 29946
rect 94024 29872 97888 29894
rect 1673 29631 1731 29637
rect 1673 29597 1685 29631
rect 1719 29628 1731 29631
rect 8294 29628 8300 29640
rect 1719 29600 8300 29628
rect 1719 29597 1731 29600
rect 1673 29591 1731 29597
rect 8294 29588 8300 29600
rect 8352 29588 8358 29640
rect 97261 29631 97319 29637
rect 97261 29597 97273 29631
rect 97307 29628 97319 29631
rect 97534 29628 97540 29640
rect 97307 29600 97540 29628
rect 97307 29597 97319 29600
rect 97261 29591 97319 29597
rect 97534 29588 97540 29600
rect 97592 29588 97598 29640
rect 842 29452 848 29504
rect 900 29492 906 29504
rect 1489 29495 1547 29501
rect 1489 29492 1501 29495
rect 900 29464 1501 29492
rect 900 29452 906 29464
rect 1489 29461 1501 29464
rect 1535 29461 1547 29495
rect 1489 29455 1547 29461
rect 97353 29495 97411 29501
rect 97353 29461 97365 29495
rect 97399 29492 97411 29495
rect 97442 29492 97448 29504
rect 97399 29464 97448 29492
rect 97399 29461 97411 29464
rect 97353 29455 97411 29461
rect 97442 29452 97448 29464
rect 97500 29452 97506 29504
rect 1104 29402 5980 29424
rect 1104 29350 4874 29402
rect 4926 29350 4938 29402
rect 4990 29350 5002 29402
rect 5054 29350 5066 29402
rect 5118 29350 5130 29402
rect 5182 29350 5980 29402
rect 1104 29328 5980 29350
rect 94024 29402 97888 29424
rect 94024 29350 97034 29402
rect 97086 29350 97098 29402
rect 97150 29350 97162 29402
rect 97214 29350 97226 29402
rect 97278 29350 97290 29402
rect 97342 29350 97888 29402
rect 94024 29328 97888 29350
rect 1104 28858 5980 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 5980 28858
rect 1104 28784 5980 28806
rect 94024 28858 97888 28880
rect 94024 28806 96374 28858
rect 96426 28806 96438 28858
rect 96490 28806 96502 28858
rect 96554 28806 96566 28858
rect 96618 28806 96630 28858
rect 96682 28806 97888 28858
rect 94024 28784 97888 28806
rect 1104 28314 5980 28336
rect 1104 28262 4874 28314
rect 4926 28262 4938 28314
rect 4990 28262 5002 28314
rect 5054 28262 5066 28314
rect 5118 28262 5130 28314
rect 5182 28262 5980 28314
rect 1104 28240 5980 28262
rect 94024 28314 97888 28336
rect 94024 28262 97034 28314
rect 97086 28262 97098 28314
rect 97150 28262 97162 28314
rect 97214 28262 97226 28314
rect 97278 28262 97290 28314
rect 97342 28262 97888 28314
rect 94024 28240 97888 28262
rect 1581 28203 1639 28209
rect 1581 28169 1593 28203
rect 1627 28200 1639 28203
rect 8294 28200 8300 28212
rect 1627 28172 8300 28200
rect 1627 28169 1639 28172
rect 1581 28163 1639 28169
rect 8294 28160 8300 28172
rect 8352 28160 8358 28212
rect 1302 28024 1308 28076
rect 1360 28064 1366 28076
rect 1397 28067 1455 28073
rect 1397 28064 1409 28067
rect 1360 28036 1409 28064
rect 1360 28024 1366 28036
rect 1397 28033 1409 28036
rect 1443 28064 1455 28067
rect 1673 28067 1731 28073
rect 1673 28064 1685 28067
rect 1443 28036 1685 28064
rect 1443 28033 1455 28036
rect 1397 28027 1455 28033
rect 1673 28033 1685 28036
rect 1719 28033 1731 28067
rect 1673 28027 1731 28033
rect 97258 28024 97264 28076
rect 97316 28024 97322 28076
rect 97442 27888 97448 27940
rect 97500 27888 97506 27940
rect 1104 27770 5980 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 5980 27770
rect 1104 27696 5980 27718
rect 94024 27770 97888 27792
rect 94024 27718 96374 27770
rect 96426 27718 96438 27770
rect 96490 27718 96502 27770
rect 96554 27718 96566 27770
rect 96618 27718 96630 27770
rect 96682 27718 97888 27770
rect 94024 27696 97888 27718
rect 1104 27226 5980 27248
rect 1104 27174 4874 27226
rect 4926 27174 4938 27226
rect 4990 27174 5002 27226
rect 5054 27174 5066 27226
rect 5118 27174 5130 27226
rect 5182 27174 5980 27226
rect 1104 27152 5980 27174
rect 94024 27226 97888 27248
rect 94024 27174 97034 27226
rect 97086 27174 97098 27226
rect 97150 27174 97162 27226
rect 97214 27174 97226 27226
rect 97278 27174 97290 27226
rect 97342 27174 97888 27226
rect 94024 27152 97888 27174
rect 1302 26936 1308 26988
rect 1360 26976 1366 26988
rect 1489 26979 1547 26985
rect 1489 26976 1501 26979
rect 1360 26948 1501 26976
rect 1360 26936 1366 26948
rect 1489 26945 1501 26948
rect 1535 26945 1547 26979
rect 1489 26939 1547 26945
rect 1673 26979 1731 26985
rect 1673 26945 1685 26979
rect 1719 26976 1731 26979
rect 8294 26976 8300 26988
rect 1719 26948 8300 26976
rect 1719 26945 1731 26948
rect 1673 26939 1731 26945
rect 1504 26908 1532 26939
rect 8294 26936 8300 26948
rect 8352 26936 8358 26988
rect 97258 26936 97264 26988
rect 97316 26936 97322 26988
rect 1765 26911 1823 26917
rect 1765 26908 1777 26911
rect 1504 26880 1777 26908
rect 1765 26877 1777 26880
rect 1811 26877 1823 26911
rect 1765 26871 1823 26877
rect 97442 26732 97448 26784
rect 97500 26732 97506 26784
rect 1104 26682 5980 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 5980 26682
rect 1104 26608 5980 26630
rect 94024 26682 97888 26704
rect 94024 26630 96374 26682
rect 96426 26630 96438 26682
rect 96490 26630 96502 26682
rect 96554 26630 96566 26682
rect 96618 26630 96630 26682
rect 96682 26630 97888 26682
rect 94024 26608 97888 26630
rect 97442 26460 97448 26512
rect 97500 26460 97506 26512
rect 1302 26324 1308 26376
rect 1360 26364 1366 26376
rect 1489 26367 1547 26373
rect 1489 26364 1501 26367
rect 1360 26336 1501 26364
rect 1360 26324 1366 26336
rect 1489 26333 1501 26336
rect 1535 26364 1547 26367
rect 1765 26367 1823 26373
rect 1765 26364 1777 26367
rect 1535 26336 1777 26364
rect 1535 26333 1547 26336
rect 1489 26327 1547 26333
rect 1765 26333 1777 26336
rect 1811 26333 1823 26367
rect 1765 26327 1823 26333
rect 96890 26324 96896 26376
rect 96948 26364 96954 26376
rect 97261 26367 97319 26373
rect 97261 26364 97273 26367
rect 96948 26336 97273 26364
rect 96948 26324 96954 26336
rect 97261 26333 97273 26336
rect 97307 26333 97319 26367
rect 97261 26327 97319 26333
rect 1670 26256 1676 26308
rect 1728 26256 1734 26308
rect 1104 26138 5980 26160
rect 1104 26086 4874 26138
rect 4926 26086 4938 26138
rect 4990 26086 5002 26138
rect 5054 26086 5066 26138
rect 5118 26086 5130 26138
rect 5182 26086 5980 26138
rect 1104 26064 5980 26086
rect 94024 26138 97888 26160
rect 94024 26086 97034 26138
rect 97086 26086 97098 26138
rect 97150 26086 97162 26138
rect 97214 26086 97226 26138
rect 97278 26086 97290 26138
rect 97342 26086 97888 26138
rect 94024 26064 97888 26086
rect 1104 25594 5980 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 5980 25594
rect 1104 25520 5980 25542
rect 94024 25594 97888 25616
rect 94024 25542 96374 25594
rect 96426 25542 96438 25594
rect 96490 25542 96502 25594
rect 96554 25542 96566 25594
rect 96618 25542 96630 25594
rect 96682 25542 97888 25594
rect 94024 25520 97888 25542
rect 1104 25050 5980 25072
rect 1104 24998 4874 25050
rect 4926 24998 4938 25050
rect 4990 24998 5002 25050
rect 5054 24998 5066 25050
rect 5118 24998 5130 25050
rect 5182 24998 5980 25050
rect 1104 24976 5980 24998
rect 94024 25050 97888 25072
rect 94024 24998 97034 25050
rect 97086 24998 97098 25050
rect 97150 24998 97162 25050
rect 97214 24998 97226 25050
rect 97278 24998 97290 25050
rect 97342 24998 97888 25050
rect 94024 24976 97888 24998
rect 1302 24760 1308 24812
rect 1360 24800 1366 24812
rect 1489 24803 1547 24809
rect 1489 24800 1501 24803
rect 1360 24772 1501 24800
rect 1360 24760 1366 24772
rect 1489 24769 1501 24772
rect 1535 24769 1547 24803
rect 1489 24763 1547 24769
rect 1673 24803 1731 24809
rect 1673 24769 1685 24803
rect 1719 24800 1731 24803
rect 8294 24800 8300 24812
rect 1719 24772 8300 24800
rect 1719 24769 1731 24772
rect 1673 24763 1731 24769
rect 1504 24732 1532 24763
rect 8294 24760 8300 24772
rect 8352 24760 8358 24812
rect 97258 24760 97264 24812
rect 97316 24760 97322 24812
rect 1765 24735 1823 24741
rect 1765 24732 1777 24735
rect 1504 24704 1777 24732
rect 1765 24701 1777 24704
rect 1811 24701 1823 24735
rect 1765 24695 1823 24701
rect 97442 24556 97448 24608
rect 97500 24556 97506 24608
rect 1104 24506 5980 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 5980 24506
rect 1104 24432 5980 24454
rect 94024 24506 97888 24528
rect 94024 24454 96374 24506
rect 96426 24454 96438 24506
rect 96490 24454 96502 24506
rect 96554 24454 96566 24506
rect 96618 24454 96630 24506
rect 96682 24454 97888 24506
rect 94024 24432 97888 24454
rect 96614 24148 96620 24200
rect 96672 24188 96678 24200
rect 97261 24191 97319 24197
rect 97261 24188 97273 24191
rect 96672 24160 97273 24188
rect 96672 24148 96678 24160
rect 97261 24157 97273 24160
rect 97307 24157 97319 24191
rect 97261 24151 97319 24157
rect 1302 24080 1308 24132
rect 1360 24120 1366 24132
rect 1489 24123 1547 24129
rect 1489 24120 1501 24123
rect 1360 24092 1501 24120
rect 1360 24080 1366 24092
rect 1489 24089 1501 24092
rect 1535 24089 1547 24123
rect 1489 24083 1547 24089
rect 1673 24123 1731 24129
rect 1673 24089 1685 24123
rect 1719 24120 1731 24123
rect 8294 24120 8300 24132
rect 1719 24092 8300 24120
rect 1719 24089 1731 24092
rect 1673 24083 1731 24089
rect 1504 24052 1532 24083
rect 8294 24080 8300 24092
rect 8352 24080 8358 24132
rect 1765 24055 1823 24061
rect 1765 24052 1777 24055
rect 1504 24024 1777 24052
rect 1765 24021 1777 24024
rect 1811 24021 1823 24055
rect 1765 24015 1823 24021
rect 97442 24012 97448 24064
rect 97500 24012 97506 24064
rect 1104 23962 5980 23984
rect 1104 23910 4874 23962
rect 4926 23910 4938 23962
rect 4990 23910 5002 23962
rect 5054 23910 5066 23962
rect 5118 23910 5130 23962
rect 5182 23910 5980 23962
rect 1104 23888 5980 23910
rect 94024 23962 97888 23984
rect 94024 23910 97034 23962
rect 97086 23910 97098 23962
rect 97150 23910 97162 23962
rect 97214 23910 97226 23962
rect 97278 23910 97290 23962
rect 97342 23910 97888 23962
rect 94024 23888 97888 23910
rect 1104 23418 5980 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 5980 23418
rect 1104 23344 5980 23366
rect 94024 23418 97888 23440
rect 94024 23366 96374 23418
rect 96426 23366 96438 23418
rect 96490 23366 96502 23418
rect 96554 23366 96566 23418
rect 96618 23366 96630 23418
rect 96682 23366 97888 23418
rect 94024 23344 97888 23366
rect 1104 22874 5980 22896
rect 1104 22822 4874 22874
rect 4926 22822 4938 22874
rect 4990 22822 5002 22874
rect 5054 22822 5066 22874
rect 5118 22822 5130 22874
rect 5182 22822 5980 22874
rect 1104 22800 5980 22822
rect 94024 22874 97888 22896
rect 94024 22822 97034 22874
rect 97086 22822 97098 22874
rect 97150 22822 97162 22874
rect 97214 22822 97226 22874
rect 97278 22822 97290 22874
rect 97342 22822 97888 22874
rect 94024 22800 97888 22822
rect 1118 22584 1124 22636
rect 1176 22624 1182 22636
rect 1489 22627 1547 22633
rect 1489 22624 1501 22627
rect 1176 22596 1501 22624
rect 1176 22584 1182 22596
rect 1489 22593 1501 22596
rect 1535 22593 1547 22627
rect 1489 22587 1547 22593
rect 1673 22627 1731 22633
rect 1673 22593 1685 22627
rect 1719 22624 1731 22627
rect 8294 22624 8300 22636
rect 1719 22596 8300 22624
rect 1719 22593 1731 22596
rect 1673 22587 1731 22593
rect 1504 22556 1532 22587
rect 8294 22584 8300 22596
rect 8352 22584 8358 22636
rect 97258 22584 97264 22636
rect 97316 22584 97322 22636
rect 1765 22559 1823 22565
rect 1765 22556 1777 22559
rect 1504 22528 1777 22556
rect 1765 22525 1777 22528
rect 1811 22525 1823 22559
rect 1765 22519 1823 22525
rect 97442 22448 97448 22500
rect 97500 22448 97506 22500
rect 1104 22330 5980 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 5980 22330
rect 1104 22256 5980 22278
rect 94024 22330 97888 22352
rect 94024 22278 96374 22330
rect 96426 22278 96438 22330
rect 96490 22278 96502 22330
rect 96554 22278 96566 22330
rect 96618 22278 96630 22330
rect 96682 22278 97888 22330
rect 94024 22256 97888 22278
rect 1104 21786 5980 21808
rect 1104 21734 4874 21786
rect 4926 21734 4938 21786
rect 4990 21734 5002 21786
rect 5054 21734 5066 21786
rect 5118 21734 5130 21786
rect 5182 21734 5980 21786
rect 1104 21712 5980 21734
rect 94024 21786 97888 21808
rect 94024 21734 97034 21786
rect 97086 21734 97098 21786
rect 97150 21734 97162 21786
rect 97214 21734 97226 21786
rect 97278 21734 97290 21786
rect 97342 21734 97888 21786
rect 94024 21712 97888 21734
rect 1302 21496 1308 21548
rect 1360 21536 1366 21548
rect 1489 21539 1547 21545
rect 1489 21536 1501 21539
rect 1360 21508 1501 21536
rect 1360 21496 1366 21508
rect 1489 21505 1501 21508
rect 1535 21505 1547 21539
rect 1489 21499 1547 21505
rect 1673 21539 1731 21545
rect 1673 21505 1685 21539
rect 1719 21536 1731 21539
rect 8294 21536 8300 21548
rect 1719 21508 8300 21536
rect 1719 21505 1731 21508
rect 1673 21499 1731 21505
rect 1504 21468 1532 21499
rect 8294 21496 8300 21508
rect 8352 21496 8358 21548
rect 97258 21496 97264 21548
rect 97316 21496 97322 21548
rect 1765 21471 1823 21477
rect 1765 21468 1777 21471
rect 1504 21440 1777 21468
rect 1765 21437 1777 21440
rect 1811 21437 1823 21471
rect 1765 21431 1823 21437
rect 97442 21292 97448 21344
rect 97500 21292 97506 21344
rect 1104 21242 5980 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 5980 21242
rect 1104 21168 5980 21190
rect 94024 21242 97888 21264
rect 94024 21190 96374 21242
rect 96426 21190 96438 21242
rect 96490 21190 96502 21242
rect 96554 21190 96566 21242
rect 96618 21190 96630 21242
rect 96682 21190 97888 21242
rect 94024 21168 97888 21190
rect 96614 20884 96620 20936
rect 96672 20924 96678 20936
rect 97261 20927 97319 20933
rect 97261 20924 97273 20927
rect 96672 20896 97273 20924
rect 96672 20884 96678 20896
rect 97261 20893 97273 20896
rect 97307 20893 97319 20927
rect 97261 20887 97319 20893
rect 1302 20816 1308 20868
rect 1360 20856 1366 20868
rect 1489 20859 1547 20865
rect 1489 20856 1501 20859
rect 1360 20828 1501 20856
rect 1360 20816 1366 20828
rect 1489 20825 1501 20828
rect 1535 20825 1547 20859
rect 1489 20819 1547 20825
rect 1504 20788 1532 20819
rect 1854 20816 1860 20868
rect 1912 20816 1918 20868
rect 1949 20791 2007 20797
rect 1949 20788 1961 20791
rect 1504 20760 1961 20788
rect 1949 20757 1961 20760
rect 1995 20757 2007 20791
rect 1949 20751 2007 20757
rect 97442 20748 97448 20800
rect 97500 20748 97506 20800
rect 1104 20698 5980 20720
rect 1104 20646 4874 20698
rect 4926 20646 4938 20698
rect 4990 20646 5002 20698
rect 5054 20646 5066 20698
rect 5118 20646 5130 20698
rect 5182 20646 5980 20698
rect 1104 20624 5980 20646
rect 94024 20698 97888 20720
rect 94024 20646 97034 20698
rect 97086 20646 97098 20698
rect 97150 20646 97162 20698
rect 97214 20646 97226 20698
rect 97278 20646 97290 20698
rect 97342 20646 97888 20698
rect 94024 20624 97888 20646
rect 1104 20154 5980 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 5980 20154
rect 1104 20080 5980 20102
rect 94024 20154 97888 20176
rect 94024 20102 96374 20154
rect 96426 20102 96438 20154
rect 96490 20102 96502 20154
rect 96554 20102 96566 20154
rect 96618 20102 96630 20154
rect 96682 20102 97888 20154
rect 94024 20080 97888 20102
rect 1104 19610 5980 19632
rect 1104 19558 4874 19610
rect 4926 19558 4938 19610
rect 4990 19558 5002 19610
rect 5054 19558 5066 19610
rect 5118 19558 5130 19610
rect 5182 19558 5980 19610
rect 1104 19536 5980 19558
rect 94024 19610 97888 19632
rect 94024 19558 97034 19610
rect 97086 19558 97098 19610
rect 97150 19558 97162 19610
rect 97214 19558 97226 19610
rect 97278 19558 97290 19610
rect 97342 19558 97888 19610
rect 94024 19536 97888 19558
rect 97442 19456 97448 19508
rect 97500 19456 97506 19508
rect 1486 19320 1492 19372
rect 1544 19360 1550 19372
rect 1765 19363 1823 19369
rect 1765 19360 1777 19363
rect 1544 19332 1777 19360
rect 1544 19320 1550 19332
rect 1765 19329 1777 19332
rect 1811 19329 1823 19363
rect 1765 19323 1823 19329
rect 97258 19320 97264 19372
rect 97316 19320 97322 19372
rect 1673 19227 1731 19233
rect 1673 19193 1685 19227
rect 1719 19224 1731 19227
rect 8294 19224 8300 19236
rect 1719 19196 8300 19224
rect 1719 19193 1731 19196
rect 1673 19187 1731 19193
rect 8294 19184 8300 19196
rect 8352 19184 8358 19236
rect 1104 19066 5980 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 5980 19066
rect 1104 18992 5980 19014
rect 94024 19066 97888 19088
rect 94024 19014 96374 19066
rect 96426 19014 96438 19066
rect 96490 19014 96502 19066
rect 96554 19014 96566 19066
rect 96618 19014 96630 19066
rect 96682 19014 97888 19066
rect 94024 18992 97888 19014
rect 96614 18708 96620 18760
rect 96672 18748 96678 18760
rect 97261 18751 97319 18757
rect 97261 18748 97273 18751
rect 96672 18720 97273 18748
rect 96672 18708 96678 18720
rect 97261 18717 97273 18720
rect 97307 18717 97319 18751
rect 97261 18711 97319 18717
rect 1302 18640 1308 18692
rect 1360 18680 1366 18692
rect 1489 18683 1547 18689
rect 1489 18680 1501 18683
rect 1360 18652 1501 18680
rect 1360 18640 1366 18652
rect 1489 18649 1501 18652
rect 1535 18649 1547 18683
rect 1489 18643 1547 18649
rect 1857 18683 1915 18689
rect 1857 18649 1869 18683
rect 1903 18680 1915 18683
rect 8294 18680 8300 18692
rect 1903 18652 8300 18680
rect 1903 18649 1915 18652
rect 1857 18643 1915 18649
rect 1504 18612 1532 18643
rect 8294 18640 8300 18652
rect 8352 18640 8358 18692
rect 1949 18615 2007 18621
rect 1949 18612 1961 18615
rect 1504 18584 1961 18612
rect 1949 18581 1961 18584
rect 1995 18581 2007 18615
rect 1949 18575 2007 18581
rect 97442 18572 97448 18624
rect 97500 18572 97506 18624
rect 1104 18522 5980 18544
rect 1104 18470 4874 18522
rect 4926 18470 4938 18522
rect 4990 18470 5002 18522
rect 5054 18470 5066 18522
rect 5118 18470 5130 18522
rect 5182 18470 5980 18522
rect 1104 18448 5980 18470
rect 94024 18522 97888 18544
rect 94024 18470 97034 18522
rect 97086 18470 97098 18522
rect 97150 18470 97162 18522
rect 97214 18470 97226 18522
rect 97278 18470 97290 18522
rect 97342 18470 97888 18522
rect 94024 18448 97888 18470
rect 1104 17978 5980 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 5980 17978
rect 1104 17904 5980 17926
rect 94024 17978 97888 18000
rect 94024 17926 96374 17978
rect 96426 17926 96438 17978
rect 96490 17926 96502 17978
rect 96554 17926 96566 17978
rect 96618 17926 96630 17978
rect 96682 17926 97888 17978
rect 94024 17904 97888 17926
rect 1104 17434 5980 17456
rect 1104 17382 4874 17434
rect 4926 17382 4938 17434
rect 4990 17382 5002 17434
rect 5054 17382 5066 17434
rect 5118 17382 5130 17434
rect 5182 17382 5980 17434
rect 1104 17360 5980 17382
rect 94024 17434 97888 17456
rect 94024 17382 97034 17434
rect 97086 17382 97098 17434
rect 97150 17382 97162 17434
rect 97214 17382 97226 17434
rect 97278 17382 97290 17434
rect 97342 17382 97888 17434
rect 94024 17360 97888 17382
rect 1581 17323 1639 17329
rect 1581 17289 1593 17323
rect 1627 17320 1639 17323
rect 8294 17320 8300 17332
rect 1627 17292 8300 17320
rect 1627 17289 1639 17292
rect 1581 17283 1639 17289
rect 8294 17280 8300 17292
rect 8352 17280 8358 17332
rect 1118 17144 1124 17196
rect 1176 17184 1182 17196
rect 1397 17187 1455 17193
rect 1397 17184 1409 17187
rect 1176 17156 1409 17184
rect 1176 17144 1182 17156
rect 1397 17153 1409 17156
rect 1443 17184 1455 17187
rect 1765 17187 1823 17193
rect 1765 17184 1777 17187
rect 1443 17156 1777 17184
rect 1443 17153 1455 17156
rect 1397 17147 1455 17153
rect 1765 17153 1777 17156
rect 1811 17153 1823 17187
rect 1765 17147 1823 17153
rect 97258 17144 97264 17196
rect 97316 17144 97322 17196
rect 97442 17008 97448 17060
rect 97500 17008 97506 17060
rect 1104 16890 5980 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 5980 16890
rect 1104 16816 5980 16838
rect 94024 16890 97888 16912
rect 94024 16838 96374 16890
rect 96426 16838 96438 16890
rect 96490 16838 96502 16890
rect 96554 16838 96566 16890
rect 96618 16838 96630 16890
rect 96682 16838 97888 16890
rect 94024 16816 97888 16838
rect 1104 16346 5980 16368
rect 1104 16294 4874 16346
rect 4926 16294 4938 16346
rect 4990 16294 5002 16346
rect 5054 16294 5066 16346
rect 5118 16294 5130 16346
rect 5182 16294 5980 16346
rect 1104 16272 5980 16294
rect 94024 16346 97888 16368
rect 94024 16294 97034 16346
rect 97086 16294 97098 16346
rect 97150 16294 97162 16346
rect 97214 16294 97226 16346
rect 97278 16294 97290 16346
rect 97342 16294 97888 16346
rect 94024 16272 97888 16294
rect 1581 16235 1639 16241
rect 1581 16201 1593 16235
rect 1627 16232 1639 16235
rect 8294 16232 8300 16244
rect 1627 16204 8300 16232
rect 1627 16201 1639 16204
rect 1581 16195 1639 16201
rect 8294 16192 8300 16204
rect 8352 16192 8358 16244
rect 1210 16056 1216 16108
rect 1268 16096 1274 16108
rect 1397 16099 1455 16105
rect 1397 16096 1409 16099
rect 1268 16068 1409 16096
rect 1268 16056 1274 16068
rect 1397 16065 1409 16068
rect 1443 16096 1455 16099
rect 1765 16099 1823 16105
rect 1765 16096 1777 16099
rect 1443 16068 1777 16096
rect 1443 16065 1455 16068
rect 1397 16059 1455 16065
rect 1765 16065 1777 16068
rect 1811 16065 1823 16099
rect 1765 16059 1823 16065
rect 97258 16056 97264 16108
rect 97316 16056 97322 16108
rect 97442 15852 97448 15904
rect 97500 15852 97506 15904
rect 1104 15802 5980 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 5980 15802
rect 1104 15728 5980 15750
rect 94024 15802 97888 15824
rect 94024 15750 96374 15802
rect 96426 15750 96438 15802
rect 96490 15750 96502 15802
rect 96554 15750 96566 15802
rect 96618 15750 96630 15802
rect 96682 15750 97888 15802
rect 94024 15728 97888 15750
rect 96614 15444 96620 15496
rect 96672 15484 96678 15496
rect 97261 15487 97319 15493
rect 97261 15484 97273 15487
rect 96672 15456 97273 15484
rect 96672 15444 96678 15456
rect 97261 15453 97273 15456
rect 97307 15453 97319 15487
rect 97261 15447 97319 15453
rect 1302 15376 1308 15428
rect 1360 15416 1366 15428
rect 1489 15419 1547 15425
rect 1489 15416 1501 15419
rect 1360 15388 1501 15416
rect 1360 15376 1366 15388
rect 1489 15385 1501 15388
rect 1535 15385 1547 15419
rect 1489 15379 1547 15385
rect 1504 15348 1532 15379
rect 1854 15376 1860 15428
rect 1912 15376 1918 15428
rect 1949 15351 2007 15357
rect 1949 15348 1961 15351
rect 1504 15320 1961 15348
rect 1949 15317 1961 15320
rect 1995 15317 2007 15351
rect 1949 15311 2007 15317
rect 97442 15308 97448 15360
rect 97500 15308 97506 15360
rect 1104 15258 5980 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 5980 15258
rect 1104 15184 5980 15206
rect 94024 15258 97888 15280
rect 94024 15206 97034 15258
rect 97086 15206 97098 15258
rect 97150 15206 97162 15258
rect 97214 15206 97226 15258
rect 97278 15206 97290 15258
rect 97342 15206 97888 15258
rect 94024 15184 97888 15206
rect 1104 14714 5980 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 5980 14714
rect 1104 14640 5980 14662
rect 94024 14714 97888 14736
rect 94024 14662 96374 14714
rect 96426 14662 96438 14714
rect 96490 14662 96502 14714
rect 96554 14662 96566 14714
rect 96618 14662 96630 14714
rect 96682 14662 97888 14714
rect 94024 14640 97888 14662
rect 1104 14170 5980 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 5980 14170
rect 1104 14096 5980 14118
rect 94024 14170 97888 14192
rect 94024 14118 97034 14170
rect 97086 14118 97098 14170
rect 97150 14118 97162 14170
rect 97214 14118 97226 14170
rect 97278 14118 97290 14170
rect 97342 14118 97888 14170
rect 94024 14096 97888 14118
rect 97442 14016 97448 14068
rect 97500 14016 97506 14068
rect 1302 13880 1308 13932
rect 1360 13920 1366 13932
rect 1489 13923 1547 13929
rect 1489 13920 1501 13923
rect 1360 13892 1501 13920
rect 1360 13880 1366 13892
rect 1489 13889 1501 13892
rect 1535 13889 1547 13923
rect 1489 13883 1547 13889
rect 1857 13923 1915 13929
rect 1857 13889 1869 13923
rect 1903 13920 1915 13923
rect 8294 13920 8300 13932
rect 1903 13892 8300 13920
rect 1903 13889 1915 13892
rect 1857 13883 1915 13889
rect 1504 13852 1532 13883
rect 8294 13880 8300 13892
rect 8352 13880 8358 13932
rect 97258 13880 97264 13932
rect 97316 13880 97322 13932
rect 1949 13855 2007 13861
rect 1949 13852 1961 13855
rect 1504 13824 1961 13852
rect 1949 13821 1961 13824
rect 1995 13821 2007 13855
rect 1949 13815 2007 13821
rect 1104 13626 5980 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 5980 13626
rect 1104 13552 5980 13574
rect 94024 13626 97888 13648
rect 94024 13574 96374 13626
rect 96426 13574 96438 13626
rect 96490 13574 96502 13626
rect 96554 13574 96566 13626
rect 96618 13574 96630 13626
rect 96682 13574 97888 13626
rect 94024 13552 97888 13574
rect 1581 13447 1639 13453
rect 1581 13413 1593 13447
rect 1627 13444 1639 13447
rect 8294 13444 8300 13456
rect 1627 13416 8300 13444
rect 1627 13413 1639 13416
rect 1581 13407 1639 13413
rect 8294 13404 8300 13416
rect 8352 13404 8358 13456
rect 1302 13268 1308 13320
rect 1360 13308 1366 13320
rect 1397 13311 1455 13317
rect 1397 13308 1409 13311
rect 1360 13280 1409 13308
rect 1360 13268 1366 13280
rect 1397 13277 1409 13280
rect 1443 13308 1455 13311
rect 1765 13311 1823 13317
rect 1765 13308 1777 13311
rect 1443 13280 1777 13308
rect 1443 13277 1455 13280
rect 1397 13271 1455 13277
rect 1765 13277 1777 13280
rect 1811 13277 1823 13311
rect 1765 13271 1823 13277
rect 96614 13268 96620 13320
rect 96672 13308 96678 13320
rect 97261 13311 97319 13317
rect 97261 13308 97273 13311
rect 96672 13280 97273 13308
rect 96672 13268 96678 13280
rect 97261 13277 97273 13280
rect 97307 13277 97319 13311
rect 97261 13271 97319 13277
rect 97442 13132 97448 13184
rect 97500 13132 97506 13184
rect 1104 13082 5980 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 5980 13082
rect 1104 13008 5980 13030
rect 94024 13082 97888 13104
rect 94024 13030 97034 13082
rect 97086 13030 97098 13082
rect 97150 13030 97162 13082
rect 97214 13030 97226 13082
rect 97278 13030 97290 13082
rect 97342 13030 97888 13082
rect 94024 13008 97888 13030
rect 1104 12538 5980 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 5980 12538
rect 1104 12464 5980 12486
rect 94024 12538 97888 12560
rect 94024 12486 96374 12538
rect 96426 12486 96438 12538
rect 96490 12486 96502 12538
rect 96554 12486 96566 12538
rect 96618 12486 96630 12538
rect 96682 12486 97888 12538
rect 94024 12464 97888 12486
rect 1104 11994 5980 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 5980 11994
rect 1104 11920 5980 11942
rect 94024 11994 97888 12016
rect 94024 11942 97034 11994
rect 97086 11942 97098 11994
rect 97150 11942 97162 11994
rect 97214 11942 97226 11994
rect 97278 11942 97290 11994
rect 97342 11942 97888 11994
rect 94024 11920 97888 11942
rect 1581 11883 1639 11889
rect 1581 11849 1593 11883
rect 1627 11880 1639 11883
rect 8294 11880 8300 11892
rect 1627 11852 8300 11880
rect 1627 11849 1639 11852
rect 1581 11843 1639 11849
rect 8294 11840 8300 11852
rect 8352 11840 8358 11892
rect 1118 11704 1124 11756
rect 1176 11744 1182 11756
rect 1397 11747 1455 11753
rect 1397 11744 1409 11747
rect 1176 11716 1409 11744
rect 1176 11704 1182 11716
rect 1397 11713 1409 11716
rect 1443 11744 1455 11747
rect 1765 11747 1823 11753
rect 1765 11744 1777 11747
rect 1443 11716 1777 11744
rect 1443 11713 1455 11716
rect 1397 11707 1455 11713
rect 1765 11713 1777 11716
rect 1811 11713 1823 11747
rect 1765 11707 1823 11713
rect 97258 11704 97264 11756
rect 97316 11704 97322 11756
rect 97442 11568 97448 11620
rect 97500 11568 97506 11620
rect 1104 11450 5980 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 5980 11450
rect 1104 11376 5980 11398
rect 94024 11450 97888 11472
rect 94024 11398 96374 11450
rect 96426 11398 96438 11450
rect 96490 11398 96502 11450
rect 96554 11398 96566 11450
rect 96618 11398 96630 11450
rect 96682 11398 97888 11450
rect 94024 11376 97888 11398
rect 1104 10906 5980 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 5980 10906
rect 1104 10832 5980 10854
rect 94024 10906 97888 10928
rect 94024 10854 97034 10906
rect 97086 10854 97098 10906
rect 97150 10854 97162 10906
rect 97214 10854 97226 10906
rect 97278 10854 97290 10906
rect 97342 10854 97888 10906
rect 94024 10832 97888 10854
rect 1104 10362 5980 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 5980 10362
rect 1104 10288 5980 10310
rect 94024 10362 97888 10384
rect 94024 10310 96374 10362
rect 96426 10310 96438 10362
rect 96490 10310 96502 10362
rect 96554 10310 96566 10362
rect 96618 10310 96630 10362
rect 96682 10310 97888 10362
rect 94024 10288 97888 10310
rect 1104 9818 5980 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 5980 9818
rect 1104 9744 5980 9766
rect 94024 9818 97888 9840
rect 94024 9766 97034 9818
rect 97086 9766 97098 9818
rect 97150 9766 97162 9818
rect 97214 9766 97226 9818
rect 97278 9766 97290 9818
rect 97342 9766 97888 9818
rect 94024 9744 97888 9766
rect 1104 9274 5980 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 5980 9274
rect 1104 9200 5980 9222
rect 94024 9274 97888 9296
rect 94024 9222 96374 9274
rect 96426 9222 96438 9274
rect 96490 9222 96502 9274
rect 96554 9222 96566 9274
rect 96618 9222 96630 9274
rect 96682 9222 97888 9274
rect 94024 9200 97888 9222
rect 1104 8730 5980 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 5980 8730
rect 1104 8656 5980 8678
rect 94024 8730 97888 8752
rect 94024 8678 97034 8730
rect 97086 8678 97098 8730
rect 97150 8678 97162 8730
rect 97214 8678 97226 8730
rect 97278 8678 97290 8730
rect 97342 8678 97888 8730
rect 94024 8656 97888 8678
rect 9122 8576 9128 8628
rect 9180 8616 9186 8628
rect 50338 8616 50344 8628
rect 9180 8588 50344 8616
rect 9180 8576 9186 8588
rect 50338 8576 50344 8588
rect 50396 8576 50402 8628
rect 97169 8483 97227 8489
rect 97169 8449 97181 8483
rect 97215 8480 97227 8483
rect 97534 8480 97540 8492
rect 97215 8452 97540 8480
rect 97215 8449 97227 8452
rect 97169 8443 97227 8449
rect 97534 8440 97540 8452
rect 97592 8440 97598 8492
rect 90910 8304 90916 8356
rect 90968 8344 90974 8356
rect 97353 8347 97411 8353
rect 97353 8344 97365 8347
rect 90968 8316 97365 8344
rect 90968 8304 90974 8316
rect 97353 8313 97365 8316
rect 97399 8313 97411 8347
rect 97353 8307 97411 8313
rect 8202 8236 8208 8288
rect 8260 8276 8266 8288
rect 9674 8276 9680 8288
rect 8260 8248 9680 8276
rect 8260 8236 8266 8248
rect 9674 8236 9680 8248
rect 9732 8236 9738 8288
rect 1104 8186 5980 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 5980 8186
rect 8110 8168 8116 8220
rect 8168 8208 8174 8220
rect 11146 8208 11152 8220
rect 8168 8180 11152 8208
rect 8168 8168 8174 8180
rect 11146 8168 11152 8180
rect 11204 8168 11210 8220
rect 94024 8186 97888 8208
rect 1104 8112 5980 8134
rect 8018 8100 8024 8152
rect 8076 8140 8082 8152
rect 11790 8140 11796 8152
rect 8076 8112 11796 8140
rect 8076 8100 8082 8112
rect 11790 8100 11796 8112
rect 11848 8100 11854 8152
rect 54478 8100 54484 8152
rect 54536 8140 54542 8152
rect 91922 8140 91928 8152
rect 54536 8112 91928 8140
rect 54536 8100 54542 8112
rect 91922 8100 91928 8112
rect 91980 8100 91986 8152
rect 94024 8134 96374 8186
rect 96426 8134 96438 8186
rect 96490 8134 96502 8186
rect 96554 8134 96566 8186
rect 96618 8134 96630 8186
rect 96682 8134 97888 8186
rect 94024 8112 97888 8134
rect 1104 7642 5980 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 5980 7642
rect 1104 7568 5980 7590
rect 94024 7642 97888 7664
rect 94024 7590 97034 7642
rect 97086 7590 97098 7642
rect 97150 7590 97162 7642
rect 97214 7590 97226 7642
rect 97278 7590 97290 7642
rect 97342 7590 97888 7642
rect 94024 7568 97888 7590
rect 1104 7098 5980 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 5980 7098
rect 1104 7024 5980 7046
rect 94024 7098 97888 7120
rect 94024 7046 96374 7098
rect 96426 7046 96438 7098
rect 96490 7046 96502 7098
rect 96554 7046 96566 7098
rect 96618 7046 96630 7098
rect 96682 7046 97888 7098
rect 94024 7024 97888 7046
rect 1104 6554 5980 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 5980 6554
rect 1104 6480 5980 6502
rect 94024 6554 97888 6576
rect 94024 6502 97034 6554
rect 97086 6502 97098 6554
rect 97150 6502 97162 6554
rect 97214 6502 97226 6554
rect 97278 6502 97290 6554
rect 97342 6502 97888 6554
rect 94024 6480 97888 6502
rect 1104 6010 97888 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 65654 6010
rect 65706 5958 65718 6010
rect 65770 5958 65782 6010
rect 65834 5958 65846 6010
rect 65898 5958 65910 6010
rect 65962 5958 96374 6010
rect 96426 5958 96438 6010
rect 96490 5958 96502 6010
rect 96554 5958 96566 6010
rect 96618 5958 96630 6010
rect 96682 5958 97888 6010
rect 1104 5936 97888 5958
rect 8938 5856 8944 5908
rect 8996 5856 9002 5908
rect 12158 5856 12164 5908
rect 12216 5896 12222 5908
rect 12802 5896 12808 5908
rect 12216 5868 12808 5896
rect 12216 5856 12222 5868
rect 12802 5856 12808 5868
rect 12860 5856 12866 5908
rect 50614 5856 50620 5908
rect 50672 5896 50678 5908
rect 50893 5899 50951 5905
rect 50893 5896 50905 5899
rect 50672 5868 50905 5896
rect 50672 5856 50678 5868
rect 50893 5865 50905 5868
rect 50939 5865 50951 5899
rect 50893 5859 50951 5865
rect 51074 5856 51080 5908
rect 51132 5856 51138 5908
rect 10042 5720 10048 5772
rect 10100 5760 10106 5772
rect 10962 5760 10968 5772
rect 10100 5732 10968 5760
rect 10100 5720 10106 5732
rect 10962 5720 10968 5732
rect 11020 5760 11026 5772
rect 51994 5760 52000 5772
rect 11020 5732 52000 5760
rect 11020 5720 11026 5732
rect 51994 5720 52000 5732
rect 52052 5720 52058 5772
rect 11146 5652 11152 5704
rect 11204 5692 11210 5704
rect 13170 5692 13176 5704
rect 11204 5664 13176 5692
rect 11204 5652 11210 5664
rect 13170 5652 13176 5664
rect 13228 5692 13234 5704
rect 53098 5692 53104 5704
rect 13228 5664 53104 5692
rect 13228 5652 13234 5664
rect 53098 5652 53104 5664
rect 53156 5652 53162 5704
rect 12802 5584 12808 5636
rect 12860 5624 12866 5636
rect 54110 5624 54116 5636
rect 12860 5596 54116 5624
rect 12860 5584 12866 5596
rect 54110 5584 54116 5596
rect 54168 5624 54174 5636
rect 54205 5627 54263 5633
rect 54205 5624 54217 5627
rect 54168 5596 54217 5624
rect 54168 5584 54174 5596
rect 54205 5593 54217 5596
rect 54251 5593 54263 5627
rect 54205 5587 54263 5593
rect 1104 5466 97888 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 35594 5466
rect 35646 5414 35658 5466
rect 35710 5414 35722 5466
rect 35774 5414 35786 5466
rect 35838 5414 35850 5466
rect 35902 5414 66314 5466
rect 66366 5414 66378 5466
rect 66430 5414 66442 5466
rect 66494 5414 66506 5466
rect 66558 5414 66570 5466
rect 66622 5414 97034 5466
rect 97086 5414 97098 5466
rect 97150 5414 97162 5466
rect 97214 5414 97226 5466
rect 97278 5414 97290 5466
rect 97342 5414 97888 5466
rect 1104 5392 97888 5414
rect 1104 4922 97888 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 65654 4922
rect 65706 4870 65718 4922
rect 65770 4870 65782 4922
rect 65834 4870 65846 4922
rect 65898 4870 65910 4922
rect 65962 4870 96374 4922
rect 96426 4870 96438 4922
rect 96490 4870 96502 4922
rect 96554 4870 96566 4922
rect 96618 4870 96630 4922
rect 96682 4870 97888 4922
rect 1104 4848 97888 4870
rect 1104 4378 97888 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 35594 4378
rect 35646 4326 35658 4378
rect 35710 4326 35722 4378
rect 35774 4326 35786 4378
rect 35838 4326 35850 4378
rect 35902 4326 66314 4378
rect 66366 4326 66378 4378
rect 66430 4326 66442 4378
rect 66494 4326 66506 4378
rect 66558 4326 66570 4378
rect 66622 4326 97034 4378
rect 97086 4326 97098 4378
rect 97150 4326 97162 4378
rect 97214 4326 97226 4378
rect 97278 4326 97290 4378
rect 97342 4326 97888 4378
rect 1104 4304 97888 4326
rect 1104 3834 97888 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 65654 3834
rect 65706 3782 65718 3834
rect 65770 3782 65782 3834
rect 65834 3782 65846 3834
rect 65898 3782 65910 3834
rect 65962 3782 96374 3834
rect 96426 3782 96438 3834
rect 96490 3782 96502 3834
rect 96554 3782 96566 3834
rect 96618 3782 96630 3834
rect 96682 3782 97888 3834
rect 1104 3760 97888 3782
rect 1104 3290 97888 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 35594 3290
rect 35646 3238 35658 3290
rect 35710 3238 35722 3290
rect 35774 3238 35786 3290
rect 35838 3238 35850 3290
rect 35902 3238 66314 3290
rect 66366 3238 66378 3290
rect 66430 3238 66442 3290
rect 66494 3238 66506 3290
rect 66558 3238 66570 3290
rect 66622 3238 97034 3290
rect 97086 3238 97098 3290
rect 97150 3238 97162 3290
rect 97214 3238 97226 3290
rect 97278 3238 97290 3290
rect 97342 3238 97888 3290
rect 1104 3216 97888 3238
rect 13170 3176 13176 3188
rect 12912 3148 13176 3176
rect 12912 3117 12940 3148
rect 13170 3136 13176 3148
rect 13228 3136 13234 3188
rect 12897 3111 12955 3117
rect 12897 3077 12909 3111
rect 12943 3077 12955 3111
rect 12897 3071 12955 3077
rect 11606 3000 11612 3052
rect 11664 3040 11670 3052
rect 11701 3043 11759 3049
rect 11701 3040 11713 3043
rect 11664 3012 11713 3040
rect 11664 3000 11670 3012
rect 11701 3009 11713 3012
rect 11747 3009 11759 3043
rect 11701 3003 11759 3009
rect 11606 2796 11612 2848
rect 11664 2796 11670 2848
rect 89530 2796 89536 2848
rect 89588 2796 89594 2848
rect 1104 2746 97888 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 65654 2746
rect 65706 2694 65718 2746
rect 65770 2694 65782 2746
rect 65834 2694 65846 2746
rect 65898 2694 65910 2746
rect 65962 2694 96374 2746
rect 96426 2694 96438 2746
rect 96490 2694 96502 2746
rect 96554 2694 96566 2746
rect 96618 2694 96630 2746
rect 96682 2694 97888 2746
rect 1104 2672 97888 2694
rect 10962 2632 10968 2644
rect 10888 2604 10968 2632
rect 10888 2505 10916 2604
rect 10962 2592 10968 2604
rect 11020 2632 11026 2644
rect 11609 2635 11667 2641
rect 11609 2632 11621 2635
rect 11020 2604 11621 2632
rect 11020 2592 11026 2604
rect 11609 2601 11621 2604
rect 11655 2601 11667 2635
rect 11609 2595 11667 2601
rect 32306 2592 32312 2644
rect 32364 2592 32370 2644
rect 33134 2592 33140 2644
rect 33192 2592 33198 2644
rect 34238 2592 34244 2644
rect 34296 2592 34302 2644
rect 35342 2592 35348 2644
rect 35400 2632 35406 2644
rect 35529 2635 35587 2641
rect 35529 2632 35541 2635
rect 35400 2604 35541 2632
rect 35400 2592 35406 2604
rect 35529 2601 35541 2604
rect 35575 2601 35587 2635
rect 35529 2595 35587 2601
rect 36446 2592 36452 2644
rect 36504 2632 36510 2644
rect 36817 2635 36875 2641
rect 36817 2632 36829 2635
rect 36504 2604 36829 2632
rect 36504 2592 36510 2604
rect 36817 2601 36829 2604
rect 36863 2601 36875 2635
rect 36817 2595 36875 2601
rect 37642 2592 37648 2644
rect 37700 2592 37706 2644
rect 38746 2592 38752 2644
rect 38804 2592 38810 2644
rect 40034 2592 40040 2644
rect 40092 2592 40098 2644
rect 40862 2592 40868 2644
rect 40920 2592 40926 2644
rect 41966 2592 41972 2644
rect 42024 2592 42030 2644
rect 43254 2592 43260 2644
rect 43312 2592 43318 2644
rect 48774 2592 48780 2644
rect 48832 2592 48838 2644
rect 74166 2592 74172 2644
rect 74224 2592 74230 2644
rect 75454 2592 75460 2644
rect 75512 2592 75518 2644
rect 76282 2592 76288 2644
rect 76340 2592 76346 2644
rect 77386 2592 77392 2644
rect 77444 2592 77450 2644
rect 78674 2592 78680 2644
rect 78732 2592 78738 2644
rect 79502 2592 79508 2644
rect 79560 2592 79566 2644
rect 80790 2592 80796 2644
rect 80848 2592 80854 2644
rect 81894 2592 81900 2644
rect 81952 2592 81958 2644
rect 83182 2592 83188 2644
rect 83240 2592 83246 2644
rect 84010 2592 84016 2644
rect 84068 2592 84074 2644
rect 85114 2592 85120 2644
rect 85172 2592 85178 2644
rect 44174 2524 44180 2576
rect 44232 2564 44238 2576
rect 44545 2567 44603 2573
rect 44545 2564 44557 2567
rect 44232 2536 44557 2564
rect 44232 2524 44238 2536
rect 44545 2533 44557 2536
rect 44591 2533 44603 2567
rect 44545 2527 44603 2533
rect 86402 2524 86408 2576
rect 86460 2524 86466 2576
rect 10873 2499 10931 2505
rect 10873 2465 10885 2499
rect 10919 2465 10931 2499
rect 10873 2459 10931 2465
rect 12802 2456 12808 2508
rect 12860 2496 12866 2508
rect 13817 2499 13875 2505
rect 13817 2496 13829 2499
rect 12860 2468 13829 2496
rect 12860 2456 12866 2468
rect 13817 2465 13829 2468
rect 13863 2465 13875 2499
rect 13817 2459 13875 2465
rect 45462 2456 45468 2508
rect 45520 2456 45526 2508
rect 46382 2456 46388 2508
rect 46440 2496 46446 2508
rect 46753 2499 46811 2505
rect 46753 2496 46765 2499
rect 46440 2468 46765 2496
rect 46440 2456 46446 2468
rect 46753 2465 46765 2468
rect 46799 2465 46811 2499
rect 46753 2459 46811 2465
rect 47486 2456 47492 2508
rect 47544 2496 47550 2508
rect 48041 2499 48099 2505
rect 48041 2496 48053 2499
rect 47544 2468 48053 2496
rect 47544 2456 47550 2468
rect 48041 2465 48053 2468
rect 48087 2465 48099 2499
rect 48041 2459 48099 2465
rect 87322 2456 87328 2508
rect 87380 2456 87386 2508
rect 88702 2456 88708 2508
rect 88760 2496 88766 2508
rect 89073 2499 89131 2505
rect 89073 2496 89085 2499
rect 88760 2468 89085 2496
rect 88760 2456 88766 2468
rect 89073 2465 89085 2468
rect 89119 2465 89131 2499
rect 89073 2459 89131 2465
rect 89806 2456 89812 2508
rect 89864 2496 89870 2508
rect 89993 2499 90051 2505
rect 89993 2496 90005 2499
rect 89864 2468 90005 2496
rect 89864 2456 89870 2468
rect 89993 2465 90005 2468
rect 90039 2465 90051 2499
rect 89993 2459 90051 2465
rect 10318 2388 10324 2440
rect 10376 2428 10382 2440
rect 11149 2431 11207 2437
rect 11149 2428 11161 2431
rect 10376 2400 11161 2428
rect 10376 2388 10382 2400
rect 11149 2397 11161 2400
rect 11195 2428 11207 2431
rect 11793 2431 11851 2437
rect 11793 2428 11805 2431
rect 11195 2400 11805 2428
rect 11195 2397 11207 2400
rect 11149 2391 11207 2397
rect 11793 2397 11805 2400
rect 11839 2397 11851 2431
rect 12345 2431 12403 2437
rect 12345 2428 12357 2431
rect 11793 2391 11851 2397
rect 12268 2400 12357 2428
rect 12268 2304 12296 2400
rect 12345 2397 12357 2400
rect 12391 2397 12403 2431
rect 12345 2391 12403 2397
rect 14550 2388 14556 2440
rect 14608 2388 14614 2440
rect 15562 2388 15568 2440
rect 15620 2388 15626 2440
rect 16850 2388 16856 2440
rect 16908 2388 16914 2440
rect 17770 2388 17776 2440
rect 17828 2388 17834 2440
rect 18782 2388 18788 2440
rect 18840 2388 18846 2440
rect 20070 2388 20076 2440
rect 20128 2388 20134 2440
rect 20990 2388 20996 2440
rect 21048 2428 21054 2440
rect 21361 2431 21419 2437
rect 21361 2428 21373 2431
rect 21048 2400 21373 2428
rect 21048 2388 21054 2400
rect 21361 2397 21373 2400
rect 21407 2397 21419 2431
rect 21361 2391 21419 2397
rect 22278 2388 22284 2440
rect 22336 2388 22342 2440
rect 23290 2388 23296 2440
rect 23348 2388 23354 2440
rect 24578 2388 24584 2440
rect 24636 2388 24642 2440
rect 25498 2388 25504 2440
rect 25556 2388 25562 2440
rect 26510 2388 26516 2440
rect 26568 2388 26574 2440
rect 27798 2388 27804 2440
rect 27856 2388 27862 2440
rect 29086 2388 29092 2440
rect 29144 2388 29150 2440
rect 30006 2388 30012 2440
rect 30064 2388 30070 2440
rect 31018 2388 31024 2440
rect 31076 2388 31082 2440
rect 32493 2431 32551 2437
rect 32493 2428 32505 2431
rect 32232 2400 32505 2428
rect 32232 2304 32260 2400
rect 32493 2397 32505 2400
rect 32539 2397 32551 2431
rect 32953 2431 33011 2437
rect 32953 2428 32965 2431
rect 32493 2391 32551 2397
rect 32876 2400 32965 2428
rect 32876 2304 32904 2400
rect 32953 2397 32965 2400
rect 32999 2397 33011 2431
rect 34425 2431 34483 2437
rect 34425 2428 34437 2431
rect 32953 2391 33011 2397
rect 34164 2400 34437 2428
rect 34164 2304 34192 2400
rect 34425 2397 34437 2400
rect 34471 2397 34483 2431
rect 35713 2431 35771 2437
rect 35713 2428 35725 2431
rect 34425 2391 34483 2397
rect 35452 2400 35725 2428
rect 35452 2304 35480 2400
rect 35713 2397 35725 2400
rect 35759 2397 35771 2431
rect 37001 2431 37059 2437
rect 37001 2428 37013 2431
rect 35713 2391 35771 2397
rect 36740 2400 37013 2428
rect 36740 2304 36768 2400
rect 37001 2397 37013 2400
rect 37047 2397 37059 2431
rect 37461 2431 37519 2437
rect 37461 2428 37473 2431
rect 37001 2391 37059 2397
rect 37384 2400 37473 2428
rect 37384 2304 37412 2400
rect 37461 2397 37473 2400
rect 37507 2397 37519 2431
rect 38933 2431 38991 2437
rect 38933 2428 38945 2431
rect 37461 2391 37519 2397
rect 38672 2400 38945 2428
rect 38672 2304 38700 2400
rect 38933 2397 38945 2400
rect 38979 2397 38991 2431
rect 40221 2431 40279 2437
rect 40221 2428 40233 2431
rect 38933 2391 38991 2397
rect 39960 2400 40233 2428
rect 39960 2304 39988 2400
rect 40221 2397 40233 2400
rect 40267 2397 40279 2431
rect 40681 2431 40739 2437
rect 40681 2428 40693 2431
rect 40221 2391 40279 2397
rect 40604 2400 40693 2428
rect 40604 2304 40632 2400
rect 40681 2397 40693 2400
rect 40727 2397 40739 2431
rect 42153 2431 42211 2437
rect 42153 2428 42165 2431
rect 40681 2391 40739 2397
rect 41892 2400 42165 2428
rect 41892 2304 41920 2400
rect 42153 2397 42165 2400
rect 42199 2397 42211 2431
rect 43441 2431 43499 2437
rect 43441 2428 43453 2431
rect 42153 2391 42211 2397
rect 43180 2400 43453 2428
rect 43180 2304 43208 2400
rect 43441 2397 43453 2400
rect 43487 2397 43499 2431
rect 45189 2431 45247 2437
rect 45189 2428 45201 2431
rect 43441 2391 43499 2397
rect 45112 2400 45201 2428
rect 44729 2363 44787 2369
rect 44729 2329 44741 2363
rect 44775 2329 44787 2363
rect 44729 2323 44787 2329
rect 12250 2252 12256 2304
rect 12308 2252 12314 2304
rect 14182 2252 14188 2304
rect 14240 2292 14246 2304
rect 14369 2295 14427 2301
rect 14369 2292 14381 2295
rect 14240 2264 14381 2292
rect 14240 2252 14246 2264
rect 14369 2261 14381 2264
rect 14415 2261 14427 2295
rect 14369 2255 14427 2261
rect 15470 2252 15476 2304
rect 15528 2292 15534 2304
rect 15749 2295 15807 2301
rect 15749 2292 15761 2295
rect 15528 2264 15761 2292
rect 15528 2252 15534 2264
rect 15749 2261 15761 2264
rect 15795 2261 15807 2295
rect 15749 2255 15807 2261
rect 16758 2252 16764 2304
rect 16816 2292 16822 2304
rect 17037 2295 17095 2301
rect 17037 2292 17049 2295
rect 16816 2264 17049 2292
rect 16816 2252 16822 2264
rect 17037 2261 17049 2264
rect 17083 2261 17095 2295
rect 17037 2255 17095 2261
rect 17402 2252 17408 2304
rect 17460 2292 17466 2304
rect 17589 2295 17647 2301
rect 17589 2292 17601 2295
rect 17460 2264 17601 2292
rect 17460 2252 17466 2264
rect 17589 2261 17601 2264
rect 17635 2261 17647 2295
rect 17589 2255 17647 2261
rect 18690 2252 18696 2304
rect 18748 2292 18754 2304
rect 18969 2295 19027 2301
rect 18969 2292 18981 2295
rect 18748 2264 18981 2292
rect 18748 2252 18754 2264
rect 18969 2261 18981 2264
rect 19015 2261 19027 2295
rect 18969 2255 19027 2261
rect 19978 2252 19984 2304
rect 20036 2292 20042 2304
rect 20257 2295 20315 2301
rect 20257 2292 20269 2295
rect 20036 2264 20269 2292
rect 20036 2252 20042 2264
rect 20257 2261 20269 2264
rect 20303 2261 20315 2295
rect 20257 2255 20315 2261
rect 21266 2252 21272 2304
rect 21324 2292 21330 2304
rect 21545 2295 21603 2301
rect 21545 2292 21557 2295
rect 21324 2264 21557 2292
rect 21324 2252 21330 2264
rect 21545 2261 21557 2264
rect 21591 2261 21603 2295
rect 21545 2255 21603 2261
rect 21910 2252 21916 2304
rect 21968 2292 21974 2304
rect 22097 2295 22155 2301
rect 22097 2292 22109 2295
rect 21968 2264 22109 2292
rect 21968 2252 21974 2264
rect 22097 2261 22109 2264
rect 22143 2261 22155 2295
rect 22097 2255 22155 2261
rect 23198 2252 23204 2304
rect 23256 2292 23262 2304
rect 23477 2295 23535 2301
rect 23477 2292 23489 2295
rect 23256 2264 23489 2292
rect 23256 2252 23262 2264
rect 23477 2261 23489 2264
rect 23523 2261 23535 2295
rect 23477 2255 23535 2261
rect 24486 2252 24492 2304
rect 24544 2292 24550 2304
rect 24765 2295 24823 2301
rect 24765 2292 24777 2295
rect 24544 2264 24777 2292
rect 24544 2252 24550 2264
rect 24765 2261 24777 2264
rect 24811 2261 24823 2295
rect 24765 2255 24823 2261
rect 25130 2252 25136 2304
rect 25188 2292 25194 2304
rect 25317 2295 25375 2301
rect 25317 2292 25329 2295
rect 25188 2264 25329 2292
rect 25188 2252 25194 2264
rect 25317 2261 25329 2264
rect 25363 2261 25375 2295
rect 25317 2255 25375 2261
rect 26418 2252 26424 2304
rect 26476 2292 26482 2304
rect 26697 2295 26755 2301
rect 26697 2292 26709 2295
rect 26476 2264 26709 2292
rect 26476 2252 26482 2264
rect 26697 2261 26709 2264
rect 26743 2261 26755 2295
rect 26697 2255 26755 2261
rect 27706 2252 27712 2304
rect 27764 2292 27770 2304
rect 27985 2295 28043 2301
rect 27985 2292 27997 2295
rect 27764 2264 27997 2292
rect 27764 2252 27770 2264
rect 27985 2261 27997 2264
rect 28031 2261 28043 2295
rect 27985 2255 28043 2261
rect 28994 2252 29000 2304
rect 29052 2292 29058 2304
rect 29273 2295 29331 2301
rect 29273 2292 29285 2295
rect 29052 2264 29285 2292
rect 29052 2252 29058 2264
rect 29273 2261 29285 2264
rect 29319 2261 29331 2295
rect 29273 2255 29331 2261
rect 29638 2252 29644 2304
rect 29696 2292 29702 2304
rect 29825 2295 29883 2301
rect 29825 2292 29837 2295
rect 29696 2264 29837 2292
rect 29696 2252 29702 2264
rect 29825 2261 29837 2264
rect 29871 2261 29883 2295
rect 29825 2255 29883 2261
rect 30926 2252 30932 2304
rect 30984 2292 30990 2304
rect 31205 2295 31263 2301
rect 31205 2292 31217 2295
rect 30984 2264 31217 2292
rect 30984 2252 30990 2264
rect 31205 2261 31217 2264
rect 31251 2261 31263 2295
rect 31205 2255 31263 2261
rect 32214 2252 32220 2304
rect 32272 2252 32278 2304
rect 32858 2252 32864 2304
rect 32916 2252 32922 2304
rect 34146 2252 34152 2304
rect 34204 2252 34210 2304
rect 35434 2252 35440 2304
rect 35492 2252 35498 2304
rect 36722 2252 36728 2304
rect 36780 2252 36786 2304
rect 37366 2252 37372 2304
rect 37424 2252 37430 2304
rect 38654 2252 38660 2304
rect 38712 2252 38718 2304
rect 39942 2252 39948 2304
rect 40000 2252 40006 2304
rect 40586 2252 40592 2304
rect 40644 2252 40650 2304
rect 41874 2252 41880 2304
rect 41932 2252 41938 2304
rect 43162 2252 43168 2304
rect 43220 2252 43226 2304
rect 44450 2252 44456 2304
rect 44508 2292 44514 2304
rect 44744 2292 44772 2323
rect 45112 2304 45140 2400
rect 45189 2397 45201 2400
rect 45235 2397 45247 2431
rect 46477 2431 46535 2437
rect 46477 2428 46489 2431
rect 45189 2391 45247 2397
rect 46400 2400 46489 2428
rect 46400 2304 46428 2400
rect 46477 2397 46489 2400
rect 46523 2397 46535 2431
rect 47765 2431 47823 2437
rect 47765 2428 47777 2431
rect 46477 2391 46535 2397
rect 47688 2400 47777 2428
rect 47688 2304 47716 2400
rect 47765 2397 47777 2400
rect 47811 2397 47823 2431
rect 47765 2391 47823 2397
rect 48961 2431 49019 2437
rect 48961 2397 48973 2431
rect 49007 2397 49019 2431
rect 48961 2391 49019 2397
rect 44508 2264 44772 2292
rect 44508 2252 44514 2264
rect 45094 2252 45100 2304
rect 45152 2252 45158 2304
rect 46382 2252 46388 2304
rect 46440 2252 46446 2304
rect 47670 2252 47676 2304
rect 47728 2252 47734 2304
rect 48314 2252 48320 2304
rect 48372 2292 48378 2304
rect 48976 2292 49004 2391
rect 56410 2388 56416 2440
rect 56468 2388 56474 2440
rect 57422 2388 57428 2440
rect 57480 2388 57486 2440
rect 58710 2388 58716 2440
rect 58768 2388 58774 2440
rect 59998 2388 60004 2440
rect 60056 2388 60062 2440
rect 60918 2388 60924 2440
rect 60976 2388 60982 2440
rect 61930 2388 61936 2440
rect 61988 2388 61994 2440
rect 63218 2388 63224 2440
rect 63276 2388 63282 2440
rect 64138 2388 64144 2440
rect 64196 2388 64202 2440
rect 65150 2388 65156 2440
rect 65208 2388 65214 2440
rect 66441 2431 66499 2437
rect 66441 2397 66453 2431
rect 66487 2428 66499 2431
rect 66714 2428 66720 2440
rect 66487 2400 66720 2428
rect 66487 2397 66499 2400
rect 66441 2391 66499 2397
rect 66714 2388 66720 2400
rect 66772 2388 66778 2440
rect 67726 2388 67732 2440
rect 67784 2388 67790 2440
rect 68646 2388 68652 2440
rect 68704 2388 68710 2440
rect 69658 2388 69664 2440
rect 69716 2388 69722 2440
rect 70946 2388 70952 2440
rect 71004 2388 71010 2440
rect 71866 2388 71872 2440
rect 71924 2388 71930 2440
rect 72878 2388 72884 2440
rect 72936 2388 72942 2440
rect 74353 2431 74411 2437
rect 74353 2428 74365 2431
rect 74092 2400 74365 2428
rect 74092 2304 74120 2400
rect 74353 2397 74365 2400
rect 74399 2397 74411 2431
rect 75641 2431 75699 2437
rect 75641 2428 75653 2431
rect 74353 2391 74411 2397
rect 75380 2400 75653 2428
rect 75380 2304 75408 2400
rect 75641 2397 75653 2400
rect 75687 2397 75699 2431
rect 76101 2431 76159 2437
rect 76101 2428 76113 2431
rect 75641 2391 75699 2397
rect 76024 2400 76113 2428
rect 76024 2304 76052 2400
rect 76101 2397 76113 2400
rect 76147 2397 76159 2431
rect 77573 2431 77631 2437
rect 77573 2428 77585 2431
rect 76101 2391 76159 2397
rect 77312 2400 77585 2428
rect 77312 2304 77340 2400
rect 77573 2397 77585 2400
rect 77619 2397 77631 2431
rect 78861 2431 78919 2437
rect 78861 2428 78873 2431
rect 77573 2391 77631 2397
rect 78600 2400 78873 2428
rect 78600 2304 78628 2400
rect 78861 2397 78873 2400
rect 78907 2397 78919 2431
rect 79321 2431 79379 2437
rect 79321 2428 79333 2431
rect 78861 2391 78919 2397
rect 79244 2400 79333 2428
rect 79244 2304 79272 2400
rect 79321 2397 79333 2400
rect 79367 2397 79379 2431
rect 80609 2431 80667 2437
rect 80609 2428 80621 2431
rect 79321 2391 79379 2397
rect 80532 2400 80621 2428
rect 80532 2304 80560 2400
rect 80609 2397 80621 2400
rect 80655 2397 80667 2431
rect 82081 2431 82139 2437
rect 82081 2428 82093 2431
rect 80609 2391 80667 2397
rect 81820 2400 82093 2428
rect 81820 2304 81848 2400
rect 82081 2397 82093 2400
rect 82127 2397 82139 2431
rect 83369 2431 83427 2437
rect 83369 2428 83381 2431
rect 82081 2391 82139 2397
rect 83108 2400 83381 2428
rect 83108 2304 83136 2400
rect 83369 2397 83381 2400
rect 83415 2397 83427 2431
rect 83829 2431 83887 2437
rect 83829 2428 83841 2431
rect 83369 2391 83427 2397
rect 83752 2400 83841 2428
rect 83752 2304 83780 2400
rect 83829 2397 83841 2400
rect 83875 2397 83887 2431
rect 85301 2431 85359 2437
rect 85301 2428 85313 2431
rect 83829 2391 83887 2397
rect 85040 2400 85313 2428
rect 85040 2304 85068 2400
rect 85301 2397 85313 2400
rect 85347 2397 85359 2431
rect 87049 2431 87107 2437
rect 87049 2428 87061 2431
rect 85301 2391 85359 2397
rect 86972 2400 87061 2428
rect 86589 2363 86647 2369
rect 86589 2329 86601 2363
rect 86635 2329 86647 2363
rect 86589 2323 86647 2329
rect 49053 2295 49111 2301
rect 49053 2292 49065 2295
rect 48372 2264 49065 2292
rect 48372 2252 48378 2264
rect 49053 2261 49065 2264
rect 49099 2261 49111 2295
rect 49053 2255 49111 2261
rect 56042 2252 56048 2304
rect 56100 2292 56106 2304
rect 56229 2295 56287 2301
rect 56229 2292 56241 2295
rect 56100 2264 56241 2292
rect 56100 2252 56106 2264
rect 56229 2261 56241 2264
rect 56275 2261 56287 2295
rect 56229 2255 56287 2261
rect 57330 2252 57336 2304
rect 57388 2292 57394 2304
rect 57609 2295 57667 2301
rect 57609 2292 57621 2295
rect 57388 2264 57621 2292
rect 57388 2252 57394 2264
rect 57609 2261 57621 2264
rect 57655 2261 57667 2295
rect 57609 2255 57667 2261
rect 58618 2252 58624 2304
rect 58676 2292 58682 2304
rect 58897 2295 58955 2301
rect 58897 2292 58909 2295
rect 58676 2264 58909 2292
rect 58676 2252 58682 2264
rect 58897 2261 58909 2264
rect 58943 2261 58955 2295
rect 58897 2255 58955 2261
rect 59906 2252 59912 2304
rect 59964 2292 59970 2304
rect 60185 2295 60243 2301
rect 60185 2292 60197 2295
rect 59964 2264 60197 2292
rect 59964 2252 59970 2264
rect 60185 2261 60197 2264
rect 60231 2261 60243 2295
rect 60185 2255 60243 2261
rect 60550 2252 60556 2304
rect 60608 2292 60614 2304
rect 60737 2295 60795 2301
rect 60737 2292 60749 2295
rect 60608 2264 60749 2292
rect 60608 2252 60614 2264
rect 60737 2261 60749 2264
rect 60783 2261 60795 2295
rect 60737 2255 60795 2261
rect 61838 2252 61844 2304
rect 61896 2292 61902 2304
rect 62117 2295 62175 2301
rect 62117 2292 62129 2295
rect 61896 2264 62129 2292
rect 61896 2252 61902 2264
rect 62117 2261 62129 2264
rect 62163 2261 62175 2295
rect 62117 2255 62175 2261
rect 63126 2252 63132 2304
rect 63184 2292 63190 2304
rect 63405 2295 63463 2301
rect 63405 2292 63417 2295
rect 63184 2264 63417 2292
rect 63184 2252 63190 2264
rect 63405 2261 63417 2264
rect 63451 2261 63463 2295
rect 63405 2255 63463 2261
rect 63770 2252 63776 2304
rect 63828 2292 63834 2304
rect 63957 2295 64015 2301
rect 63957 2292 63969 2295
rect 63828 2264 63969 2292
rect 63828 2252 63834 2264
rect 63957 2261 63969 2264
rect 64003 2261 64015 2295
rect 63957 2255 64015 2261
rect 65058 2252 65064 2304
rect 65116 2292 65122 2304
rect 65337 2295 65395 2301
rect 65337 2292 65349 2295
rect 65116 2264 65349 2292
rect 65116 2252 65122 2264
rect 65337 2261 65349 2264
rect 65383 2261 65395 2295
rect 65337 2255 65395 2261
rect 66625 2295 66683 2301
rect 66625 2261 66637 2295
rect 66671 2292 66683 2295
rect 66714 2292 66720 2304
rect 66671 2264 66720 2292
rect 66671 2261 66683 2264
rect 66625 2255 66683 2261
rect 66714 2252 66720 2264
rect 66772 2252 66778 2304
rect 67634 2252 67640 2304
rect 67692 2292 67698 2304
rect 67913 2295 67971 2301
rect 67913 2292 67925 2295
rect 67692 2264 67925 2292
rect 67692 2252 67698 2264
rect 67913 2261 67925 2264
rect 67959 2261 67971 2295
rect 67913 2255 67971 2261
rect 68278 2252 68284 2304
rect 68336 2292 68342 2304
rect 68465 2295 68523 2301
rect 68465 2292 68477 2295
rect 68336 2264 68477 2292
rect 68336 2252 68342 2264
rect 68465 2261 68477 2264
rect 68511 2261 68523 2295
rect 68465 2255 68523 2261
rect 69566 2252 69572 2304
rect 69624 2292 69630 2304
rect 69845 2295 69903 2301
rect 69845 2292 69857 2295
rect 69624 2264 69857 2292
rect 69624 2252 69630 2264
rect 69845 2261 69857 2264
rect 69891 2261 69903 2295
rect 69845 2255 69903 2261
rect 70854 2252 70860 2304
rect 70912 2292 70918 2304
rect 71133 2295 71191 2301
rect 71133 2292 71145 2295
rect 70912 2264 71145 2292
rect 70912 2252 70918 2264
rect 71133 2261 71145 2264
rect 71179 2261 71191 2295
rect 71133 2255 71191 2261
rect 71498 2252 71504 2304
rect 71556 2292 71562 2304
rect 71685 2295 71743 2301
rect 71685 2292 71697 2295
rect 71556 2264 71697 2292
rect 71556 2252 71562 2264
rect 71685 2261 71697 2264
rect 71731 2261 71743 2295
rect 71685 2255 71743 2261
rect 72786 2252 72792 2304
rect 72844 2292 72850 2304
rect 73065 2295 73123 2301
rect 73065 2292 73077 2295
rect 72844 2264 73077 2292
rect 72844 2252 72850 2264
rect 73065 2261 73077 2264
rect 73111 2261 73123 2295
rect 73065 2255 73123 2261
rect 74074 2252 74080 2304
rect 74132 2252 74138 2304
rect 75362 2252 75368 2304
rect 75420 2252 75426 2304
rect 76006 2252 76012 2304
rect 76064 2252 76070 2304
rect 77294 2252 77300 2304
rect 77352 2252 77358 2304
rect 78582 2252 78588 2304
rect 78640 2252 78646 2304
rect 79226 2252 79232 2304
rect 79284 2252 79290 2304
rect 80514 2252 80520 2304
rect 80572 2252 80578 2304
rect 81802 2252 81808 2304
rect 81860 2252 81866 2304
rect 83090 2252 83096 2304
rect 83148 2252 83154 2304
rect 83734 2252 83740 2304
rect 83792 2252 83798 2304
rect 85022 2252 85028 2304
rect 85080 2252 85086 2304
rect 86310 2252 86316 2304
rect 86368 2292 86374 2304
rect 86604 2292 86632 2323
rect 86972 2304 87000 2400
rect 87049 2397 87061 2400
rect 87095 2397 87107 2431
rect 88797 2431 88855 2437
rect 88797 2428 88809 2431
rect 87049 2391 87107 2397
rect 88536 2400 88809 2428
rect 86368 2264 86632 2292
rect 86368 2252 86374 2264
rect 86954 2252 86960 2304
rect 87012 2252 87018 2304
rect 88242 2252 88248 2304
rect 88300 2292 88306 2304
rect 88536 2301 88564 2400
rect 88797 2397 88809 2400
rect 88843 2397 88855 2431
rect 88797 2391 88855 2397
rect 89530 2388 89536 2440
rect 89588 2428 89594 2440
rect 89717 2431 89775 2437
rect 89717 2428 89729 2431
rect 89588 2400 89729 2428
rect 89588 2388 89594 2400
rect 89717 2397 89729 2400
rect 89763 2397 89775 2431
rect 89717 2391 89775 2397
rect 88521 2295 88579 2301
rect 88521 2292 88533 2295
rect 88300 2264 88533 2292
rect 88300 2252 88306 2264
rect 88521 2261 88533 2264
rect 88567 2261 88579 2295
rect 88521 2255 88579 2261
rect 1104 2202 97888 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 35594 2202
rect 35646 2150 35658 2202
rect 35710 2150 35722 2202
rect 35774 2150 35786 2202
rect 35838 2150 35850 2202
rect 35902 2150 66314 2202
rect 66366 2150 66378 2202
rect 66430 2150 66442 2202
rect 66494 2150 66506 2202
rect 66558 2150 66570 2202
rect 66622 2150 97034 2202
rect 97086 2150 97098 2202
rect 97150 2150 97162 2202
rect 97214 2150 97226 2202
rect 97278 2150 97290 2202
rect 97342 2150 97888 2202
rect 1104 2128 97888 2150
<< via1 >>
rect 4874 95718 4926 95770
rect 4938 95718 4990 95770
rect 5002 95718 5054 95770
rect 5066 95718 5118 95770
rect 5130 95718 5182 95770
rect 35594 95718 35646 95770
rect 35658 95718 35710 95770
rect 35722 95718 35774 95770
rect 35786 95718 35838 95770
rect 35850 95718 35902 95770
rect 66314 95718 66366 95770
rect 66378 95718 66430 95770
rect 66442 95718 66494 95770
rect 66506 95718 66558 95770
rect 66570 95718 66622 95770
rect 97034 95718 97086 95770
rect 97098 95718 97150 95770
rect 97162 95718 97214 95770
rect 97226 95718 97278 95770
rect 97290 95718 97342 95770
rect 14096 95659 14148 95668
rect 14096 95625 14105 95659
rect 14105 95625 14139 95659
rect 14139 95625 14148 95659
rect 14096 95616 14148 95625
rect 15384 95659 15436 95668
rect 15384 95625 15393 95659
rect 15393 95625 15427 95659
rect 15427 95625 15436 95659
rect 15384 95616 15436 95625
rect 16672 95659 16724 95668
rect 16672 95625 16681 95659
rect 16681 95625 16715 95659
rect 16715 95625 16724 95659
rect 16672 95616 16724 95625
rect 17316 95659 17368 95668
rect 17316 95625 17325 95659
rect 17325 95625 17359 95659
rect 17359 95625 17368 95659
rect 17316 95616 17368 95625
rect 18604 95659 18656 95668
rect 18604 95625 18613 95659
rect 18613 95625 18647 95659
rect 18647 95625 18656 95659
rect 18604 95616 18656 95625
rect 19892 95659 19944 95668
rect 19892 95625 19901 95659
rect 19901 95625 19935 95659
rect 19935 95625 19944 95659
rect 19892 95616 19944 95625
rect 21180 95659 21232 95668
rect 21180 95625 21189 95659
rect 21189 95625 21223 95659
rect 21223 95625 21232 95659
rect 21180 95616 21232 95625
rect 21824 95659 21876 95668
rect 21824 95625 21833 95659
rect 21833 95625 21867 95659
rect 21867 95625 21876 95659
rect 21824 95616 21876 95625
rect 23112 95659 23164 95668
rect 23112 95625 23121 95659
rect 23121 95625 23155 95659
rect 23155 95625 23164 95659
rect 23112 95616 23164 95625
rect 25044 95659 25096 95668
rect 25044 95625 25053 95659
rect 25053 95625 25087 95659
rect 25087 95625 25096 95659
rect 25044 95616 25096 95625
rect 26332 95659 26384 95668
rect 26332 95625 26341 95659
rect 26341 95625 26375 95659
rect 26375 95625 26384 95659
rect 26332 95616 26384 95625
rect 27620 95659 27672 95668
rect 27620 95625 27629 95659
rect 27629 95625 27663 95659
rect 27663 95625 27672 95659
rect 27620 95616 27672 95625
rect 29092 95616 29144 95668
rect 29552 95659 29604 95668
rect 29552 95625 29561 95659
rect 29561 95625 29595 95659
rect 29595 95625 29604 95659
rect 29552 95616 29604 95625
rect 30840 95659 30892 95668
rect 30840 95625 30849 95659
rect 30849 95625 30883 95659
rect 30883 95625 30892 95659
rect 30840 95616 30892 95625
rect 32496 95659 32548 95668
rect 32496 95625 32505 95659
rect 32505 95625 32539 95659
rect 32539 95625 32548 95659
rect 32496 95616 32548 95625
rect 33048 95659 33100 95668
rect 33048 95625 33057 95659
rect 33057 95625 33091 95659
rect 33091 95625 33100 95659
rect 33048 95616 33100 95625
rect 34428 95659 34480 95668
rect 34428 95625 34437 95659
rect 34437 95625 34471 95659
rect 34471 95625 34480 95659
rect 34428 95616 34480 95625
rect 35348 95616 35400 95668
rect 37004 95659 37056 95668
rect 37004 95625 37013 95659
rect 37013 95625 37047 95659
rect 37047 95625 37056 95659
rect 37004 95616 37056 95625
rect 37556 95659 37608 95668
rect 37556 95625 37565 95659
rect 37565 95625 37599 95659
rect 37599 95625 37608 95659
rect 37556 95616 37608 95625
rect 38936 95659 38988 95668
rect 38936 95625 38945 95659
rect 38945 95625 38979 95659
rect 38979 95625 38988 95659
rect 38936 95616 38988 95625
rect 39856 95616 39908 95668
rect 40776 95659 40828 95668
rect 40776 95625 40785 95659
rect 40785 95625 40819 95659
rect 40819 95625 40828 95659
rect 40776 95616 40828 95625
rect 42156 95659 42208 95668
rect 42156 95625 42165 95659
rect 42165 95625 42199 95659
rect 42199 95625 42208 95659
rect 42156 95616 42208 95625
rect 43444 95659 43496 95668
rect 43444 95625 43453 95659
rect 43453 95625 43487 95659
rect 43487 95625 43496 95659
rect 43444 95616 43496 95625
rect 44732 95659 44784 95668
rect 44732 95625 44741 95659
rect 44741 95625 44775 95659
rect 44775 95625 44784 95659
rect 44732 95616 44784 95625
rect 45284 95659 45336 95668
rect 45284 95625 45293 95659
rect 45293 95625 45327 95659
rect 45327 95625 45336 95659
rect 45284 95616 45336 95625
rect 46664 95659 46716 95668
rect 46664 95625 46673 95659
rect 46673 95625 46707 95659
rect 46707 95625 46716 95659
rect 46664 95616 46716 95625
rect 47952 95659 48004 95668
rect 47952 95625 47961 95659
rect 47961 95625 47995 95659
rect 47995 95625 48004 95659
rect 47952 95616 48004 95625
rect 48504 95659 48556 95668
rect 48504 95625 48513 95659
rect 48513 95625 48547 95659
rect 48547 95625 48556 95659
rect 48504 95616 48556 95625
rect 50988 95616 51040 95668
rect 54392 95616 54444 95668
rect 32312 95523 32364 95532
rect 32312 95489 32321 95523
rect 32321 95489 32355 95523
rect 32355 95489 32364 95523
rect 32312 95480 32364 95489
rect 33232 95523 33284 95532
rect 33232 95489 33241 95523
rect 33241 95489 33275 95523
rect 33275 95489 33284 95523
rect 33232 95480 33284 95489
rect 34244 95523 34296 95532
rect 34244 95489 34253 95523
rect 34253 95489 34287 95523
rect 34287 95489 34296 95523
rect 34244 95480 34296 95489
rect 35348 95480 35400 95532
rect 36452 95480 36504 95532
rect 37740 95523 37792 95532
rect 37740 95489 37749 95523
rect 37749 95489 37783 95523
rect 37783 95489 37792 95523
rect 37740 95480 37792 95489
rect 38752 95523 38804 95532
rect 38752 95489 38761 95523
rect 38761 95489 38795 95523
rect 38795 95489 38804 95523
rect 38752 95480 38804 95489
rect 39764 95480 39816 95532
rect 40960 95523 41012 95532
rect 40960 95489 40969 95523
rect 40969 95489 41003 95523
rect 41003 95489 41012 95523
rect 40960 95480 41012 95489
rect 41972 95523 42024 95532
rect 41972 95489 41981 95523
rect 41981 95489 42015 95523
rect 42015 95489 42024 95523
rect 41972 95480 42024 95489
rect 43260 95523 43312 95532
rect 43260 95489 43269 95523
rect 43269 95489 43303 95523
rect 43303 95489 43312 95523
rect 43260 95480 43312 95489
rect 44180 95480 44232 95532
rect 45468 95523 45520 95532
rect 45468 95489 45477 95523
rect 45477 95489 45511 95523
rect 45511 95489 45520 95523
rect 45468 95480 45520 95489
rect 46480 95523 46532 95532
rect 46480 95489 46489 95523
rect 46489 95489 46523 95523
rect 46523 95489 46532 95523
rect 46480 95480 46532 95489
rect 47768 95523 47820 95532
rect 47768 95489 47777 95523
rect 47777 95489 47811 95523
rect 47811 95489 47820 95523
rect 47768 95480 47820 95489
rect 48688 95523 48740 95532
rect 48688 95489 48697 95523
rect 48697 95489 48731 95523
rect 48731 95489 48740 95523
rect 48688 95480 48740 95489
rect 51080 95523 51132 95532
rect 51080 95489 51089 95523
rect 51089 95489 51123 95523
rect 51123 95489 51132 95523
rect 51080 95480 51132 95489
rect 51816 95480 51868 95532
rect 52920 95523 52972 95532
rect 52920 95489 52929 95523
rect 52929 95489 52963 95523
rect 52963 95489 52972 95523
rect 52920 95480 52972 95489
rect 56416 95616 56468 95668
rect 58532 95659 58584 95668
rect 58532 95625 58541 95659
rect 58541 95625 58575 95659
rect 58575 95625 58584 95659
rect 58532 95616 58584 95625
rect 59820 95659 59872 95668
rect 59820 95625 59829 95659
rect 59829 95625 59863 95659
rect 59863 95625 59872 95659
rect 59820 95616 59872 95625
rect 57704 95523 57756 95532
rect 57704 95489 57713 95523
rect 57713 95489 57747 95523
rect 57747 95489 57756 95523
rect 57704 95480 57756 95489
rect 60464 95659 60516 95668
rect 60464 95625 60473 95659
rect 60473 95625 60507 95659
rect 60507 95625 60516 95659
rect 60464 95616 60516 95625
rect 61752 95659 61804 95668
rect 61752 95625 61761 95659
rect 61761 95625 61795 95659
rect 61795 95625 61804 95659
rect 61752 95616 61804 95625
rect 63040 95659 63092 95668
rect 63040 95625 63049 95659
rect 63049 95625 63083 95659
rect 63083 95625 63092 95659
rect 63040 95616 63092 95625
rect 63684 95659 63736 95668
rect 63684 95625 63693 95659
rect 63693 95625 63727 95659
rect 63727 95625 63736 95659
rect 63684 95616 63736 95625
rect 64972 95659 65024 95668
rect 64972 95625 64981 95659
rect 64981 95625 65015 95659
rect 65015 95625 65024 95659
rect 64972 95616 65024 95625
rect 66720 95616 66772 95668
rect 67916 95659 67968 95668
rect 67916 95625 67925 95659
rect 67925 95625 67959 95659
rect 67959 95625 67968 95659
rect 67916 95616 67968 95625
rect 68560 95616 68612 95668
rect 69848 95616 69900 95668
rect 70768 95659 70820 95668
rect 70768 95625 70777 95659
rect 70777 95625 70811 95659
rect 70811 95625 70820 95659
rect 70768 95616 70820 95625
rect 71412 95659 71464 95668
rect 71412 95625 71421 95659
rect 71421 95625 71455 95659
rect 71455 95625 71464 95659
rect 71412 95616 71464 95625
rect 72700 95659 72752 95668
rect 72700 95625 72709 95659
rect 72709 95625 72743 95659
rect 72743 95625 72752 95659
rect 72700 95616 72752 95625
rect 74356 95659 74408 95668
rect 74356 95625 74365 95659
rect 74365 95625 74399 95659
rect 74399 95625 74408 95659
rect 74356 95616 74408 95625
rect 75644 95659 75696 95668
rect 75644 95625 75653 95659
rect 75653 95625 75687 95659
rect 75687 95625 75696 95659
rect 75644 95616 75696 95625
rect 76196 95659 76248 95668
rect 76196 95625 76205 95659
rect 76205 95625 76239 95659
rect 76239 95625 76248 95659
rect 76196 95616 76248 95625
rect 77576 95659 77628 95668
rect 77576 95625 77585 95659
rect 77585 95625 77619 95659
rect 77619 95625 77628 95659
rect 77576 95616 77628 95625
rect 78496 95616 78548 95668
rect 79416 95659 79468 95668
rect 79416 95625 79425 95659
rect 79425 95625 79459 95659
rect 79459 95625 79468 95659
rect 79416 95616 79468 95625
rect 80796 95659 80848 95668
rect 80796 95625 80805 95659
rect 80805 95625 80839 95659
rect 80839 95625 80848 95659
rect 80796 95616 80848 95625
rect 82084 95659 82136 95668
rect 82084 95625 82093 95659
rect 82093 95625 82127 95659
rect 82127 95625 82136 95659
rect 82084 95616 82136 95625
rect 83372 95659 83424 95668
rect 83372 95625 83381 95659
rect 83381 95625 83415 95659
rect 83415 95625 83424 95659
rect 83372 95616 83424 95625
rect 83924 95659 83976 95668
rect 83924 95625 83933 95659
rect 83933 95625 83967 95659
rect 83967 95625 83976 95659
rect 83924 95616 83976 95625
rect 85304 95659 85356 95668
rect 85304 95625 85313 95659
rect 85313 95625 85347 95659
rect 85347 95625 85356 95659
rect 85304 95616 85356 95625
rect 86592 95659 86644 95668
rect 86592 95625 86601 95659
rect 86601 95625 86635 95659
rect 86635 95625 86644 95659
rect 86592 95616 86644 95625
rect 87144 95659 87196 95668
rect 87144 95625 87153 95659
rect 87153 95625 87187 95659
rect 87187 95625 87196 95659
rect 87144 95616 87196 95625
rect 88156 95616 88208 95668
rect 89628 95616 89680 95668
rect 91008 95616 91060 95668
rect 74172 95523 74224 95532
rect 74172 95489 74181 95523
rect 74181 95489 74215 95523
rect 74215 95489 74224 95523
rect 74172 95480 74224 95489
rect 75460 95523 75512 95532
rect 75460 95489 75469 95523
rect 75469 95489 75503 95523
rect 75503 95489 75512 95523
rect 75460 95480 75512 95489
rect 76380 95523 76432 95532
rect 76380 95489 76389 95523
rect 76389 95489 76423 95523
rect 76423 95489 76432 95523
rect 76380 95480 76432 95489
rect 77392 95523 77444 95532
rect 77392 95489 77401 95523
rect 77401 95489 77435 95523
rect 77435 95489 77444 95523
rect 77392 95480 77444 95489
rect 78588 95480 78640 95532
rect 79600 95523 79652 95532
rect 79600 95489 79609 95523
rect 79609 95489 79643 95523
rect 79643 95489 79652 95523
rect 79600 95480 79652 95489
rect 80612 95523 80664 95532
rect 80612 95489 80621 95523
rect 80621 95489 80655 95523
rect 80655 95489 80664 95523
rect 80612 95480 80664 95489
rect 81900 95523 81952 95532
rect 81900 95489 81909 95523
rect 81909 95489 81943 95523
rect 81943 95489 81952 95523
rect 81900 95480 81952 95489
rect 83188 95523 83240 95532
rect 83188 95489 83197 95523
rect 83197 95489 83231 95523
rect 83231 95489 83240 95523
rect 83188 95480 83240 95489
rect 84108 95523 84160 95532
rect 84108 95489 84117 95523
rect 84117 95489 84151 95523
rect 84151 95489 84160 95523
rect 84108 95480 84160 95489
rect 85120 95523 85172 95532
rect 85120 95489 85129 95523
rect 85129 95489 85163 95523
rect 85163 95489 85172 95523
rect 85120 95480 85172 95489
rect 86408 95523 86460 95532
rect 86408 95489 86417 95523
rect 86417 95489 86451 95523
rect 86451 95489 86460 95523
rect 86408 95480 86460 95489
rect 87328 95523 87380 95532
rect 87328 95489 87337 95523
rect 87337 95489 87371 95523
rect 87371 95489 87380 95523
rect 87328 95480 87380 95489
rect 88340 95523 88392 95532
rect 88340 95489 88349 95523
rect 88349 95489 88383 95523
rect 88383 95489 88392 95523
rect 88340 95480 88392 95489
rect 89628 95523 89680 95532
rect 89628 95489 89637 95523
rect 89637 95489 89671 95523
rect 89671 95489 89680 95523
rect 89628 95480 89680 95489
rect 90916 95523 90968 95532
rect 90916 95489 90925 95523
rect 90925 95489 90959 95523
rect 90959 95489 90968 95523
rect 90916 95480 90968 95489
rect 25504 95455 25556 95464
rect 25504 95421 25513 95455
rect 25513 95421 25547 95455
rect 25547 95421 25556 95455
rect 25504 95412 25556 95421
rect 52368 95412 52420 95464
rect 54116 95455 54168 95464
rect 54116 95421 54125 95455
rect 54125 95421 54159 95455
rect 54159 95421 54168 95455
rect 54116 95412 54168 95421
rect 56784 95412 56836 95464
rect 66720 95455 66772 95464
rect 66720 95421 66729 95455
rect 66729 95421 66763 95455
rect 66763 95421 66772 95455
rect 66720 95412 66772 95421
rect 67456 95412 67508 95464
rect 18788 95387 18840 95396
rect 18788 95353 18797 95387
rect 18797 95353 18831 95387
rect 18831 95353 18840 95387
rect 18788 95344 18840 95353
rect 20076 95387 20128 95396
rect 20076 95353 20085 95387
rect 20085 95353 20119 95387
rect 20119 95353 20128 95387
rect 20076 95344 20128 95353
rect 20996 95344 21048 95396
rect 23296 95387 23348 95396
rect 23296 95353 23305 95387
rect 23305 95353 23339 95387
rect 23339 95353 23348 95387
rect 23296 95344 23348 95353
rect 28724 95344 28776 95396
rect 60004 95387 60056 95396
rect 60004 95353 60013 95387
rect 60013 95353 60047 95387
rect 60047 95353 60056 95387
rect 60004 95344 60056 95353
rect 61936 95387 61988 95396
rect 61936 95353 61945 95387
rect 61945 95353 61979 95387
rect 61979 95353 61988 95387
rect 61936 95344 61988 95353
rect 63224 95387 63276 95396
rect 63224 95353 63233 95387
rect 63233 95353 63267 95387
rect 63267 95353 63276 95387
rect 63224 95344 63276 95353
rect 14464 95319 14516 95328
rect 14464 95285 14473 95319
rect 14473 95285 14507 95319
rect 14507 95285 14516 95319
rect 14464 95276 14516 95285
rect 15752 95319 15804 95328
rect 15752 95285 15761 95319
rect 15761 95285 15795 95319
rect 15795 95285 15804 95319
rect 15752 95276 15804 95285
rect 16580 95276 16632 95328
rect 17684 95319 17736 95328
rect 17684 95285 17693 95319
rect 17693 95285 17727 95319
rect 17727 95285 17736 95319
rect 17684 95276 17736 95285
rect 22192 95319 22244 95328
rect 22192 95285 22201 95319
rect 22201 95285 22235 95319
rect 22235 95285 22244 95319
rect 22192 95276 22244 95285
rect 26516 95319 26568 95328
rect 26516 95285 26525 95319
rect 26525 95285 26559 95319
rect 26559 95285 26568 95319
rect 26516 95276 26568 95285
rect 27804 95319 27856 95328
rect 27804 95285 27813 95319
rect 27813 95285 27847 95319
rect 27847 95285 27856 95319
rect 27804 95276 27856 95285
rect 29920 95319 29972 95328
rect 29920 95285 29929 95319
rect 29929 95285 29963 95319
rect 29963 95285 29972 95319
rect 29920 95276 29972 95285
rect 31024 95319 31076 95328
rect 31024 95285 31033 95319
rect 31033 95285 31067 95319
rect 31067 95285 31076 95319
rect 31024 95276 31076 95285
rect 56508 95276 56560 95328
rect 57520 95319 57572 95328
rect 57520 95285 57529 95319
rect 57529 95285 57563 95319
rect 57563 95285 57572 95319
rect 57520 95276 57572 95285
rect 58900 95319 58952 95328
rect 58900 95285 58909 95319
rect 58909 95285 58943 95319
rect 58943 95285 58952 95319
rect 58900 95276 58952 95285
rect 60832 95319 60884 95328
rect 60832 95285 60841 95319
rect 60841 95285 60875 95319
rect 60875 95285 60884 95319
rect 60832 95276 60884 95285
rect 64052 95319 64104 95328
rect 64052 95285 64061 95319
rect 64061 95285 64095 95319
rect 64095 95285 64104 95319
rect 64052 95276 64104 95285
rect 65248 95319 65300 95328
rect 65248 95285 65257 95319
rect 65257 95285 65291 95319
rect 65291 95285 65300 95319
rect 65248 95276 65300 95285
rect 68836 95276 68888 95328
rect 69664 95319 69716 95328
rect 69664 95285 69673 95319
rect 69673 95285 69707 95319
rect 69707 95285 69716 95319
rect 69664 95276 69716 95285
rect 70952 95319 71004 95328
rect 70952 95285 70961 95319
rect 70961 95285 70995 95319
rect 70995 95285 71004 95319
rect 70952 95276 71004 95285
rect 71780 95319 71832 95328
rect 71780 95285 71789 95319
rect 71789 95285 71823 95319
rect 71823 95285 71832 95319
rect 71780 95276 71832 95285
rect 73068 95319 73120 95328
rect 73068 95285 73077 95319
rect 73077 95285 73111 95319
rect 73111 95285 73120 95319
rect 73068 95276 73120 95285
rect 4214 95174 4266 95226
rect 4278 95174 4330 95226
rect 4342 95174 4394 95226
rect 4406 95174 4458 95226
rect 4470 95174 4522 95226
rect 34934 95174 34986 95226
rect 34998 95174 35050 95226
rect 35062 95174 35114 95226
rect 35126 95174 35178 95226
rect 35190 95174 35242 95226
rect 65654 95174 65706 95226
rect 65718 95174 65770 95226
rect 65782 95174 65834 95226
rect 65846 95174 65898 95226
rect 65910 95174 65962 95226
rect 96374 95174 96426 95226
rect 96438 95174 96490 95226
rect 96502 95174 96554 95226
rect 96566 95174 96618 95226
rect 96630 95174 96682 95226
rect 24400 95115 24452 95124
rect 24400 95081 24409 95115
rect 24409 95081 24443 95115
rect 24443 95081 24452 95115
rect 24400 95072 24452 95081
rect 52920 95072 52972 95124
rect 56784 95115 56836 95124
rect 56784 95081 56793 95115
rect 56793 95081 56827 95115
rect 56827 95081 56836 95115
rect 56784 95072 56836 95081
rect 52460 94936 52512 94988
rect 52920 94979 52972 94988
rect 52920 94945 52929 94979
rect 52929 94945 52963 94979
rect 52963 94945 52972 94979
rect 52920 94936 52972 94945
rect 24308 94868 24360 94920
rect 51080 94732 51132 94784
rect 4874 94630 4926 94682
rect 4938 94630 4990 94682
rect 5002 94630 5054 94682
rect 5066 94630 5118 94682
rect 5130 94630 5182 94682
rect 35594 94630 35646 94682
rect 35658 94630 35710 94682
rect 35722 94630 35774 94682
rect 35786 94630 35838 94682
rect 35850 94630 35902 94682
rect 66314 94630 66366 94682
rect 66378 94630 66430 94682
rect 66442 94630 66494 94682
rect 66506 94630 66558 94682
rect 66570 94630 66622 94682
rect 97034 94630 97086 94682
rect 97098 94630 97150 94682
rect 97162 94630 97214 94682
rect 97226 94630 97278 94682
rect 97290 94630 97342 94682
rect 4214 94086 4266 94138
rect 4278 94086 4330 94138
rect 4342 94086 4394 94138
rect 4406 94086 4458 94138
rect 4470 94086 4522 94138
rect 34934 94086 34986 94138
rect 34998 94086 35050 94138
rect 35062 94086 35114 94138
rect 35126 94086 35178 94138
rect 35190 94086 35242 94138
rect 65654 94086 65706 94138
rect 65718 94086 65770 94138
rect 65782 94086 65834 94138
rect 65846 94086 65898 94138
rect 65910 94086 65962 94138
rect 96374 94086 96426 94138
rect 96438 94086 96490 94138
rect 96502 94086 96554 94138
rect 96566 94086 96618 94138
rect 96630 94086 96682 94138
rect 54116 93984 54168 94036
rect 52552 93780 52604 93832
rect 54116 93848 54168 93900
rect 91652 93848 91704 93900
rect 4874 93542 4926 93594
rect 4938 93542 4990 93594
rect 5002 93542 5054 93594
rect 5066 93542 5118 93594
rect 5130 93542 5182 93594
rect 35594 93542 35646 93594
rect 35658 93542 35710 93594
rect 35722 93542 35774 93594
rect 35786 93542 35838 93594
rect 35850 93542 35902 93594
rect 66314 93542 66366 93594
rect 66378 93542 66430 93594
rect 66442 93542 66494 93594
rect 66506 93542 66558 93594
rect 66570 93542 66622 93594
rect 97034 93542 97086 93594
rect 97098 93542 97150 93594
rect 97162 93542 97214 93594
rect 97226 93542 97278 93594
rect 97290 93542 97342 93594
rect 56784 93483 56836 93492
rect 31852 93304 31904 93356
rect 5540 93168 5592 93220
rect 8944 93143 8996 93152
rect 8944 93109 8953 93143
rect 8953 93109 8987 93143
rect 8987 93109 8996 93143
rect 8944 93100 8996 93109
rect 10048 93143 10100 93152
rect 10048 93109 10057 93143
rect 10057 93109 10091 93143
rect 10091 93109 10100 93143
rect 10048 93100 10100 93109
rect 11152 93143 11204 93152
rect 11152 93109 11161 93143
rect 11161 93109 11195 93143
rect 11195 93109 11204 93143
rect 11152 93100 11204 93109
rect 12256 93143 12308 93152
rect 12256 93109 12265 93143
rect 12265 93109 12299 93143
rect 12299 93109 12308 93143
rect 12256 93100 12308 93109
rect 13268 93143 13320 93152
rect 13268 93109 13277 93143
rect 13277 93109 13311 93143
rect 13311 93109 13320 93143
rect 13268 93100 13320 93109
rect 50712 93236 50764 93288
rect 52920 93304 52972 93356
rect 54208 93304 54260 93356
rect 56784 93449 56793 93483
rect 56793 93449 56827 93483
rect 56827 93449 56836 93483
rect 56784 93440 56836 93449
rect 57060 93236 57112 93288
rect 31852 93143 31904 93152
rect 31852 93109 31861 93143
rect 31861 93109 31895 93143
rect 31895 93109 31904 93143
rect 31852 93100 31904 93109
rect 49884 93100 49936 93152
rect 51080 93143 51132 93152
rect 51080 93109 51089 93143
rect 51089 93109 51123 93143
rect 51123 93109 51132 93143
rect 51080 93100 51132 93109
rect 52000 93143 52052 93152
rect 52000 93109 52009 93143
rect 52009 93109 52043 93143
rect 52043 93109 52052 93143
rect 52000 93100 52052 93109
rect 52552 93100 52604 93152
rect 54208 93143 54260 93152
rect 54208 93109 54217 93143
rect 54217 93109 54251 93143
rect 54251 93109 54260 93143
rect 54208 93100 54260 93109
rect 55128 93143 55180 93152
rect 55128 93109 55137 93143
rect 55137 93109 55171 93143
rect 55171 93109 55180 93143
rect 55128 93100 55180 93109
rect 57060 93143 57112 93152
rect 57060 93109 57069 93143
rect 57069 93109 57103 93143
rect 57103 93109 57112 93143
rect 57060 93100 57112 93109
rect 91744 93100 91796 93152
rect 4214 92998 4266 93050
rect 4278 92998 4330 93050
rect 4342 92998 4394 93050
rect 4406 92998 4458 93050
rect 4470 92998 4522 93050
rect 34934 92998 34986 93050
rect 34998 92998 35050 93050
rect 35062 92998 35114 93050
rect 35126 92998 35178 93050
rect 35190 92998 35242 93050
rect 65654 92998 65706 93050
rect 65718 92998 65770 93050
rect 65782 92998 65834 93050
rect 65846 92998 65898 93050
rect 65910 92998 65962 93050
rect 96374 92998 96426 93050
rect 96438 92998 96490 93050
rect 96502 92998 96554 93050
rect 96566 92998 96618 93050
rect 96630 92998 96682 93050
rect 57060 92896 57112 92948
rect 91836 92896 91888 92948
rect 10048 92828 10100 92880
rect 52000 92828 52052 92880
rect 12256 92760 12308 92812
rect 54208 92760 54260 92812
rect 11152 92692 11204 92744
rect 52552 92692 52604 92744
rect 4874 92454 4926 92506
rect 4938 92454 4990 92506
rect 5002 92454 5054 92506
rect 5066 92454 5118 92506
rect 5130 92454 5182 92506
rect 50528 92420 50580 92472
rect 51080 92420 51132 92472
rect 97034 92454 97086 92506
rect 97098 92454 97150 92506
rect 97162 92454 97214 92506
rect 97226 92454 97278 92506
rect 97290 92454 97342 92506
rect 4214 91910 4266 91962
rect 4278 91910 4330 91962
rect 4342 91910 4394 91962
rect 4406 91910 4458 91962
rect 4470 91910 4522 91962
rect 96374 91910 96426 91962
rect 96438 91910 96490 91962
rect 96502 91910 96554 91962
rect 96566 91910 96618 91962
rect 96630 91910 96682 91962
rect 4874 91366 4926 91418
rect 4938 91366 4990 91418
rect 5002 91366 5054 91418
rect 5066 91366 5118 91418
rect 5130 91366 5182 91418
rect 97034 91366 97086 91418
rect 97098 91366 97150 91418
rect 97162 91366 97214 91418
rect 97226 91366 97278 91418
rect 97290 91366 97342 91418
rect 4214 90822 4266 90874
rect 4278 90822 4330 90874
rect 4342 90822 4394 90874
rect 4406 90822 4458 90874
rect 4470 90822 4522 90874
rect 96374 90822 96426 90874
rect 96438 90822 96490 90874
rect 96502 90822 96554 90874
rect 96566 90822 96618 90874
rect 96630 90822 96682 90874
rect 5724 90448 5776 90500
rect 55128 90448 55180 90500
rect 4874 90278 4926 90330
rect 4938 90278 4990 90330
rect 5002 90278 5054 90330
rect 5066 90278 5118 90330
rect 5130 90278 5182 90330
rect 97034 90278 97086 90330
rect 97098 90278 97150 90330
rect 97162 90278 97214 90330
rect 97226 90278 97278 90330
rect 97290 90278 97342 90330
rect 5632 90108 5684 90160
rect 8484 90108 8536 90160
rect 4214 89734 4266 89786
rect 4278 89734 4330 89786
rect 4342 89734 4394 89786
rect 4406 89734 4458 89786
rect 4470 89734 4522 89786
rect 96374 89734 96426 89786
rect 96438 89734 96490 89786
rect 96502 89734 96554 89786
rect 96566 89734 96618 89786
rect 96630 89734 96682 89786
rect 4874 89190 4926 89242
rect 4938 89190 4990 89242
rect 5002 89190 5054 89242
rect 5066 89190 5118 89242
rect 5130 89190 5182 89242
rect 97034 89190 97086 89242
rect 97098 89190 97150 89242
rect 97162 89190 97214 89242
rect 97226 89190 97278 89242
rect 97290 89190 97342 89242
rect 4214 88646 4266 88698
rect 4278 88646 4330 88698
rect 4342 88646 4394 88698
rect 4406 88646 4458 88698
rect 4470 88646 4522 88698
rect 96374 88646 96426 88698
rect 96438 88646 96490 88698
rect 96502 88646 96554 88698
rect 96566 88646 96618 88698
rect 96630 88646 96682 88698
rect 4874 88102 4926 88154
rect 4938 88102 4990 88154
rect 5002 88102 5054 88154
rect 5066 88102 5118 88154
rect 5130 88102 5182 88154
rect 97034 88102 97086 88154
rect 97098 88102 97150 88154
rect 97162 88102 97214 88154
rect 97226 88102 97278 88154
rect 97290 88102 97342 88154
rect 4214 87558 4266 87610
rect 4278 87558 4330 87610
rect 4342 87558 4394 87610
rect 4406 87558 4458 87610
rect 4470 87558 4522 87610
rect 96374 87558 96426 87610
rect 96438 87558 96490 87610
rect 96502 87558 96554 87610
rect 96566 87558 96618 87610
rect 96630 87558 96682 87610
rect 97356 87431 97408 87440
rect 97356 87397 97365 87431
rect 97365 87397 97399 87431
rect 97399 87397 97408 87431
rect 97356 87388 97408 87397
rect 8300 87252 8352 87304
rect 97540 87295 97592 87304
rect 97540 87261 97549 87295
rect 97549 87261 97583 87295
rect 97583 87261 97592 87295
rect 97540 87252 97592 87261
rect 848 87116 900 87168
rect 4874 87014 4926 87066
rect 4938 87014 4990 87066
rect 5002 87014 5054 87066
rect 5066 87014 5118 87066
rect 5130 87014 5182 87066
rect 97034 87014 97086 87066
rect 97098 87014 97150 87066
rect 97162 87014 97214 87066
rect 97226 87014 97278 87066
rect 97290 87014 97342 87066
rect 8300 86776 8352 86828
rect 97540 86819 97592 86828
rect 97540 86785 97549 86819
rect 97549 86785 97583 86819
rect 97583 86785 97592 86819
rect 97540 86776 97592 86785
rect 848 86572 900 86624
rect 97356 86615 97408 86624
rect 97356 86581 97365 86615
rect 97365 86581 97399 86615
rect 97399 86581 97408 86615
rect 97356 86572 97408 86581
rect 4214 86470 4266 86522
rect 4278 86470 4330 86522
rect 4342 86470 4394 86522
rect 4406 86470 4458 86522
rect 4470 86470 4522 86522
rect 96374 86470 96426 86522
rect 96438 86470 96490 86522
rect 96502 86470 96554 86522
rect 96566 86470 96618 86522
rect 96630 86470 96682 86522
rect 4874 85926 4926 85978
rect 4938 85926 4990 85978
rect 5002 85926 5054 85978
rect 5066 85926 5118 85978
rect 5130 85926 5182 85978
rect 97034 85926 97086 85978
rect 97098 85926 97150 85978
rect 97162 85926 97214 85978
rect 97226 85926 97278 85978
rect 97290 85926 97342 85978
rect 4214 85382 4266 85434
rect 4278 85382 4330 85434
rect 4342 85382 4394 85434
rect 4406 85382 4458 85434
rect 4470 85382 4522 85434
rect 96374 85382 96426 85434
rect 96438 85382 96490 85434
rect 96502 85382 96554 85434
rect 96566 85382 96618 85434
rect 96630 85382 96682 85434
rect 97356 85255 97408 85264
rect 97356 85221 97365 85255
rect 97365 85221 97399 85255
rect 97399 85221 97408 85255
rect 97356 85212 97408 85221
rect 8300 85076 8352 85128
rect 97540 85119 97592 85128
rect 97540 85085 97549 85119
rect 97549 85085 97583 85119
rect 97583 85085 97592 85119
rect 97540 85076 97592 85085
rect 848 84940 900 84992
rect 4874 84838 4926 84890
rect 4938 84838 4990 84890
rect 5002 84838 5054 84890
rect 5066 84838 5118 84890
rect 5130 84838 5182 84890
rect 97034 84838 97086 84890
rect 97098 84838 97150 84890
rect 97162 84838 97214 84890
rect 97226 84838 97278 84890
rect 97290 84838 97342 84890
rect 1676 84643 1728 84652
rect 1676 84609 1685 84643
rect 1685 84609 1719 84643
rect 1719 84609 1728 84643
rect 1676 84600 1728 84609
rect 97540 84643 97592 84652
rect 97540 84609 97549 84643
rect 97549 84609 97583 84643
rect 97583 84609 97592 84643
rect 97540 84600 97592 84609
rect 848 84464 900 84516
rect 97356 84439 97408 84448
rect 97356 84405 97365 84439
rect 97365 84405 97399 84439
rect 97399 84405 97408 84439
rect 97356 84396 97408 84405
rect 4214 84294 4266 84346
rect 4278 84294 4330 84346
rect 4342 84294 4394 84346
rect 4406 84294 4458 84346
rect 4470 84294 4522 84346
rect 96374 84294 96426 84346
rect 96438 84294 96490 84346
rect 96502 84294 96554 84346
rect 96566 84294 96618 84346
rect 96630 84294 96682 84346
rect 4874 83750 4926 83802
rect 4938 83750 4990 83802
rect 5002 83750 5054 83802
rect 5066 83750 5118 83802
rect 5130 83750 5182 83802
rect 97034 83750 97086 83802
rect 97098 83750 97150 83802
rect 97162 83750 97214 83802
rect 97226 83750 97278 83802
rect 97290 83750 97342 83802
rect 8300 83512 8352 83564
rect 97540 83555 97592 83564
rect 97540 83521 97549 83555
rect 97549 83521 97583 83555
rect 97583 83521 97592 83555
rect 97540 83512 97592 83521
rect 848 83308 900 83360
rect 97356 83351 97408 83360
rect 97356 83317 97365 83351
rect 97365 83317 97399 83351
rect 97399 83317 97408 83351
rect 97356 83308 97408 83317
rect 4214 83206 4266 83258
rect 4278 83206 4330 83258
rect 4342 83206 4394 83258
rect 4406 83206 4458 83258
rect 4470 83206 4522 83258
rect 96374 83206 96426 83258
rect 96438 83206 96490 83258
rect 96502 83206 96554 83258
rect 96566 83206 96618 83258
rect 96630 83206 96682 83258
rect 4874 82662 4926 82714
rect 4938 82662 4990 82714
rect 5002 82662 5054 82714
rect 5066 82662 5118 82714
rect 5130 82662 5182 82714
rect 97034 82662 97086 82714
rect 97098 82662 97150 82714
rect 97162 82662 97214 82714
rect 97226 82662 97278 82714
rect 97290 82662 97342 82714
rect 4214 82118 4266 82170
rect 4278 82118 4330 82170
rect 4342 82118 4394 82170
rect 4406 82118 4458 82170
rect 4470 82118 4522 82170
rect 96374 82118 96426 82170
rect 96438 82118 96490 82170
rect 96502 82118 96554 82170
rect 96566 82118 96618 82170
rect 96630 82118 96682 82170
rect 97356 81991 97408 82000
rect 97356 81957 97365 81991
rect 97365 81957 97399 81991
rect 97399 81957 97408 81991
rect 97356 81948 97408 81957
rect 8300 81812 8352 81864
rect 97540 81855 97592 81864
rect 97540 81821 97549 81855
rect 97549 81821 97583 81855
rect 97583 81821 97592 81855
rect 97540 81812 97592 81821
rect 848 81676 900 81728
rect 4874 81574 4926 81626
rect 4938 81574 4990 81626
rect 5002 81574 5054 81626
rect 5066 81574 5118 81626
rect 5130 81574 5182 81626
rect 97034 81574 97086 81626
rect 97098 81574 97150 81626
rect 97162 81574 97214 81626
rect 97226 81574 97278 81626
rect 97290 81574 97342 81626
rect 8300 81336 8352 81388
rect 97540 81379 97592 81388
rect 97540 81345 97549 81379
rect 97549 81345 97583 81379
rect 97583 81345 97592 81379
rect 97540 81336 97592 81345
rect 848 81132 900 81184
rect 97356 81175 97408 81184
rect 97356 81141 97365 81175
rect 97365 81141 97399 81175
rect 97399 81141 97408 81175
rect 97356 81132 97408 81141
rect 4214 81030 4266 81082
rect 4278 81030 4330 81082
rect 4342 81030 4394 81082
rect 4406 81030 4458 81082
rect 4470 81030 4522 81082
rect 96374 81030 96426 81082
rect 96438 81030 96490 81082
rect 96502 81030 96554 81082
rect 96566 81030 96618 81082
rect 96630 81030 96682 81082
rect 4874 80486 4926 80538
rect 4938 80486 4990 80538
rect 5002 80486 5054 80538
rect 5066 80486 5118 80538
rect 5130 80486 5182 80538
rect 97034 80486 97086 80538
rect 97098 80486 97150 80538
rect 97162 80486 97214 80538
rect 97226 80486 97278 80538
rect 97290 80486 97342 80538
rect 4214 79942 4266 79994
rect 4278 79942 4330 79994
rect 4342 79942 4394 79994
rect 4406 79942 4458 79994
rect 4470 79942 4522 79994
rect 96374 79942 96426 79994
rect 96438 79942 96490 79994
rect 96502 79942 96554 79994
rect 96566 79942 96618 79994
rect 96630 79942 96682 79994
rect 97356 79815 97408 79824
rect 97356 79781 97365 79815
rect 97365 79781 97399 79815
rect 97399 79781 97408 79815
rect 97356 79772 97408 79781
rect 8300 79636 8352 79688
rect 97540 79679 97592 79688
rect 97540 79645 97549 79679
rect 97549 79645 97583 79679
rect 97583 79645 97592 79679
rect 97540 79636 97592 79645
rect 848 79500 900 79552
rect 4874 79398 4926 79450
rect 4938 79398 4990 79450
rect 5002 79398 5054 79450
rect 5066 79398 5118 79450
rect 5130 79398 5182 79450
rect 97034 79398 97086 79450
rect 97098 79398 97150 79450
rect 97162 79398 97214 79450
rect 97226 79398 97278 79450
rect 97290 79398 97342 79450
rect 8300 79160 8352 79212
rect 97448 79203 97500 79212
rect 97448 79169 97457 79203
rect 97457 79169 97491 79203
rect 97491 79169 97500 79203
rect 97448 79160 97500 79169
rect 848 79024 900 79076
rect 97264 79067 97316 79076
rect 97264 79033 97273 79067
rect 97273 79033 97307 79067
rect 97307 79033 97316 79067
rect 97264 79024 97316 79033
rect 4214 78854 4266 78906
rect 4278 78854 4330 78906
rect 4342 78854 4394 78906
rect 4406 78854 4458 78906
rect 4470 78854 4522 78906
rect 96374 78854 96426 78906
rect 96438 78854 96490 78906
rect 96502 78854 96554 78906
rect 96566 78854 96618 78906
rect 96630 78854 96682 78906
rect 4874 78310 4926 78362
rect 4938 78310 4990 78362
rect 5002 78310 5054 78362
rect 5066 78310 5118 78362
rect 5130 78310 5182 78362
rect 97034 78310 97086 78362
rect 97098 78310 97150 78362
rect 97162 78310 97214 78362
rect 97226 78310 97278 78362
rect 97290 78310 97342 78362
rect 8300 78072 8352 78124
rect 97540 78115 97592 78124
rect 97540 78081 97549 78115
rect 97549 78081 97583 78115
rect 97583 78081 97592 78115
rect 97540 78072 97592 78081
rect 848 77868 900 77920
rect 97356 77911 97408 77920
rect 97356 77877 97365 77911
rect 97365 77877 97399 77911
rect 97399 77877 97408 77911
rect 97356 77868 97408 77877
rect 4214 77766 4266 77818
rect 4278 77766 4330 77818
rect 4342 77766 4394 77818
rect 4406 77766 4458 77818
rect 4470 77766 4522 77818
rect 96374 77766 96426 77818
rect 96438 77766 96490 77818
rect 96502 77766 96554 77818
rect 96566 77766 96618 77818
rect 96630 77766 96682 77818
rect 4874 77222 4926 77274
rect 4938 77222 4990 77274
rect 5002 77222 5054 77274
rect 5066 77222 5118 77274
rect 5130 77222 5182 77274
rect 97034 77222 97086 77274
rect 97098 77222 97150 77274
rect 97162 77222 97214 77274
rect 97226 77222 97278 77274
rect 97290 77222 97342 77274
rect 4214 76678 4266 76730
rect 4278 76678 4330 76730
rect 4342 76678 4394 76730
rect 4406 76678 4458 76730
rect 4470 76678 4522 76730
rect 96374 76678 96426 76730
rect 96438 76678 96490 76730
rect 96502 76678 96554 76730
rect 96566 76678 96618 76730
rect 96630 76678 96682 76730
rect 97356 76551 97408 76560
rect 97356 76517 97365 76551
rect 97365 76517 97399 76551
rect 97399 76517 97408 76551
rect 97356 76508 97408 76517
rect 8300 76372 8352 76424
rect 97540 76415 97592 76424
rect 97540 76381 97549 76415
rect 97549 76381 97583 76415
rect 97583 76381 97592 76415
rect 97540 76372 97592 76381
rect 848 76236 900 76288
rect 4874 76134 4926 76186
rect 4938 76134 4990 76186
rect 5002 76134 5054 76186
rect 5066 76134 5118 76186
rect 5130 76134 5182 76186
rect 97034 76134 97086 76186
rect 97098 76134 97150 76186
rect 97162 76134 97214 76186
rect 97226 76134 97278 76186
rect 97290 76134 97342 76186
rect 848 76032 900 76084
rect 1676 75939 1728 75948
rect 1676 75905 1685 75939
rect 1685 75905 1719 75939
rect 1719 75905 1728 75939
rect 1676 75896 1728 75905
rect 97540 75939 97592 75948
rect 97540 75905 97549 75939
rect 97549 75905 97583 75939
rect 97583 75905 97592 75939
rect 97540 75896 97592 75905
rect 97356 75735 97408 75744
rect 97356 75701 97365 75735
rect 97365 75701 97399 75735
rect 97399 75701 97408 75735
rect 97356 75692 97408 75701
rect 4214 75590 4266 75642
rect 4278 75590 4330 75642
rect 4342 75590 4394 75642
rect 4406 75590 4458 75642
rect 4470 75590 4522 75642
rect 96374 75590 96426 75642
rect 96438 75590 96490 75642
rect 96502 75590 96554 75642
rect 96566 75590 96618 75642
rect 96630 75590 96682 75642
rect 4874 75046 4926 75098
rect 4938 75046 4990 75098
rect 5002 75046 5054 75098
rect 5066 75046 5118 75098
rect 5130 75046 5182 75098
rect 97034 75046 97086 75098
rect 97098 75046 97150 75098
rect 97162 75046 97214 75098
rect 97226 75046 97278 75098
rect 97290 75046 97342 75098
rect 4214 74502 4266 74554
rect 4278 74502 4330 74554
rect 4342 74502 4394 74554
rect 4406 74502 4458 74554
rect 4470 74502 4522 74554
rect 96374 74502 96426 74554
rect 96438 74502 96490 74554
rect 96502 74502 96554 74554
rect 96566 74502 96618 74554
rect 96630 74502 96682 74554
rect 97264 74375 97316 74384
rect 97264 74341 97273 74375
rect 97273 74341 97307 74375
rect 97307 74341 97316 74375
rect 97264 74332 97316 74341
rect 8300 74196 8352 74248
rect 97448 74171 97500 74180
rect 97448 74137 97457 74171
rect 97457 74137 97491 74171
rect 97491 74137 97500 74171
rect 97448 74128 97500 74137
rect 848 74060 900 74112
rect 4874 73958 4926 74010
rect 4938 73958 4990 74010
rect 5002 73958 5054 74010
rect 5066 73958 5118 74010
rect 5130 73958 5182 74010
rect 97034 73958 97086 74010
rect 97098 73958 97150 74010
rect 97162 73958 97214 74010
rect 97226 73958 97278 74010
rect 97290 73958 97342 74010
rect 8300 73720 8352 73772
rect 97540 73763 97592 73772
rect 97540 73729 97549 73763
rect 97549 73729 97583 73763
rect 97583 73729 97592 73763
rect 97540 73720 97592 73729
rect 848 73584 900 73636
rect 97356 73559 97408 73568
rect 97356 73525 97365 73559
rect 97365 73525 97399 73559
rect 97399 73525 97408 73559
rect 97356 73516 97408 73525
rect 4214 73414 4266 73466
rect 4278 73414 4330 73466
rect 4342 73414 4394 73466
rect 4406 73414 4458 73466
rect 4470 73414 4522 73466
rect 96374 73414 96426 73466
rect 96438 73414 96490 73466
rect 96502 73414 96554 73466
rect 96566 73414 96618 73466
rect 96630 73414 96682 73466
rect 4874 72870 4926 72922
rect 4938 72870 4990 72922
rect 5002 72870 5054 72922
rect 5066 72870 5118 72922
rect 5130 72870 5182 72922
rect 97034 72870 97086 72922
rect 97098 72870 97150 72922
rect 97162 72870 97214 72922
rect 97226 72870 97278 72922
rect 97290 72870 97342 72922
rect 8300 72632 8352 72684
rect 97264 72607 97316 72616
rect 97264 72573 97273 72607
rect 97273 72573 97307 72607
rect 97307 72573 97316 72607
rect 97264 72564 97316 72573
rect 97540 72607 97592 72616
rect 97540 72573 97549 72607
rect 97549 72573 97583 72607
rect 97583 72573 97592 72607
rect 97540 72564 97592 72573
rect 848 72428 900 72480
rect 4214 72326 4266 72378
rect 4278 72326 4330 72378
rect 4342 72326 4394 72378
rect 4406 72326 4458 72378
rect 4470 72326 4522 72378
rect 96374 72326 96426 72378
rect 96438 72326 96490 72378
rect 96502 72326 96554 72378
rect 96566 72326 96618 72378
rect 96630 72326 96682 72378
rect 97540 72199 97592 72208
rect 97540 72165 97549 72199
rect 97549 72165 97583 72199
rect 97583 72165 97592 72199
rect 97540 72156 97592 72165
rect 4874 71782 4926 71834
rect 4938 71782 4990 71834
rect 5002 71782 5054 71834
rect 5066 71782 5118 71834
rect 5130 71782 5182 71834
rect 97034 71782 97086 71834
rect 97098 71782 97150 71834
rect 97162 71782 97214 71834
rect 97226 71782 97278 71834
rect 97290 71782 97342 71834
rect 4214 71238 4266 71290
rect 4278 71238 4330 71290
rect 4342 71238 4394 71290
rect 4406 71238 4458 71290
rect 4470 71238 4522 71290
rect 96374 71238 96426 71290
rect 96438 71238 96490 71290
rect 96502 71238 96554 71290
rect 96566 71238 96618 71290
rect 96630 71238 96682 71290
rect 97356 71111 97408 71120
rect 97356 71077 97365 71111
rect 97365 71077 97399 71111
rect 97399 71077 97408 71111
rect 97356 71068 97408 71077
rect 8300 70932 8352 70984
rect 97540 70975 97592 70984
rect 97540 70941 97549 70975
rect 97549 70941 97583 70975
rect 97583 70941 97592 70975
rect 97540 70932 97592 70941
rect 848 70796 900 70848
rect 4874 70694 4926 70746
rect 4938 70694 4990 70746
rect 5002 70694 5054 70746
rect 5066 70694 5118 70746
rect 5130 70694 5182 70746
rect 97034 70694 97086 70746
rect 97098 70694 97150 70746
rect 97162 70694 97214 70746
rect 97226 70694 97278 70746
rect 97290 70694 97342 70746
rect 5540 70635 5592 70644
rect 5540 70601 5549 70635
rect 5549 70601 5583 70635
rect 5583 70601 5592 70635
rect 5540 70592 5592 70601
rect 97448 70635 97500 70644
rect 97448 70601 97457 70635
rect 97457 70601 97491 70635
rect 97491 70601 97500 70635
rect 97448 70592 97500 70601
rect 1308 70456 1360 70508
rect 97264 70499 97316 70508
rect 97264 70465 97273 70499
rect 97273 70465 97307 70499
rect 97307 70465 97316 70499
rect 97264 70456 97316 70465
rect 1584 70295 1636 70304
rect 1584 70261 1593 70295
rect 1593 70261 1627 70295
rect 1627 70261 1636 70295
rect 1584 70252 1636 70261
rect 4214 70150 4266 70202
rect 4278 70150 4330 70202
rect 4342 70150 4394 70202
rect 4406 70150 4458 70202
rect 4470 70150 4522 70202
rect 96374 70150 96426 70202
rect 96438 70150 96490 70202
rect 96502 70150 96554 70202
rect 96566 70150 96618 70202
rect 96630 70150 96682 70202
rect 5540 69844 5592 69896
rect 5632 69708 5684 69760
rect 4874 69606 4926 69658
rect 4938 69606 4990 69658
rect 5002 69606 5054 69658
rect 5066 69606 5118 69658
rect 5130 69606 5182 69658
rect 97034 69606 97086 69658
rect 97098 69606 97150 69658
rect 97162 69606 97214 69658
rect 97226 69606 97278 69658
rect 97290 69606 97342 69658
rect 5632 69547 5684 69556
rect 5632 69513 5641 69547
rect 5641 69513 5675 69547
rect 5675 69513 5684 69547
rect 5632 69504 5684 69513
rect 4214 69062 4266 69114
rect 4278 69062 4330 69114
rect 4342 69062 4394 69114
rect 4406 69062 4458 69114
rect 4470 69062 4522 69114
rect 96374 69062 96426 69114
rect 96438 69062 96490 69114
rect 96502 69062 96554 69114
rect 96566 69062 96618 69114
rect 96630 69062 96682 69114
rect 97264 68799 97316 68808
rect 97264 68765 97273 68799
rect 97273 68765 97307 68799
rect 97307 68765 97316 68799
rect 97264 68756 97316 68765
rect 1124 68688 1176 68740
rect 8300 68688 8352 68740
rect 97448 68663 97500 68672
rect 97448 68629 97457 68663
rect 97457 68629 97491 68663
rect 97491 68629 97500 68663
rect 97448 68620 97500 68629
rect 4874 68518 4926 68570
rect 4938 68518 4990 68570
rect 5002 68518 5054 68570
rect 5066 68518 5118 68570
rect 5130 68518 5182 68570
rect 97034 68518 97086 68570
rect 97098 68518 97150 68570
rect 97162 68518 97214 68570
rect 97226 68518 97278 68570
rect 97290 68518 97342 68570
rect 1308 68280 1360 68332
rect 97264 68323 97316 68332
rect 97264 68289 97273 68323
rect 97273 68289 97307 68323
rect 97307 68289 97316 68323
rect 97264 68280 97316 68289
rect 8300 68144 8352 68196
rect 97448 68119 97500 68128
rect 97448 68085 97457 68119
rect 97457 68085 97491 68119
rect 97491 68085 97500 68119
rect 97448 68076 97500 68085
rect 4214 67974 4266 68026
rect 4278 67974 4330 68026
rect 4342 67974 4394 68026
rect 4406 67974 4458 68026
rect 4470 67974 4522 68026
rect 96374 67974 96426 68026
rect 96438 67974 96490 68026
rect 96502 67974 96554 68026
rect 96566 67974 96618 68026
rect 96630 67974 96682 68026
rect 4874 67430 4926 67482
rect 4938 67430 4990 67482
rect 5002 67430 5054 67482
rect 5066 67430 5118 67482
rect 5130 67430 5182 67482
rect 97034 67430 97086 67482
rect 97098 67430 97150 67482
rect 97162 67430 97214 67482
rect 97226 67430 97278 67482
rect 97290 67430 97342 67482
rect 1308 67192 1360 67244
rect 97264 67235 97316 67244
rect 97264 67201 97273 67235
rect 97273 67201 97307 67235
rect 97307 67201 97316 67235
rect 97264 67192 97316 67201
rect 8300 67056 8352 67108
rect 97448 67031 97500 67040
rect 97448 66997 97457 67031
rect 97457 66997 97491 67031
rect 97491 66997 97500 67031
rect 97448 66988 97500 66997
rect 4214 66886 4266 66938
rect 4278 66886 4330 66938
rect 4342 66886 4394 66938
rect 4406 66886 4458 66938
rect 4470 66886 4522 66938
rect 96374 66886 96426 66938
rect 96438 66886 96490 66938
rect 96502 66886 96554 66938
rect 96566 66886 96618 66938
rect 96630 66886 96682 66938
rect 4874 66342 4926 66394
rect 4938 66342 4990 66394
rect 5002 66342 5054 66394
rect 5066 66342 5118 66394
rect 5130 66342 5182 66394
rect 97034 66342 97086 66394
rect 97098 66342 97150 66394
rect 97162 66342 97214 66394
rect 97226 66342 97278 66394
rect 97290 66342 97342 66394
rect 4214 65798 4266 65850
rect 4278 65798 4330 65850
rect 4342 65798 4394 65850
rect 4406 65798 4458 65850
rect 4470 65798 4522 65850
rect 96374 65798 96426 65850
rect 96438 65798 96490 65850
rect 96502 65798 96554 65850
rect 96566 65798 96618 65850
rect 96630 65798 96682 65850
rect 8300 65628 8352 65680
rect 97264 65535 97316 65544
rect 97264 65501 97273 65535
rect 97273 65501 97307 65535
rect 97307 65501 97316 65535
rect 97264 65492 97316 65501
rect 1124 65424 1176 65476
rect 97448 65399 97500 65408
rect 97448 65365 97457 65399
rect 97457 65365 97491 65399
rect 97491 65365 97500 65399
rect 97448 65356 97500 65365
rect 4874 65254 4926 65306
rect 4938 65254 4990 65306
rect 5002 65254 5054 65306
rect 5066 65254 5118 65306
rect 5130 65254 5182 65306
rect 97034 65254 97086 65306
rect 97098 65254 97150 65306
rect 97162 65254 97214 65306
rect 97226 65254 97278 65306
rect 97290 65254 97342 65306
rect 1308 65016 1360 65068
rect 97264 65059 97316 65068
rect 97264 65025 97273 65059
rect 97273 65025 97307 65059
rect 97307 65025 97316 65059
rect 97264 65016 97316 65025
rect 1676 64923 1728 64932
rect 1676 64889 1685 64923
rect 1685 64889 1719 64923
rect 1719 64889 1728 64923
rect 1676 64880 1728 64889
rect 97448 64923 97500 64932
rect 97448 64889 97457 64923
rect 97457 64889 97491 64923
rect 97491 64889 97500 64923
rect 97448 64880 97500 64889
rect 4214 64710 4266 64762
rect 4278 64710 4330 64762
rect 4342 64710 4394 64762
rect 4406 64710 4458 64762
rect 4470 64710 4522 64762
rect 96374 64710 96426 64762
rect 96438 64710 96490 64762
rect 96502 64710 96554 64762
rect 96566 64710 96618 64762
rect 96630 64710 96682 64762
rect 4874 64166 4926 64218
rect 4938 64166 4990 64218
rect 5002 64166 5054 64218
rect 5066 64166 5118 64218
rect 5130 64166 5182 64218
rect 97034 64166 97086 64218
rect 97098 64166 97150 64218
rect 97162 64166 97214 64218
rect 97226 64166 97278 64218
rect 97290 64166 97342 64218
rect 4214 63622 4266 63674
rect 4278 63622 4330 63674
rect 4342 63622 4394 63674
rect 4406 63622 4458 63674
rect 4470 63622 4522 63674
rect 96374 63622 96426 63674
rect 96438 63622 96490 63674
rect 96502 63622 96554 63674
rect 96566 63622 96618 63674
rect 96630 63622 96682 63674
rect 97264 63359 97316 63368
rect 97264 63325 97273 63359
rect 97273 63325 97307 63359
rect 97307 63325 97316 63359
rect 97264 63316 97316 63325
rect 1124 63248 1176 63300
rect 8300 63248 8352 63300
rect 97448 63223 97500 63232
rect 97448 63189 97457 63223
rect 97457 63189 97491 63223
rect 97491 63189 97500 63223
rect 97448 63180 97500 63189
rect 4874 63078 4926 63130
rect 4938 63078 4990 63130
rect 5002 63078 5054 63130
rect 5066 63078 5118 63130
rect 5130 63078 5182 63130
rect 97034 63078 97086 63130
rect 97098 63078 97150 63130
rect 97162 63078 97214 63130
rect 97226 63078 97278 63130
rect 97290 63078 97342 63130
rect 1308 62840 1360 62892
rect 97264 62883 97316 62892
rect 97264 62849 97273 62883
rect 97273 62849 97307 62883
rect 97307 62849 97316 62883
rect 97264 62840 97316 62849
rect 8300 62704 8352 62756
rect 97448 62679 97500 62688
rect 97448 62645 97457 62679
rect 97457 62645 97491 62679
rect 97491 62645 97500 62679
rect 97448 62636 97500 62645
rect 4214 62534 4266 62586
rect 4278 62534 4330 62586
rect 4342 62534 4394 62586
rect 4406 62534 4458 62586
rect 4470 62534 4522 62586
rect 96374 62534 96426 62586
rect 96438 62534 96490 62586
rect 96502 62534 96554 62586
rect 96566 62534 96618 62586
rect 96630 62534 96682 62586
rect 4874 61990 4926 62042
rect 4938 61990 4990 62042
rect 5002 61990 5054 62042
rect 5066 61990 5118 62042
rect 5130 61990 5182 62042
rect 97034 61990 97086 62042
rect 97098 61990 97150 62042
rect 97162 61990 97214 62042
rect 97226 61990 97278 62042
rect 97290 61990 97342 62042
rect 1308 61752 1360 61804
rect 97264 61795 97316 61804
rect 97264 61761 97273 61795
rect 97273 61761 97307 61795
rect 97307 61761 97316 61795
rect 97264 61752 97316 61761
rect 8300 61616 8352 61668
rect 97448 61591 97500 61600
rect 97448 61557 97457 61591
rect 97457 61557 97491 61591
rect 97491 61557 97500 61591
rect 97448 61548 97500 61557
rect 4214 61446 4266 61498
rect 4278 61446 4330 61498
rect 4342 61446 4394 61498
rect 4406 61446 4458 61498
rect 4470 61446 4522 61498
rect 96374 61446 96426 61498
rect 96438 61446 96490 61498
rect 96502 61446 96554 61498
rect 96566 61446 96618 61498
rect 96630 61446 96682 61498
rect 4874 60902 4926 60954
rect 4938 60902 4990 60954
rect 5002 60902 5054 60954
rect 5066 60902 5118 60954
rect 5130 60902 5182 60954
rect 97034 60902 97086 60954
rect 97098 60902 97150 60954
rect 97162 60902 97214 60954
rect 97226 60902 97278 60954
rect 97290 60902 97342 60954
rect 4214 60358 4266 60410
rect 4278 60358 4330 60410
rect 4342 60358 4394 60410
rect 4406 60358 4458 60410
rect 4470 60358 4522 60410
rect 96374 60358 96426 60410
rect 96438 60358 96490 60410
rect 96502 60358 96554 60410
rect 96566 60358 96618 60410
rect 96630 60358 96682 60410
rect 8300 60256 8352 60308
rect 97264 60095 97316 60104
rect 97264 60061 97273 60095
rect 97273 60061 97307 60095
rect 97307 60061 97316 60095
rect 97264 60052 97316 60061
rect 1216 59984 1268 60036
rect 50436 59984 50488 60036
rect 50620 59984 50672 60036
rect 97448 59959 97500 59968
rect 97448 59925 97457 59959
rect 97457 59925 97491 59959
rect 97491 59925 97500 59959
rect 97448 59916 97500 59925
rect 4874 59814 4926 59866
rect 4938 59814 4990 59866
rect 5002 59814 5054 59866
rect 5066 59814 5118 59866
rect 5130 59814 5182 59866
rect 97034 59814 97086 59866
rect 97098 59814 97150 59866
rect 97162 59814 97214 59866
rect 97226 59814 97278 59866
rect 97290 59814 97342 59866
rect 1216 59576 1268 59628
rect 97264 59619 97316 59628
rect 97264 59585 97273 59619
rect 97273 59585 97307 59619
rect 97307 59585 97316 59619
rect 97264 59576 97316 59585
rect 1584 59415 1636 59424
rect 1584 59381 1593 59415
rect 1593 59381 1627 59415
rect 1627 59381 1636 59415
rect 1584 59372 1636 59381
rect 97448 59415 97500 59424
rect 97448 59381 97457 59415
rect 97457 59381 97491 59415
rect 97491 59381 97500 59415
rect 97448 59372 97500 59381
rect 4214 59270 4266 59322
rect 4278 59270 4330 59322
rect 4342 59270 4394 59322
rect 4406 59270 4458 59322
rect 4470 59270 4522 59322
rect 96374 59270 96426 59322
rect 96438 59270 96490 59322
rect 96502 59270 96554 59322
rect 96566 59270 96618 59322
rect 96630 59270 96682 59322
rect 4874 58726 4926 58778
rect 4938 58726 4990 58778
rect 5002 58726 5054 58778
rect 5066 58726 5118 58778
rect 5130 58726 5182 58778
rect 97034 58726 97086 58778
rect 97098 58726 97150 58778
rect 97162 58726 97214 58778
rect 97226 58726 97278 58778
rect 97290 58726 97342 58778
rect 4214 58182 4266 58234
rect 4278 58182 4330 58234
rect 4342 58182 4394 58234
rect 4406 58182 4458 58234
rect 4470 58182 4522 58234
rect 96374 58182 96426 58234
rect 96438 58182 96490 58234
rect 96502 58182 96554 58234
rect 96566 58182 96618 58234
rect 96630 58182 96682 58234
rect 1308 57876 1360 57928
rect 97264 57919 97316 57928
rect 97264 57885 97273 57919
rect 97273 57885 97307 57919
rect 97307 57885 97316 57919
rect 97264 57876 97316 57885
rect 1584 57783 1636 57792
rect 1584 57749 1593 57783
rect 1593 57749 1627 57783
rect 1627 57749 1636 57783
rect 1584 57740 1636 57749
rect 97448 57783 97500 57792
rect 97448 57749 97457 57783
rect 97457 57749 97491 57783
rect 97491 57749 97500 57783
rect 97448 57740 97500 57749
rect 4874 57638 4926 57690
rect 4938 57638 4990 57690
rect 5002 57638 5054 57690
rect 5066 57638 5118 57690
rect 5130 57638 5182 57690
rect 97034 57638 97086 57690
rect 97098 57638 97150 57690
rect 97162 57638 97214 57690
rect 97226 57638 97278 57690
rect 97290 57638 97342 57690
rect 1308 57400 1360 57452
rect 97264 57443 97316 57452
rect 97264 57409 97273 57443
rect 97273 57409 97307 57443
rect 97307 57409 97316 57443
rect 97264 57400 97316 57409
rect 8300 57264 8352 57316
rect 97448 57239 97500 57248
rect 97448 57205 97457 57239
rect 97457 57205 97491 57239
rect 97491 57205 97500 57239
rect 97448 57196 97500 57205
rect 4214 57094 4266 57146
rect 4278 57094 4330 57146
rect 4342 57094 4394 57146
rect 4406 57094 4458 57146
rect 4470 57094 4522 57146
rect 96374 57094 96426 57146
rect 96438 57094 96490 57146
rect 96502 57094 96554 57146
rect 96566 57094 96618 57146
rect 96630 57094 96682 57146
rect 4874 56550 4926 56602
rect 4938 56550 4990 56602
rect 5002 56550 5054 56602
rect 5066 56550 5118 56602
rect 5130 56550 5182 56602
rect 97034 56550 97086 56602
rect 97098 56550 97150 56602
rect 97162 56550 97214 56602
rect 97226 56550 97278 56602
rect 97290 56550 97342 56602
rect 1308 56312 1360 56364
rect 97264 56355 97316 56364
rect 97264 56321 97273 56355
rect 97273 56321 97307 56355
rect 97307 56321 97316 56355
rect 97264 56312 97316 56321
rect 8300 56176 8352 56228
rect 97448 56151 97500 56160
rect 97448 56117 97457 56151
rect 97457 56117 97491 56151
rect 97491 56117 97500 56151
rect 97448 56108 97500 56117
rect 4214 56006 4266 56058
rect 4278 56006 4330 56058
rect 4342 56006 4394 56058
rect 4406 56006 4458 56058
rect 4470 56006 4522 56058
rect 96374 56006 96426 56058
rect 96438 56006 96490 56058
rect 96502 56006 96554 56058
rect 96566 56006 96618 56058
rect 96630 56006 96682 56058
rect 4874 55462 4926 55514
rect 4938 55462 4990 55514
rect 5002 55462 5054 55514
rect 5066 55462 5118 55514
rect 5130 55462 5182 55514
rect 97034 55462 97086 55514
rect 97098 55462 97150 55514
rect 97162 55462 97214 55514
rect 97226 55462 97278 55514
rect 97290 55462 97342 55514
rect 4214 54918 4266 54970
rect 4278 54918 4330 54970
rect 4342 54918 4394 54970
rect 4406 54918 4458 54970
rect 4470 54918 4522 54970
rect 96374 54918 96426 54970
rect 96438 54918 96490 54970
rect 96502 54918 96554 54970
rect 96566 54918 96618 54970
rect 96630 54918 96682 54970
rect 8300 54816 8352 54868
rect 1308 54612 1360 54664
rect 97264 54655 97316 54664
rect 97264 54621 97273 54655
rect 97273 54621 97307 54655
rect 97307 54621 97316 54655
rect 97264 54612 97316 54621
rect 97448 54519 97500 54528
rect 97448 54485 97457 54519
rect 97457 54485 97491 54519
rect 97491 54485 97500 54519
rect 97448 54476 97500 54485
rect 4874 54374 4926 54426
rect 4938 54374 4990 54426
rect 5002 54374 5054 54426
rect 5066 54374 5118 54426
rect 5130 54374 5182 54426
rect 97034 54374 97086 54426
rect 97098 54374 97150 54426
rect 97162 54374 97214 54426
rect 97226 54374 97278 54426
rect 97290 54374 97342 54426
rect 1216 54136 1268 54188
rect 97264 54179 97316 54188
rect 97264 54145 97273 54179
rect 97273 54145 97307 54179
rect 97307 54145 97316 54179
rect 97264 54136 97316 54145
rect 1584 53975 1636 53984
rect 1584 53941 1593 53975
rect 1593 53941 1627 53975
rect 1627 53941 1636 53975
rect 1584 53932 1636 53941
rect 97448 53975 97500 53984
rect 97448 53941 97457 53975
rect 97457 53941 97491 53975
rect 97491 53941 97500 53975
rect 97448 53932 97500 53941
rect 4214 53830 4266 53882
rect 4278 53830 4330 53882
rect 4342 53830 4394 53882
rect 4406 53830 4458 53882
rect 4470 53830 4522 53882
rect 96374 53830 96426 53882
rect 96438 53830 96490 53882
rect 96502 53830 96554 53882
rect 96566 53830 96618 53882
rect 96630 53830 96682 53882
rect 4874 53286 4926 53338
rect 4938 53286 4990 53338
rect 5002 53286 5054 53338
rect 5066 53286 5118 53338
rect 5130 53286 5182 53338
rect 97034 53286 97086 53338
rect 97098 53286 97150 53338
rect 97162 53286 97214 53338
rect 97226 53286 97278 53338
rect 97290 53286 97342 53338
rect 4214 52742 4266 52794
rect 4278 52742 4330 52794
rect 4342 52742 4394 52794
rect 4406 52742 4458 52794
rect 4470 52742 4522 52794
rect 96374 52742 96426 52794
rect 96438 52742 96490 52794
rect 96502 52742 96554 52794
rect 96566 52742 96618 52794
rect 96630 52742 96682 52794
rect 4874 52198 4926 52250
rect 4938 52198 4990 52250
rect 5002 52198 5054 52250
rect 5066 52198 5118 52250
rect 5130 52198 5182 52250
rect 97034 52198 97086 52250
rect 97098 52198 97150 52250
rect 97162 52198 97214 52250
rect 97226 52198 97278 52250
rect 97290 52198 97342 52250
rect 4214 51654 4266 51706
rect 4278 51654 4330 51706
rect 4342 51654 4394 51706
rect 4406 51654 4458 51706
rect 4470 51654 4522 51706
rect 96374 51654 96426 51706
rect 96438 51654 96490 51706
rect 96502 51654 96554 51706
rect 96566 51654 96618 51706
rect 96630 51654 96682 51706
rect 4874 51110 4926 51162
rect 4938 51110 4990 51162
rect 5002 51110 5054 51162
rect 5066 51110 5118 51162
rect 5130 51110 5182 51162
rect 97034 51110 97086 51162
rect 97098 51110 97150 51162
rect 97162 51110 97214 51162
rect 97226 51110 97278 51162
rect 97290 51110 97342 51162
rect 5724 51008 5776 51060
rect 8484 51008 8536 51060
rect 7472 50804 7524 50856
rect 92112 50804 92164 50856
rect 4214 50566 4266 50618
rect 4278 50566 4330 50618
rect 4342 50566 4394 50618
rect 4406 50566 4458 50618
rect 4470 50566 4522 50618
rect 8208 50600 8260 50652
rect 9864 50600 9916 50652
rect 10232 50192 10284 50244
rect 8024 50124 8076 50176
rect 11796 50124 11848 50176
rect 53380 50192 53432 50244
rect 52276 50124 52328 50176
rect 96374 50566 96426 50618
rect 96438 50566 96490 50618
rect 96502 50566 96554 50618
rect 96566 50566 96618 50618
rect 96630 50566 96682 50618
rect 4874 50022 4926 50074
rect 4938 50022 4990 50074
rect 5002 50022 5054 50074
rect 5066 50022 5118 50074
rect 5130 50022 5182 50074
rect 7472 50056 7524 50108
rect 8116 50056 8168 50108
rect 11152 50056 11204 50108
rect 52920 50056 52972 50108
rect 54484 49988 54536 50040
rect 91928 49988 91980 50040
rect 92112 49988 92164 50040
rect 97034 50022 97086 50074
rect 97098 50022 97150 50074
rect 97162 50022 97214 50074
rect 97226 50022 97278 50074
rect 97290 50022 97342 50074
rect 4214 49478 4266 49530
rect 4278 49478 4330 49530
rect 4342 49478 4394 49530
rect 4406 49478 4458 49530
rect 4470 49478 4522 49530
rect 96374 49478 96426 49530
rect 96438 49478 96490 49530
rect 96502 49478 96554 49530
rect 96566 49478 96618 49530
rect 96630 49478 96682 49530
rect 4874 48934 4926 48986
rect 4938 48934 4990 48986
rect 5002 48934 5054 48986
rect 5066 48934 5118 48986
rect 5130 48934 5182 48986
rect 97034 48934 97086 48986
rect 97098 48934 97150 48986
rect 97162 48934 97214 48986
rect 97226 48934 97278 48986
rect 97290 48934 97342 48986
rect 5540 48875 5592 48884
rect 5540 48841 5549 48875
rect 5549 48841 5583 48875
rect 5583 48841 5592 48875
rect 5540 48832 5592 48841
rect 8484 48832 8536 48884
rect 12900 48764 12952 48816
rect 52276 48764 52328 48816
rect 91744 48764 91796 48816
rect 1216 48696 1268 48748
rect 5632 48696 5684 48748
rect 11152 48696 11204 48748
rect 55588 48696 55640 48748
rect 10232 48628 10284 48680
rect 51816 48628 51868 48680
rect 54484 48628 54536 48680
rect 91836 48628 91888 48680
rect 11888 48560 11940 48612
rect 54024 48560 54076 48612
rect 50344 48492 50396 48544
rect 55404 48492 55456 48544
rect 4214 48390 4266 48442
rect 4278 48390 4330 48442
rect 4342 48390 4394 48442
rect 4406 48390 4458 48442
rect 4470 48390 4522 48442
rect 11336 48424 11388 48476
rect 53380 48424 53432 48476
rect 91652 48492 91704 48544
rect 96374 48390 96426 48442
rect 96438 48390 96490 48442
rect 96502 48390 96554 48442
rect 96566 48390 96618 48442
rect 96630 48390 96682 48442
rect 5632 48263 5684 48272
rect 5632 48229 5641 48263
rect 5641 48229 5675 48263
rect 5675 48229 5684 48263
rect 5632 48220 5684 48229
rect 4874 47846 4926 47898
rect 4938 47846 4990 47898
rect 5002 47846 5054 47898
rect 5066 47846 5118 47898
rect 5130 47846 5182 47898
rect 97034 47846 97086 47898
rect 97098 47846 97150 47898
rect 97162 47846 97214 47898
rect 97226 47846 97278 47898
rect 97290 47846 97342 47898
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 96374 47302 96426 47354
rect 96438 47302 96490 47354
rect 96502 47302 96554 47354
rect 96566 47302 96618 47354
rect 96630 47302 96682 47354
rect 4874 46758 4926 46810
rect 4938 46758 4990 46810
rect 5002 46758 5054 46810
rect 5066 46758 5118 46810
rect 5130 46758 5182 46810
rect 97034 46758 97086 46810
rect 97098 46758 97150 46810
rect 97162 46758 97214 46810
rect 97226 46758 97278 46810
rect 97290 46758 97342 46810
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 96374 46214 96426 46266
rect 96438 46214 96490 46266
rect 96502 46214 96554 46266
rect 96566 46214 96618 46266
rect 96630 46214 96682 46266
rect 1676 45951 1728 45960
rect 1676 45917 1685 45951
rect 1685 45917 1719 45951
rect 1719 45917 1728 45951
rect 1676 45908 1728 45917
rect 97540 45951 97592 45960
rect 97540 45917 97549 45951
rect 97549 45917 97583 45951
rect 97583 45917 97592 45951
rect 97540 45908 97592 45917
rect 848 45772 900 45824
rect 97448 45772 97500 45824
rect 4874 45670 4926 45722
rect 4938 45670 4990 45722
rect 5002 45670 5054 45722
rect 5066 45670 5118 45722
rect 5130 45670 5182 45722
rect 97034 45670 97086 45722
rect 97098 45670 97150 45722
rect 97162 45670 97214 45722
rect 97226 45670 97278 45722
rect 97290 45670 97342 45722
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 96374 45126 96426 45178
rect 96438 45126 96490 45178
rect 96502 45126 96554 45178
rect 96566 45126 96618 45178
rect 96630 45126 96682 45178
rect 4874 44582 4926 44634
rect 4938 44582 4990 44634
rect 5002 44582 5054 44634
rect 5066 44582 5118 44634
rect 5130 44582 5182 44634
rect 97034 44582 97086 44634
rect 97098 44582 97150 44634
rect 97162 44582 97214 44634
rect 97226 44582 97278 44634
rect 97290 44582 97342 44634
rect 848 44480 900 44532
rect 8300 44344 8352 44396
rect 97540 44387 97592 44396
rect 97540 44353 97549 44387
rect 97549 44353 97583 44387
rect 97583 44353 97592 44387
rect 97540 44344 97592 44353
rect 97356 44251 97408 44260
rect 97356 44217 97365 44251
rect 97365 44217 97399 44251
rect 97399 44217 97408 44251
rect 97356 44208 97408 44217
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 96374 44038 96426 44090
rect 96438 44038 96490 44090
rect 96502 44038 96554 44090
rect 96566 44038 96618 44090
rect 96630 44038 96682 44090
rect 4874 43494 4926 43546
rect 4938 43494 4990 43546
rect 5002 43494 5054 43546
rect 5066 43494 5118 43546
rect 5130 43494 5182 43546
rect 97034 43494 97086 43546
rect 97098 43494 97150 43546
rect 97162 43494 97214 43546
rect 97226 43494 97278 43546
rect 97290 43494 97342 43546
rect 8300 43256 8352 43308
rect 97540 43299 97592 43308
rect 97540 43265 97549 43299
rect 97549 43265 97583 43299
rect 97583 43265 97592 43299
rect 97540 43256 97592 43265
rect 97356 43163 97408 43172
rect 97356 43129 97365 43163
rect 97365 43129 97399 43163
rect 97399 43129 97408 43163
rect 97356 43120 97408 43129
rect 848 43052 900 43104
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 96374 42950 96426 43002
rect 96438 42950 96490 43002
rect 96502 42950 96554 43002
rect 96566 42950 96618 43002
rect 96630 42950 96682 43002
rect 8300 42644 8352 42696
rect 97540 42687 97592 42696
rect 97540 42653 97549 42687
rect 97549 42653 97583 42687
rect 97583 42653 97592 42687
rect 97540 42644 97592 42653
rect 848 42508 900 42560
rect 97448 42508 97500 42560
rect 4874 42406 4926 42458
rect 4938 42406 4990 42458
rect 5002 42406 5054 42458
rect 5066 42406 5118 42458
rect 5130 42406 5182 42458
rect 97034 42406 97086 42458
rect 97098 42406 97150 42458
rect 97162 42406 97214 42458
rect 97226 42406 97278 42458
rect 97290 42406 97342 42458
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 96374 41862 96426 41914
rect 96438 41862 96490 41914
rect 96502 41862 96554 41914
rect 96566 41862 96618 41914
rect 96630 41862 96682 41914
rect 4874 41318 4926 41370
rect 4938 41318 4990 41370
rect 5002 41318 5054 41370
rect 5066 41318 5118 41370
rect 5130 41318 5182 41370
rect 97034 41318 97086 41370
rect 97098 41318 97150 41370
rect 97162 41318 97214 41370
rect 97226 41318 97278 41370
rect 97290 41318 97342 41370
rect 97356 41259 97408 41268
rect 97356 41225 97365 41259
rect 97365 41225 97399 41259
rect 97399 41225 97408 41259
rect 97356 41216 97408 41225
rect 8300 41080 8352 41132
rect 97540 41123 97592 41132
rect 97540 41089 97549 41123
rect 97549 41089 97583 41123
rect 97583 41089 97592 41123
rect 97540 41080 97592 41089
rect 848 40944 900 40996
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 96374 40774 96426 40826
rect 96438 40774 96490 40826
rect 96502 40774 96554 40826
rect 96566 40774 96618 40826
rect 96630 40774 96682 40826
rect 1676 40511 1728 40520
rect 1676 40477 1685 40511
rect 1685 40477 1719 40511
rect 1719 40477 1728 40511
rect 1676 40468 1728 40477
rect 97540 40511 97592 40520
rect 97540 40477 97549 40511
rect 97549 40477 97583 40511
rect 97583 40477 97592 40511
rect 97540 40468 97592 40477
rect 848 40332 900 40384
rect 97448 40332 97500 40384
rect 4874 40230 4926 40282
rect 4938 40230 4990 40282
rect 5002 40230 5054 40282
rect 5066 40230 5118 40282
rect 5130 40230 5182 40282
rect 97034 40230 97086 40282
rect 97098 40230 97150 40282
rect 97162 40230 97214 40282
rect 97226 40230 97278 40282
rect 97290 40230 97342 40282
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 96374 39686 96426 39738
rect 96438 39686 96490 39738
rect 96502 39686 96554 39738
rect 96566 39686 96618 39738
rect 96630 39686 96682 39738
rect 4874 39142 4926 39194
rect 4938 39142 4990 39194
rect 5002 39142 5054 39194
rect 5066 39142 5118 39194
rect 5130 39142 5182 39194
rect 97034 39142 97086 39194
rect 97098 39142 97150 39194
rect 97162 39142 97214 39194
rect 97226 39142 97278 39194
rect 97290 39142 97342 39194
rect 97356 39083 97408 39092
rect 97356 39049 97365 39083
rect 97365 39049 97399 39083
rect 97399 39049 97408 39083
rect 97356 39040 97408 39049
rect 8300 38904 8352 38956
rect 97540 38947 97592 38956
rect 97540 38913 97549 38947
rect 97549 38913 97583 38947
rect 97583 38913 97592 38947
rect 97540 38904 97592 38913
rect 848 38700 900 38752
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 96374 38598 96426 38650
rect 96438 38598 96490 38650
rect 96502 38598 96554 38650
rect 96566 38598 96618 38650
rect 96630 38598 96682 38650
rect 4874 38054 4926 38106
rect 4938 38054 4990 38106
rect 5002 38054 5054 38106
rect 5066 38054 5118 38106
rect 5130 38054 5182 38106
rect 97034 38054 97086 38106
rect 97098 38054 97150 38106
rect 97162 38054 97214 38106
rect 97226 38054 97278 38106
rect 97290 38054 97342 38106
rect 97356 37995 97408 38004
rect 97356 37961 97365 37995
rect 97365 37961 97399 37995
rect 97399 37961 97408 37995
rect 97356 37952 97408 37961
rect 8300 37816 8352 37868
rect 97540 37859 97592 37868
rect 97540 37825 97549 37859
rect 97549 37825 97583 37859
rect 97583 37825 97592 37859
rect 97540 37816 97592 37825
rect 848 37612 900 37664
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 96374 37510 96426 37562
rect 96438 37510 96490 37562
rect 96502 37510 96554 37562
rect 96566 37510 96618 37562
rect 96630 37510 96682 37562
rect 96620 37272 96672 37324
rect 8300 37204 8352 37256
rect 97448 37179 97500 37188
rect 97448 37145 97457 37179
rect 97457 37145 97491 37179
rect 97491 37145 97500 37179
rect 97448 37136 97500 37145
rect 848 37068 900 37120
rect 4874 36966 4926 37018
rect 4938 36966 4990 37018
rect 5002 36966 5054 37018
rect 5066 36966 5118 37018
rect 5130 36966 5182 37018
rect 97034 36966 97086 37018
rect 97098 36966 97150 37018
rect 97162 36966 97214 37018
rect 97226 36966 97278 37018
rect 97290 36966 97342 37018
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 96374 36422 96426 36474
rect 96438 36422 96490 36474
rect 96502 36422 96554 36474
rect 96566 36422 96618 36474
rect 96630 36422 96682 36474
rect 4874 35878 4926 35930
rect 4938 35878 4990 35930
rect 5002 35878 5054 35930
rect 5066 35878 5118 35930
rect 5130 35878 5182 35930
rect 97034 35878 97086 35930
rect 97098 35878 97150 35930
rect 97162 35878 97214 35930
rect 97226 35878 97278 35930
rect 97290 35878 97342 35930
rect 97356 35819 97408 35828
rect 97356 35785 97365 35819
rect 97365 35785 97399 35819
rect 97399 35785 97408 35819
rect 97356 35776 97408 35785
rect 8300 35640 8352 35692
rect 97540 35683 97592 35692
rect 97540 35649 97549 35683
rect 97549 35649 97583 35683
rect 97583 35649 97592 35683
rect 97540 35640 97592 35649
rect 848 35504 900 35556
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 96374 35334 96426 35386
rect 96438 35334 96490 35386
rect 96502 35334 96554 35386
rect 96566 35334 96618 35386
rect 96630 35334 96682 35386
rect 1676 35071 1728 35080
rect 1676 35037 1685 35071
rect 1685 35037 1719 35071
rect 1719 35037 1728 35071
rect 1676 35028 1728 35037
rect 97540 35071 97592 35080
rect 97540 35037 97549 35071
rect 97549 35037 97583 35071
rect 97583 35037 97592 35071
rect 97540 35028 97592 35037
rect 848 34892 900 34944
rect 97448 34892 97500 34944
rect 4874 34790 4926 34842
rect 4938 34790 4990 34842
rect 5002 34790 5054 34842
rect 5066 34790 5118 34842
rect 5130 34790 5182 34842
rect 97034 34790 97086 34842
rect 97098 34790 97150 34842
rect 97162 34790 97214 34842
rect 97226 34790 97278 34842
rect 97290 34790 97342 34842
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 96374 34246 96426 34298
rect 96438 34246 96490 34298
rect 96502 34246 96554 34298
rect 96566 34246 96618 34298
rect 96630 34246 96682 34298
rect 4874 33702 4926 33754
rect 4938 33702 4990 33754
rect 5002 33702 5054 33754
rect 5066 33702 5118 33754
rect 5130 33702 5182 33754
rect 97034 33702 97086 33754
rect 97098 33702 97150 33754
rect 97162 33702 97214 33754
rect 97226 33702 97278 33754
rect 97290 33702 97342 33754
rect 97356 33643 97408 33652
rect 97356 33609 97365 33643
rect 97365 33609 97399 33643
rect 97399 33609 97408 33643
rect 97356 33600 97408 33609
rect 8300 33464 8352 33516
rect 97540 33507 97592 33516
rect 97540 33473 97549 33507
rect 97549 33473 97583 33507
rect 97583 33473 97592 33507
rect 97540 33464 97592 33473
rect 848 33260 900 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 96374 33158 96426 33210
rect 96438 33158 96490 33210
rect 96502 33158 96554 33210
rect 96566 33158 96618 33210
rect 96630 33158 96682 33210
rect 4874 32614 4926 32666
rect 4938 32614 4990 32666
rect 5002 32614 5054 32666
rect 5066 32614 5118 32666
rect 5130 32614 5182 32666
rect 97034 32614 97086 32666
rect 97098 32614 97150 32666
rect 97162 32614 97214 32666
rect 97226 32614 97278 32666
rect 97290 32614 97342 32666
rect 97264 32487 97316 32496
rect 97264 32453 97273 32487
rect 97273 32453 97307 32487
rect 97307 32453 97316 32487
rect 97264 32444 97316 32453
rect 8300 32376 8352 32428
rect 97448 32419 97500 32428
rect 97448 32385 97457 32419
rect 97457 32385 97491 32419
rect 97491 32385 97500 32419
rect 97448 32376 97500 32385
rect 848 32172 900 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 96374 32070 96426 32122
rect 96438 32070 96490 32122
rect 96502 32070 96554 32122
rect 96566 32070 96618 32122
rect 96630 32070 96682 32122
rect 848 31900 900 31952
rect 96620 31900 96672 31952
rect 1676 31807 1728 31816
rect 1676 31773 1685 31807
rect 1685 31773 1719 31807
rect 1719 31773 1728 31807
rect 1676 31764 1728 31773
rect 97540 31807 97592 31816
rect 97540 31773 97549 31807
rect 97549 31773 97583 31807
rect 97583 31773 97592 31807
rect 97540 31764 97592 31773
rect 4874 31526 4926 31578
rect 4938 31526 4990 31578
rect 5002 31526 5054 31578
rect 5066 31526 5118 31578
rect 5130 31526 5182 31578
rect 97034 31526 97086 31578
rect 97098 31526 97150 31578
rect 97162 31526 97214 31578
rect 97226 31526 97278 31578
rect 97290 31526 97342 31578
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 96374 30982 96426 31034
rect 96438 30982 96490 31034
rect 96502 30982 96554 31034
rect 96566 30982 96618 31034
rect 96630 30982 96682 31034
rect 97540 30583 97592 30592
rect 97540 30549 97549 30583
rect 97549 30549 97583 30583
rect 97583 30549 97592 30583
rect 97540 30540 97592 30549
rect 4874 30438 4926 30490
rect 4938 30438 4990 30490
rect 5002 30438 5054 30490
rect 5066 30438 5118 30490
rect 5130 30438 5182 30490
rect 97034 30438 97086 30490
rect 97098 30438 97150 30490
rect 97162 30438 97214 30490
rect 97226 30438 97278 30490
rect 97290 30438 97342 30490
rect 8300 30200 8352 30252
rect 97264 30243 97316 30252
rect 97264 30209 97273 30243
rect 97273 30209 97307 30243
rect 97307 30209 97316 30243
rect 97264 30200 97316 30209
rect 97540 30175 97592 30184
rect 97540 30141 97549 30175
rect 97549 30141 97583 30175
rect 97583 30141 97592 30175
rect 97540 30132 97592 30141
rect 848 30064 900 30116
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 96374 29894 96426 29946
rect 96438 29894 96490 29946
rect 96502 29894 96554 29946
rect 96566 29894 96618 29946
rect 96630 29894 96682 29946
rect 8300 29588 8352 29640
rect 97540 29631 97592 29640
rect 97540 29597 97549 29631
rect 97549 29597 97583 29631
rect 97583 29597 97592 29631
rect 97540 29588 97592 29597
rect 848 29452 900 29504
rect 97448 29452 97500 29504
rect 4874 29350 4926 29402
rect 4938 29350 4990 29402
rect 5002 29350 5054 29402
rect 5066 29350 5118 29402
rect 5130 29350 5182 29402
rect 97034 29350 97086 29402
rect 97098 29350 97150 29402
rect 97162 29350 97214 29402
rect 97226 29350 97278 29402
rect 97290 29350 97342 29402
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 96374 28806 96426 28858
rect 96438 28806 96490 28858
rect 96502 28806 96554 28858
rect 96566 28806 96618 28858
rect 96630 28806 96682 28858
rect 4874 28262 4926 28314
rect 4938 28262 4990 28314
rect 5002 28262 5054 28314
rect 5066 28262 5118 28314
rect 5130 28262 5182 28314
rect 97034 28262 97086 28314
rect 97098 28262 97150 28314
rect 97162 28262 97214 28314
rect 97226 28262 97278 28314
rect 97290 28262 97342 28314
rect 8300 28160 8352 28212
rect 1308 28024 1360 28076
rect 97264 28067 97316 28076
rect 97264 28033 97273 28067
rect 97273 28033 97307 28067
rect 97307 28033 97316 28067
rect 97264 28024 97316 28033
rect 97448 27931 97500 27940
rect 97448 27897 97457 27931
rect 97457 27897 97491 27931
rect 97491 27897 97500 27931
rect 97448 27888 97500 27897
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 96374 27718 96426 27770
rect 96438 27718 96490 27770
rect 96502 27718 96554 27770
rect 96566 27718 96618 27770
rect 96630 27718 96682 27770
rect 4874 27174 4926 27226
rect 4938 27174 4990 27226
rect 5002 27174 5054 27226
rect 5066 27174 5118 27226
rect 5130 27174 5182 27226
rect 97034 27174 97086 27226
rect 97098 27174 97150 27226
rect 97162 27174 97214 27226
rect 97226 27174 97278 27226
rect 97290 27174 97342 27226
rect 1308 26936 1360 26988
rect 8300 26936 8352 26988
rect 97264 26979 97316 26988
rect 97264 26945 97273 26979
rect 97273 26945 97307 26979
rect 97307 26945 97316 26979
rect 97264 26936 97316 26945
rect 97448 26775 97500 26784
rect 97448 26741 97457 26775
rect 97457 26741 97491 26775
rect 97491 26741 97500 26775
rect 97448 26732 97500 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 96374 26630 96426 26682
rect 96438 26630 96490 26682
rect 96502 26630 96554 26682
rect 96566 26630 96618 26682
rect 96630 26630 96682 26682
rect 97448 26503 97500 26512
rect 97448 26469 97457 26503
rect 97457 26469 97491 26503
rect 97491 26469 97500 26503
rect 97448 26460 97500 26469
rect 1308 26324 1360 26376
rect 96896 26324 96948 26376
rect 1676 26299 1728 26308
rect 1676 26265 1685 26299
rect 1685 26265 1719 26299
rect 1719 26265 1728 26299
rect 1676 26256 1728 26265
rect 4874 26086 4926 26138
rect 4938 26086 4990 26138
rect 5002 26086 5054 26138
rect 5066 26086 5118 26138
rect 5130 26086 5182 26138
rect 97034 26086 97086 26138
rect 97098 26086 97150 26138
rect 97162 26086 97214 26138
rect 97226 26086 97278 26138
rect 97290 26086 97342 26138
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 96374 25542 96426 25594
rect 96438 25542 96490 25594
rect 96502 25542 96554 25594
rect 96566 25542 96618 25594
rect 96630 25542 96682 25594
rect 4874 24998 4926 25050
rect 4938 24998 4990 25050
rect 5002 24998 5054 25050
rect 5066 24998 5118 25050
rect 5130 24998 5182 25050
rect 97034 24998 97086 25050
rect 97098 24998 97150 25050
rect 97162 24998 97214 25050
rect 97226 24998 97278 25050
rect 97290 24998 97342 25050
rect 1308 24760 1360 24812
rect 8300 24760 8352 24812
rect 97264 24803 97316 24812
rect 97264 24769 97273 24803
rect 97273 24769 97307 24803
rect 97307 24769 97316 24803
rect 97264 24760 97316 24769
rect 97448 24599 97500 24608
rect 97448 24565 97457 24599
rect 97457 24565 97491 24599
rect 97491 24565 97500 24599
rect 97448 24556 97500 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 96374 24454 96426 24506
rect 96438 24454 96490 24506
rect 96502 24454 96554 24506
rect 96566 24454 96618 24506
rect 96630 24454 96682 24506
rect 96620 24148 96672 24200
rect 1308 24080 1360 24132
rect 8300 24080 8352 24132
rect 97448 24055 97500 24064
rect 97448 24021 97457 24055
rect 97457 24021 97491 24055
rect 97491 24021 97500 24055
rect 97448 24012 97500 24021
rect 4874 23910 4926 23962
rect 4938 23910 4990 23962
rect 5002 23910 5054 23962
rect 5066 23910 5118 23962
rect 5130 23910 5182 23962
rect 97034 23910 97086 23962
rect 97098 23910 97150 23962
rect 97162 23910 97214 23962
rect 97226 23910 97278 23962
rect 97290 23910 97342 23962
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 96374 23366 96426 23418
rect 96438 23366 96490 23418
rect 96502 23366 96554 23418
rect 96566 23366 96618 23418
rect 96630 23366 96682 23418
rect 4874 22822 4926 22874
rect 4938 22822 4990 22874
rect 5002 22822 5054 22874
rect 5066 22822 5118 22874
rect 5130 22822 5182 22874
rect 97034 22822 97086 22874
rect 97098 22822 97150 22874
rect 97162 22822 97214 22874
rect 97226 22822 97278 22874
rect 97290 22822 97342 22874
rect 1124 22584 1176 22636
rect 8300 22584 8352 22636
rect 97264 22627 97316 22636
rect 97264 22593 97273 22627
rect 97273 22593 97307 22627
rect 97307 22593 97316 22627
rect 97264 22584 97316 22593
rect 97448 22491 97500 22500
rect 97448 22457 97457 22491
rect 97457 22457 97491 22491
rect 97491 22457 97500 22491
rect 97448 22448 97500 22457
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 96374 22278 96426 22330
rect 96438 22278 96490 22330
rect 96502 22278 96554 22330
rect 96566 22278 96618 22330
rect 96630 22278 96682 22330
rect 4874 21734 4926 21786
rect 4938 21734 4990 21786
rect 5002 21734 5054 21786
rect 5066 21734 5118 21786
rect 5130 21734 5182 21786
rect 97034 21734 97086 21786
rect 97098 21734 97150 21786
rect 97162 21734 97214 21786
rect 97226 21734 97278 21786
rect 97290 21734 97342 21786
rect 1308 21496 1360 21548
rect 8300 21496 8352 21548
rect 97264 21539 97316 21548
rect 97264 21505 97273 21539
rect 97273 21505 97307 21539
rect 97307 21505 97316 21539
rect 97264 21496 97316 21505
rect 97448 21335 97500 21344
rect 97448 21301 97457 21335
rect 97457 21301 97491 21335
rect 97491 21301 97500 21335
rect 97448 21292 97500 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 96374 21190 96426 21242
rect 96438 21190 96490 21242
rect 96502 21190 96554 21242
rect 96566 21190 96618 21242
rect 96630 21190 96682 21242
rect 96620 20884 96672 20936
rect 1308 20816 1360 20868
rect 1860 20859 1912 20868
rect 1860 20825 1869 20859
rect 1869 20825 1903 20859
rect 1903 20825 1912 20859
rect 1860 20816 1912 20825
rect 97448 20791 97500 20800
rect 97448 20757 97457 20791
rect 97457 20757 97491 20791
rect 97491 20757 97500 20791
rect 97448 20748 97500 20757
rect 4874 20646 4926 20698
rect 4938 20646 4990 20698
rect 5002 20646 5054 20698
rect 5066 20646 5118 20698
rect 5130 20646 5182 20698
rect 97034 20646 97086 20698
rect 97098 20646 97150 20698
rect 97162 20646 97214 20698
rect 97226 20646 97278 20698
rect 97290 20646 97342 20698
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 96374 20102 96426 20154
rect 96438 20102 96490 20154
rect 96502 20102 96554 20154
rect 96566 20102 96618 20154
rect 96630 20102 96682 20154
rect 4874 19558 4926 19610
rect 4938 19558 4990 19610
rect 5002 19558 5054 19610
rect 5066 19558 5118 19610
rect 5130 19558 5182 19610
rect 97034 19558 97086 19610
rect 97098 19558 97150 19610
rect 97162 19558 97214 19610
rect 97226 19558 97278 19610
rect 97290 19558 97342 19610
rect 97448 19499 97500 19508
rect 97448 19465 97457 19499
rect 97457 19465 97491 19499
rect 97491 19465 97500 19499
rect 97448 19456 97500 19465
rect 1492 19363 1544 19372
rect 1492 19329 1501 19363
rect 1501 19329 1535 19363
rect 1535 19329 1544 19363
rect 1492 19320 1544 19329
rect 97264 19363 97316 19372
rect 97264 19329 97273 19363
rect 97273 19329 97307 19363
rect 97307 19329 97316 19363
rect 97264 19320 97316 19329
rect 8300 19184 8352 19236
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 96374 19014 96426 19066
rect 96438 19014 96490 19066
rect 96502 19014 96554 19066
rect 96566 19014 96618 19066
rect 96630 19014 96682 19066
rect 96620 18708 96672 18760
rect 1308 18640 1360 18692
rect 8300 18640 8352 18692
rect 97448 18615 97500 18624
rect 97448 18581 97457 18615
rect 97457 18581 97491 18615
rect 97491 18581 97500 18615
rect 97448 18572 97500 18581
rect 4874 18470 4926 18522
rect 4938 18470 4990 18522
rect 5002 18470 5054 18522
rect 5066 18470 5118 18522
rect 5130 18470 5182 18522
rect 97034 18470 97086 18522
rect 97098 18470 97150 18522
rect 97162 18470 97214 18522
rect 97226 18470 97278 18522
rect 97290 18470 97342 18522
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 96374 17926 96426 17978
rect 96438 17926 96490 17978
rect 96502 17926 96554 17978
rect 96566 17926 96618 17978
rect 96630 17926 96682 17978
rect 4874 17382 4926 17434
rect 4938 17382 4990 17434
rect 5002 17382 5054 17434
rect 5066 17382 5118 17434
rect 5130 17382 5182 17434
rect 97034 17382 97086 17434
rect 97098 17382 97150 17434
rect 97162 17382 97214 17434
rect 97226 17382 97278 17434
rect 97290 17382 97342 17434
rect 8300 17280 8352 17332
rect 1124 17144 1176 17196
rect 97264 17187 97316 17196
rect 97264 17153 97273 17187
rect 97273 17153 97307 17187
rect 97307 17153 97316 17187
rect 97264 17144 97316 17153
rect 97448 17051 97500 17060
rect 97448 17017 97457 17051
rect 97457 17017 97491 17051
rect 97491 17017 97500 17051
rect 97448 17008 97500 17017
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 96374 16838 96426 16890
rect 96438 16838 96490 16890
rect 96502 16838 96554 16890
rect 96566 16838 96618 16890
rect 96630 16838 96682 16890
rect 4874 16294 4926 16346
rect 4938 16294 4990 16346
rect 5002 16294 5054 16346
rect 5066 16294 5118 16346
rect 5130 16294 5182 16346
rect 97034 16294 97086 16346
rect 97098 16294 97150 16346
rect 97162 16294 97214 16346
rect 97226 16294 97278 16346
rect 97290 16294 97342 16346
rect 8300 16192 8352 16244
rect 1216 16056 1268 16108
rect 97264 16099 97316 16108
rect 97264 16065 97273 16099
rect 97273 16065 97307 16099
rect 97307 16065 97316 16099
rect 97264 16056 97316 16065
rect 97448 15895 97500 15904
rect 97448 15861 97457 15895
rect 97457 15861 97491 15895
rect 97491 15861 97500 15895
rect 97448 15852 97500 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 96374 15750 96426 15802
rect 96438 15750 96490 15802
rect 96502 15750 96554 15802
rect 96566 15750 96618 15802
rect 96630 15750 96682 15802
rect 96620 15444 96672 15496
rect 1308 15376 1360 15428
rect 1860 15419 1912 15428
rect 1860 15385 1869 15419
rect 1869 15385 1903 15419
rect 1903 15385 1912 15419
rect 1860 15376 1912 15385
rect 97448 15351 97500 15360
rect 97448 15317 97457 15351
rect 97457 15317 97491 15351
rect 97491 15317 97500 15351
rect 97448 15308 97500 15317
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 97034 15206 97086 15258
rect 97098 15206 97150 15258
rect 97162 15206 97214 15258
rect 97226 15206 97278 15258
rect 97290 15206 97342 15258
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 96374 14662 96426 14714
rect 96438 14662 96490 14714
rect 96502 14662 96554 14714
rect 96566 14662 96618 14714
rect 96630 14662 96682 14714
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 97034 14118 97086 14170
rect 97098 14118 97150 14170
rect 97162 14118 97214 14170
rect 97226 14118 97278 14170
rect 97290 14118 97342 14170
rect 97448 14059 97500 14068
rect 97448 14025 97457 14059
rect 97457 14025 97491 14059
rect 97491 14025 97500 14059
rect 97448 14016 97500 14025
rect 1308 13880 1360 13932
rect 8300 13880 8352 13932
rect 97264 13923 97316 13932
rect 97264 13889 97273 13923
rect 97273 13889 97307 13923
rect 97307 13889 97316 13923
rect 97264 13880 97316 13889
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 96374 13574 96426 13626
rect 96438 13574 96490 13626
rect 96502 13574 96554 13626
rect 96566 13574 96618 13626
rect 96630 13574 96682 13626
rect 8300 13404 8352 13456
rect 1308 13268 1360 13320
rect 96620 13268 96672 13320
rect 97448 13175 97500 13184
rect 97448 13141 97457 13175
rect 97457 13141 97491 13175
rect 97491 13141 97500 13175
rect 97448 13132 97500 13141
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 97034 13030 97086 13082
rect 97098 13030 97150 13082
rect 97162 13030 97214 13082
rect 97226 13030 97278 13082
rect 97290 13030 97342 13082
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 96374 12486 96426 12538
rect 96438 12486 96490 12538
rect 96502 12486 96554 12538
rect 96566 12486 96618 12538
rect 96630 12486 96682 12538
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 97034 11942 97086 11994
rect 97098 11942 97150 11994
rect 97162 11942 97214 11994
rect 97226 11942 97278 11994
rect 97290 11942 97342 11994
rect 8300 11840 8352 11892
rect 1124 11704 1176 11756
rect 97264 11747 97316 11756
rect 97264 11713 97273 11747
rect 97273 11713 97307 11747
rect 97307 11713 97316 11747
rect 97264 11704 97316 11713
rect 97448 11611 97500 11620
rect 97448 11577 97457 11611
rect 97457 11577 97491 11611
rect 97491 11577 97500 11611
rect 97448 11568 97500 11577
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 96374 11398 96426 11450
rect 96438 11398 96490 11450
rect 96502 11398 96554 11450
rect 96566 11398 96618 11450
rect 96630 11398 96682 11450
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 97034 10854 97086 10906
rect 97098 10854 97150 10906
rect 97162 10854 97214 10906
rect 97226 10854 97278 10906
rect 97290 10854 97342 10906
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 96374 10310 96426 10362
rect 96438 10310 96490 10362
rect 96502 10310 96554 10362
rect 96566 10310 96618 10362
rect 96630 10310 96682 10362
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 97034 9766 97086 9818
rect 97098 9766 97150 9818
rect 97162 9766 97214 9818
rect 97226 9766 97278 9818
rect 97290 9766 97342 9818
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 96374 9222 96426 9274
rect 96438 9222 96490 9274
rect 96502 9222 96554 9274
rect 96566 9222 96618 9274
rect 96630 9222 96682 9274
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 97034 8678 97086 8730
rect 97098 8678 97150 8730
rect 97162 8678 97214 8730
rect 97226 8678 97278 8730
rect 97290 8678 97342 8730
rect 9128 8576 9180 8628
rect 50344 8576 50396 8628
rect 97540 8483 97592 8492
rect 97540 8449 97549 8483
rect 97549 8449 97583 8483
rect 97583 8449 97592 8483
rect 97540 8440 97592 8449
rect 90916 8304 90968 8356
rect 8208 8236 8260 8288
rect 9680 8236 9732 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 8116 8168 8168 8220
rect 11152 8168 11204 8220
rect 8024 8100 8076 8152
rect 11796 8100 11848 8152
rect 54484 8100 54536 8152
rect 91928 8100 91980 8152
rect 96374 8134 96426 8186
rect 96438 8134 96490 8186
rect 96502 8134 96554 8186
rect 96566 8134 96618 8186
rect 96630 8134 96682 8186
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 97034 7590 97086 7642
rect 97098 7590 97150 7642
rect 97162 7590 97214 7642
rect 97226 7590 97278 7642
rect 97290 7590 97342 7642
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 96374 7046 96426 7098
rect 96438 7046 96490 7098
rect 96502 7046 96554 7098
rect 96566 7046 96618 7098
rect 96630 7046 96682 7098
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 97034 6502 97086 6554
rect 97098 6502 97150 6554
rect 97162 6502 97214 6554
rect 97226 6502 97278 6554
rect 97290 6502 97342 6554
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 65654 5958 65706 6010
rect 65718 5958 65770 6010
rect 65782 5958 65834 6010
rect 65846 5958 65898 6010
rect 65910 5958 65962 6010
rect 96374 5958 96426 6010
rect 96438 5958 96490 6010
rect 96502 5958 96554 6010
rect 96566 5958 96618 6010
rect 96630 5958 96682 6010
rect 8944 5899 8996 5908
rect 8944 5865 8953 5899
rect 8953 5865 8987 5899
rect 8987 5865 8996 5899
rect 8944 5856 8996 5865
rect 12164 5899 12216 5908
rect 12164 5865 12173 5899
rect 12173 5865 12207 5899
rect 12207 5865 12216 5899
rect 12164 5856 12216 5865
rect 12808 5856 12860 5908
rect 50620 5856 50672 5908
rect 51080 5899 51132 5908
rect 51080 5865 51089 5899
rect 51089 5865 51123 5899
rect 51123 5865 51132 5899
rect 51080 5856 51132 5865
rect 10048 5763 10100 5772
rect 10048 5729 10057 5763
rect 10057 5729 10091 5763
rect 10091 5729 10100 5763
rect 10048 5720 10100 5729
rect 10968 5720 11020 5772
rect 52000 5763 52052 5772
rect 52000 5729 52009 5763
rect 52009 5729 52043 5763
rect 52043 5729 52052 5763
rect 52000 5720 52052 5729
rect 11152 5695 11204 5704
rect 11152 5661 11161 5695
rect 11161 5661 11195 5695
rect 11195 5661 11204 5695
rect 11152 5652 11204 5661
rect 13176 5652 13228 5704
rect 53104 5695 53156 5704
rect 53104 5661 53113 5695
rect 53113 5661 53147 5695
rect 53147 5661 53156 5695
rect 53104 5652 53156 5661
rect 12808 5584 12860 5636
rect 54116 5584 54168 5636
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 35594 5414 35646 5466
rect 35658 5414 35710 5466
rect 35722 5414 35774 5466
rect 35786 5414 35838 5466
rect 35850 5414 35902 5466
rect 66314 5414 66366 5466
rect 66378 5414 66430 5466
rect 66442 5414 66494 5466
rect 66506 5414 66558 5466
rect 66570 5414 66622 5466
rect 97034 5414 97086 5466
rect 97098 5414 97150 5466
rect 97162 5414 97214 5466
rect 97226 5414 97278 5466
rect 97290 5414 97342 5466
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 65654 4870 65706 4922
rect 65718 4870 65770 4922
rect 65782 4870 65834 4922
rect 65846 4870 65898 4922
rect 65910 4870 65962 4922
rect 96374 4870 96426 4922
rect 96438 4870 96490 4922
rect 96502 4870 96554 4922
rect 96566 4870 96618 4922
rect 96630 4870 96682 4922
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 35594 4326 35646 4378
rect 35658 4326 35710 4378
rect 35722 4326 35774 4378
rect 35786 4326 35838 4378
rect 35850 4326 35902 4378
rect 66314 4326 66366 4378
rect 66378 4326 66430 4378
rect 66442 4326 66494 4378
rect 66506 4326 66558 4378
rect 66570 4326 66622 4378
rect 97034 4326 97086 4378
rect 97098 4326 97150 4378
rect 97162 4326 97214 4378
rect 97226 4326 97278 4378
rect 97290 4326 97342 4378
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 65654 3782 65706 3834
rect 65718 3782 65770 3834
rect 65782 3782 65834 3834
rect 65846 3782 65898 3834
rect 65910 3782 65962 3834
rect 96374 3782 96426 3834
rect 96438 3782 96490 3834
rect 96502 3782 96554 3834
rect 96566 3782 96618 3834
rect 96630 3782 96682 3834
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 35594 3238 35646 3290
rect 35658 3238 35710 3290
rect 35722 3238 35774 3290
rect 35786 3238 35838 3290
rect 35850 3238 35902 3290
rect 66314 3238 66366 3290
rect 66378 3238 66430 3290
rect 66442 3238 66494 3290
rect 66506 3238 66558 3290
rect 66570 3238 66622 3290
rect 97034 3238 97086 3290
rect 97098 3238 97150 3290
rect 97162 3238 97214 3290
rect 97226 3238 97278 3290
rect 97290 3238 97342 3290
rect 13176 3179 13228 3188
rect 13176 3145 13185 3179
rect 13185 3145 13219 3179
rect 13219 3145 13228 3179
rect 13176 3136 13228 3145
rect 11612 3000 11664 3052
rect 11612 2839 11664 2848
rect 11612 2805 11621 2839
rect 11621 2805 11655 2839
rect 11655 2805 11664 2839
rect 11612 2796 11664 2805
rect 89536 2839 89588 2848
rect 89536 2805 89545 2839
rect 89545 2805 89579 2839
rect 89579 2805 89588 2839
rect 89536 2796 89588 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 65654 2694 65706 2746
rect 65718 2694 65770 2746
rect 65782 2694 65834 2746
rect 65846 2694 65898 2746
rect 65910 2694 65962 2746
rect 96374 2694 96426 2746
rect 96438 2694 96490 2746
rect 96502 2694 96554 2746
rect 96566 2694 96618 2746
rect 96630 2694 96682 2746
rect 10968 2592 11020 2644
rect 32312 2635 32364 2644
rect 32312 2601 32321 2635
rect 32321 2601 32355 2635
rect 32355 2601 32364 2635
rect 32312 2592 32364 2601
rect 33140 2635 33192 2644
rect 33140 2601 33149 2635
rect 33149 2601 33183 2635
rect 33183 2601 33192 2635
rect 33140 2592 33192 2601
rect 34244 2635 34296 2644
rect 34244 2601 34253 2635
rect 34253 2601 34287 2635
rect 34287 2601 34296 2635
rect 34244 2592 34296 2601
rect 35348 2592 35400 2644
rect 36452 2592 36504 2644
rect 37648 2635 37700 2644
rect 37648 2601 37657 2635
rect 37657 2601 37691 2635
rect 37691 2601 37700 2635
rect 37648 2592 37700 2601
rect 38752 2635 38804 2644
rect 38752 2601 38761 2635
rect 38761 2601 38795 2635
rect 38795 2601 38804 2635
rect 38752 2592 38804 2601
rect 40040 2635 40092 2644
rect 40040 2601 40049 2635
rect 40049 2601 40083 2635
rect 40083 2601 40092 2635
rect 40040 2592 40092 2601
rect 40868 2635 40920 2644
rect 40868 2601 40877 2635
rect 40877 2601 40911 2635
rect 40911 2601 40920 2635
rect 40868 2592 40920 2601
rect 41972 2635 42024 2644
rect 41972 2601 41981 2635
rect 41981 2601 42015 2635
rect 42015 2601 42024 2635
rect 41972 2592 42024 2601
rect 43260 2635 43312 2644
rect 43260 2601 43269 2635
rect 43269 2601 43303 2635
rect 43303 2601 43312 2635
rect 43260 2592 43312 2601
rect 48780 2635 48832 2644
rect 48780 2601 48789 2635
rect 48789 2601 48823 2635
rect 48823 2601 48832 2635
rect 48780 2592 48832 2601
rect 74172 2635 74224 2644
rect 74172 2601 74181 2635
rect 74181 2601 74215 2635
rect 74215 2601 74224 2635
rect 74172 2592 74224 2601
rect 75460 2635 75512 2644
rect 75460 2601 75469 2635
rect 75469 2601 75503 2635
rect 75503 2601 75512 2635
rect 75460 2592 75512 2601
rect 76288 2635 76340 2644
rect 76288 2601 76297 2635
rect 76297 2601 76331 2635
rect 76331 2601 76340 2635
rect 76288 2592 76340 2601
rect 77392 2635 77444 2644
rect 77392 2601 77401 2635
rect 77401 2601 77435 2635
rect 77435 2601 77444 2635
rect 77392 2592 77444 2601
rect 78680 2635 78732 2644
rect 78680 2601 78689 2635
rect 78689 2601 78723 2635
rect 78723 2601 78732 2635
rect 78680 2592 78732 2601
rect 79508 2635 79560 2644
rect 79508 2601 79517 2635
rect 79517 2601 79551 2635
rect 79551 2601 79560 2635
rect 79508 2592 79560 2601
rect 80796 2635 80848 2644
rect 80796 2601 80805 2635
rect 80805 2601 80839 2635
rect 80839 2601 80848 2635
rect 80796 2592 80848 2601
rect 81900 2635 81952 2644
rect 81900 2601 81909 2635
rect 81909 2601 81943 2635
rect 81943 2601 81952 2635
rect 81900 2592 81952 2601
rect 83188 2635 83240 2644
rect 83188 2601 83197 2635
rect 83197 2601 83231 2635
rect 83231 2601 83240 2635
rect 83188 2592 83240 2601
rect 84016 2635 84068 2644
rect 84016 2601 84025 2635
rect 84025 2601 84059 2635
rect 84059 2601 84068 2635
rect 84016 2592 84068 2601
rect 85120 2635 85172 2644
rect 85120 2601 85129 2635
rect 85129 2601 85163 2635
rect 85163 2601 85172 2635
rect 85120 2592 85172 2601
rect 44180 2524 44232 2576
rect 86408 2567 86460 2576
rect 86408 2533 86417 2567
rect 86417 2533 86451 2567
rect 86451 2533 86460 2567
rect 86408 2524 86460 2533
rect 12808 2499 12860 2508
rect 12808 2465 12817 2499
rect 12817 2465 12851 2499
rect 12851 2465 12860 2499
rect 12808 2456 12860 2465
rect 45468 2499 45520 2508
rect 45468 2465 45477 2499
rect 45477 2465 45511 2499
rect 45511 2465 45520 2499
rect 45468 2456 45520 2465
rect 46388 2456 46440 2508
rect 47492 2456 47544 2508
rect 87328 2499 87380 2508
rect 87328 2465 87337 2499
rect 87337 2465 87371 2499
rect 87371 2465 87380 2499
rect 87328 2456 87380 2465
rect 88708 2456 88760 2508
rect 89812 2456 89864 2508
rect 10324 2388 10376 2440
rect 14556 2431 14608 2440
rect 14556 2397 14565 2431
rect 14565 2397 14599 2431
rect 14599 2397 14608 2431
rect 14556 2388 14608 2397
rect 15568 2431 15620 2440
rect 15568 2397 15577 2431
rect 15577 2397 15611 2431
rect 15611 2397 15620 2431
rect 15568 2388 15620 2397
rect 16856 2431 16908 2440
rect 16856 2397 16865 2431
rect 16865 2397 16899 2431
rect 16899 2397 16908 2431
rect 16856 2388 16908 2397
rect 17776 2431 17828 2440
rect 17776 2397 17785 2431
rect 17785 2397 17819 2431
rect 17819 2397 17828 2431
rect 17776 2388 17828 2397
rect 18788 2431 18840 2440
rect 18788 2397 18797 2431
rect 18797 2397 18831 2431
rect 18831 2397 18840 2431
rect 18788 2388 18840 2397
rect 20076 2431 20128 2440
rect 20076 2397 20085 2431
rect 20085 2397 20119 2431
rect 20119 2397 20128 2431
rect 20076 2388 20128 2397
rect 20996 2388 21048 2440
rect 22284 2431 22336 2440
rect 22284 2397 22293 2431
rect 22293 2397 22327 2431
rect 22327 2397 22336 2431
rect 22284 2388 22336 2397
rect 23296 2431 23348 2440
rect 23296 2397 23305 2431
rect 23305 2397 23339 2431
rect 23339 2397 23348 2431
rect 23296 2388 23348 2397
rect 24584 2431 24636 2440
rect 24584 2397 24593 2431
rect 24593 2397 24627 2431
rect 24627 2397 24636 2431
rect 24584 2388 24636 2397
rect 25504 2431 25556 2440
rect 25504 2397 25513 2431
rect 25513 2397 25547 2431
rect 25547 2397 25556 2431
rect 25504 2388 25556 2397
rect 26516 2431 26568 2440
rect 26516 2397 26525 2431
rect 26525 2397 26559 2431
rect 26559 2397 26568 2431
rect 26516 2388 26568 2397
rect 27804 2431 27856 2440
rect 27804 2397 27813 2431
rect 27813 2397 27847 2431
rect 27847 2397 27856 2431
rect 27804 2388 27856 2397
rect 29092 2431 29144 2440
rect 29092 2397 29101 2431
rect 29101 2397 29135 2431
rect 29135 2397 29144 2431
rect 29092 2388 29144 2397
rect 30012 2431 30064 2440
rect 30012 2397 30021 2431
rect 30021 2397 30055 2431
rect 30055 2397 30064 2431
rect 30012 2388 30064 2397
rect 31024 2431 31076 2440
rect 31024 2397 31033 2431
rect 31033 2397 31067 2431
rect 31067 2397 31076 2431
rect 31024 2388 31076 2397
rect 12256 2295 12308 2304
rect 12256 2261 12265 2295
rect 12265 2261 12299 2295
rect 12299 2261 12308 2295
rect 12256 2252 12308 2261
rect 14188 2252 14240 2304
rect 15476 2252 15528 2304
rect 16764 2252 16816 2304
rect 17408 2252 17460 2304
rect 18696 2252 18748 2304
rect 19984 2252 20036 2304
rect 21272 2252 21324 2304
rect 21916 2252 21968 2304
rect 23204 2252 23256 2304
rect 24492 2252 24544 2304
rect 25136 2252 25188 2304
rect 26424 2252 26476 2304
rect 27712 2252 27764 2304
rect 29000 2252 29052 2304
rect 29644 2252 29696 2304
rect 30932 2252 30984 2304
rect 32220 2295 32272 2304
rect 32220 2261 32229 2295
rect 32229 2261 32263 2295
rect 32263 2261 32272 2295
rect 32220 2252 32272 2261
rect 32864 2295 32916 2304
rect 32864 2261 32873 2295
rect 32873 2261 32907 2295
rect 32907 2261 32916 2295
rect 32864 2252 32916 2261
rect 34152 2295 34204 2304
rect 34152 2261 34161 2295
rect 34161 2261 34195 2295
rect 34195 2261 34204 2295
rect 34152 2252 34204 2261
rect 35440 2295 35492 2304
rect 35440 2261 35449 2295
rect 35449 2261 35483 2295
rect 35483 2261 35492 2295
rect 35440 2252 35492 2261
rect 36728 2295 36780 2304
rect 36728 2261 36737 2295
rect 36737 2261 36771 2295
rect 36771 2261 36780 2295
rect 36728 2252 36780 2261
rect 37372 2295 37424 2304
rect 37372 2261 37381 2295
rect 37381 2261 37415 2295
rect 37415 2261 37424 2295
rect 37372 2252 37424 2261
rect 38660 2295 38712 2304
rect 38660 2261 38669 2295
rect 38669 2261 38703 2295
rect 38703 2261 38712 2295
rect 38660 2252 38712 2261
rect 39948 2295 40000 2304
rect 39948 2261 39957 2295
rect 39957 2261 39991 2295
rect 39991 2261 40000 2295
rect 39948 2252 40000 2261
rect 40592 2295 40644 2304
rect 40592 2261 40601 2295
rect 40601 2261 40635 2295
rect 40635 2261 40644 2295
rect 40592 2252 40644 2261
rect 41880 2295 41932 2304
rect 41880 2261 41889 2295
rect 41889 2261 41923 2295
rect 41923 2261 41932 2295
rect 41880 2252 41932 2261
rect 43168 2295 43220 2304
rect 43168 2261 43177 2295
rect 43177 2261 43211 2295
rect 43211 2261 43220 2295
rect 43168 2252 43220 2261
rect 44456 2295 44508 2304
rect 44456 2261 44465 2295
rect 44465 2261 44499 2295
rect 44499 2261 44508 2295
rect 44456 2252 44508 2261
rect 45100 2295 45152 2304
rect 45100 2261 45109 2295
rect 45109 2261 45143 2295
rect 45143 2261 45152 2295
rect 45100 2252 45152 2261
rect 46388 2295 46440 2304
rect 46388 2261 46397 2295
rect 46397 2261 46431 2295
rect 46431 2261 46440 2295
rect 46388 2252 46440 2261
rect 47676 2295 47728 2304
rect 47676 2261 47685 2295
rect 47685 2261 47719 2295
rect 47719 2261 47728 2295
rect 47676 2252 47728 2261
rect 48320 2252 48372 2304
rect 56416 2431 56468 2440
rect 56416 2397 56425 2431
rect 56425 2397 56459 2431
rect 56459 2397 56468 2431
rect 56416 2388 56468 2397
rect 57428 2431 57480 2440
rect 57428 2397 57437 2431
rect 57437 2397 57471 2431
rect 57471 2397 57480 2431
rect 57428 2388 57480 2397
rect 58716 2431 58768 2440
rect 58716 2397 58725 2431
rect 58725 2397 58759 2431
rect 58759 2397 58768 2431
rect 58716 2388 58768 2397
rect 60004 2431 60056 2440
rect 60004 2397 60013 2431
rect 60013 2397 60047 2431
rect 60047 2397 60056 2431
rect 60004 2388 60056 2397
rect 60924 2431 60976 2440
rect 60924 2397 60933 2431
rect 60933 2397 60967 2431
rect 60967 2397 60976 2431
rect 60924 2388 60976 2397
rect 61936 2431 61988 2440
rect 61936 2397 61945 2431
rect 61945 2397 61979 2431
rect 61979 2397 61988 2431
rect 61936 2388 61988 2397
rect 63224 2431 63276 2440
rect 63224 2397 63233 2431
rect 63233 2397 63267 2431
rect 63267 2397 63276 2431
rect 63224 2388 63276 2397
rect 64144 2431 64196 2440
rect 64144 2397 64153 2431
rect 64153 2397 64187 2431
rect 64187 2397 64196 2431
rect 64144 2388 64196 2397
rect 65156 2431 65208 2440
rect 65156 2397 65165 2431
rect 65165 2397 65199 2431
rect 65199 2397 65208 2431
rect 65156 2388 65208 2397
rect 66720 2388 66772 2440
rect 67732 2431 67784 2440
rect 67732 2397 67741 2431
rect 67741 2397 67775 2431
rect 67775 2397 67784 2431
rect 67732 2388 67784 2397
rect 68652 2431 68704 2440
rect 68652 2397 68661 2431
rect 68661 2397 68695 2431
rect 68695 2397 68704 2431
rect 68652 2388 68704 2397
rect 69664 2431 69716 2440
rect 69664 2397 69673 2431
rect 69673 2397 69707 2431
rect 69707 2397 69716 2431
rect 69664 2388 69716 2397
rect 70952 2431 71004 2440
rect 70952 2397 70961 2431
rect 70961 2397 70995 2431
rect 70995 2397 71004 2431
rect 70952 2388 71004 2397
rect 71872 2431 71924 2440
rect 71872 2397 71881 2431
rect 71881 2397 71915 2431
rect 71915 2397 71924 2431
rect 71872 2388 71924 2397
rect 72884 2431 72936 2440
rect 72884 2397 72893 2431
rect 72893 2397 72927 2431
rect 72927 2397 72936 2431
rect 72884 2388 72936 2397
rect 56048 2252 56100 2304
rect 57336 2252 57388 2304
rect 58624 2252 58676 2304
rect 59912 2252 59964 2304
rect 60556 2252 60608 2304
rect 61844 2252 61896 2304
rect 63132 2252 63184 2304
rect 63776 2252 63828 2304
rect 65064 2252 65116 2304
rect 66720 2252 66772 2304
rect 67640 2252 67692 2304
rect 68284 2252 68336 2304
rect 69572 2252 69624 2304
rect 70860 2252 70912 2304
rect 71504 2252 71556 2304
rect 72792 2252 72844 2304
rect 74080 2295 74132 2304
rect 74080 2261 74089 2295
rect 74089 2261 74123 2295
rect 74123 2261 74132 2295
rect 74080 2252 74132 2261
rect 75368 2295 75420 2304
rect 75368 2261 75377 2295
rect 75377 2261 75411 2295
rect 75411 2261 75420 2295
rect 75368 2252 75420 2261
rect 76012 2295 76064 2304
rect 76012 2261 76021 2295
rect 76021 2261 76055 2295
rect 76055 2261 76064 2295
rect 76012 2252 76064 2261
rect 77300 2295 77352 2304
rect 77300 2261 77309 2295
rect 77309 2261 77343 2295
rect 77343 2261 77352 2295
rect 77300 2252 77352 2261
rect 78588 2295 78640 2304
rect 78588 2261 78597 2295
rect 78597 2261 78631 2295
rect 78631 2261 78640 2295
rect 78588 2252 78640 2261
rect 79232 2295 79284 2304
rect 79232 2261 79241 2295
rect 79241 2261 79275 2295
rect 79275 2261 79284 2295
rect 79232 2252 79284 2261
rect 80520 2295 80572 2304
rect 80520 2261 80529 2295
rect 80529 2261 80563 2295
rect 80563 2261 80572 2295
rect 80520 2252 80572 2261
rect 81808 2295 81860 2304
rect 81808 2261 81817 2295
rect 81817 2261 81851 2295
rect 81851 2261 81860 2295
rect 81808 2252 81860 2261
rect 83096 2295 83148 2304
rect 83096 2261 83105 2295
rect 83105 2261 83139 2295
rect 83139 2261 83148 2295
rect 83096 2252 83148 2261
rect 83740 2295 83792 2304
rect 83740 2261 83749 2295
rect 83749 2261 83783 2295
rect 83783 2261 83792 2295
rect 83740 2252 83792 2261
rect 85028 2295 85080 2304
rect 85028 2261 85037 2295
rect 85037 2261 85071 2295
rect 85071 2261 85080 2295
rect 85028 2252 85080 2261
rect 86316 2295 86368 2304
rect 86316 2261 86325 2295
rect 86325 2261 86359 2295
rect 86359 2261 86368 2295
rect 86316 2252 86368 2261
rect 86960 2295 87012 2304
rect 86960 2261 86969 2295
rect 86969 2261 87003 2295
rect 87003 2261 87012 2295
rect 86960 2252 87012 2261
rect 88248 2252 88300 2304
rect 89536 2388 89588 2440
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
rect 35594 2150 35646 2202
rect 35658 2150 35710 2202
rect 35722 2150 35774 2202
rect 35786 2150 35838 2202
rect 35850 2150 35902 2202
rect 66314 2150 66366 2202
rect 66378 2150 66430 2202
rect 66442 2150 66494 2202
rect 66506 2150 66558 2202
rect 66570 2150 66622 2202
rect 97034 2150 97086 2202
rect 97098 2150 97150 2202
rect 97162 2150 97214 2202
rect 97226 2150 97278 2202
rect 97290 2150 97342 2202
<< metal2 >>
rect 14186 97322 14242 98000
rect 15474 97322 15530 98000
rect 16762 97322 16818 98000
rect 17406 97322 17462 98000
rect 18694 97322 18750 98000
rect 19982 97322 20038 98000
rect 21270 97322 21326 98000
rect 21914 97322 21970 98000
rect 23202 97322 23258 98000
rect 24490 97322 24546 98000
rect 25134 97322 25190 98000
rect 26422 97322 26478 98000
rect 27710 97322 27766 98000
rect 14108 97294 14242 97322
rect 4874 95772 5182 95781
rect 4874 95770 4880 95772
rect 4936 95770 4960 95772
rect 5016 95770 5040 95772
rect 5096 95770 5120 95772
rect 5176 95770 5182 95772
rect 4936 95718 4938 95770
rect 5118 95718 5120 95770
rect 4874 95716 4880 95718
rect 4936 95716 4960 95718
rect 5016 95716 5040 95718
rect 5096 95716 5120 95718
rect 5176 95716 5182 95718
rect 4874 95707 5182 95716
rect 14108 95674 14136 97294
rect 14186 97200 14242 97294
rect 15396 97294 15530 97322
rect 15396 95674 15424 97294
rect 15474 97200 15530 97294
rect 16684 97294 16818 97322
rect 16684 95674 16712 97294
rect 16762 97200 16818 97294
rect 17328 97294 17462 97322
rect 17328 95674 17356 97294
rect 17406 97200 17462 97294
rect 18616 97294 18750 97322
rect 18616 95674 18644 97294
rect 18694 97200 18750 97294
rect 19904 97294 20038 97322
rect 19904 95674 19932 97294
rect 19982 97200 20038 97294
rect 21192 97294 21326 97322
rect 21192 95674 21220 97294
rect 21270 97200 21326 97294
rect 21836 97294 21970 97322
rect 21836 95674 21864 97294
rect 21914 97200 21970 97294
rect 23124 97294 23258 97322
rect 23124 95674 23152 97294
rect 23202 97200 23258 97294
rect 24412 97294 24546 97322
rect 14096 95668 14148 95674
rect 14096 95610 14148 95616
rect 15384 95668 15436 95674
rect 15384 95610 15436 95616
rect 16672 95668 16724 95674
rect 16672 95610 16724 95616
rect 17316 95668 17368 95674
rect 17316 95610 17368 95616
rect 18604 95668 18656 95674
rect 18604 95610 18656 95616
rect 19892 95668 19944 95674
rect 19892 95610 19944 95616
rect 21180 95668 21232 95674
rect 21180 95610 21232 95616
rect 21824 95668 21876 95674
rect 21824 95610 21876 95616
rect 23112 95668 23164 95674
rect 23112 95610 23164 95616
rect 18788 95396 18840 95402
rect 18788 95338 18840 95344
rect 20076 95396 20128 95402
rect 20076 95338 20128 95344
rect 20996 95396 21048 95402
rect 20996 95338 21048 95344
rect 23296 95396 23348 95402
rect 23296 95338 23348 95344
rect 14464 95328 14516 95334
rect 14464 95270 14516 95276
rect 15752 95328 15804 95334
rect 15752 95270 15804 95276
rect 16580 95328 16632 95334
rect 16580 95270 16632 95276
rect 17684 95328 17736 95334
rect 17684 95270 17736 95276
rect 4214 95228 4522 95237
rect 4214 95226 4220 95228
rect 4276 95226 4300 95228
rect 4356 95226 4380 95228
rect 4436 95226 4460 95228
rect 4516 95226 4522 95228
rect 4276 95174 4278 95226
rect 4458 95174 4460 95226
rect 4214 95172 4220 95174
rect 4276 95172 4300 95174
rect 4356 95172 4380 95174
rect 4436 95172 4460 95174
rect 4516 95172 4522 95174
rect 4214 95163 4522 95172
rect 4874 94684 5182 94693
rect 4874 94682 4880 94684
rect 4936 94682 4960 94684
rect 5016 94682 5040 94684
rect 5096 94682 5120 94684
rect 5176 94682 5182 94684
rect 4936 94630 4938 94682
rect 5118 94630 5120 94682
rect 4874 94628 4880 94630
rect 4936 94628 4960 94630
rect 5016 94628 5040 94630
rect 5096 94628 5120 94630
rect 5176 94628 5182 94630
rect 4874 94619 5182 94628
rect 4214 94140 4522 94149
rect 4214 94138 4220 94140
rect 4276 94138 4300 94140
rect 4356 94138 4380 94140
rect 4436 94138 4460 94140
rect 4516 94138 4522 94140
rect 4276 94086 4278 94138
rect 4458 94086 4460 94138
rect 4214 94084 4220 94086
rect 4276 94084 4300 94086
rect 4356 94084 4380 94086
rect 4436 94084 4460 94086
rect 4516 94084 4522 94086
rect 4214 94075 4522 94084
rect 4874 93596 5182 93605
rect 4874 93594 4880 93596
rect 4936 93594 4960 93596
rect 5016 93594 5040 93596
rect 5096 93594 5120 93596
rect 5176 93594 5182 93596
rect 4936 93542 4938 93594
rect 5118 93542 5120 93594
rect 4874 93540 4880 93542
rect 4936 93540 4960 93542
rect 5016 93540 5040 93542
rect 5096 93540 5120 93542
rect 5176 93540 5182 93542
rect 4874 93531 5182 93540
rect 5540 93220 5592 93226
rect 5540 93162 5592 93168
rect 4214 93052 4522 93061
rect 4214 93050 4220 93052
rect 4276 93050 4300 93052
rect 4356 93050 4380 93052
rect 4436 93050 4460 93052
rect 4516 93050 4522 93052
rect 4276 92998 4278 93050
rect 4458 92998 4460 93050
rect 4214 92996 4220 92998
rect 4276 92996 4300 92998
rect 4356 92996 4380 92998
rect 4436 92996 4460 92998
rect 4516 92996 4522 92998
rect 4214 92987 4522 92996
rect 4874 92508 5182 92517
rect 4874 92506 4880 92508
rect 4936 92506 4960 92508
rect 5016 92506 5040 92508
rect 5096 92506 5120 92508
rect 5176 92506 5182 92508
rect 4936 92454 4938 92506
rect 5118 92454 5120 92506
rect 4874 92452 4880 92454
rect 4936 92452 4960 92454
rect 5016 92452 5040 92454
rect 5096 92452 5120 92454
rect 5176 92452 5182 92454
rect 4874 92443 5182 92452
rect 4214 91964 4522 91973
rect 4214 91962 4220 91964
rect 4276 91962 4300 91964
rect 4356 91962 4380 91964
rect 4436 91962 4460 91964
rect 4516 91962 4522 91964
rect 4276 91910 4278 91962
rect 4458 91910 4460 91962
rect 4214 91908 4220 91910
rect 4276 91908 4300 91910
rect 4356 91908 4380 91910
rect 4436 91908 4460 91910
rect 4516 91908 4522 91910
rect 4214 91899 4522 91908
rect 4874 91420 5182 91429
rect 4874 91418 4880 91420
rect 4936 91418 4960 91420
rect 5016 91418 5040 91420
rect 5096 91418 5120 91420
rect 5176 91418 5182 91420
rect 4936 91366 4938 91418
rect 5118 91366 5120 91418
rect 4874 91364 4880 91366
rect 4936 91364 4960 91366
rect 5016 91364 5040 91366
rect 5096 91364 5120 91366
rect 5176 91364 5182 91366
rect 4874 91355 5182 91364
rect 4214 90876 4522 90885
rect 4214 90874 4220 90876
rect 4276 90874 4300 90876
rect 4356 90874 4380 90876
rect 4436 90874 4460 90876
rect 4516 90874 4522 90876
rect 4276 90822 4278 90874
rect 4458 90822 4460 90874
rect 4214 90820 4220 90822
rect 4276 90820 4300 90822
rect 4356 90820 4380 90822
rect 4436 90820 4460 90822
rect 4516 90820 4522 90822
rect 4214 90811 4522 90820
rect 4874 90332 5182 90341
rect 4874 90330 4880 90332
rect 4936 90330 4960 90332
rect 5016 90330 5040 90332
rect 5096 90330 5120 90332
rect 5176 90330 5182 90332
rect 4936 90278 4938 90330
rect 5118 90278 5120 90330
rect 4874 90276 4880 90278
rect 4936 90276 4960 90278
rect 5016 90276 5040 90278
rect 5096 90276 5120 90278
rect 5176 90276 5182 90278
rect 4874 90267 5182 90276
rect 4214 89788 4522 89797
rect 4214 89786 4220 89788
rect 4276 89786 4300 89788
rect 4356 89786 4380 89788
rect 4436 89786 4460 89788
rect 4516 89786 4522 89788
rect 4276 89734 4278 89786
rect 4458 89734 4460 89786
rect 4214 89732 4220 89734
rect 4276 89732 4300 89734
rect 4356 89732 4380 89734
rect 4436 89732 4460 89734
rect 4516 89732 4522 89734
rect 4214 89723 4522 89732
rect 4874 89244 5182 89253
rect 4874 89242 4880 89244
rect 4936 89242 4960 89244
rect 5016 89242 5040 89244
rect 5096 89242 5120 89244
rect 5176 89242 5182 89244
rect 4936 89190 4938 89242
rect 5118 89190 5120 89242
rect 4874 89188 4880 89190
rect 4936 89188 4960 89190
rect 5016 89188 5040 89190
rect 5096 89188 5120 89190
rect 5176 89188 5182 89190
rect 4874 89179 5182 89188
rect 4214 88700 4522 88709
rect 4214 88698 4220 88700
rect 4276 88698 4300 88700
rect 4356 88698 4380 88700
rect 4436 88698 4460 88700
rect 4516 88698 4522 88700
rect 4276 88646 4278 88698
rect 4458 88646 4460 88698
rect 4214 88644 4220 88646
rect 4276 88644 4300 88646
rect 4356 88644 4380 88646
rect 4436 88644 4460 88646
rect 4516 88644 4522 88646
rect 4214 88635 4522 88644
rect 4874 88156 5182 88165
rect 4874 88154 4880 88156
rect 4936 88154 4960 88156
rect 5016 88154 5040 88156
rect 5096 88154 5120 88156
rect 5176 88154 5182 88156
rect 4936 88102 4938 88154
rect 5118 88102 5120 88154
rect 4874 88100 4880 88102
rect 4936 88100 4960 88102
rect 5016 88100 5040 88102
rect 5096 88100 5120 88102
rect 5176 88100 5182 88102
rect 4874 88091 5182 88100
rect 4214 87612 4522 87621
rect 4214 87610 4220 87612
rect 4276 87610 4300 87612
rect 4356 87610 4380 87612
rect 4436 87610 4460 87612
rect 4516 87610 4522 87612
rect 4276 87558 4278 87610
rect 4458 87558 4460 87610
rect 4214 87556 4220 87558
rect 4276 87556 4300 87558
rect 4356 87556 4380 87558
rect 4436 87556 4460 87558
rect 4516 87556 4522 87558
rect 4214 87547 4522 87556
rect 846 87272 902 87281
rect 846 87207 902 87216
rect 860 87174 888 87207
rect 848 87168 900 87174
rect 848 87110 900 87116
rect 4874 87068 5182 87077
rect 4874 87066 4880 87068
rect 4936 87066 4960 87068
rect 5016 87066 5040 87068
rect 5096 87066 5120 87068
rect 5176 87066 5182 87068
rect 4936 87014 4938 87066
rect 5118 87014 5120 87066
rect 4874 87012 4880 87014
rect 4936 87012 4960 87014
rect 5016 87012 5040 87014
rect 5096 87012 5120 87014
rect 5176 87012 5182 87014
rect 4874 87003 5182 87012
rect 848 86624 900 86630
rect 846 86592 848 86601
rect 900 86592 902 86601
rect 846 86527 902 86536
rect 4214 86524 4522 86533
rect 4214 86522 4220 86524
rect 4276 86522 4300 86524
rect 4356 86522 4380 86524
rect 4436 86522 4460 86524
rect 4516 86522 4522 86524
rect 4276 86470 4278 86522
rect 4458 86470 4460 86522
rect 4214 86468 4220 86470
rect 4276 86468 4300 86470
rect 4356 86468 4380 86470
rect 4436 86468 4460 86470
rect 4516 86468 4522 86470
rect 4214 86459 4522 86468
rect 4874 85980 5182 85989
rect 4874 85978 4880 85980
rect 4936 85978 4960 85980
rect 5016 85978 5040 85980
rect 5096 85978 5120 85980
rect 5176 85978 5182 85980
rect 4936 85926 4938 85978
rect 5118 85926 5120 85978
rect 4874 85924 4880 85926
rect 4936 85924 4960 85926
rect 5016 85924 5040 85926
rect 5096 85924 5120 85926
rect 5176 85924 5182 85926
rect 4874 85915 5182 85924
rect 4214 85436 4522 85445
rect 4214 85434 4220 85436
rect 4276 85434 4300 85436
rect 4356 85434 4380 85436
rect 4436 85434 4460 85436
rect 4516 85434 4522 85436
rect 4276 85382 4278 85434
rect 4458 85382 4460 85434
rect 4214 85380 4220 85382
rect 4276 85380 4300 85382
rect 4356 85380 4380 85382
rect 4436 85380 4460 85382
rect 4516 85380 4522 85382
rect 4214 85371 4522 85380
rect 848 84992 900 84998
rect 846 84960 848 84969
rect 900 84960 902 84969
rect 846 84895 902 84904
rect 4874 84892 5182 84901
rect 4874 84890 4880 84892
rect 4936 84890 4960 84892
rect 5016 84890 5040 84892
rect 5096 84890 5120 84892
rect 5176 84890 5182 84892
rect 4936 84838 4938 84890
rect 5118 84838 5120 84890
rect 4874 84836 4880 84838
rect 4936 84836 4960 84838
rect 5016 84836 5040 84838
rect 5096 84836 5120 84838
rect 5176 84836 5182 84838
rect 4874 84827 5182 84836
rect 1676 84652 1728 84658
rect 1676 84594 1728 84600
rect 846 84552 902 84561
rect 846 84487 848 84496
rect 900 84487 902 84496
rect 848 84458 900 84464
rect 1688 84153 1716 84594
rect 4214 84348 4522 84357
rect 4214 84346 4220 84348
rect 4276 84346 4300 84348
rect 4356 84346 4380 84348
rect 4436 84346 4460 84348
rect 4516 84346 4522 84348
rect 4276 84294 4278 84346
rect 4458 84294 4460 84346
rect 4214 84292 4220 84294
rect 4276 84292 4300 84294
rect 4356 84292 4380 84294
rect 4436 84292 4460 84294
rect 4516 84292 4522 84294
rect 4214 84283 4522 84292
rect 1674 84144 1730 84153
rect 1674 84079 1730 84088
rect 4874 83804 5182 83813
rect 4874 83802 4880 83804
rect 4936 83802 4960 83804
rect 5016 83802 5040 83804
rect 5096 83802 5120 83804
rect 5176 83802 5182 83804
rect 4936 83750 4938 83802
rect 5118 83750 5120 83802
rect 4874 83748 4880 83750
rect 4936 83748 4960 83750
rect 5016 83748 5040 83750
rect 5096 83748 5120 83750
rect 5176 83748 5182 83750
rect 4874 83739 5182 83748
rect 848 83360 900 83366
rect 848 83302 900 83308
rect 860 83201 888 83302
rect 4214 83260 4522 83269
rect 4214 83258 4220 83260
rect 4276 83258 4300 83260
rect 4356 83258 4380 83260
rect 4436 83258 4460 83260
rect 4516 83258 4522 83260
rect 4276 83206 4278 83258
rect 4458 83206 4460 83258
rect 4214 83204 4220 83206
rect 4276 83204 4300 83206
rect 4356 83204 4380 83206
rect 4436 83204 4460 83206
rect 4516 83204 4522 83206
rect 846 83192 902 83201
rect 4214 83195 4522 83204
rect 846 83127 902 83136
rect 4874 82716 5182 82725
rect 4874 82714 4880 82716
rect 4936 82714 4960 82716
rect 5016 82714 5040 82716
rect 5096 82714 5120 82716
rect 5176 82714 5182 82716
rect 4936 82662 4938 82714
rect 5118 82662 5120 82714
rect 4874 82660 4880 82662
rect 4936 82660 4960 82662
rect 5016 82660 5040 82662
rect 5096 82660 5120 82662
rect 5176 82660 5182 82662
rect 4874 82651 5182 82660
rect 4214 82172 4522 82181
rect 4214 82170 4220 82172
rect 4276 82170 4300 82172
rect 4356 82170 4380 82172
rect 4436 82170 4460 82172
rect 4516 82170 4522 82172
rect 4276 82118 4278 82170
rect 4458 82118 4460 82170
rect 4214 82116 4220 82118
rect 4276 82116 4300 82118
rect 4356 82116 4380 82118
rect 4436 82116 4460 82118
rect 4516 82116 4522 82118
rect 4214 82107 4522 82116
rect 846 81832 902 81841
rect 846 81767 902 81776
rect 860 81734 888 81767
rect 848 81728 900 81734
rect 848 81670 900 81676
rect 4874 81628 5182 81637
rect 4874 81626 4880 81628
rect 4936 81626 4960 81628
rect 5016 81626 5040 81628
rect 5096 81626 5120 81628
rect 5176 81626 5182 81628
rect 4936 81574 4938 81626
rect 5118 81574 5120 81626
rect 4874 81572 4880 81574
rect 4936 81572 4960 81574
rect 5016 81572 5040 81574
rect 5096 81572 5120 81574
rect 5176 81572 5182 81574
rect 4874 81563 5182 81572
rect 848 81184 900 81190
rect 846 81152 848 81161
rect 900 81152 902 81161
rect 846 81087 902 81096
rect 4214 81084 4522 81093
rect 4214 81082 4220 81084
rect 4276 81082 4300 81084
rect 4356 81082 4380 81084
rect 4436 81082 4460 81084
rect 4516 81082 4522 81084
rect 4276 81030 4278 81082
rect 4458 81030 4460 81082
rect 4214 81028 4220 81030
rect 4276 81028 4300 81030
rect 4356 81028 4380 81030
rect 4436 81028 4460 81030
rect 4516 81028 4522 81030
rect 4214 81019 4522 81028
rect 4874 80540 5182 80549
rect 4874 80538 4880 80540
rect 4936 80538 4960 80540
rect 5016 80538 5040 80540
rect 5096 80538 5120 80540
rect 5176 80538 5182 80540
rect 4936 80486 4938 80538
rect 5118 80486 5120 80538
rect 4874 80484 4880 80486
rect 4936 80484 4960 80486
rect 5016 80484 5040 80486
rect 5096 80484 5120 80486
rect 5176 80484 5182 80486
rect 4874 80475 5182 80484
rect 4214 79996 4522 80005
rect 4214 79994 4220 79996
rect 4276 79994 4300 79996
rect 4356 79994 4380 79996
rect 4436 79994 4460 79996
rect 4516 79994 4522 79996
rect 4276 79942 4278 79994
rect 4458 79942 4460 79994
rect 4214 79940 4220 79942
rect 4276 79940 4300 79942
rect 4356 79940 4380 79942
rect 4436 79940 4460 79942
rect 4516 79940 4522 79942
rect 4214 79931 4522 79940
rect 848 79552 900 79558
rect 846 79520 848 79529
rect 900 79520 902 79529
rect 846 79455 902 79464
rect 4874 79452 5182 79461
rect 4874 79450 4880 79452
rect 4936 79450 4960 79452
rect 5016 79450 5040 79452
rect 5096 79450 5120 79452
rect 5176 79450 5182 79452
rect 4936 79398 4938 79450
rect 5118 79398 5120 79450
rect 4874 79396 4880 79398
rect 4936 79396 4960 79398
rect 5016 79396 5040 79398
rect 5096 79396 5120 79398
rect 5176 79396 5182 79398
rect 4874 79387 5182 79396
rect 846 79112 902 79121
rect 846 79047 848 79056
rect 900 79047 902 79056
rect 848 79018 900 79024
rect 4214 78908 4522 78917
rect 4214 78906 4220 78908
rect 4276 78906 4300 78908
rect 4356 78906 4380 78908
rect 4436 78906 4460 78908
rect 4516 78906 4522 78908
rect 4276 78854 4278 78906
rect 4458 78854 4460 78906
rect 4214 78852 4220 78854
rect 4276 78852 4300 78854
rect 4356 78852 4380 78854
rect 4436 78852 4460 78854
rect 4516 78852 4522 78854
rect 4214 78843 4522 78852
rect 4874 78364 5182 78373
rect 4874 78362 4880 78364
rect 4936 78362 4960 78364
rect 5016 78362 5040 78364
rect 5096 78362 5120 78364
rect 5176 78362 5182 78364
rect 4936 78310 4938 78362
rect 5118 78310 5120 78362
rect 4874 78308 4880 78310
rect 4936 78308 4960 78310
rect 5016 78308 5040 78310
rect 5096 78308 5120 78310
rect 5176 78308 5182 78310
rect 4874 78299 5182 78308
rect 848 77920 900 77926
rect 848 77862 900 77868
rect 860 77761 888 77862
rect 4214 77820 4522 77829
rect 4214 77818 4220 77820
rect 4276 77818 4300 77820
rect 4356 77818 4380 77820
rect 4436 77818 4460 77820
rect 4516 77818 4522 77820
rect 4276 77766 4278 77818
rect 4458 77766 4460 77818
rect 4214 77764 4220 77766
rect 4276 77764 4300 77766
rect 4356 77764 4380 77766
rect 4436 77764 4460 77766
rect 4516 77764 4522 77766
rect 846 77752 902 77761
rect 4214 77755 4522 77764
rect 846 77687 902 77696
rect 4874 77276 5182 77285
rect 4874 77274 4880 77276
rect 4936 77274 4960 77276
rect 5016 77274 5040 77276
rect 5096 77274 5120 77276
rect 5176 77274 5182 77276
rect 4936 77222 4938 77274
rect 5118 77222 5120 77274
rect 4874 77220 4880 77222
rect 4936 77220 4960 77222
rect 5016 77220 5040 77222
rect 5096 77220 5120 77222
rect 5176 77220 5182 77222
rect 4874 77211 5182 77220
rect 4214 76732 4522 76741
rect 4214 76730 4220 76732
rect 4276 76730 4300 76732
rect 4356 76730 4380 76732
rect 4436 76730 4460 76732
rect 4516 76730 4522 76732
rect 4276 76678 4278 76730
rect 4458 76678 4460 76730
rect 4214 76676 4220 76678
rect 4276 76676 4300 76678
rect 4356 76676 4380 76678
rect 4436 76676 4460 76678
rect 4516 76676 4522 76678
rect 4214 76667 4522 76676
rect 846 76392 902 76401
rect 846 76327 902 76336
rect 860 76294 888 76327
rect 848 76288 900 76294
rect 848 76230 900 76236
rect 4874 76188 5182 76197
rect 4874 76186 4880 76188
rect 4936 76186 4960 76188
rect 5016 76186 5040 76188
rect 5096 76186 5120 76188
rect 5176 76186 5182 76188
rect 4936 76134 4938 76186
rect 5118 76134 5120 76186
rect 4874 76132 4880 76134
rect 4936 76132 4960 76134
rect 5016 76132 5040 76134
rect 5096 76132 5120 76134
rect 5176 76132 5182 76134
rect 4874 76123 5182 76132
rect 848 76084 900 76090
rect 848 76026 900 76032
rect 860 75721 888 76026
rect 1676 75948 1728 75954
rect 1676 75890 1728 75896
rect 846 75712 902 75721
rect 846 75647 902 75656
rect 1688 75449 1716 75890
rect 4214 75644 4522 75653
rect 4214 75642 4220 75644
rect 4276 75642 4300 75644
rect 4356 75642 4380 75644
rect 4436 75642 4460 75644
rect 4516 75642 4522 75644
rect 4276 75590 4278 75642
rect 4458 75590 4460 75642
rect 4214 75588 4220 75590
rect 4276 75588 4300 75590
rect 4356 75588 4380 75590
rect 4436 75588 4460 75590
rect 4516 75588 4522 75590
rect 4214 75579 4522 75588
rect 1674 75440 1730 75449
rect 1674 75375 1730 75384
rect 4874 75100 5182 75109
rect 4874 75098 4880 75100
rect 4936 75098 4960 75100
rect 5016 75098 5040 75100
rect 5096 75098 5120 75100
rect 5176 75098 5182 75100
rect 4936 75046 4938 75098
rect 5118 75046 5120 75098
rect 4874 75044 4880 75046
rect 4936 75044 4960 75046
rect 5016 75044 5040 75046
rect 5096 75044 5120 75046
rect 5176 75044 5182 75046
rect 4874 75035 5182 75044
rect 4214 74556 4522 74565
rect 4214 74554 4220 74556
rect 4276 74554 4300 74556
rect 4356 74554 4380 74556
rect 4436 74554 4460 74556
rect 4516 74554 4522 74556
rect 4276 74502 4278 74554
rect 4458 74502 4460 74554
rect 4214 74500 4220 74502
rect 4276 74500 4300 74502
rect 4356 74500 4380 74502
rect 4436 74500 4460 74502
rect 4516 74500 4522 74502
rect 4214 74491 4522 74500
rect 848 74112 900 74118
rect 846 74080 848 74089
rect 900 74080 902 74089
rect 846 74015 902 74024
rect 4874 74012 5182 74021
rect 4874 74010 4880 74012
rect 4936 74010 4960 74012
rect 5016 74010 5040 74012
rect 5096 74010 5120 74012
rect 5176 74010 5182 74012
rect 4936 73958 4938 74010
rect 5118 73958 5120 74010
rect 4874 73956 4880 73958
rect 4936 73956 4960 73958
rect 5016 73956 5040 73958
rect 5096 73956 5120 73958
rect 5176 73956 5182 73958
rect 4874 73947 5182 73956
rect 846 73672 902 73681
rect 846 73607 848 73616
rect 900 73607 902 73616
rect 848 73578 900 73584
rect 4214 73468 4522 73477
rect 4214 73466 4220 73468
rect 4276 73466 4300 73468
rect 4356 73466 4380 73468
rect 4436 73466 4460 73468
rect 4516 73466 4522 73468
rect 4276 73414 4278 73466
rect 4458 73414 4460 73466
rect 4214 73412 4220 73414
rect 4276 73412 4300 73414
rect 4356 73412 4380 73414
rect 4436 73412 4460 73414
rect 4516 73412 4522 73414
rect 4214 73403 4522 73412
rect 4874 72924 5182 72933
rect 4874 72922 4880 72924
rect 4936 72922 4960 72924
rect 5016 72922 5040 72924
rect 5096 72922 5120 72924
rect 5176 72922 5182 72924
rect 4936 72870 4938 72922
rect 5118 72870 5120 72922
rect 4874 72868 4880 72870
rect 4936 72868 4960 72870
rect 5016 72868 5040 72870
rect 5096 72868 5120 72870
rect 5176 72868 5182 72870
rect 4874 72859 5182 72868
rect 848 72480 900 72486
rect 848 72422 900 72428
rect 860 72321 888 72422
rect 4214 72380 4522 72389
rect 4214 72378 4220 72380
rect 4276 72378 4300 72380
rect 4356 72378 4380 72380
rect 4436 72378 4460 72380
rect 4516 72378 4522 72380
rect 4276 72326 4278 72378
rect 4458 72326 4460 72378
rect 4214 72324 4220 72326
rect 4276 72324 4300 72326
rect 4356 72324 4380 72326
rect 4436 72324 4460 72326
rect 4516 72324 4522 72326
rect 846 72312 902 72321
rect 4214 72315 4522 72324
rect 846 72247 902 72256
rect 4874 71836 5182 71845
rect 4874 71834 4880 71836
rect 4936 71834 4960 71836
rect 5016 71834 5040 71836
rect 5096 71834 5120 71836
rect 5176 71834 5182 71836
rect 4936 71782 4938 71834
rect 5118 71782 5120 71834
rect 4874 71780 4880 71782
rect 4936 71780 4960 71782
rect 5016 71780 5040 71782
rect 5096 71780 5120 71782
rect 5176 71780 5182 71782
rect 4874 71771 5182 71780
rect 4214 71292 4522 71301
rect 4214 71290 4220 71292
rect 4276 71290 4300 71292
rect 4356 71290 4380 71292
rect 4436 71290 4460 71292
rect 4516 71290 4522 71292
rect 4276 71238 4278 71290
rect 4458 71238 4460 71290
rect 4214 71236 4220 71238
rect 4276 71236 4300 71238
rect 4356 71236 4380 71238
rect 4436 71236 4460 71238
rect 4516 71236 4522 71238
rect 4214 71227 4522 71236
rect 846 70952 902 70961
rect 846 70887 902 70896
rect 860 70854 888 70887
rect 848 70848 900 70854
rect 848 70790 900 70796
rect 4874 70748 5182 70757
rect 4874 70746 4880 70748
rect 4936 70746 4960 70748
rect 5016 70746 5040 70748
rect 5096 70746 5120 70748
rect 5176 70746 5182 70748
rect 4936 70694 4938 70746
rect 5118 70694 5120 70746
rect 4874 70692 4880 70694
rect 4936 70692 4960 70694
rect 5016 70692 5040 70694
rect 5096 70692 5120 70694
rect 5176 70692 5182 70694
rect 4874 70683 5182 70692
rect 5552 70650 5580 93162
rect 8944 93152 8996 93158
rect 8944 93094 8996 93100
rect 10048 93152 10100 93158
rect 10048 93094 10100 93100
rect 11152 93152 11204 93158
rect 11152 93094 11204 93100
rect 12256 93152 12308 93158
rect 12256 93094 12308 93100
rect 13268 93152 13320 93158
rect 13268 93094 13320 93100
rect 8956 90930 8984 93094
rect 10060 92886 10088 93094
rect 10048 92880 10100 92886
rect 10048 92822 10100 92828
rect 10060 90930 10088 92822
rect 11164 92750 11192 93094
rect 12268 92818 12296 93094
rect 12256 92812 12308 92818
rect 12256 92754 12308 92760
rect 11152 92744 11204 92750
rect 11152 92686 11204 92692
rect 11164 90930 11192 92686
rect 12268 90930 12296 92754
rect 8496 90902 8984 90930
rect 9982 90902 10088 90930
rect 11086 90902 11192 90930
rect 12190 90902 12296 90930
rect 5724 90500 5776 90506
rect 5724 90442 5776 90448
rect 5632 90160 5684 90166
rect 5632 90102 5684 90108
rect 5540 70644 5592 70650
rect 5540 70586 5592 70592
rect 1308 70508 1360 70514
rect 1308 70450 1360 70456
rect 1320 70145 1348 70450
rect 1584 70304 1636 70310
rect 1584 70246 1636 70252
rect 1306 70136 1362 70145
rect 1306 70071 1362 70080
rect 1596 70009 1624 70246
rect 4214 70204 4522 70213
rect 4214 70202 4220 70204
rect 4276 70202 4300 70204
rect 4356 70202 4380 70204
rect 4436 70202 4460 70204
rect 4516 70202 4522 70204
rect 4276 70150 4278 70202
rect 4458 70150 4460 70202
rect 4214 70148 4220 70150
rect 4276 70148 4300 70150
rect 4356 70148 4380 70150
rect 4436 70148 4460 70150
rect 4516 70148 4522 70150
rect 4214 70139 4522 70148
rect 1582 70000 1638 70009
rect 1582 69935 1638 69944
rect 5552 69902 5580 70586
rect 5540 69896 5592 69902
rect 5540 69838 5592 69844
rect 5644 69766 5672 90102
rect 5632 69760 5684 69766
rect 5632 69702 5684 69708
rect 4874 69660 5182 69669
rect 4874 69658 4880 69660
rect 4936 69658 4960 69660
rect 5016 69658 5040 69660
rect 5096 69658 5120 69660
rect 5176 69658 5182 69660
rect 4936 69606 4938 69658
rect 5118 69606 5120 69658
rect 4874 69604 4880 69606
rect 4936 69604 4960 69606
rect 5016 69604 5040 69606
rect 5096 69604 5120 69606
rect 5176 69604 5182 69606
rect 4874 69595 5182 69604
rect 5644 69562 5672 69702
rect 5632 69556 5684 69562
rect 5632 69498 5684 69504
rect 4214 69116 4522 69125
rect 4214 69114 4220 69116
rect 4276 69114 4300 69116
rect 4356 69114 4380 69116
rect 4436 69114 4460 69116
rect 4516 69114 4522 69116
rect 4276 69062 4278 69114
rect 4458 69062 4460 69114
rect 4214 69060 4220 69062
rect 4276 69060 4300 69062
rect 4356 69060 4380 69062
rect 4436 69060 4460 69062
rect 4516 69060 4522 69062
rect 4214 69051 4522 69060
rect 1122 68776 1178 68785
rect 1122 68711 1124 68720
rect 1176 68711 1178 68720
rect 1124 68682 1176 68688
rect 4874 68572 5182 68581
rect 4874 68570 4880 68572
rect 4936 68570 4960 68572
rect 5016 68570 5040 68572
rect 5096 68570 5120 68572
rect 5176 68570 5182 68572
rect 4936 68518 4938 68570
rect 5118 68518 5120 68570
rect 4874 68516 4880 68518
rect 4936 68516 4960 68518
rect 5016 68516 5040 68518
rect 5096 68516 5120 68518
rect 5176 68516 5182 68518
rect 4874 68507 5182 68516
rect 1308 68332 1360 68338
rect 1308 68274 1360 68280
rect 1320 68105 1348 68274
rect 1306 68096 1362 68105
rect 1306 68031 1362 68040
rect 4214 68028 4522 68037
rect 4214 68026 4220 68028
rect 4276 68026 4300 68028
rect 4356 68026 4380 68028
rect 4436 68026 4460 68028
rect 4516 68026 4522 68028
rect 4276 67974 4278 68026
rect 4458 67974 4460 68026
rect 4214 67972 4220 67974
rect 4276 67972 4300 67974
rect 4356 67972 4380 67974
rect 4436 67972 4460 67974
rect 4516 67972 4522 67974
rect 4214 67963 4522 67972
rect 4874 67484 5182 67493
rect 4874 67482 4880 67484
rect 4936 67482 4960 67484
rect 5016 67482 5040 67484
rect 5096 67482 5120 67484
rect 5176 67482 5182 67484
rect 4936 67430 4938 67482
rect 5118 67430 5120 67482
rect 4874 67428 4880 67430
rect 4936 67428 4960 67430
rect 5016 67428 5040 67430
rect 5096 67428 5120 67430
rect 5176 67428 5182 67430
rect 4874 67419 5182 67428
rect 1308 67244 1360 67250
rect 1308 67186 1360 67192
rect 1320 66745 1348 67186
rect 4214 66940 4522 66949
rect 4214 66938 4220 66940
rect 4276 66938 4300 66940
rect 4356 66938 4380 66940
rect 4436 66938 4460 66940
rect 4516 66938 4522 66940
rect 4276 66886 4278 66938
rect 4458 66886 4460 66938
rect 4214 66884 4220 66886
rect 4276 66884 4300 66886
rect 4356 66884 4380 66886
rect 4436 66884 4460 66886
rect 4516 66884 4522 66886
rect 4214 66875 4522 66884
rect 1306 66736 1362 66745
rect 1306 66671 1362 66680
rect 4874 66396 5182 66405
rect 4874 66394 4880 66396
rect 4936 66394 4960 66396
rect 5016 66394 5040 66396
rect 5096 66394 5120 66396
rect 5176 66394 5182 66396
rect 4936 66342 4938 66394
rect 5118 66342 5120 66394
rect 4874 66340 4880 66342
rect 4936 66340 4960 66342
rect 5016 66340 5040 66342
rect 5096 66340 5120 66342
rect 5176 66340 5182 66342
rect 4874 66331 5182 66340
rect 4214 65852 4522 65861
rect 4214 65850 4220 65852
rect 4276 65850 4300 65852
rect 4356 65850 4380 65852
rect 4436 65850 4460 65852
rect 4516 65850 4522 65852
rect 4276 65798 4278 65850
rect 4458 65798 4460 65850
rect 4214 65796 4220 65798
rect 4276 65796 4300 65798
rect 4356 65796 4380 65798
rect 4436 65796 4460 65798
rect 4516 65796 4522 65798
rect 4214 65787 4522 65796
rect 1124 65476 1176 65482
rect 1124 65418 1176 65424
rect 1136 65385 1164 65418
rect 1122 65376 1178 65385
rect 1122 65311 1178 65320
rect 4874 65308 5182 65317
rect 4874 65306 4880 65308
rect 4936 65306 4960 65308
rect 5016 65306 5040 65308
rect 5096 65306 5120 65308
rect 5176 65306 5182 65308
rect 4936 65254 4938 65306
rect 5118 65254 5120 65306
rect 4874 65252 4880 65254
rect 4936 65252 4960 65254
rect 5016 65252 5040 65254
rect 5096 65252 5120 65254
rect 5176 65252 5182 65254
rect 4874 65243 5182 65252
rect 1308 65068 1360 65074
rect 1308 65010 1360 65016
rect 1320 64705 1348 65010
rect 1676 64932 1728 64938
rect 1676 64874 1728 64880
rect 5644 64874 5672 69498
rect 1306 64696 1362 64705
rect 1306 64631 1362 64640
rect 1688 64569 1716 64874
rect 5552 64846 5672 64874
rect 4214 64764 4522 64773
rect 4214 64762 4220 64764
rect 4276 64762 4300 64764
rect 4356 64762 4380 64764
rect 4436 64762 4460 64764
rect 4516 64762 4522 64764
rect 4276 64710 4278 64762
rect 4458 64710 4460 64762
rect 4214 64708 4220 64710
rect 4276 64708 4300 64710
rect 4356 64708 4380 64710
rect 4436 64708 4460 64710
rect 4516 64708 4522 64710
rect 4214 64699 4522 64708
rect 1674 64560 1730 64569
rect 1674 64495 1730 64504
rect 4874 64220 5182 64229
rect 4874 64218 4880 64220
rect 4936 64218 4960 64220
rect 5016 64218 5040 64220
rect 5096 64218 5120 64220
rect 5176 64218 5182 64220
rect 4936 64166 4938 64218
rect 5118 64166 5120 64218
rect 4874 64164 4880 64166
rect 4936 64164 4960 64166
rect 5016 64164 5040 64166
rect 5096 64164 5120 64166
rect 5176 64164 5182 64166
rect 4874 64155 5182 64164
rect 4214 63676 4522 63685
rect 4214 63674 4220 63676
rect 4276 63674 4300 63676
rect 4356 63674 4380 63676
rect 4436 63674 4460 63676
rect 4516 63674 4522 63676
rect 4276 63622 4278 63674
rect 4458 63622 4460 63674
rect 4214 63620 4220 63622
rect 4276 63620 4300 63622
rect 4356 63620 4380 63622
rect 4436 63620 4460 63622
rect 4516 63620 4522 63622
rect 4214 63611 4522 63620
rect 1122 63336 1178 63345
rect 1122 63271 1124 63280
rect 1176 63271 1178 63280
rect 1124 63242 1176 63248
rect 4874 63132 5182 63141
rect 4874 63130 4880 63132
rect 4936 63130 4960 63132
rect 5016 63130 5040 63132
rect 5096 63130 5120 63132
rect 5176 63130 5182 63132
rect 4936 63078 4938 63130
rect 5118 63078 5120 63130
rect 4874 63076 4880 63078
rect 4936 63076 4960 63078
rect 5016 63076 5040 63078
rect 5096 63076 5120 63078
rect 5176 63076 5182 63078
rect 4874 63067 5182 63076
rect 1308 62892 1360 62898
rect 1308 62834 1360 62840
rect 1320 62665 1348 62834
rect 1306 62656 1362 62665
rect 1306 62591 1362 62600
rect 4214 62588 4522 62597
rect 4214 62586 4220 62588
rect 4276 62586 4300 62588
rect 4356 62586 4380 62588
rect 4436 62586 4460 62588
rect 4516 62586 4522 62588
rect 4276 62534 4278 62586
rect 4458 62534 4460 62586
rect 4214 62532 4220 62534
rect 4276 62532 4300 62534
rect 4356 62532 4380 62534
rect 4436 62532 4460 62534
rect 4516 62532 4522 62534
rect 4214 62523 4522 62532
rect 4874 62044 5182 62053
rect 4874 62042 4880 62044
rect 4936 62042 4960 62044
rect 5016 62042 5040 62044
rect 5096 62042 5120 62044
rect 5176 62042 5182 62044
rect 4936 61990 4938 62042
rect 5118 61990 5120 62042
rect 4874 61988 4880 61990
rect 4936 61988 4960 61990
rect 5016 61988 5040 61990
rect 5096 61988 5120 61990
rect 5176 61988 5182 61990
rect 4874 61979 5182 61988
rect 1308 61804 1360 61810
rect 1308 61746 1360 61752
rect 1320 61305 1348 61746
rect 4214 61500 4522 61509
rect 4214 61498 4220 61500
rect 4276 61498 4300 61500
rect 4356 61498 4380 61500
rect 4436 61498 4460 61500
rect 4516 61498 4522 61500
rect 4276 61446 4278 61498
rect 4458 61446 4460 61498
rect 4214 61444 4220 61446
rect 4276 61444 4300 61446
rect 4356 61444 4380 61446
rect 4436 61444 4460 61446
rect 4516 61444 4522 61446
rect 4214 61435 4522 61444
rect 1306 61296 1362 61305
rect 1306 61231 1362 61240
rect 4874 60956 5182 60965
rect 4874 60954 4880 60956
rect 4936 60954 4960 60956
rect 5016 60954 5040 60956
rect 5096 60954 5120 60956
rect 5176 60954 5182 60956
rect 4936 60902 4938 60954
rect 5118 60902 5120 60954
rect 4874 60900 4880 60902
rect 4936 60900 4960 60902
rect 5016 60900 5040 60902
rect 5096 60900 5120 60902
rect 5176 60900 5182 60902
rect 4874 60891 5182 60900
rect 4214 60412 4522 60421
rect 4214 60410 4220 60412
rect 4276 60410 4300 60412
rect 4356 60410 4380 60412
rect 4436 60410 4460 60412
rect 4516 60410 4522 60412
rect 4276 60358 4278 60410
rect 4458 60358 4460 60410
rect 4214 60356 4220 60358
rect 4276 60356 4300 60358
rect 4356 60356 4380 60358
rect 4436 60356 4460 60358
rect 4516 60356 4522 60358
rect 4214 60347 4522 60356
rect 1216 60036 1268 60042
rect 1216 59978 1268 59984
rect 1228 59945 1256 59978
rect 1214 59936 1270 59945
rect 1214 59871 1270 59880
rect 4874 59868 5182 59877
rect 4874 59866 4880 59868
rect 4936 59866 4960 59868
rect 5016 59866 5040 59868
rect 5096 59866 5120 59868
rect 5176 59866 5182 59868
rect 4936 59814 4938 59866
rect 5118 59814 5120 59866
rect 4874 59812 4880 59814
rect 4936 59812 4960 59814
rect 5016 59812 5040 59814
rect 5096 59812 5120 59814
rect 5176 59812 5182 59814
rect 4874 59803 5182 59812
rect 1216 59628 1268 59634
rect 1216 59570 1268 59576
rect 1228 59265 1256 59570
rect 1584 59424 1636 59430
rect 1584 59366 1636 59372
rect 1214 59256 1270 59265
rect 1214 59191 1270 59200
rect 1596 59129 1624 59366
rect 4214 59324 4522 59333
rect 4214 59322 4220 59324
rect 4276 59322 4300 59324
rect 4356 59322 4380 59324
rect 4436 59322 4460 59324
rect 4516 59322 4522 59324
rect 4276 59270 4278 59322
rect 4458 59270 4460 59322
rect 4214 59268 4220 59270
rect 4276 59268 4300 59270
rect 4356 59268 4380 59270
rect 4436 59268 4460 59270
rect 4516 59268 4522 59270
rect 4214 59259 4522 59268
rect 1582 59120 1638 59129
rect 1582 59055 1638 59064
rect 4874 58780 5182 58789
rect 4874 58778 4880 58780
rect 4936 58778 4960 58780
rect 5016 58778 5040 58780
rect 5096 58778 5120 58780
rect 5176 58778 5182 58780
rect 4936 58726 4938 58778
rect 5118 58726 5120 58778
rect 4874 58724 4880 58726
rect 4936 58724 4960 58726
rect 5016 58724 5040 58726
rect 5096 58724 5120 58726
rect 5176 58724 5182 58726
rect 4874 58715 5182 58724
rect 4214 58236 4522 58245
rect 4214 58234 4220 58236
rect 4276 58234 4300 58236
rect 4356 58234 4380 58236
rect 4436 58234 4460 58236
rect 4516 58234 4522 58236
rect 4276 58182 4278 58234
rect 4458 58182 4460 58234
rect 4214 58180 4220 58182
rect 4276 58180 4300 58182
rect 4356 58180 4380 58182
rect 4436 58180 4460 58182
rect 4516 58180 4522 58182
rect 4214 58171 4522 58180
rect 1582 58032 1638 58041
rect 1582 57967 1638 57976
rect 1308 57928 1360 57934
rect 1306 57896 1308 57905
rect 1360 57896 1362 57905
rect 1306 57831 1362 57840
rect 1596 57798 1624 57967
rect 1584 57792 1636 57798
rect 1584 57734 1636 57740
rect 4874 57692 5182 57701
rect 4874 57690 4880 57692
rect 4936 57690 4960 57692
rect 5016 57690 5040 57692
rect 5096 57690 5120 57692
rect 5176 57690 5182 57692
rect 4936 57638 4938 57690
rect 5118 57638 5120 57690
rect 4874 57636 4880 57638
rect 4936 57636 4960 57638
rect 5016 57636 5040 57638
rect 5096 57636 5120 57638
rect 5176 57636 5182 57638
rect 4874 57627 5182 57636
rect 1308 57452 1360 57458
rect 1308 57394 1360 57400
rect 1320 57225 1348 57394
rect 1306 57216 1362 57225
rect 1306 57151 1362 57160
rect 4214 57148 4522 57157
rect 4214 57146 4220 57148
rect 4276 57146 4300 57148
rect 4356 57146 4380 57148
rect 4436 57146 4460 57148
rect 4516 57146 4522 57148
rect 4276 57094 4278 57146
rect 4458 57094 4460 57146
rect 4214 57092 4220 57094
rect 4276 57092 4300 57094
rect 4356 57092 4380 57094
rect 4436 57092 4460 57094
rect 4516 57092 4522 57094
rect 4214 57083 4522 57092
rect 4874 56604 5182 56613
rect 4874 56602 4880 56604
rect 4936 56602 4960 56604
rect 5016 56602 5040 56604
rect 5096 56602 5120 56604
rect 5176 56602 5182 56604
rect 4936 56550 4938 56602
rect 5118 56550 5120 56602
rect 4874 56548 4880 56550
rect 4936 56548 4960 56550
rect 5016 56548 5040 56550
rect 5096 56548 5120 56550
rect 5176 56548 5182 56550
rect 4874 56539 5182 56548
rect 1308 56364 1360 56370
rect 1308 56306 1360 56312
rect 1320 55865 1348 56306
rect 4214 56060 4522 56069
rect 4214 56058 4220 56060
rect 4276 56058 4300 56060
rect 4356 56058 4380 56060
rect 4436 56058 4460 56060
rect 4516 56058 4522 56060
rect 4276 56006 4278 56058
rect 4458 56006 4460 56058
rect 4214 56004 4220 56006
rect 4276 56004 4300 56006
rect 4356 56004 4380 56006
rect 4436 56004 4460 56006
rect 4516 56004 4522 56006
rect 4214 55995 4522 56004
rect 1306 55856 1362 55865
rect 1306 55791 1362 55800
rect 4874 55516 5182 55525
rect 4874 55514 4880 55516
rect 4936 55514 4960 55516
rect 5016 55514 5040 55516
rect 5096 55514 5120 55516
rect 5176 55514 5182 55516
rect 4936 55462 4938 55514
rect 5118 55462 5120 55514
rect 4874 55460 4880 55462
rect 4936 55460 4960 55462
rect 5016 55460 5040 55462
rect 5096 55460 5120 55462
rect 5176 55460 5182 55462
rect 4874 55451 5182 55460
rect 4214 54972 4522 54981
rect 4214 54970 4220 54972
rect 4276 54970 4300 54972
rect 4356 54970 4380 54972
rect 4436 54970 4460 54972
rect 4516 54970 4522 54972
rect 4276 54918 4278 54970
rect 4458 54918 4460 54970
rect 4214 54916 4220 54918
rect 4276 54916 4300 54918
rect 4356 54916 4380 54918
rect 4436 54916 4460 54918
rect 4516 54916 4522 54918
rect 4214 54907 4522 54916
rect 1308 54664 1360 54670
rect 1308 54606 1360 54612
rect 1320 54505 1348 54606
rect 1306 54496 1362 54505
rect 1306 54431 1362 54440
rect 4874 54428 5182 54437
rect 4874 54426 4880 54428
rect 4936 54426 4960 54428
rect 5016 54426 5040 54428
rect 5096 54426 5120 54428
rect 5176 54426 5182 54428
rect 4936 54374 4938 54426
rect 5118 54374 5120 54426
rect 4874 54372 4880 54374
rect 4936 54372 4960 54374
rect 5016 54372 5040 54374
rect 5096 54372 5120 54374
rect 5176 54372 5182 54374
rect 4874 54363 5182 54372
rect 1216 54188 1268 54194
rect 1216 54130 1268 54136
rect 1228 53825 1256 54130
rect 1584 53984 1636 53990
rect 1584 53926 1636 53932
rect 1214 53816 1270 53825
rect 1214 53751 1270 53760
rect 1596 53689 1624 53926
rect 4214 53884 4522 53893
rect 4214 53882 4220 53884
rect 4276 53882 4300 53884
rect 4356 53882 4380 53884
rect 4436 53882 4460 53884
rect 4516 53882 4522 53884
rect 4276 53830 4278 53882
rect 4458 53830 4460 53882
rect 4214 53828 4220 53830
rect 4276 53828 4300 53830
rect 4356 53828 4380 53830
rect 4436 53828 4460 53830
rect 4516 53828 4522 53830
rect 4214 53819 4522 53828
rect 1582 53680 1638 53689
rect 1582 53615 1638 53624
rect 4874 53340 5182 53349
rect 4874 53338 4880 53340
rect 4936 53338 4960 53340
rect 5016 53338 5040 53340
rect 5096 53338 5120 53340
rect 5176 53338 5182 53340
rect 4936 53286 4938 53338
rect 5118 53286 5120 53338
rect 4874 53284 4880 53286
rect 4936 53284 4960 53286
rect 5016 53284 5040 53286
rect 5096 53284 5120 53286
rect 5176 53284 5182 53286
rect 4874 53275 5182 53284
rect 4214 52796 4522 52805
rect 4214 52794 4220 52796
rect 4276 52794 4300 52796
rect 4356 52794 4380 52796
rect 4436 52794 4460 52796
rect 4516 52794 4522 52796
rect 4276 52742 4278 52794
rect 4458 52742 4460 52794
rect 4214 52740 4220 52742
rect 4276 52740 4300 52742
rect 4356 52740 4380 52742
rect 4436 52740 4460 52742
rect 4516 52740 4522 52742
rect 4214 52731 4522 52740
rect 4874 52252 5182 52261
rect 4874 52250 4880 52252
rect 4936 52250 4960 52252
rect 5016 52250 5040 52252
rect 5096 52250 5120 52252
rect 5176 52250 5182 52252
rect 4936 52198 4938 52250
rect 5118 52198 5120 52250
rect 4874 52196 4880 52198
rect 4936 52196 4960 52198
rect 5016 52196 5040 52198
rect 5096 52196 5120 52198
rect 5176 52196 5182 52198
rect 4874 52187 5182 52196
rect 4214 51708 4522 51717
rect 4214 51706 4220 51708
rect 4276 51706 4300 51708
rect 4356 51706 4380 51708
rect 4436 51706 4460 51708
rect 4516 51706 4522 51708
rect 4276 51654 4278 51706
rect 4458 51654 4460 51706
rect 4214 51652 4220 51654
rect 4276 51652 4300 51654
rect 4356 51652 4380 51654
rect 4436 51652 4460 51654
rect 4516 51652 4522 51654
rect 4214 51643 4522 51652
rect 4874 51164 5182 51173
rect 4874 51162 4880 51164
rect 4936 51162 4960 51164
rect 5016 51162 5040 51164
rect 5096 51162 5120 51164
rect 5176 51162 5182 51164
rect 4936 51110 4938 51162
rect 5118 51110 5120 51162
rect 4874 51108 4880 51110
rect 4936 51108 4960 51110
rect 5016 51108 5040 51110
rect 5096 51108 5120 51110
rect 5176 51108 5182 51110
rect 4874 51099 5182 51108
rect 4214 50620 4522 50629
rect 4214 50618 4220 50620
rect 4276 50618 4300 50620
rect 4356 50618 4380 50620
rect 4436 50618 4460 50620
rect 4516 50618 4522 50620
rect 4276 50566 4278 50618
rect 4458 50566 4460 50618
rect 4214 50564 4220 50566
rect 4276 50564 4300 50566
rect 4356 50564 4380 50566
rect 4436 50564 4460 50566
rect 4516 50564 4522 50566
rect 4214 50555 4522 50564
rect 4874 50076 5182 50085
rect 4874 50074 4880 50076
rect 4936 50074 4960 50076
rect 5016 50074 5040 50076
rect 5096 50074 5120 50076
rect 5176 50074 5182 50076
rect 4936 50022 4938 50074
rect 5118 50022 5120 50074
rect 4874 50020 4880 50022
rect 4936 50020 4960 50022
rect 5016 50020 5040 50022
rect 5096 50020 5120 50022
rect 5176 50020 5182 50022
rect 4874 50011 5182 50020
rect 4214 49532 4522 49541
rect 4214 49530 4220 49532
rect 4276 49530 4300 49532
rect 4356 49530 4380 49532
rect 4436 49530 4460 49532
rect 4516 49530 4522 49532
rect 4276 49478 4278 49530
rect 4458 49478 4460 49530
rect 4214 49476 4220 49478
rect 4276 49476 4300 49478
rect 4356 49476 4380 49478
rect 4436 49476 4460 49478
rect 4516 49476 4522 49478
rect 4214 49467 4522 49476
rect 4874 48988 5182 48997
rect 4874 48986 4880 48988
rect 4936 48986 4960 48988
rect 5016 48986 5040 48988
rect 5096 48986 5120 48988
rect 5176 48986 5182 48988
rect 4936 48934 4938 48986
rect 5118 48934 5120 48986
rect 4874 48932 4880 48934
rect 4936 48932 4960 48934
rect 5016 48932 5040 48934
rect 5096 48932 5120 48934
rect 5176 48932 5182 48934
rect 4874 48923 5182 48932
rect 5552 48890 5580 64846
rect 5736 51066 5764 90442
rect 8496 90166 8524 90902
rect 13280 90545 13308 93094
rect 14476 90930 14504 95270
rect 15764 90930 15792 95270
rect 14398 90902 14504 90930
rect 15502 90902 15792 90930
rect 16592 90916 16620 95270
rect 17696 90916 17724 95270
rect 18800 90916 18828 95338
rect 20088 90930 20116 95338
rect 19918 90902 20116 90930
rect 21008 90916 21036 95338
rect 22192 95328 22244 95334
rect 22192 95270 22244 95276
rect 22204 90930 22232 95270
rect 23308 90930 23336 95338
rect 24412 95130 24440 97294
rect 24490 97200 24546 97294
rect 25056 97294 25190 97322
rect 25056 95674 25084 97294
rect 25134 97200 25190 97294
rect 26344 97294 26478 97322
rect 26344 95674 26372 97294
rect 26422 97200 26478 97294
rect 27632 97294 27766 97322
rect 27632 95674 27660 97294
rect 27710 97200 27766 97294
rect 28998 97322 29054 98000
rect 29642 97322 29698 98000
rect 30930 97322 30986 98000
rect 28998 97294 29132 97322
rect 28998 97200 29054 97294
rect 29104 95674 29132 97294
rect 29564 97294 29698 97322
rect 29564 95674 29592 97294
rect 29642 97200 29698 97294
rect 30852 97294 30986 97322
rect 30852 95674 30880 97294
rect 30930 97200 30986 97294
rect 32218 97322 32274 98000
rect 32862 97322 32918 98000
rect 34150 97322 34206 98000
rect 35438 97322 35494 98000
rect 32218 97294 32536 97322
rect 32218 97200 32274 97294
rect 32508 95674 32536 97294
rect 32862 97294 33088 97322
rect 32862 97200 32918 97294
rect 33060 95674 33088 97294
rect 34150 97294 34468 97322
rect 34150 97200 34206 97294
rect 34440 95674 34468 97294
rect 35360 97294 35494 97322
rect 35360 95674 35388 97294
rect 35438 97200 35494 97294
rect 36726 97322 36782 98000
rect 37370 97322 37426 98000
rect 38658 97322 38714 98000
rect 39946 97322 40002 98000
rect 36726 97294 37044 97322
rect 36726 97200 36782 97294
rect 35594 95772 35902 95781
rect 35594 95770 35600 95772
rect 35656 95770 35680 95772
rect 35736 95770 35760 95772
rect 35816 95770 35840 95772
rect 35896 95770 35902 95772
rect 35656 95718 35658 95770
rect 35838 95718 35840 95770
rect 35594 95716 35600 95718
rect 35656 95716 35680 95718
rect 35736 95716 35760 95718
rect 35816 95716 35840 95718
rect 35896 95716 35902 95718
rect 35594 95707 35902 95716
rect 37016 95674 37044 97294
rect 37370 97294 37596 97322
rect 37370 97200 37426 97294
rect 37568 95674 37596 97294
rect 38658 97294 38976 97322
rect 38658 97200 38714 97294
rect 38948 95674 38976 97294
rect 39868 97294 40002 97322
rect 39868 95674 39896 97294
rect 39946 97200 40002 97294
rect 40590 97322 40646 98000
rect 41878 97322 41934 98000
rect 43166 97322 43222 98000
rect 44454 97322 44510 98000
rect 45098 97322 45154 98000
rect 46386 97322 46442 98000
rect 47674 97322 47730 98000
rect 48318 97322 48374 98000
rect 50250 97322 50306 98000
rect 40590 97294 40816 97322
rect 40590 97200 40646 97294
rect 40788 95674 40816 97294
rect 41878 97294 42196 97322
rect 41878 97200 41934 97294
rect 42168 95674 42196 97294
rect 43166 97294 43484 97322
rect 43166 97200 43222 97294
rect 43456 95674 43484 97294
rect 44454 97294 44772 97322
rect 44454 97200 44510 97294
rect 44744 95674 44772 97294
rect 45098 97294 45324 97322
rect 45098 97200 45154 97294
rect 45296 95674 45324 97294
rect 46386 97294 46704 97322
rect 46386 97200 46442 97294
rect 46676 95674 46704 97294
rect 47674 97294 47992 97322
rect 47674 97200 47730 97294
rect 47964 95674 47992 97294
rect 48318 97294 48544 97322
rect 48318 97200 48374 97294
rect 48516 95674 48544 97294
rect 49896 97294 50306 97322
rect 25044 95668 25096 95674
rect 25044 95610 25096 95616
rect 26332 95668 26384 95674
rect 26332 95610 26384 95616
rect 27620 95668 27672 95674
rect 27620 95610 27672 95616
rect 29092 95668 29144 95674
rect 29092 95610 29144 95616
rect 29552 95668 29604 95674
rect 29552 95610 29604 95616
rect 30840 95668 30892 95674
rect 30840 95610 30892 95616
rect 32496 95668 32548 95674
rect 32496 95610 32548 95616
rect 33048 95668 33100 95674
rect 33048 95610 33100 95616
rect 34428 95668 34480 95674
rect 34428 95610 34480 95616
rect 35348 95668 35400 95674
rect 35348 95610 35400 95616
rect 37004 95668 37056 95674
rect 37004 95610 37056 95616
rect 37556 95668 37608 95674
rect 37556 95610 37608 95616
rect 38936 95668 38988 95674
rect 38936 95610 38988 95616
rect 39856 95668 39908 95674
rect 39856 95610 39908 95616
rect 40776 95668 40828 95674
rect 40776 95610 40828 95616
rect 42156 95668 42208 95674
rect 42156 95610 42208 95616
rect 43444 95668 43496 95674
rect 43444 95610 43496 95616
rect 44732 95668 44784 95674
rect 44732 95610 44784 95616
rect 45284 95668 45336 95674
rect 45284 95610 45336 95616
rect 46664 95668 46716 95674
rect 46664 95610 46716 95616
rect 47952 95668 48004 95674
rect 47952 95610 48004 95616
rect 48504 95668 48556 95674
rect 48504 95610 48556 95616
rect 32312 95532 32364 95538
rect 32312 95474 32364 95480
rect 33232 95532 33284 95538
rect 33232 95474 33284 95480
rect 34244 95532 34296 95538
rect 34244 95474 34296 95480
rect 35348 95532 35400 95538
rect 35348 95474 35400 95480
rect 36452 95532 36504 95538
rect 36452 95474 36504 95480
rect 37740 95532 37792 95538
rect 37740 95474 37792 95480
rect 38752 95532 38804 95538
rect 38752 95474 38804 95480
rect 39764 95532 39816 95538
rect 39764 95474 39816 95480
rect 40960 95532 41012 95538
rect 40960 95474 41012 95480
rect 41972 95532 42024 95538
rect 41972 95474 42024 95480
rect 43260 95532 43312 95538
rect 43260 95474 43312 95480
rect 44180 95532 44232 95538
rect 44180 95474 44232 95480
rect 45468 95532 45520 95538
rect 45468 95474 45520 95480
rect 46480 95532 46532 95538
rect 46480 95474 46532 95480
rect 47768 95532 47820 95538
rect 47768 95474 47820 95480
rect 48688 95532 48740 95538
rect 48688 95474 48740 95480
rect 25504 95464 25556 95470
rect 25504 95406 25556 95412
rect 24400 95124 24452 95130
rect 24400 95066 24452 95072
rect 24308 94920 24360 94926
rect 24308 94862 24360 94868
rect 22126 90902 22232 90930
rect 23230 90902 23336 90930
rect 24320 90916 24348 94862
rect 25516 90930 25544 95406
rect 28724 95396 28776 95402
rect 28724 95338 28776 95344
rect 26516 95328 26568 95334
rect 26516 95270 26568 95276
rect 27804 95328 27856 95334
rect 27804 95270 27856 95276
rect 25438 90902 25544 90930
rect 26528 90916 26556 95270
rect 27816 90930 27844 95270
rect 27646 90902 27844 90930
rect 28736 90916 28764 95338
rect 29920 95328 29972 95334
rect 29920 95270 29972 95276
rect 31024 95328 31076 95334
rect 31024 95270 31076 95276
rect 29932 90930 29960 95270
rect 31036 90930 31064 95270
rect 31852 93356 31904 93362
rect 31852 93298 31904 93304
rect 31864 93158 31892 93298
rect 31852 93152 31904 93158
rect 31852 93094 31904 93100
rect 32324 90930 32352 95474
rect 33244 90930 33272 95474
rect 29854 90902 29960 90930
rect 30958 90902 31064 90930
rect 32062 90902 32352 90930
rect 33166 90902 33272 90930
rect 34256 90916 34284 95474
rect 34934 95228 35242 95237
rect 34934 95226 34940 95228
rect 34996 95226 35020 95228
rect 35076 95226 35100 95228
rect 35156 95226 35180 95228
rect 35236 95226 35242 95228
rect 34996 95174 34998 95226
rect 35178 95174 35180 95226
rect 34934 95172 34940 95174
rect 34996 95172 35020 95174
rect 35076 95172 35100 95174
rect 35156 95172 35180 95174
rect 35236 95172 35242 95174
rect 34934 95163 35242 95172
rect 34934 94140 35242 94149
rect 34934 94138 34940 94140
rect 34996 94138 35020 94140
rect 35076 94138 35100 94140
rect 35156 94138 35180 94140
rect 35236 94138 35242 94140
rect 34996 94086 34998 94138
rect 35178 94086 35180 94138
rect 34934 94084 34940 94086
rect 34996 94084 35020 94086
rect 35076 94084 35100 94086
rect 35156 94084 35180 94086
rect 35236 94084 35242 94086
rect 34934 94075 35242 94084
rect 34934 93052 35242 93061
rect 34934 93050 34940 93052
rect 34996 93050 35020 93052
rect 35076 93050 35100 93052
rect 35156 93050 35180 93052
rect 35236 93050 35242 93052
rect 34996 92998 34998 93050
rect 35178 92998 35180 93050
rect 34934 92996 34940 92998
rect 34996 92996 35020 92998
rect 35076 92996 35100 92998
rect 35156 92996 35180 92998
rect 35236 92996 35242 92998
rect 34934 92987 35242 92996
rect 35360 90916 35388 95474
rect 35594 94684 35902 94693
rect 35594 94682 35600 94684
rect 35656 94682 35680 94684
rect 35736 94682 35760 94684
rect 35816 94682 35840 94684
rect 35896 94682 35902 94684
rect 35656 94630 35658 94682
rect 35838 94630 35840 94682
rect 35594 94628 35600 94630
rect 35656 94628 35680 94630
rect 35736 94628 35760 94630
rect 35816 94628 35840 94630
rect 35896 94628 35902 94630
rect 35594 94619 35902 94628
rect 35594 93596 35902 93605
rect 35594 93594 35600 93596
rect 35656 93594 35680 93596
rect 35736 93594 35760 93596
rect 35816 93594 35840 93596
rect 35896 93594 35902 93596
rect 35656 93542 35658 93594
rect 35838 93542 35840 93594
rect 35594 93540 35600 93542
rect 35656 93540 35680 93542
rect 35736 93540 35760 93542
rect 35816 93540 35840 93542
rect 35896 93540 35902 93542
rect 35594 93531 35902 93540
rect 36464 90916 36492 95474
rect 37752 90930 37780 95474
rect 38764 90930 38792 95474
rect 37582 90902 37780 90930
rect 38686 90902 38792 90930
rect 39776 90916 39804 95474
rect 40972 90930 41000 95474
rect 40894 90902 41000 90930
rect 41984 90916 42012 95474
rect 43272 90930 43300 95474
rect 43102 90902 43300 90930
rect 44192 90916 44220 95474
rect 45480 90930 45508 95474
rect 46492 90930 46520 95474
rect 47780 90930 47808 95474
rect 48700 90930 48728 95474
rect 49896 93158 49924 97294
rect 50250 97200 50306 97294
rect 50894 97322 50950 98000
rect 51538 97322 51594 98000
rect 52826 97322 52882 98000
rect 54114 97322 54170 98000
rect 56046 97322 56102 98000
rect 57334 97322 57390 98000
rect 58622 97322 58678 98000
rect 59910 97322 59966 98000
rect 60554 97322 60610 98000
rect 61842 97322 61898 98000
rect 63130 97322 63186 98000
rect 63774 97322 63830 98000
rect 65062 97322 65118 98000
rect 50894 97294 51028 97322
rect 50894 97200 50950 97294
rect 51000 95674 51028 97294
rect 51538 97294 51856 97322
rect 51538 97200 51594 97294
rect 50988 95668 51040 95674
rect 50988 95610 51040 95616
rect 51828 95538 51856 97294
rect 52826 97294 52960 97322
rect 52826 97200 52882 97294
rect 52932 95538 52960 97294
rect 54114 97294 54432 97322
rect 54114 97200 54170 97294
rect 54404 95674 54432 97294
rect 56046 97294 56456 97322
rect 56046 97200 56102 97294
rect 56428 95674 56456 97294
rect 57334 97294 57744 97322
rect 57334 97200 57390 97294
rect 54392 95668 54444 95674
rect 54392 95610 54444 95616
rect 56416 95668 56468 95674
rect 56416 95610 56468 95616
rect 57716 95538 57744 97294
rect 58544 97294 58678 97322
rect 58544 95674 58572 97294
rect 58622 97200 58678 97294
rect 59832 97294 59966 97322
rect 59832 95674 59860 97294
rect 59910 97200 59966 97294
rect 60476 97294 60610 97322
rect 60476 95674 60504 97294
rect 60554 97200 60610 97294
rect 61764 97294 61898 97322
rect 61764 95674 61792 97294
rect 61842 97200 61898 97294
rect 63052 97294 63186 97322
rect 63052 95674 63080 97294
rect 63130 97200 63186 97294
rect 63696 97294 63830 97322
rect 63696 95674 63724 97294
rect 63774 97200 63830 97294
rect 64984 97294 65118 97322
rect 64984 95674 65012 97294
rect 65062 97200 65118 97294
rect 66350 97322 66406 98000
rect 67638 97322 67694 98000
rect 68282 97322 68338 98000
rect 69570 97322 69626 98000
rect 70858 97322 70914 98000
rect 71502 97322 71558 98000
rect 72790 97322 72846 98000
rect 66350 97294 66760 97322
rect 66350 97200 66406 97294
rect 66314 95772 66622 95781
rect 66314 95770 66320 95772
rect 66376 95770 66400 95772
rect 66456 95770 66480 95772
rect 66536 95770 66560 95772
rect 66616 95770 66622 95772
rect 66376 95718 66378 95770
rect 66558 95718 66560 95770
rect 66314 95716 66320 95718
rect 66376 95716 66400 95718
rect 66456 95716 66480 95718
rect 66536 95716 66560 95718
rect 66616 95716 66622 95718
rect 66314 95707 66622 95716
rect 66732 95674 66760 97294
rect 67638 97294 67956 97322
rect 67638 97200 67694 97294
rect 67928 95674 67956 97294
rect 68282 97294 68600 97322
rect 68282 97200 68338 97294
rect 68572 95674 68600 97294
rect 69570 97294 69888 97322
rect 69570 97200 69626 97294
rect 69860 95674 69888 97294
rect 70780 97294 70914 97322
rect 70780 95674 70808 97294
rect 70858 97200 70914 97294
rect 71424 97294 71558 97322
rect 71424 95674 71452 97294
rect 71502 97200 71558 97294
rect 72712 97294 72846 97322
rect 72712 95674 72740 97294
rect 72790 97200 72846 97294
rect 74078 97322 74134 98000
rect 75366 97322 75422 98000
rect 76010 97322 76066 98000
rect 77298 97322 77354 98000
rect 78586 97322 78642 98000
rect 74078 97294 74396 97322
rect 74078 97200 74134 97294
rect 74368 95674 74396 97294
rect 75366 97294 75684 97322
rect 75366 97200 75422 97294
rect 75656 95674 75684 97294
rect 76010 97294 76236 97322
rect 76010 97200 76066 97294
rect 76208 95674 76236 97294
rect 77298 97294 77616 97322
rect 77298 97200 77354 97294
rect 77588 95674 77616 97294
rect 78508 97294 78642 97322
rect 78508 95674 78536 97294
rect 78586 97200 78642 97294
rect 79230 97322 79286 98000
rect 80518 97322 80574 98000
rect 81806 97322 81862 98000
rect 83094 97322 83150 98000
rect 83738 97322 83794 98000
rect 85026 97322 85082 98000
rect 86314 97322 86370 98000
rect 86958 97322 87014 98000
rect 88246 97322 88302 98000
rect 79230 97294 79456 97322
rect 79230 97200 79286 97294
rect 79428 95674 79456 97294
rect 80518 97294 80836 97322
rect 80518 97200 80574 97294
rect 80808 95674 80836 97294
rect 81806 97294 82124 97322
rect 81806 97200 81862 97294
rect 82096 95674 82124 97294
rect 83094 97294 83412 97322
rect 83094 97200 83150 97294
rect 83384 95674 83412 97294
rect 83738 97294 83964 97322
rect 83738 97200 83794 97294
rect 83936 95674 83964 97294
rect 85026 97294 85344 97322
rect 85026 97200 85082 97294
rect 85316 95674 85344 97294
rect 86314 97294 86632 97322
rect 86314 97200 86370 97294
rect 86604 95674 86632 97294
rect 86958 97294 87184 97322
rect 86958 97200 87014 97294
rect 87156 95674 87184 97294
rect 88168 97294 88302 97322
rect 88168 95674 88196 97294
rect 88246 97200 88302 97294
rect 89534 97322 89590 98000
rect 90822 97322 90878 98000
rect 89534 97294 89668 97322
rect 89534 97200 89590 97294
rect 89640 95674 89668 97294
rect 90822 97294 91048 97322
rect 90822 97200 90878 97294
rect 91020 95674 91048 97294
rect 97034 95772 97342 95781
rect 97034 95770 97040 95772
rect 97096 95770 97120 95772
rect 97176 95770 97200 95772
rect 97256 95770 97280 95772
rect 97336 95770 97342 95772
rect 97096 95718 97098 95770
rect 97278 95718 97280 95770
rect 97034 95716 97040 95718
rect 97096 95716 97120 95718
rect 97176 95716 97200 95718
rect 97256 95716 97280 95718
rect 97336 95716 97342 95718
rect 97034 95707 97342 95716
rect 58532 95668 58584 95674
rect 58532 95610 58584 95616
rect 59820 95668 59872 95674
rect 59820 95610 59872 95616
rect 60464 95668 60516 95674
rect 60464 95610 60516 95616
rect 61752 95668 61804 95674
rect 61752 95610 61804 95616
rect 63040 95668 63092 95674
rect 63040 95610 63092 95616
rect 63684 95668 63736 95674
rect 63684 95610 63736 95616
rect 64972 95668 65024 95674
rect 64972 95610 65024 95616
rect 66720 95668 66772 95674
rect 66720 95610 66772 95616
rect 67916 95668 67968 95674
rect 67916 95610 67968 95616
rect 68560 95668 68612 95674
rect 68560 95610 68612 95616
rect 69848 95668 69900 95674
rect 69848 95610 69900 95616
rect 70768 95668 70820 95674
rect 70768 95610 70820 95616
rect 71412 95668 71464 95674
rect 71412 95610 71464 95616
rect 72700 95668 72752 95674
rect 72700 95610 72752 95616
rect 74356 95668 74408 95674
rect 74356 95610 74408 95616
rect 75644 95668 75696 95674
rect 75644 95610 75696 95616
rect 76196 95668 76248 95674
rect 76196 95610 76248 95616
rect 77576 95668 77628 95674
rect 77576 95610 77628 95616
rect 78496 95668 78548 95674
rect 78496 95610 78548 95616
rect 79416 95668 79468 95674
rect 79416 95610 79468 95616
rect 80796 95668 80848 95674
rect 80796 95610 80848 95616
rect 82084 95668 82136 95674
rect 82084 95610 82136 95616
rect 83372 95668 83424 95674
rect 83372 95610 83424 95616
rect 83924 95668 83976 95674
rect 83924 95610 83976 95616
rect 85304 95668 85356 95674
rect 85304 95610 85356 95616
rect 86592 95668 86644 95674
rect 86592 95610 86644 95616
rect 87144 95668 87196 95674
rect 87144 95610 87196 95616
rect 88156 95668 88208 95674
rect 88156 95610 88208 95616
rect 89628 95668 89680 95674
rect 89628 95610 89680 95616
rect 91008 95668 91060 95674
rect 91008 95610 91060 95616
rect 51080 95532 51132 95538
rect 51080 95474 51132 95480
rect 51816 95532 51868 95538
rect 51816 95474 51868 95480
rect 52920 95532 52972 95538
rect 52920 95474 52972 95480
rect 57704 95532 57756 95538
rect 57704 95474 57756 95480
rect 74172 95532 74224 95538
rect 74172 95474 74224 95480
rect 75460 95532 75512 95538
rect 75460 95474 75512 95480
rect 76380 95532 76432 95538
rect 76380 95474 76432 95480
rect 77392 95532 77444 95538
rect 77392 95474 77444 95480
rect 78588 95532 78640 95538
rect 78588 95474 78640 95480
rect 79600 95532 79652 95538
rect 79600 95474 79652 95480
rect 80612 95532 80664 95538
rect 80612 95474 80664 95480
rect 81900 95532 81952 95538
rect 81900 95474 81952 95480
rect 83188 95532 83240 95538
rect 83188 95474 83240 95480
rect 84108 95532 84160 95538
rect 84108 95474 84160 95480
rect 85120 95532 85172 95538
rect 85120 95474 85172 95480
rect 86408 95532 86460 95538
rect 86408 95474 86460 95480
rect 87328 95532 87380 95538
rect 87328 95474 87380 95480
rect 88340 95532 88392 95538
rect 88340 95474 88392 95480
rect 89628 95532 89680 95538
rect 89628 95474 89680 95480
rect 90916 95532 90968 95538
rect 90916 95474 90968 95480
rect 51092 94790 51120 95474
rect 52368 95464 52420 95470
rect 52368 95406 52420 95412
rect 52380 95010 52408 95406
rect 52932 95130 52960 95474
rect 54116 95464 54168 95470
rect 54116 95406 54168 95412
rect 56784 95464 56836 95470
rect 56784 95406 56836 95412
rect 66720 95464 66772 95470
rect 66720 95406 66772 95412
rect 67456 95464 67508 95470
rect 67456 95406 67508 95412
rect 52920 95124 52972 95130
rect 52920 95066 52972 95072
rect 52380 94994 52500 95010
rect 52380 94988 52512 94994
rect 52380 94982 52460 94988
rect 52460 94930 52512 94936
rect 52920 94988 52972 94994
rect 52920 94930 52972 94936
rect 51080 94784 51132 94790
rect 51080 94726 51132 94732
rect 50712 93288 50764 93294
rect 50712 93230 50764 93236
rect 49884 93152 49936 93158
rect 49884 93094 49936 93100
rect 50528 92472 50580 92478
rect 50528 92414 50580 92420
rect 45310 90902 45508 90930
rect 46414 90902 46520 90930
rect 47518 90902 47808 90930
rect 48622 90902 48728 90930
rect 13266 90536 13322 90545
rect 13266 90471 13322 90480
rect 8484 90160 8536 90166
rect 8484 90102 8536 90108
rect 8298 87544 8354 87553
rect 8298 87479 8354 87488
rect 8312 87310 8340 87479
rect 8300 87304 8352 87310
rect 8300 87246 8352 87252
rect 8300 86828 8352 86834
rect 8300 86770 8352 86776
rect 8312 86737 8340 86770
rect 8298 86728 8354 86737
rect 8298 86663 8354 86672
rect 8298 85368 8354 85377
rect 8298 85303 8354 85312
rect 8312 85134 8340 85303
rect 8300 85128 8352 85134
rect 8300 85070 8352 85076
rect 8300 83564 8352 83570
rect 8300 83506 8352 83512
rect 8312 83473 8340 83506
rect 8298 83464 8354 83473
rect 8298 83399 8354 83408
rect 8298 82104 8354 82113
rect 8298 82039 8354 82048
rect 8312 81870 8340 82039
rect 8300 81864 8352 81870
rect 8300 81806 8352 81812
rect 8300 81388 8352 81394
rect 8300 81330 8352 81336
rect 8312 81297 8340 81330
rect 8298 81288 8354 81297
rect 8298 81223 8354 81232
rect 8298 79928 8354 79937
rect 8298 79863 8354 79872
rect 8312 79694 8340 79863
rect 8300 79688 8352 79694
rect 8300 79630 8352 79636
rect 8300 79212 8352 79218
rect 8300 79154 8352 79160
rect 8312 79121 8340 79154
rect 8298 79112 8354 79121
rect 8298 79047 8354 79056
rect 8300 78124 8352 78130
rect 8300 78066 8352 78072
rect 8312 78033 8340 78066
rect 8298 78024 8354 78033
rect 8298 77959 8354 77968
rect 8298 76664 8354 76673
rect 8298 76599 8354 76608
rect 8312 76430 8340 76599
rect 8300 76424 8352 76430
rect 8300 76366 8352 76372
rect 8298 74488 8354 74497
rect 8298 74423 8354 74432
rect 8312 74254 8340 74423
rect 8300 74248 8352 74254
rect 8300 74190 8352 74196
rect 8300 73772 8352 73778
rect 8300 73714 8352 73720
rect 8312 73681 8340 73714
rect 8298 73672 8354 73681
rect 8298 73607 8354 73616
rect 8300 72684 8352 72690
rect 8300 72626 8352 72632
rect 8312 72593 8340 72626
rect 8298 72584 8354 72593
rect 8298 72519 8354 72528
rect 8298 71224 8354 71233
rect 8298 71159 8354 71168
rect 8312 70990 8340 71159
rect 8300 70984 8352 70990
rect 8300 70926 8352 70932
rect 8300 68740 8352 68746
rect 8300 68682 8352 68688
rect 8312 68649 8340 68682
rect 8298 68640 8354 68649
rect 8298 68575 8354 68584
rect 8300 68196 8352 68202
rect 8300 68138 8352 68144
rect 8312 68105 8340 68138
rect 8298 68096 8354 68105
rect 8298 68031 8354 68040
rect 8300 67108 8352 67114
rect 8300 67050 8352 67056
rect 8312 67017 8340 67050
rect 8298 67008 8354 67017
rect 8298 66943 8354 66952
rect 8298 65784 8354 65793
rect 8298 65719 8354 65728
rect 8312 65686 8340 65719
rect 8300 65680 8352 65686
rect 8300 65622 8352 65628
rect 8300 63300 8352 63306
rect 8300 63242 8352 63248
rect 8312 63209 8340 63242
rect 8298 63200 8354 63209
rect 8298 63135 8354 63144
rect 8300 62756 8352 62762
rect 8300 62698 8352 62704
rect 8312 62665 8340 62698
rect 8298 62656 8354 62665
rect 8298 62591 8354 62600
rect 8300 61668 8352 61674
rect 8300 61610 8352 61616
rect 8312 61577 8340 61610
rect 8298 61568 8354 61577
rect 8298 61503 8354 61512
rect 8298 60344 8354 60353
rect 8298 60279 8300 60288
rect 8352 60279 8354 60288
rect 8300 60250 8352 60256
rect 50436 60036 50488 60042
rect 50436 59978 50488 59984
rect 8300 57316 8352 57322
rect 8300 57258 8352 57264
rect 8312 57225 8340 57258
rect 8298 57216 8354 57225
rect 8298 57151 8354 57160
rect 8300 56228 8352 56234
rect 8300 56170 8352 56176
rect 8312 56137 8340 56170
rect 8298 56128 8354 56137
rect 8298 56063 8354 56072
rect 8298 54904 8354 54913
rect 8298 54839 8300 54848
rect 8352 54839 8354 54848
rect 8300 54810 8352 54816
rect 5724 51060 5776 51066
rect 5724 51002 5776 51008
rect 8484 51060 8536 51066
rect 8484 51002 8536 51008
rect 7472 50856 7524 50862
rect 7472 50798 7524 50804
rect 7484 50114 7512 50798
rect 8496 50674 8524 51002
rect 8208 50652 8260 50658
rect 8496 50646 8878 50674
rect 9864 50652 9916 50658
rect 8208 50594 8260 50600
rect 9864 50594 9916 50600
rect 8024 50176 8076 50182
rect 8024 50118 8076 50124
rect 7472 50108 7524 50114
rect 7472 50050 7524 50056
rect 5540 48884 5592 48890
rect 5540 48826 5592 48832
rect 1216 48748 1268 48754
rect 1216 48690 1268 48696
rect 5632 48748 5684 48754
rect 5632 48690 5684 48696
rect 1228 48385 1256 48690
rect 4214 48444 4522 48453
rect 4214 48442 4220 48444
rect 4276 48442 4300 48444
rect 4356 48442 4380 48444
rect 4436 48442 4460 48444
rect 4516 48442 4522 48444
rect 4276 48390 4278 48442
rect 4458 48390 4460 48442
rect 4214 48388 4220 48390
rect 4276 48388 4300 48390
rect 4356 48388 4380 48390
rect 4436 48388 4460 48390
rect 4516 48388 4522 48390
rect 1214 48376 1270 48385
rect 4214 48379 4522 48388
rect 1214 48311 1270 48320
rect 5644 48278 5672 48690
rect 5632 48272 5684 48278
rect 5632 48214 5684 48220
rect 4874 47900 5182 47909
rect 4874 47898 4880 47900
rect 4936 47898 4960 47900
rect 5016 47898 5040 47900
rect 5096 47898 5120 47900
rect 5176 47898 5182 47900
rect 4936 47846 4938 47898
rect 5118 47846 5120 47898
rect 4874 47844 4880 47846
rect 4936 47844 4960 47846
rect 5016 47844 5040 47846
rect 5096 47844 5120 47846
rect 5176 47844 5182 47846
rect 4874 47835 5182 47844
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 4874 46812 5182 46821
rect 4874 46810 4880 46812
rect 4936 46810 4960 46812
rect 5016 46810 5040 46812
rect 5096 46810 5120 46812
rect 5176 46810 5182 46812
rect 4936 46758 4938 46810
rect 5118 46758 5120 46810
rect 4874 46756 4880 46758
rect 4936 46756 4960 46758
rect 5016 46756 5040 46758
rect 5096 46756 5120 46758
rect 5176 46756 5182 46758
rect 4874 46747 5182 46756
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 1676 45960 1728 45966
rect 1676 45902 1728 45908
rect 848 45824 900 45830
rect 846 45792 848 45801
rect 900 45792 902 45801
rect 846 45727 902 45736
rect 1688 45393 1716 45902
rect 4874 45724 5182 45733
rect 4874 45722 4880 45724
rect 4936 45722 4960 45724
rect 5016 45722 5040 45724
rect 5096 45722 5120 45724
rect 5176 45722 5182 45724
rect 4936 45670 4938 45722
rect 5118 45670 5120 45722
rect 4874 45668 4880 45670
rect 4936 45668 4960 45670
rect 5016 45668 5040 45670
rect 5096 45668 5120 45670
rect 5176 45668 5182 45670
rect 4874 45659 5182 45668
rect 1674 45384 1730 45393
rect 1674 45319 1730 45328
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 4874 44636 5182 44645
rect 4874 44634 4880 44636
rect 4936 44634 4960 44636
rect 5016 44634 5040 44636
rect 5096 44634 5120 44636
rect 5176 44634 5182 44636
rect 4936 44582 4938 44634
rect 5118 44582 5120 44634
rect 4874 44580 4880 44582
rect 4936 44580 4960 44582
rect 5016 44580 5040 44582
rect 5096 44580 5120 44582
rect 5176 44580 5182 44582
rect 4874 44571 5182 44580
rect 848 44532 900 44538
rect 848 44474 900 44480
rect 860 44441 888 44474
rect 846 44432 902 44441
rect 846 44367 902 44376
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 4874 43548 5182 43557
rect 4874 43546 4880 43548
rect 4936 43546 4960 43548
rect 5016 43546 5040 43548
rect 5096 43546 5120 43548
rect 5176 43546 5182 43548
rect 4936 43494 4938 43546
rect 5118 43494 5120 43546
rect 4874 43492 4880 43494
rect 4936 43492 4960 43494
rect 5016 43492 5040 43494
rect 5096 43492 5120 43494
rect 5176 43492 5182 43494
rect 4874 43483 5182 43492
rect 848 43104 900 43110
rect 846 43072 848 43081
rect 900 43072 902 43081
rect 846 43007 902 43016
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 848 42560 900 42566
rect 848 42502 900 42508
rect 860 42401 888 42502
rect 4874 42460 5182 42469
rect 4874 42458 4880 42460
rect 4936 42458 4960 42460
rect 5016 42458 5040 42460
rect 5096 42458 5120 42460
rect 5176 42458 5182 42460
rect 4936 42406 4938 42458
rect 5118 42406 5120 42458
rect 4874 42404 4880 42406
rect 4936 42404 4960 42406
rect 5016 42404 5040 42406
rect 5096 42404 5120 42406
rect 5176 42404 5182 42406
rect 846 42392 902 42401
rect 4874 42395 5182 42404
rect 846 42327 902 42336
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 4874 41372 5182 41381
rect 4874 41370 4880 41372
rect 4936 41370 4960 41372
rect 5016 41370 5040 41372
rect 5096 41370 5120 41372
rect 5176 41370 5182 41372
rect 4936 41318 4938 41370
rect 5118 41318 5120 41370
rect 4874 41316 4880 41318
rect 4936 41316 4960 41318
rect 5016 41316 5040 41318
rect 5096 41316 5120 41318
rect 5176 41316 5182 41318
rect 4874 41307 5182 41316
rect 846 41032 902 41041
rect 846 40967 848 40976
rect 900 40967 902 40976
rect 848 40938 900 40944
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 1676 40520 1728 40526
rect 1676 40462 1728 40468
rect 848 40384 900 40390
rect 846 40352 848 40361
rect 900 40352 902 40361
rect 846 40287 902 40296
rect 1688 39953 1716 40462
rect 4874 40284 5182 40293
rect 4874 40282 4880 40284
rect 4936 40282 4960 40284
rect 5016 40282 5040 40284
rect 5096 40282 5120 40284
rect 5176 40282 5182 40284
rect 4936 40230 4938 40282
rect 5118 40230 5120 40282
rect 4874 40228 4880 40230
rect 4936 40228 4960 40230
rect 5016 40228 5040 40230
rect 5096 40228 5120 40230
rect 5176 40228 5182 40230
rect 4874 40219 5182 40228
rect 1674 39944 1730 39953
rect 1674 39879 1730 39888
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 4874 39196 5182 39205
rect 4874 39194 4880 39196
rect 4936 39194 4960 39196
rect 5016 39194 5040 39196
rect 5096 39194 5120 39196
rect 5176 39194 5182 39196
rect 4936 39142 4938 39194
rect 5118 39142 5120 39194
rect 4874 39140 4880 39142
rect 4936 39140 4960 39142
rect 5016 39140 5040 39142
rect 5096 39140 5120 39142
rect 5176 39140 5182 39142
rect 4874 39131 5182 39140
rect 848 38752 900 38758
rect 846 38720 848 38729
rect 900 38720 902 38729
rect 846 38655 902 38664
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 4874 38108 5182 38117
rect 4874 38106 4880 38108
rect 4936 38106 4960 38108
rect 5016 38106 5040 38108
rect 5096 38106 5120 38108
rect 5176 38106 5182 38108
rect 4936 38054 4938 38106
rect 5118 38054 5120 38106
rect 4874 38052 4880 38054
rect 4936 38052 4960 38054
rect 5016 38052 5040 38054
rect 5096 38052 5120 38054
rect 5176 38052 5182 38054
rect 4874 38043 5182 38052
rect 848 37664 900 37670
rect 846 37632 848 37641
rect 900 37632 902 37641
rect 846 37567 902 37576
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 848 37120 900 37126
rect 848 37062 900 37068
rect 860 36961 888 37062
rect 4874 37020 5182 37029
rect 4874 37018 4880 37020
rect 4936 37018 4960 37020
rect 5016 37018 5040 37020
rect 5096 37018 5120 37020
rect 5176 37018 5182 37020
rect 4936 36966 4938 37018
rect 5118 36966 5120 37018
rect 4874 36964 4880 36966
rect 4936 36964 4960 36966
rect 5016 36964 5040 36966
rect 5096 36964 5120 36966
rect 5176 36964 5182 36966
rect 846 36952 902 36961
rect 4874 36955 5182 36964
rect 846 36887 902 36896
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4874 35932 5182 35941
rect 4874 35930 4880 35932
rect 4936 35930 4960 35932
rect 5016 35930 5040 35932
rect 5096 35930 5120 35932
rect 5176 35930 5182 35932
rect 4936 35878 4938 35930
rect 5118 35878 5120 35930
rect 4874 35876 4880 35878
rect 4936 35876 4960 35878
rect 5016 35876 5040 35878
rect 5096 35876 5120 35878
rect 5176 35876 5182 35878
rect 4874 35867 5182 35876
rect 846 35592 902 35601
rect 846 35527 848 35536
rect 900 35527 902 35536
rect 848 35498 900 35504
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 1676 35080 1728 35086
rect 1676 35022 1728 35028
rect 848 34944 900 34950
rect 846 34912 848 34921
rect 900 34912 902 34921
rect 846 34847 902 34856
rect 1688 34513 1716 35022
rect 4874 34844 5182 34853
rect 4874 34842 4880 34844
rect 4936 34842 4960 34844
rect 5016 34842 5040 34844
rect 5096 34842 5120 34844
rect 5176 34842 5182 34844
rect 4936 34790 4938 34842
rect 5118 34790 5120 34842
rect 4874 34788 4880 34790
rect 4936 34788 4960 34790
rect 5016 34788 5040 34790
rect 5096 34788 5120 34790
rect 5176 34788 5182 34790
rect 4874 34779 5182 34788
rect 1674 34504 1730 34513
rect 1674 34439 1730 34448
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4874 33756 5182 33765
rect 4874 33754 4880 33756
rect 4936 33754 4960 33756
rect 5016 33754 5040 33756
rect 5096 33754 5120 33756
rect 5176 33754 5182 33756
rect 4936 33702 4938 33754
rect 5118 33702 5120 33754
rect 4874 33700 4880 33702
rect 4936 33700 4960 33702
rect 5016 33700 5040 33702
rect 5096 33700 5120 33702
rect 5176 33700 5182 33702
rect 4874 33691 5182 33700
rect 848 33312 900 33318
rect 846 33280 848 33289
rect 900 33280 902 33289
rect 846 33215 902 33224
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4874 32668 5182 32677
rect 4874 32666 4880 32668
rect 4936 32666 4960 32668
rect 5016 32666 5040 32668
rect 5096 32666 5120 32668
rect 5176 32666 5182 32668
rect 4936 32614 4938 32666
rect 5118 32614 5120 32666
rect 4874 32612 4880 32614
rect 4936 32612 4960 32614
rect 5016 32612 5040 32614
rect 5096 32612 5120 32614
rect 5176 32612 5182 32614
rect 4874 32603 5182 32612
rect 848 32224 900 32230
rect 846 32192 848 32201
rect 900 32192 902 32201
rect 846 32127 902 32136
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 848 31952 900 31958
rect 848 31894 900 31900
rect 860 31521 888 31894
rect 1676 31816 1728 31822
rect 1676 31758 1728 31764
rect 846 31512 902 31521
rect 846 31447 902 31456
rect 1688 31249 1716 31758
rect 4874 31580 5182 31589
rect 4874 31578 4880 31580
rect 4936 31578 4960 31580
rect 5016 31578 5040 31580
rect 5096 31578 5120 31580
rect 5176 31578 5182 31580
rect 4936 31526 4938 31578
rect 5118 31526 5120 31578
rect 4874 31524 4880 31526
rect 4936 31524 4960 31526
rect 5016 31524 5040 31526
rect 5096 31524 5120 31526
rect 5176 31524 5182 31526
rect 4874 31515 5182 31524
rect 1674 31240 1730 31249
rect 1674 31175 1730 31184
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4874 30492 5182 30501
rect 4874 30490 4880 30492
rect 4936 30490 4960 30492
rect 5016 30490 5040 30492
rect 5096 30490 5120 30492
rect 5176 30490 5182 30492
rect 4936 30438 4938 30490
rect 5118 30438 5120 30490
rect 4874 30436 4880 30438
rect 4936 30436 4960 30438
rect 5016 30436 5040 30438
rect 5096 30436 5120 30438
rect 5176 30436 5182 30438
rect 4874 30427 5182 30436
rect 846 30152 902 30161
rect 846 30087 848 30096
rect 900 30087 902 30096
rect 848 30058 900 30064
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 848 29504 900 29510
rect 846 29472 848 29481
rect 900 29472 902 29481
rect 846 29407 902 29416
rect 4874 29404 5182 29413
rect 4874 29402 4880 29404
rect 4936 29402 4960 29404
rect 5016 29402 5040 29404
rect 5096 29402 5120 29404
rect 5176 29402 5182 29404
rect 4936 29350 4938 29402
rect 5118 29350 5120 29402
rect 4874 29348 4880 29350
rect 4936 29348 4960 29350
rect 5016 29348 5040 29350
rect 5096 29348 5120 29350
rect 5176 29348 5182 29350
rect 4874 29339 5182 29348
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4874 28316 5182 28325
rect 4874 28314 4880 28316
rect 4936 28314 4960 28316
rect 5016 28314 5040 28316
rect 5096 28314 5120 28316
rect 5176 28314 5182 28316
rect 4936 28262 4938 28314
rect 5118 28262 5120 28314
rect 4874 28260 4880 28262
rect 4936 28260 4960 28262
rect 5016 28260 5040 28262
rect 5096 28260 5120 28262
rect 5176 28260 5182 28262
rect 4874 28251 5182 28260
rect 1308 28076 1360 28082
rect 1308 28018 1360 28024
rect 1320 27985 1348 28018
rect 1306 27976 1362 27985
rect 1306 27911 1362 27920
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4874 27228 5182 27237
rect 4874 27226 4880 27228
rect 4936 27226 4960 27228
rect 5016 27226 5040 27228
rect 5096 27226 5120 27228
rect 5176 27226 5182 27228
rect 4936 27174 4938 27226
rect 5118 27174 5120 27226
rect 4874 27172 4880 27174
rect 4936 27172 4960 27174
rect 5016 27172 5040 27174
rect 5096 27172 5120 27174
rect 5176 27172 5182 27174
rect 4874 27163 5182 27172
rect 1308 26988 1360 26994
rect 1308 26930 1360 26936
rect 1320 26625 1348 26930
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 1306 26616 1362 26625
rect 4214 26619 4522 26628
rect 1306 26551 1362 26560
rect 1308 26376 1360 26382
rect 1308 26318 1360 26324
rect 1320 25945 1348 26318
rect 1676 26308 1728 26314
rect 1676 26250 1728 26256
rect 1306 25936 1362 25945
rect 1306 25871 1362 25880
rect 1688 25809 1716 26250
rect 4874 26140 5182 26149
rect 4874 26138 4880 26140
rect 4936 26138 4960 26140
rect 5016 26138 5040 26140
rect 5096 26138 5120 26140
rect 5176 26138 5182 26140
rect 4936 26086 4938 26138
rect 5118 26086 5120 26138
rect 4874 26084 4880 26086
rect 4936 26084 4960 26086
rect 5016 26084 5040 26086
rect 5096 26084 5120 26086
rect 5176 26084 5182 26086
rect 4874 26075 5182 26084
rect 1674 25800 1730 25809
rect 1674 25735 1730 25744
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4874 25052 5182 25061
rect 4874 25050 4880 25052
rect 4936 25050 4960 25052
rect 5016 25050 5040 25052
rect 5096 25050 5120 25052
rect 5176 25050 5182 25052
rect 4936 24998 4938 25050
rect 5118 24998 5120 25050
rect 4874 24996 4880 24998
rect 4936 24996 4960 24998
rect 5016 24996 5040 24998
rect 5096 24996 5120 24998
rect 5176 24996 5182 24998
rect 4874 24987 5182 24996
rect 1308 24812 1360 24818
rect 1308 24754 1360 24760
rect 1320 24585 1348 24754
rect 1306 24576 1362 24585
rect 1306 24511 1362 24520
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 1308 24132 1360 24138
rect 1308 24074 1360 24080
rect 1320 23905 1348 24074
rect 4874 23964 5182 23973
rect 4874 23962 4880 23964
rect 4936 23962 4960 23964
rect 5016 23962 5040 23964
rect 5096 23962 5120 23964
rect 5176 23962 5182 23964
rect 4936 23910 4938 23962
rect 5118 23910 5120 23962
rect 4874 23908 4880 23910
rect 4936 23908 4960 23910
rect 5016 23908 5040 23910
rect 5096 23908 5120 23910
rect 5176 23908 5182 23910
rect 1306 23896 1362 23905
rect 4874 23899 5182 23908
rect 1306 23831 1362 23840
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4874 22876 5182 22885
rect 4874 22874 4880 22876
rect 4936 22874 4960 22876
rect 5016 22874 5040 22876
rect 5096 22874 5120 22876
rect 5176 22874 5182 22876
rect 4936 22822 4938 22874
rect 5118 22822 5120 22874
rect 4874 22820 4880 22822
rect 4936 22820 4960 22822
rect 5016 22820 5040 22822
rect 5096 22820 5120 22822
rect 5176 22820 5182 22822
rect 4874 22811 5182 22820
rect 1124 22636 1176 22642
rect 1124 22578 1176 22584
rect 1136 22545 1164 22578
rect 1122 22536 1178 22545
rect 1122 22471 1178 22480
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4874 21788 5182 21797
rect 4874 21786 4880 21788
rect 4936 21786 4960 21788
rect 5016 21786 5040 21788
rect 5096 21786 5120 21788
rect 5176 21786 5182 21788
rect 4936 21734 4938 21786
rect 5118 21734 5120 21786
rect 4874 21732 4880 21734
rect 4936 21732 4960 21734
rect 5016 21732 5040 21734
rect 5096 21732 5120 21734
rect 5176 21732 5182 21734
rect 4874 21723 5182 21732
rect 1308 21548 1360 21554
rect 1308 21490 1360 21496
rect 1320 21185 1348 21490
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 1306 21176 1362 21185
rect 4214 21179 4522 21188
rect 1306 21111 1362 21120
rect 1308 20868 1360 20874
rect 1308 20810 1360 20816
rect 1860 20868 1912 20874
rect 1860 20810 1912 20816
rect 1320 20505 1348 20810
rect 1306 20496 1362 20505
rect 1306 20431 1362 20440
rect 1872 20369 1900 20810
rect 4874 20700 5182 20709
rect 4874 20698 4880 20700
rect 4936 20698 4960 20700
rect 5016 20698 5040 20700
rect 5096 20698 5120 20700
rect 5176 20698 5182 20700
rect 4936 20646 4938 20698
rect 5118 20646 5120 20698
rect 4874 20644 4880 20646
rect 4936 20644 4960 20646
rect 5016 20644 5040 20646
rect 5096 20644 5120 20646
rect 5176 20644 5182 20646
rect 4874 20635 5182 20644
rect 1858 20360 1914 20369
rect 1858 20295 1914 20304
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4874 19612 5182 19621
rect 4874 19610 4880 19612
rect 4936 19610 4960 19612
rect 5016 19610 5040 19612
rect 5096 19610 5120 19612
rect 5176 19610 5182 19612
rect 4936 19558 4938 19610
rect 5118 19558 5120 19610
rect 4874 19556 4880 19558
rect 4936 19556 4960 19558
rect 5016 19556 5040 19558
rect 5096 19556 5120 19558
rect 5176 19556 5182 19558
rect 4874 19547 5182 19556
rect 1492 19372 1544 19378
rect 1492 19314 1544 19320
rect 1504 19145 1532 19314
rect 1490 19136 1546 19145
rect 1490 19071 1546 19080
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 1308 18692 1360 18698
rect 1308 18634 1360 18640
rect 1320 18465 1348 18634
rect 4874 18524 5182 18533
rect 4874 18522 4880 18524
rect 4936 18522 4960 18524
rect 5016 18522 5040 18524
rect 5096 18522 5120 18524
rect 5176 18522 5182 18524
rect 4936 18470 4938 18522
rect 5118 18470 5120 18522
rect 4874 18468 4880 18470
rect 4936 18468 4960 18470
rect 5016 18468 5040 18470
rect 5096 18468 5120 18470
rect 5176 18468 5182 18470
rect 1306 18456 1362 18465
rect 4874 18459 5182 18468
rect 1306 18391 1362 18400
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4874 17436 5182 17445
rect 4874 17434 4880 17436
rect 4936 17434 4960 17436
rect 5016 17434 5040 17436
rect 5096 17434 5120 17436
rect 5176 17434 5182 17436
rect 4936 17382 4938 17434
rect 5118 17382 5120 17434
rect 4874 17380 4880 17382
rect 4936 17380 4960 17382
rect 5016 17380 5040 17382
rect 5096 17380 5120 17382
rect 5176 17380 5182 17382
rect 4874 17371 5182 17380
rect 1124 17196 1176 17202
rect 1124 17138 1176 17144
rect 1136 17105 1164 17138
rect 1122 17096 1178 17105
rect 1122 17031 1178 17040
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4874 16348 5182 16357
rect 4874 16346 4880 16348
rect 4936 16346 4960 16348
rect 5016 16346 5040 16348
rect 5096 16346 5120 16348
rect 5176 16346 5182 16348
rect 4936 16294 4938 16346
rect 5118 16294 5120 16346
rect 4874 16292 4880 16294
rect 4936 16292 4960 16294
rect 5016 16292 5040 16294
rect 5096 16292 5120 16294
rect 5176 16292 5182 16294
rect 4874 16283 5182 16292
rect 1216 16108 1268 16114
rect 1216 16050 1268 16056
rect 1228 15745 1256 16050
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 1214 15736 1270 15745
rect 4214 15739 4522 15748
rect 1214 15671 1270 15680
rect 1308 15428 1360 15434
rect 1308 15370 1360 15376
rect 1860 15428 1912 15434
rect 1860 15370 1912 15376
rect 1320 15065 1348 15370
rect 1306 15056 1362 15065
rect 1306 14991 1362 15000
rect 1872 14929 1900 15370
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 1858 14920 1914 14929
rect 1858 14855 1914 14864
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 1308 13932 1360 13938
rect 1308 13874 1360 13880
rect 1320 13705 1348 13874
rect 1306 13696 1362 13705
rect 1306 13631 1362 13640
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 1308 13320 1360 13326
rect 1308 13262 1360 13268
rect 1320 13025 1348 13262
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 1306 13016 1362 13025
rect 4874 13019 5182 13028
rect 1306 12951 1362 12960
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 1124 11756 1176 11762
rect 1124 11698 1176 11704
rect 1136 11665 1164 11698
rect 1122 11656 1178 11665
rect 1122 11591 1178 11600
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 8036 8158 8064 50118
rect 8116 50108 8168 50114
rect 8116 50050 8168 50056
rect 8128 8226 8156 50050
rect 8220 8294 8248 50594
rect 9876 50266 9904 50594
rect 9876 50250 10272 50266
rect 9876 50244 10284 50250
rect 9876 50238 10232 50244
rect 10232 50186 10284 50192
rect 11796 50176 11848 50182
rect 11086 50114 11192 50130
rect 11848 50124 12190 50130
rect 11796 50118 12190 50124
rect 11086 50108 11204 50114
rect 11086 50102 11152 50108
rect 11808 50102 12190 50118
rect 11152 50050 11204 50056
rect 8496 48890 8878 48906
rect 14384 48892 14412 50116
rect 15488 48892 15516 50116
rect 16592 48892 16620 50116
rect 17696 48892 17724 50116
rect 18800 48892 18828 50116
rect 19904 48892 19932 50116
rect 21008 48892 21036 50116
rect 22112 48892 22140 50116
rect 23216 48892 23244 50116
rect 24320 48892 24348 50116
rect 25424 48892 25452 50116
rect 26528 48892 26556 50116
rect 27632 48892 27660 50116
rect 28736 48892 28764 50116
rect 29840 48892 29868 50116
rect 30944 48892 30972 50116
rect 32048 48892 32076 50116
rect 33152 48892 33180 50116
rect 34256 48892 34284 50116
rect 35360 48892 35388 50116
rect 36464 48892 36492 50116
rect 37568 48892 37596 50116
rect 38672 48892 38700 50116
rect 39776 48892 39804 50116
rect 40880 48892 40908 50116
rect 41984 48892 42012 50116
rect 43088 48892 43116 50116
rect 44192 48892 44220 50116
rect 45296 48892 45324 50116
rect 46400 48892 46428 50116
rect 47504 48892 47532 50116
rect 48608 48892 48636 50116
rect 50448 48906 50476 59978
rect 50540 50674 50568 92414
rect 50724 90794 50752 93230
rect 51092 93158 51120 94726
rect 52552 93832 52604 93838
rect 52552 93774 52604 93780
rect 52564 93158 52592 93774
rect 52932 93362 52960 94930
rect 54128 94042 54156 95406
rect 56508 95328 56560 95334
rect 56508 95270 56560 95276
rect 54116 94036 54168 94042
rect 54116 93978 54168 93984
rect 54128 93906 54156 93978
rect 54116 93900 54168 93906
rect 54116 93842 54168 93848
rect 52920 93356 52972 93362
rect 52920 93298 52972 93304
rect 54208 93356 54260 93362
rect 54208 93298 54260 93304
rect 54220 93158 54248 93298
rect 51080 93152 51132 93158
rect 51080 93094 51132 93100
rect 52000 93152 52052 93158
rect 52000 93094 52052 93100
rect 52552 93152 52604 93158
rect 52552 93094 52604 93100
rect 54208 93152 54260 93158
rect 54208 93094 54260 93100
rect 55128 93152 55180 93158
rect 55128 93094 55180 93100
rect 51092 92478 51120 93094
rect 52012 92886 52040 93094
rect 52000 92880 52052 92886
rect 52000 92822 52052 92828
rect 51080 92472 51132 92478
rect 51080 92414 51132 92420
rect 52012 91202 52040 92822
rect 52564 92750 52592 93094
rect 54220 92818 54248 93094
rect 54208 92812 54260 92818
rect 54208 92754 54260 92760
rect 52552 92744 52604 92750
rect 52552 92686 52604 92692
rect 51966 91174 52040 91202
rect 51966 90916 51994 91174
rect 52564 90930 52592 92686
rect 54220 91202 54248 92754
rect 54174 91174 54248 91202
rect 52564 90902 53084 90930
rect 54174 90916 54202 91174
rect 50632 90766 50876 90794
rect 50632 60042 50660 90766
rect 55140 90522 55168 93094
rect 56520 90930 56548 95270
rect 56796 95130 56824 95406
rect 60004 95396 60056 95402
rect 60004 95338 60056 95344
rect 61936 95396 61988 95402
rect 61936 95338 61988 95344
rect 63224 95396 63276 95402
rect 63224 95338 63276 95344
rect 57520 95328 57572 95334
rect 57520 95270 57572 95276
rect 58900 95328 58952 95334
rect 58900 95270 58952 95276
rect 56784 95124 56836 95130
rect 56784 95066 56836 95072
rect 56796 93498 56824 95066
rect 56784 93492 56836 93498
rect 56784 93434 56836 93440
rect 57060 93288 57112 93294
rect 57060 93230 57112 93236
rect 57072 93158 57100 93230
rect 57060 93152 57112 93158
rect 57060 93094 57112 93100
rect 57072 92954 57100 93094
rect 57060 92948 57112 92954
rect 57060 92890 57112 92896
rect 57532 91202 57560 95270
rect 56396 90902 56548 90930
rect 57486 91174 57560 91202
rect 57486 90916 57514 91174
rect 58912 90930 58940 95270
rect 60016 90930 60044 95338
rect 60832 95328 60884 95334
rect 60832 95270 60884 95276
rect 60844 91202 60872 95270
rect 61948 91202 61976 95338
rect 58604 90902 58940 90930
rect 59708 90902 60044 90930
rect 60798 91174 60872 91202
rect 61902 91174 61976 91202
rect 60798 90916 60826 91174
rect 61902 90916 61930 91174
rect 63236 90930 63264 95338
rect 64052 95328 64104 95334
rect 64052 95270 64104 95276
rect 65248 95328 65300 95334
rect 65248 95270 65300 95276
rect 64064 91202 64092 95270
rect 65260 91202 65288 95270
rect 65654 95228 65962 95237
rect 65654 95226 65660 95228
rect 65716 95226 65740 95228
rect 65796 95226 65820 95228
rect 65876 95226 65900 95228
rect 65956 95226 65962 95228
rect 65716 95174 65718 95226
rect 65898 95174 65900 95226
rect 65654 95172 65660 95174
rect 65716 95172 65740 95174
rect 65796 95172 65820 95174
rect 65876 95172 65900 95174
rect 65956 95172 65962 95174
rect 65654 95163 65962 95172
rect 66314 94684 66622 94693
rect 66314 94682 66320 94684
rect 66376 94682 66400 94684
rect 66456 94682 66480 94684
rect 66536 94682 66560 94684
rect 66616 94682 66622 94684
rect 66376 94630 66378 94682
rect 66558 94630 66560 94682
rect 66314 94628 66320 94630
rect 66376 94628 66400 94630
rect 66456 94628 66480 94630
rect 66536 94628 66560 94630
rect 66616 94628 66622 94630
rect 66314 94619 66622 94628
rect 65654 94140 65962 94149
rect 65654 94138 65660 94140
rect 65716 94138 65740 94140
rect 65796 94138 65820 94140
rect 65876 94138 65900 94140
rect 65956 94138 65962 94140
rect 65716 94086 65718 94138
rect 65898 94086 65900 94138
rect 65654 94084 65660 94086
rect 65716 94084 65740 94086
rect 65796 94084 65820 94086
rect 65876 94084 65900 94086
rect 65956 94084 65962 94086
rect 65654 94075 65962 94084
rect 66314 93596 66622 93605
rect 66314 93594 66320 93596
rect 66376 93594 66400 93596
rect 66456 93594 66480 93596
rect 66536 93594 66560 93596
rect 66616 93594 66622 93596
rect 66376 93542 66378 93594
rect 66558 93542 66560 93594
rect 66314 93540 66320 93542
rect 66376 93540 66400 93542
rect 66456 93540 66480 93542
rect 66536 93540 66560 93542
rect 66616 93540 66622 93542
rect 66314 93531 66622 93540
rect 65654 93052 65962 93061
rect 65654 93050 65660 93052
rect 65716 93050 65740 93052
rect 65796 93050 65820 93052
rect 65876 93050 65900 93052
rect 65956 93050 65962 93052
rect 65716 92998 65718 93050
rect 65898 92998 65900 93050
rect 65654 92996 65660 92998
rect 65716 92996 65740 92998
rect 65796 92996 65820 92998
rect 65876 92996 65900 92998
rect 65956 92996 65962 92998
rect 65654 92987 65962 92996
rect 64064 91174 64138 91202
rect 63020 90902 63264 90930
rect 64110 90916 64138 91174
rect 65214 91174 65288 91202
rect 65214 90916 65242 91174
rect 66732 90930 66760 95406
rect 67468 91202 67496 95406
rect 68836 95328 68888 95334
rect 68836 95270 68888 95276
rect 69664 95328 69716 95334
rect 69664 95270 69716 95276
rect 70952 95328 71004 95334
rect 70952 95270 71004 95276
rect 71780 95328 71832 95334
rect 71780 95270 71832 95276
rect 73068 95328 73120 95334
rect 73068 95270 73120 95276
rect 66332 90902 66760 90930
rect 67422 91174 67496 91202
rect 67422 90916 67450 91174
rect 68848 90930 68876 95270
rect 69676 91202 69704 95270
rect 68540 90902 68876 90930
rect 69630 91174 69704 91202
rect 69630 90916 69658 91174
rect 70964 90930 70992 95270
rect 71792 91202 71820 95270
rect 71792 91174 71866 91202
rect 70748 90902 70992 90930
rect 71838 90916 71866 91174
rect 73080 90930 73108 95270
rect 74184 90930 74212 95474
rect 75472 90930 75500 95474
rect 76392 90930 76420 95474
rect 77404 91202 77432 95474
rect 72956 90902 73108 90930
rect 74060 90902 74212 90930
rect 75164 90902 75500 90930
rect 76268 90902 76420 90930
rect 77358 91174 77432 91202
rect 77358 90916 77386 91174
rect 78600 90930 78628 95474
rect 79612 91202 79640 95474
rect 78476 90902 78628 90930
rect 79566 91174 79640 91202
rect 80624 91202 80652 95474
rect 80624 91174 80698 91202
rect 79566 90916 79594 91174
rect 80670 90916 80698 91174
rect 81912 90930 81940 95474
rect 83200 90930 83228 95474
rect 84120 90930 84148 95474
rect 85132 91202 85160 95474
rect 81788 90902 81940 90930
rect 82892 90902 83228 90930
rect 83996 90902 84148 90930
rect 85086 91174 85160 91202
rect 85086 90916 85114 91174
rect 86420 90930 86448 95474
rect 87340 91202 87368 95474
rect 86204 90902 86448 90930
rect 87294 91174 87368 91202
rect 88352 91202 88380 95474
rect 88352 91174 88426 91202
rect 87294 90916 87322 91174
rect 88398 90916 88426 91174
rect 89640 90930 89668 95474
rect 90928 90930 90956 95474
rect 96374 95228 96682 95237
rect 96374 95226 96380 95228
rect 96436 95226 96460 95228
rect 96516 95226 96540 95228
rect 96596 95226 96620 95228
rect 96676 95226 96682 95228
rect 96436 95174 96438 95226
rect 96618 95174 96620 95226
rect 96374 95172 96380 95174
rect 96436 95172 96460 95174
rect 96516 95172 96540 95174
rect 96596 95172 96620 95174
rect 96676 95172 96682 95174
rect 96374 95163 96682 95172
rect 97034 94684 97342 94693
rect 97034 94682 97040 94684
rect 97096 94682 97120 94684
rect 97176 94682 97200 94684
rect 97256 94682 97280 94684
rect 97336 94682 97342 94684
rect 97096 94630 97098 94682
rect 97278 94630 97280 94682
rect 97034 94628 97040 94630
rect 97096 94628 97120 94630
rect 97176 94628 97200 94630
rect 97256 94628 97280 94630
rect 97336 94628 97342 94630
rect 97034 94619 97342 94628
rect 96374 94140 96682 94149
rect 96374 94138 96380 94140
rect 96436 94138 96460 94140
rect 96516 94138 96540 94140
rect 96596 94138 96620 94140
rect 96676 94138 96682 94140
rect 96436 94086 96438 94138
rect 96618 94086 96620 94138
rect 96374 94084 96380 94086
rect 96436 94084 96460 94086
rect 96516 94084 96540 94086
rect 96596 94084 96620 94086
rect 96676 94084 96682 94086
rect 96374 94075 96682 94084
rect 91652 93900 91704 93906
rect 91652 93842 91704 93848
rect 89516 90902 89668 90930
rect 90620 90902 90956 90930
rect 55140 90506 55292 90522
rect 55128 90500 55292 90506
rect 55180 90494 55292 90500
rect 55128 90442 55180 90448
rect 50620 60036 50672 60042
rect 50620 59978 50672 59984
rect 50540 50646 50876 50674
rect 52932 50250 53420 50266
rect 52932 50244 53432 50250
rect 52932 50238 53380 50244
rect 52276 50176 52328 50182
rect 51980 50124 52276 50130
rect 51980 50118 52328 50124
rect 51980 50102 52316 50118
rect 52932 50114 52960 50238
rect 53380 50186 53432 50192
rect 56244 50238 56396 50266
rect 57348 50238 57500 50266
rect 58452 50238 58604 50266
rect 59556 50238 59708 50266
rect 60812 50238 60964 50266
rect 61916 50238 62068 50266
rect 63020 50238 63172 50266
rect 64124 50238 64276 50266
rect 65228 50238 65380 50266
rect 66332 50238 66484 50266
rect 67436 50238 67588 50266
rect 68540 50238 68692 50266
rect 69644 50238 69796 50266
rect 70748 50238 70900 50266
rect 71852 50238 72004 50266
rect 72956 50238 73108 50266
rect 74060 50238 74212 50266
rect 75164 50238 75316 50266
rect 76268 50238 76420 50266
rect 77372 50238 77524 50266
rect 78476 50238 78628 50266
rect 79580 50238 79732 50266
rect 80684 50238 80836 50266
rect 81788 50238 81940 50266
rect 82892 50238 83044 50266
rect 83996 50238 84148 50266
rect 85100 50238 85252 50266
rect 86204 50238 86356 50266
rect 87308 50238 87460 50266
rect 88412 50238 88564 50266
rect 52920 50108 52972 50114
rect 54188 50102 54524 50130
rect 52920 50050 52972 50056
rect 54496 50046 54524 50102
rect 54484 50040 54536 50046
rect 54484 49982 54536 49988
rect 8484 48884 8878 48890
rect 8536 48878 8878 48884
rect 50448 48878 50876 48906
rect 8484 48826 8536 48832
rect 12900 48816 12952 48822
rect 12952 48764 13294 48770
rect 12900 48758 13294 48764
rect 11152 48748 11204 48754
rect 12912 48742 13294 48758
rect 11152 48690 11204 48696
rect 10232 48680 10284 48686
rect 9982 48628 10232 48634
rect 9982 48622 10284 48628
rect 9982 48606 10272 48622
rect 11164 48498 11192 48690
rect 11900 48618 12190 48634
rect 11888 48612 12190 48618
rect 11940 48606 12190 48612
rect 11888 48554 11940 48560
rect 50344 48544 50396 48550
rect 11086 48482 11376 48498
rect 50344 48486 50396 48492
rect 11086 48476 11388 48482
rect 11086 48470 11336 48476
rect 11336 48418 11388 48424
rect 8298 44432 8354 44441
rect 8298 44367 8300 44376
rect 8352 44367 8354 44376
rect 8300 44338 8352 44344
rect 8298 43344 8354 43353
rect 8298 43279 8300 43288
rect 8352 43279 8354 43288
rect 8300 43250 8352 43256
rect 8300 42696 8352 42702
rect 8298 42664 8300 42673
rect 8352 42664 8354 42673
rect 8298 42599 8354 42608
rect 8298 41168 8354 41177
rect 8298 41103 8300 41112
rect 8352 41103 8354 41112
rect 8300 41074 8352 41080
rect 8298 38992 8354 39001
rect 8298 38927 8300 38936
rect 8352 38927 8354 38936
rect 8300 38898 8352 38904
rect 8298 37904 8354 37913
rect 8298 37839 8300 37848
rect 8352 37839 8354 37848
rect 8300 37810 8352 37816
rect 8300 37256 8352 37262
rect 8298 37224 8300 37233
rect 8352 37224 8354 37233
rect 8298 37159 8354 37168
rect 8298 35728 8354 35737
rect 8298 35663 8300 35672
rect 8352 35663 8354 35672
rect 8300 35634 8352 35640
rect 8298 33552 8354 33561
rect 8298 33487 8300 33496
rect 8352 33487 8354 33496
rect 8300 33458 8352 33464
rect 8298 32464 8354 32473
rect 8298 32399 8300 32408
rect 8352 32399 8354 32408
rect 8300 32370 8352 32376
rect 8298 30288 8354 30297
rect 8298 30223 8300 30232
rect 8352 30223 8354 30232
rect 8300 30194 8352 30200
rect 8300 29640 8352 29646
rect 8298 29608 8300 29617
rect 8352 29608 8354 29617
rect 8298 29543 8354 29552
rect 8300 28212 8352 28218
rect 8300 28154 8352 28160
rect 8312 28121 8340 28154
rect 8298 28112 8354 28121
rect 8298 28047 8354 28056
rect 8298 27024 8354 27033
rect 8298 26959 8300 26968
rect 8352 26959 8354 26968
rect 8300 26930 8352 26936
rect 8298 24848 8354 24857
rect 8298 24783 8300 24792
rect 8352 24783 8354 24792
rect 8300 24754 8352 24760
rect 8300 24132 8352 24138
rect 8300 24074 8352 24080
rect 8312 24041 8340 24074
rect 8298 24032 8354 24041
rect 8298 23967 8354 23976
rect 8298 22672 8354 22681
rect 8298 22607 8300 22616
rect 8352 22607 8354 22616
rect 8300 22578 8352 22584
rect 8298 21584 8354 21593
rect 8298 21519 8300 21528
rect 8352 21519 8354 21528
rect 8300 21490 8352 21496
rect 8300 19236 8352 19242
rect 8300 19178 8352 19184
rect 8312 19009 8340 19178
rect 8298 19000 8354 19009
rect 8298 18935 8354 18944
rect 8300 18692 8352 18698
rect 8300 18634 8352 18640
rect 8312 18601 8340 18634
rect 8298 18592 8354 18601
rect 8298 18527 8354 18536
rect 8300 17332 8352 17338
rect 8300 17274 8352 17280
rect 8312 17241 8340 17274
rect 8298 17232 8354 17241
rect 8298 17167 8354 17176
rect 8300 16244 8352 16250
rect 8300 16186 8352 16192
rect 8312 16153 8340 16186
rect 8298 16144 8354 16153
rect 8298 16079 8354 16088
rect 8298 13968 8354 13977
rect 8298 13903 8300 13912
rect 8352 13903 8354 13912
rect 8300 13874 8352 13880
rect 8300 13456 8352 13462
rect 8300 13398 8352 13404
rect 8312 13297 8340 13398
rect 8298 13288 8354 13297
rect 8298 13223 8354 13232
rect 8300 11892 8352 11898
rect 8300 11834 8352 11840
rect 8312 11801 8340 11834
rect 8298 11792 8354 11801
rect 8298 11727 8354 11736
rect 8878 8634 9168 8650
rect 50356 8634 50384 48486
rect 8878 8628 9180 8634
rect 8878 8622 9128 8628
rect 8208 8288 8260 8294
rect 8208 8230 8260 8236
rect 8116 8220 8168 8226
rect 8116 8162 8168 8168
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 8024 8152 8076 8158
rect 8024 8094 8076 8100
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 8956 5914 8984 8622
rect 9128 8570 9180 8576
rect 50344 8628 50396 8634
rect 50344 8570 50396 8576
rect 9680 8288 9732 8294
rect 9732 8236 10088 8242
rect 9680 8230 10088 8236
rect 9692 8214 10088 8230
rect 11086 8226 11192 8242
rect 11086 8220 11204 8226
rect 11086 8214 11152 8220
rect 8944 5908 8996 5914
rect 8944 5850 8996 5856
rect 10060 5778 10088 8214
rect 11152 8162 11204 8168
rect 10048 5772 10100 5778
rect 10048 5714 10100 5720
rect 10968 5772 11020 5778
rect 10968 5714 11020 5720
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 10980 2650 11008 5714
rect 11164 5710 11192 8162
rect 11796 8152 11848 8158
rect 11848 8100 12190 8106
rect 11796 8094 12190 8100
rect 11808 8092 12190 8094
rect 11808 8078 12204 8092
rect 14398 8078 14596 8106
rect 15502 8078 15608 8106
rect 16606 8078 16896 8106
rect 17710 8078 17816 8106
rect 12176 5914 12204 8078
rect 12164 5908 12216 5914
rect 12164 5850 12216 5856
rect 12808 5908 12860 5914
rect 12808 5850 12860 5856
rect 11152 5704 11204 5710
rect 11152 5646 11204 5652
rect 12820 5642 12848 5850
rect 13176 5704 13228 5710
rect 13176 5646 13228 5652
rect 12808 5636 12860 5642
rect 12808 5578 12860 5584
rect 11612 3052 11664 3058
rect 11612 2994 11664 3000
rect 11624 2854 11652 2994
rect 11612 2848 11664 2854
rect 11612 2790 11664 2796
rect 10968 2644 11020 2650
rect 10968 2586 11020 2592
rect 10324 2440 10376 2446
rect 10324 2382 10376 2388
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 10336 800 10364 2382
rect 11624 800 11652 2790
rect 12820 2514 12848 5578
rect 13188 3194 13216 5646
rect 13176 3188 13228 3194
rect 13176 3130 13228 3136
rect 12808 2508 12860 2514
rect 12808 2450 12860 2456
rect 14568 2446 14596 8078
rect 15580 2446 15608 8078
rect 16868 2446 16896 8078
rect 17788 2446 17816 8078
rect 18800 2446 18828 8092
rect 19918 8078 20116 8106
rect 20088 2446 20116 8078
rect 21008 2446 21036 8092
rect 22126 8078 22324 8106
rect 23230 8078 23336 8106
rect 24334 8078 24624 8106
rect 25438 8078 25544 8106
rect 22296 2446 22324 8078
rect 23308 2446 23336 8078
rect 24596 2446 24624 8078
rect 25516 2446 25544 8078
rect 26528 2446 26556 8092
rect 27646 8078 27844 8106
rect 28750 8078 29132 8106
rect 29854 8078 30052 8106
rect 30958 8078 31064 8106
rect 32062 8078 32352 8106
rect 27816 2446 27844 8078
rect 29104 2446 29132 8078
rect 30024 2446 30052 8078
rect 31036 2446 31064 8078
rect 32324 2650 32352 8078
rect 33152 2650 33180 8092
rect 34256 2650 34284 8092
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 35360 2650 35388 8092
rect 35594 5468 35902 5477
rect 35594 5466 35600 5468
rect 35656 5466 35680 5468
rect 35736 5466 35760 5468
rect 35816 5466 35840 5468
rect 35896 5466 35902 5468
rect 35656 5414 35658 5466
rect 35838 5414 35840 5466
rect 35594 5412 35600 5414
rect 35656 5412 35680 5414
rect 35736 5412 35760 5414
rect 35816 5412 35840 5414
rect 35896 5412 35902 5414
rect 35594 5403 35902 5412
rect 35594 4380 35902 4389
rect 35594 4378 35600 4380
rect 35656 4378 35680 4380
rect 35736 4378 35760 4380
rect 35816 4378 35840 4380
rect 35896 4378 35902 4380
rect 35656 4326 35658 4378
rect 35838 4326 35840 4378
rect 35594 4324 35600 4326
rect 35656 4324 35680 4326
rect 35736 4324 35760 4326
rect 35816 4324 35840 4326
rect 35896 4324 35902 4326
rect 35594 4315 35902 4324
rect 35594 3292 35902 3301
rect 35594 3290 35600 3292
rect 35656 3290 35680 3292
rect 35736 3290 35760 3292
rect 35816 3290 35840 3292
rect 35896 3290 35902 3292
rect 35656 3238 35658 3290
rect 35838 3238 35840 3290
rect 35594 3236 35600 3238
rect 35656 3236 35680 3238
rect 35736 3236 35760 3238
rect 35816 3236 35840 3238
rect 35896 3236 35902 3238
rect 35594 3227 35902 3236
rect 36464 2650 36492 8092
rect 37582 8078 37688 8106
rect 38686 8078 38792 8106
rect 39790 8078 40080 8106
rect 37660 2650 37688 8078
rect 38764 2650 38792 8078
rect 40052 2650 40080 8078
rect 40880 2650 40908 8092
rect 41984 2650 42012 8092
rect 43102 8078 43300 8106
rect 43272 2650 43300 8078
rect 32312 2644 32364 2650
rect 32312 2586 32364 2592
rect 33140 2644 33192 2650
rect 33140 2586 33192 2592
rect 34244 2644 34296 2650
rect 34244 2586 34296 2592
rect 35348 2644 35400 2650
rect 35348 2586 35400 2592
rect 36452 2644 36504 2650
rect 36452 2586 36504 2592
rect 37648 2644 37700 2650
rect 37648 2586 37700 2592
rect 38752 2644 38804 2650
rect 38752 2586 38804 2592
rect 40040 2644 40092 2650
rect 40040 2586 40092 2592
rect 40868 2644 40920 2650
rect 40868 2586 40920 2592
rect 41972 2644 42024 2650
rect 41972 2586 42024 2592
rect 43260 2644 43312 2650
rect 43260 2586 43312 2592
rect 44192 2582 44220 8092
rect 45310 8078 45508 8106
rect 44180 2576 44232 2582
rect 44180 2518 44232 2524
rect 45480 2514 45508 8078
rect 46400 2514 46428 8092
rect 47504 2514 47532 8092
rect 48622 8078 48820 8106
rect 48792 2650 48820 8078
rect 50632 5914 50660 48878
rect 52276 48816 52328 48822
rect 51828 48764 52276 48770
rect 56244 48770 56272 50238
rect 57348 48770 57376 50238
rect 58452 48770 58480 50238
rect 59556 48770 59584 50238
rect 51828 48758 52328 48764
rect 51828 48742 52316 48758
rect 55292 48754 55628 48770
rect 55292 48748 55640 48754
rect 55292 48742 55588 48748
rect 51828 48686 51856 48742
rect 51816 48680 51868 48686
rect 54484 48680 54536 48686
rect 51816 48622 51868 48628
rect 54036 48628 54484 48634
rect 54036 48622 54536 48628
rect 54036 48618 54524 48622
rect 54024 48612 54524 48618
rect 54076 48606 54524 48612
rect 54024 48554 54076 48560
rect 55416 48550 55444 48742
rect 56244 48742 56396 48770
rect 57348 48742 57500 48770
rect 58452 48742 58604 48770
rect 59556 48742 59708 48770
rect 55588 48690 55640 48696
rect 60936 48634 60964 50238
rect 62040 48634 62068 50238
rect 63144 48770 63172 50238
rect 64248 48770 64276 50238
rect 65352 48770 65380 50238
rect 66456 48770 66484 50238
rect 63020 48742 63172 48770
rect 64124 48742 64276 48770
rect 65228 48742 65380 48770
rect 66332 48742 66484 48770
rect 67560 48634 67588 50238
rect 68664 48770 68692 50238
rect 69768 48770 69796 50238
rect 70872 48770 70900 50238
rect 71976 48770 72004 50238
rect 73080 48770 73108 50238
rect 68540 48742 68692 48770
rect 69644 48742 69796 48770
rect 70748 48742 70900 48770
rect 71852 48742 72004 48770
rect 72956 48742 73108 48770
rect 74184 48634 74212 50238
rect 75288 48634 75316 50238
rect 76392 48770 76420 50238
rect 77496 48770 77524 50238
rect 78600 48770 78628 50238
rect 79704 48770 79732 50238
rect 80808 48770 80836 50238
rect 81912 48770 81940 50238
rect 83016 48770 83044 50238
rect 84120 48770 84148 50238
rect 76268 48742 76420 48770
rect 77372 48742 77524 48770
rect 78476 48742 78628 48770
rect 79580 48742 79732 48770
rect 80684 48742 80836 48770
rect 81788 48742 81940 48770
rect 82892 48742 83044 48770
rect 83996 48742 84148 48770
rect 85224 48634 85252 50238
rect 86328 48770 86356 50238
rect 86204 48742 86356 48770
rect 87432 48634 87460 50238
rect 88536 48634 88564 50238
rect 60812 48606 60964 48634
rect 61916 48606 62068 48634
rect 67436 48606 67588 48634
rect 74060 48606 74212 48634
rect 75164 48606 75316 48634
rect 85100 48606 85252 48634
rect 87308 48606 87460 48634
rect 88412 48606 88564 48634
rect 89364 50238 89516 50266
rect 90468 50238 90620 50266
rect 89364 48634 89392 50238
rect 90468 48770 90496 50238
rect 90468 48742 90620 48770
rect 89364 48606 89516 48634
rect 91664 48550 91692 93842
rect 97034 93596 97342 93605
rect 97034 93594 97040 93596
rect 97096 93594 97120 93596
rect 97176 93594 97200 93596
rect 97256 93594 97280 93596
rect 97336 93594 97342 93596
rect 97096 93542 97098 93594
rect 97278 93542 97280 93594
rect 97034 93540 97040 93542
rect 97096 93540 97120 93542
rect 97176 93540 97200 93542
rect 97256 93540 97280 93542
rect 97336 93540 97342 93542
rect 97034 93531 97342 93540
rect 91744 93152 91796 93158
rect 91744 93094 91796 93100
rect 91756 48822 91784 93094
rect 96374 93052 96682 93061
rect 96374 93050 96380 93052
rect 96436 93050 96460 93052
rect 96516 93050 96540 93052
rect 96596 93050 96620 93052
rect 96676 93050 96682 93052
rect 96436 92998 96438 93050
rect 96618 92998 96620 93050
rect 96374 92996 96380 92998
rect 96436 92996 96460 92998
rect 96516 92996 96540 92998
rect 96596 92996 96620 92998
rect 96676 92996 96682 92998
rect 96374 92987 96682 92996
rect 91836 92948 91888 92954
rect 91836 92890 91888 92896
rect 91744 48816 91796 48822
rect 91744 48758 91796 48764
rect 91848 48686 91876 92890
rect 97034 92508 97342 92517
rect 97034 92506 97040 92508
rect 97096 92506 97120 92508
rect 97176 92506 97200 92508
rect 97256 92506 97280 92508
rect 97336 92506 97342 92508
rect 97096 92454 97098 92506
rect 97278 92454 97280 92506
rect 97034 92452 97040 92454
rect 97096 92452 97120 92454
rect 97176 92452 97200 92454
rect 97256 92452 97280 92454
rect 97336 92452 97342 92454
rect 97034 92443 97342 92452
rect 96374 91964 96682 91973
rect 96374 91962 96380 91964
rect 96436 91962 96460 91964
rect 96516 91962 96540 91964
rect 96596 91962 96620 91964
rect 96676 91962 96682 91964
rect 96436 91910 96438 91962
rect 96618 91910 96620 91962
rect 96374 91908 96380 91910
rect 96436 91908 96460 91910
rect 96516 91908 96540 91910
rect 96596 91908 96620 91910
rect 96676 91908 96682 91910
rect 96374 91899 96682 91908
rect 97034 91420 97342 91429
rect 97034 91418 97040 91420
rect 97096 91418 97120 91420
rect 97176 91418 97200 91420
rect 97256 91418 97280 91420
rect 97336 91418 97342 91420
rect 97096 91366 97098 91418
rect 97278 91366 97280 91418
rect 97034 91364 97040 91366
rect 97096 91364 97120 91366
rect 97176 91364 97200 91366
rect 97256 91364 97280 91366
rect 97336 91364 97342 91366
rect 97034 91355 97342 91364
rect 96374 90876 96682 90885
rect 96374 90874 96380 90876
rect 96436 90874 96460 90876
rect 96516 90874 96540 90876
rect 96596 90874 96620 90876
rect 96676 90874 96682 90876
rect 96436 90822 96438 90874
rect 96618 90822 96620 90874
rect 96374 90820 96380 90822
rect 96436 90820 96460 90822
rect 96516 90820 96540 90822
rect 96596 90820 96620 90822
rect 96676 90820 96682 90822
rect 96374 90811 96682 90820
rect 97034 90332 97342 90341
rect 97034 90330 97040 90332
rect 97096 90330 97120 90332
rect 97176 90330 97200 90332
rect 97256 90330 97280 90332
rect 97336 90330 97342 90332
rect 97096 90278 97098 90330
rect 97278 90278 97280 90330
rect 97034 90276 97040 90278
rect 97096 90276 97120 90278
rect 97176 90276 97200 90278
rect 97256 90276 97280 90278
rect 97336 90276 97342 90278
rect 97034 90267 97342 90276
rect 96374 89788 96682 89797
rect 96374 89786 96380 89788
rect 96436 89786 96460 89788
rect 96516 89786 96540 89788
rect 96596 89786 96620 89788
rect 96676 89786 96682 89788
rect 96436 89734 96438 89786
rect 96618 89734 96620 89786
rect 96374 89732 96380 89734
rect 96436 89732 96460 89734
rect 96516 89732 96540 89734
rect 96596 89732 96620 89734
rect 96676 89732 96682 89734
rect 96374 89723 96682 89732
rect 97034 89244 97342 89253
rect 97034 89242 97040 89244
rect 97096 89242 97120 89244
rect 97176 89242 97200 89244
rect 97256 89242 97280 89244
rect 97336 89242 97342 89244
rect 97096 89190 97098 89242
rect 97278 89190 97280 89242
rect 97034 89188 97040 89190
rect 97096 89188 97120 89190
rect 97176 89188 97200 89190
rect 97256 89188 97280 89190
rect 97336 89188 97342 89190
rect 97034 89179 97342 89188
rect 96374 88700 96682 88709
rect 96374 88698 96380 88700
rect 96436 88698 96460 88700
rect 96516 88698 96540 88700
rect 96596 88698 96620 88700
rect 96676 88698 96682 88700
rect 96436 88646 96438 88698
rect 96618 88646 96620 88698
rect 96374 88644 96380 88646
rect 96436 88644 96460 88646
rect 96516 88644 96540 88646
rect 96596 88644 96620 88646
rect 96676 88644 96682 88646
rect 96374 88635 96682 88644
rect 97034 88156 97342 88165
rect 97034 88154 97040 88156
rect 97096 88154 97120 88156
rect 97176 88154 97200 88156
rect 97256 88154 97280 88156
rect 97336 88154 97342 88156
rect 97096 88102 97098 88154
rect 97278 88102 97280 88154
rect 97034 88100 97040 88102
rect 97096 88100 97120 88102
rect 97176 88100 97200 88102
rect 97256 88100 97280 88102
rect 97336 88100 97342 88102
rect 97034 88091 97342 88100
rect 96374 87612 96682 87621
rect 96374 87610 96380 87612
rect 96436 87610 96460 87612
rect 96516 87610 96540 87612
rect 96596 87610 96620 87612
rect 96676 87610 96682 87612
rect 96436 87558 96438 87610
rect 96618 87558 96620 87610
rect 96374 87556 96380 87558
rect 96436 87556 96460 87558
rect 96516 87556 96540 87558
rect 96596 87556 96620 87558
rect 96676 87556 96682 87558
rect 96374 87547 96682 87556
rect 97356 87440 97408 87446
rect 97354 87408 97356 87417
rect 97408 87408 97410 87417
rect 97354 87343 97410 87352
rect 97540 87304 97592 87310
rect 97540 87246 97592 87252
rect 97552 87145 97580 87246
rect 97538 87136 97594 87145
rect 97034 87068 97342 87077
rect 97538 87071 97594 87080
rect 97034 87066 97040 87068
rect 97096 87066 97120 87068
rect 97176 87066 97200 87068
rect 97256 87066 97280 87068
rect 97336 87066 97342 87068
rect 97096 87014 97098 87066
rect 97278 87014 97280 87066
rect 97034 87012 97040 87014
rect 97096 87012 97120 87014
rect 97176 87012 97200 87014
rect 97256 87012 97280 87014
rect 97336 87012 97342 87014
rect 97034 87003 97342 87012
rect 97540 86828 97592 86834
rect 97540 86770 97592 86776
rect 97356 86624 97408 86630
rect 97356 86566 97408 86572
rect 96374 86524 96682 86533
rect 96374 86522 96380 86524
rect 96436 86522 96460 86524
rect 96516 86522 96540 86524
rect 96596 86522 96620 86524
rect 96676 86522 96682 86524
rect 96436 86470 96438 86522
rect 96618 86470 96620 86522
rect 96374 86468 96380 86470
rect 96436 86468 96460 86470
rect 96516 86468 96540 86470
rect 96596 86468 96620 86470
rect 96676 86468 96682 86470
rect 96374 86459 96682 86468
rect 97368 86329 97396 86566
rect 97552 86465 97580 86770
rect 97538 86456 97594 86465
rect 97538 86391 97594 86400
rect 97354 86320 97410 86329
rect 97354 86255 97410 86264
rect 97034 85980 97342 85989
rect 97034 85978 97040 85980
rect 97096 85978 97120 85980
rect 97176 85978 97200 85980
rect 97256 85978 97280 85980
rect 97336 85978 97342 85980
rect 97096 85926 97098 85978
rect 97278 85926 97280 85978
rect 97034 85924 97040 85926
rect 97096 85924 97120 85926
rect 97176 85924 97200 85926
rect 97256 85924 97280 85926
rect 97336 85924 97342 85926
rect 97034 85915 97342 85924
rect 96374 85436 96682 85445
rect 96374 85434 96380 85436
rect 96436 85434 96460 85436
rect 96516 85434 96540 85436
rect 96596 85434 96620 85436
rect 96676 85434 96682 85436
rect 96436 85382 96438 85434
rect 96618 85382 96620 85434
rect 96374 85380 96380 85382
rect 96436 85380 96460 85382
rect 96516 85380 96540 85382
rect 96596 85380 96620 85382
rect 96676 85380 96682 85382
rect 96374 85371 96682 85380
rect 97356 85264 97408 85270
rect 97354 85232 97356 85241
rect 97408 85232 97410 85241
rect 97354 85167 97410 85176
rect 97540 85128 97592 85134
rect 97538 85096 97540 85105
rect 97592 85096 97594 85105
rect 97538 85031 97594 85040
rect 97034 84892 97342 84901
rect 97034 84890 97040 84892
rect 97096 84890 97120 84892
rect 97176 84890 97200 84892
rect 97256 84890 97280 84892
rect 97336 84890 97342 84892
rect 97096 84838 97098 84890
rect 97278 84838 97280 84890
rect 97034 84836 97040 84838
rect 97096 84836 97120 84838
rect 97176 84836 97200 84838
rect 97256 84836 97280 84838
rect 97336 84836 97342 84838
rect 97034 84827 97342 84836
rect 97540 84652 97592 84658
rect 97540 84594 97592 84600
rect 97356 84448 97408 84454
rect 97552 84425 97580 84594
rect 97356 84390 97408 84396
rect 97538 84416 97594 84425
rect 96374 84348 96682 84357
rect 96374 84346 96380 84348
rect 96436 84346 96460 84348
rect 96516 84346 96540 84348
rect 96596 84346 96620 84348
rect 96676 84346 96682 84348
rect 96436 84294 96438 84346
rect 96618 84294 96620 84346
rect 96374 84292 96380 84294
rect 96436 84292 96460 84294
rect 96516 84292 96540 84294
rect 96596 84292 96620 84294
rect 96676 84292 96682 84294
rect 96374 84283 96682 84292
rect 97368 84153 97396 84390
rect 97538 84351 97594 84360
rect 97354 84144 97410 84153
rect 97354 84079 97410 84088
rect 97034 83804 97342 83813
rect 97034 83802 97040 83804
rect 97096 83802 97120 83804
rect 97176 83802 97200 83804
rect 97256 83802 97280 83804
rect 97336 83802 97342 83804
rect 97096 83750 97098 83802
rect 97278 83750 97280 83802
rect 97034 83748 97040 83750
rect 97096 83748 97120 83750
rect 97176 83748 97200 83750
rect 97256 83748 97280 83750
rect 97336 83748 97342 83750
rect 97034 83739 97342 83748
rect 97540 83564 97592 83570
rect 97540 83506 97592 83512
rect 97356 83360 97408 83366
rect 97356 83302 97408 83308
rect 96374 83260 96682 83269
rect 96374 83258 96380 83260
rect 96436 83258 96460 83260
rect 96516 83258 96540 83260
rect 96596 83258 96620 83260
rect 96676 83258 96682 83260
rect 96436 83206 96438 83258
rect 96618 83206 96620 83258
rect 96374 83204 96380 83206
rect 96436 83204 96460 83206
rect 96516 83204 96540 83206
rect 96596 83204 96620 83206
rect 96676 83204 96682 83206
rect 96374 83195 96682 83204
rect 97368 83065 97396 83302
rect 97552 83065 97580 83506
rect 97354 83056 97410 83065
rect 97354 82991 97410 83000
rect 97538 83056 97594 83065
rect 97538 82991 97594 83000
rect 97034 82716 97342 82725
rect 97034 82714 97040 82716
rect 97096 82714 97120 82716
rect 97176 82714 97200 82716
rect 97256 82714 97280 82716
rect 97336 82714 97342 82716
rect 97096 82662 97098 82714
rect 97278 82662 97280 82714
rect 97034 82660 97040 82662
rect 97096 82660 97120 82662
rect 97176 82660 97200 82662
rect 97256 82660 97280 82662
rect 97336 82660 97342 82662
rect 97034 82651 97342 82660
rect 96374 82172 96682 82181
rect 96374 82170 96380 82172
rect 96436 82170 96460 82172
rect 96516 82170 96540 82172
rect 96596 82170 96620 82172
rect 96676 82170 96682 82172
rect 96436 82118 96438 82170
rect 96618 82118 96620 82170
rect 96374 82116 96380 82118
rect 96436 82116 96460 82118
rect 96516 82116 96540 82118
rect 96596 82116 96620 82118
rect 96676 82116 96682 82118
rect 96374 82107 96682 82116
rect 97356 82000 97408 82006
rect 97354 81968 97356 81977
rect 97408 81968 97410 81977
rect 97354 81903 97410 81912
rect 97540 81864 97592 81870
rect 97540 81806 97592 81812
rect 97552 81705 97580 81806
rect 97538 81696 97594 81705
rect 97034 81628 97342 81637
rect 97538 81631 97594 81640
rect 97034 81626 97040 81628
rect 97096 81626 97120 81628
rect 97176 81626 97200 81628
rect 97256 81626 97280 81628
rect 97336 81626 97342 81628
rect 97096 81574 97098 81626
rect 97278 81574 97280 81626
rect 97034 81572 97040 81574
rect 97096 81572 97120 81574
rect 97176 81572 97200 81574
rect 97256 81572 97280 81574
rect 97336 81572 97342 81574
rect 97034 81563 97342 81572
rect 97540 81388 97592 81394
rect 97540 81330 97592 81336
rect 97356 81184 97408 81190
rect 97356 81126 97408 81132
rect 96374 81084 96682 81093
rect 96374 81082 96380 81084
rect 96436 81082 96460 81084
rect 96516 81082 96540 81084
rect 96596 81082 96620 81084
rect 96676 81082 96682 81084
rect 96436 81030 96438 81082
rect 96618 81030 96620 81082
rect 96374 81028 96380 81030
rect 96436 81028 96460 81030
rect 96516 81028 96540 81030
rect 96596 81028 96620 81030
rect 96676 81028 96682 81030
rect 96374 81019 96682 81028
rect 97368 80889 97396 81126
rect 97552 81025 97580 81330
rect 97538 81016 97594 81025
rect 97538 80951 97594 80960
rect 97354 80880 97410 80889
rect 97354 80815 97410 80824
rect 97034 80540 97342 80549
rect 97034 80538 97040 80540
rect 97096 80538 97120 80540
rect 97176 80538 97200 80540
rect 97256 80538 97280 80540
rect 97336 80538 97342 80540
rect 97096 80486 97098 80538
rect 97278 80486 97280 80538
rect 97034 80484 97040 80486
rect 97096 80484 97120 80486
rect 97176 80484 97200 80486
rect 97256 80484 97280 80486
rect 97336 80484 97342 80486
rect 97034 80475 97342 80484
rect 96374 79996 96682 80005
rect 96374 79994 96380 79996
rect 96436 79994 96460 79996
rect 96516 79994 96540 79996
rect 96596 79994 96620 79996
rect 96676 79994 96682 79996
rect 96436 79942 96438 79994
rect 96618 79942 96620 79994
rect 96374 79940 96380 79942
rect 96436 79940 96460 79942
rect 96516 79940 96540 79942
rect 96596 79940 96620 79942
rect 96676 79940 96682 79942
rect 96374 79931 96682 79940
rect 97356 79824 97408 79830
rect 97354 79792 97356 79801
rect 97408 79792 97410 79801
rect 97354 79727 97410 79736
rect 97540 79688 97592 79694
rect 97538 79656 97540 79665
rect 97592 79656 97594 79665
rect 97538 79591 97594 79600
rect 97034 79452 97342 79461
rect 97034 79450 97040 79452
rect 97096 79450 97120 79452
rect 97176 79450 97200 79452
rect 97256 79450 97280 79452
rect 97336 79450 97342 79452
rect 97096 79398 97098 79450
rect 97278 79398 97280 79450
rect 97034 79396 97040 79398
rect 97096 79396 97120 79398
rect 97176 79396 97200 79398
rect 97256 79396 97280 79398
rect 97336 79396 97342 79398
rect 97034 79387 97342 79396
rect 97448 79212 97500 79218
rect 97448 79154 97500 79160
rect 97264 79076 97316 79082
rect 97264 79018 97316 79024
rect 96374 78908 96682 78917
rect 96374 78906 96380 78908
rect 96436 78906 96460 78908
rect 96516 78906 96540 78908
rect 96596 78906 96620 78908
rect 96676 78906 96682 78908
rect 96436 78854 96438 78906
rect 96618 78854 96620 78906
rect 96374 78852 96380 78854
rect 96436 78852 96460 78854
rect 96516 78852 96540 78854
rect 96596 78852 96620 78854
rect 96676 78852 96682 78854
rect 96374 78843 96682 78852
rect 97276 78713 97304 79018
rect 97460 78985 97488 79154
rect 97446 78976 97502 78985
rect 97446 78911 97502 78920
rect 97262 78704 97318 78713
rect 97262 78639 97318 78648
rect 97034 78364 97342 78373
rect 97034 78362 97040 78364
rect 97096 78362 97120 78364
rect 97176 78362 97200 78364
rect 97256 78362 97280 78364
rect 97336 78362 97342 78364
rect 97096 78310 97098 78362
rect 97278 78310 97280 78362
rect 97034 78308 97040 78310
rect 97096 78308 97120 78310
rect 97176 78308 97200 78310
rect 97256 78308 97280 78310
rect 97336 78308 97342 78310
rect 97034 78299 97342 78308
rect 97540 78124 97592 78130
rect 97540 78066 97592 78072
rect 97356 77920 97408 77926
rect 97356 77862 97408 77868
rect 96374 77820 96682 77829
rect 96374 77818 96380 77820
rect 96436 77818 96460 77820
rect 96516 77818 96540 77820
rect 96596 77818 96620 77820
rect 96676 77818 96682 77820
rect 96436 77766 96438 77818
rect 96618 77766 96620 77818
rect 96374 77764 96380 77766
rect 96436 77764 96460 77766
rect 96516 77764 96540 77766
rect 96596 77764 96620 77766
rect 96676 77764 96682 77766
rect 96374 77755 96682 77764
rect 97368 77625 97396 77862
rect 97552 77625 97580 78066
rect 97354 77616 97410 77625
rect 97354 77551 97410 77560
rect 97538 77616 97594 77625
rect 97538 77551 97594 77560
rect 97034 77276 97342 77285
rect 97034 77274 97040 77276
rect 97096 77274 97120 77276
rect 97176 77274 97200 77276
rect 97256 77274 97280 77276
rect 97336 77274 97342 77276
rect 97096 77222 97098 77274
rect 97278 77222 97280 77274
rect 97034 77220 97040 77222
rect 97096 77220 97120 77222
rect 97176 77220 97200 77222
rect 97256 77220 97280 77222
rect 97336 77220 97342 77222
rect 97034 77211 97342 77220
rect 96374 76732 96682 76741
rect 96374 76730 96380 76732
rect 96436 76730 96460 76732
rect 96516 76730 96540 76732
rect 96596 76730 96620 76732
rect 96676 76730 96682 76732
rect 96436 76678 96438 76730
rect 96618 76678 96620 76730
rect 96374 76676 96380 76678
rect 96436 76676 96460 76678
rect 96516 76676 96540 76678
rect 96596 76676 96620 76678
rect 96676 76676 96682 76678
rect 96374 76667 96682 76676
rect 97356 76560 97408 76566
rect 97354 76528 97356 76537
rect 97408 76528 97410 76537
rect 97354 76463 97410 76472
rect 97540 76424 97592 76430
rect 97540 76366 97592 76372
rect 97552 76265 97580 76366
rect 97538 76256 97594 76265
rect 97034 76188 97342 76197
rect 97538 76191 97594 76200
rect 97034 76186 97040 76188
rect 97096 76186 97120 76188
rect 97176 76186 97200 76188
rect 97256 76186 97280 76188
rect 97336 76186 97342 76188
rect 97096 76134 97098 76186
rect 97278 76134 97280 76186
rect 97034 76132 97040 76134
rect 97096 76132 97120 76134
rect 97176 76132 97200 76134
rect 97256 76132 97280 76134
rect 97336 76132 97342 76134
rect 97034 76123 97342 76132
rect 97540 75948 97592 75954
rect 97540 75890 97592 75896
rect 97356 75744 97408 75750
rect 97356 75686 97408 75692
rect 96374 75644 96682 75653
rect 96374 75642 96380 75644
rect 96436 75642 96460 75644
rect 96516 75642 96540 75644
rect 96596 75642 96620 75644
rect 96676 75642 96682 75644
rect 96436 75590 96438 75642
rect 96618 75590 96620 75642
rect 96374 75588 96380 75590
rect 96436 75588 96460 75590
rect 96516 75588 96540 75590
rect 96596 75588 96620 75590
rect 96676 75588 96682 75590
rect 96374 75579 96682 75588
rect 97368 75449 97396 75686
rect 97552 75585 97580 75890
rect 97538 75576 97594 75585
rect 97538 75511 97594 75520
rect 97354 75440 97410 75449
rect 97354 75375 97410 75384
rect 97034 75100 97342 75109
rect 97034 75098 97040 75100
rect 97096 75098 97120 75100
rect 97176 75098 97200 75100
rect 97256 75098 97280 75100
rect 97336 75098 97342 75100
rect 97096 75046 97098 75098
rect 97278 75046 97280 75098
rect 97034 75044 97040 75046
rect 97096 75044 97120 75046
rect 97176 75044 97200 75046
rect 97256 75044 97280 75046
rect 97336 75044 97342 75046
rect 97034 75035 97342 75044
rect 96374 74556 96682 74565
rect 96374 74554 96380 74556
rect 96436 74554 96460 74556
rect 96516 74554 96540 74556
rect 96596 74554 96620 74556
rect 96676 74554 96682 74556
rect 96436 74502 96438 74554
rect 96618 74502 96620 74554
rect 96374 74500 96380 74502
rect 96436 74500 96460 74502
rect 96516 74500 96540 74502
rect 96596 74500 96620 74502
rect 96676 74500 96682 74502
rect 96374 74491 96682 74500
rect 97264 74384 97316 74390
rect 97262 74352 97264 74361
rect 97316 74352 97318 74361
rect 97262 74287 97318 74296
rect 97446 74216 97502 74225
rect 97446 74151 97448 74160
rect 97500 74151 97502 74160
rect 97448 74122 97500 74128
rect 97034 74012 97342 74021
rect 97034 74010 97040 74012
rect 97096 74010 97120 74012
rect 97176 74010 97200 74012
rect 97256 74010 97280 74012
rect 97336 74010 97342 74012
rect 97096 73958 97098 74010
rect 97278 73958 97280 74010
rect 97034 73956 97040 73958
rect 97096 73956 97120 73958
rect 97176 73956 97200 73958
rect 97256 73956 97280 73958
rect 97336 73956 97342 73958
rect 97034 73947 97342 73956
rect 97540 73772 97592 73778
rect 97540 73714 97592 73720
rect 97356 73568 97408 73574
rect 97552 73545 97580 73714
rect 97356 73510 97408 73516
rect 97538 73536 97594 73545
rect 96374 73468 96682 73477
rect 96374 73466 96380 73468
rect 96436 73466 96460 73468
rect 96516 73466 96540 73468
rect 96596 73466 96620 73468
rect 96676 73466 96682 73468
rect 96436 73414 96438 73466
rect 96618 73414 96620 73466
rect 96374 73412 96380 73414
rect 96436 73412 96460 73414
rect 96516 73412 96540 73414
rect 96596 73412 96620 73414
rect 96676 73412 96682 73414
rect 96374 73403 96682 73412
rect 97368 73273 97396 73510
rect 97538 73471 97594 73480
rect 97354 73264 97410 73273
rect 97354 73199 97410 73208
rect 97034 72924 97342 72933
rect 97034 72922 97040 72924
rect 97096 72922 97120 72924
rect 97176 72922 97200 72924
rect 97256 72922 97280 72924
rect 97336 72922 97342 72924
rect 97096 72870 97098 72922
rect 97278 72870 97280 72922
rect 97034 72868 97040 72870
rect 97096 72868 97120 72870
rect 97176 72868 97200 72870
rect 97256 72868 97280 72870
rect 97336 72868 97342 72870
rect 97034 72859 97342 72868
rect 97264 72616 97316 72622
rect 97264 72558 97316 72564
rect 97540 72616 97592 72622
rect 97540 72558 97592 72564
rect 96374 72380 96682 72389
rect 96374 72378 96380 72380
rect 96436 72378 96460 72380
rect 96516 72378 96540 72380
rect 96596 72378 96620 72380
rect 96676 72378 96682 72380
rect 96436 72326 96438 72378
rect 96618 72326 96620 72378
rect 96374 72324 96380 72326
rect 96436 72324 96460 72326
rect 96516 72324 96540 72326
rect 96596 72324 96620 72326
rect 96676 72324 96682 72326
rect 96374 72315 96682 72324
rect 97276 72185 97304 72558
rect 97552 72214 97580 72558
rect 97540 72208 97592 72214
rect 97262 72176 97318 72185
rect 97262 72111 97318 72120
rect 97538 72176 97540 72185
rect 97592 72176 97594 72185
rect 97538 72111 97594 72120
rect 97034 71836 97342 71845
rect 97034 71834 97040 71836
rect 97096 71834 97120 71836
rect 97176 71834 97200 71836
rect 97256 71834 97280 71836
rect 97336 71834 97342 71836
rect 97096 71782 97098 71834
rect 97278 71782 97280 71834
rect 97034 71780 97040 71782
rect 97096 71780 97120 71782
rect 97176 71780 97200 71782
rect 97256 71780 97280 71782
rect 97336 71780 97342 71782
rect 97034 71771 97342 71780
rect 96374 71292 96682 71301
rect 96374 71290 96380 71292
rect 96436 71290 96460 71292
rect 96516 71290 96540 71292
rect 96596 71290 96620 71292
rect 96676 71290 96682 71292
rect 96436 71238 96438 71290
rect 96618 71238 96620 71290
rect 96374 71236 96380 71238
rect 96436 71236 96460 71238
rect 96516 71236 96540 71238
rect 96596 71236 96620 71238
rect 96676 71236 96682 71238
rect 96374 71227 96682 71236
rect 97356 71120 97408 71126
rect 97354 71088 97356 71097
rect 97408 71088 97410 71097
rect 97354 71023 97410 71032
rect 97540 70984 97592 70990
rect 97540 70926 97592 70932
rect 97552 70825 97580 70926
rect 97538 70816 97594 70825
rect 97034 70748 97342 70757
rect 97538 70751 97594 70760
rect 97034 70746 97040 70748
rect 97096 70746 97120 70748
rect 97176 70746 97200 70748
rect 97256 70746 97280 70748
rect 97336 70746 97342 70748
rect 97096 70694 97098 70746
rect 97278 70694 97280 70746
rect 97034 70692 97040 70694
rect 97096 70692 97120 70694
rect 97176 70692 97200 70694
rect 97256 70692 97280 70694
rect 97336 70692 97342 70694
rect 97034 70683 97342 70692
rect 97448 70644 97500 70650
rect 97448 70586 97500 70592
rect 97264 70508 97316 70514
rect 97264 70450 97316 70456
rect 96374 70204 96682 70213
rect 96374 70202 96380 70204
rect 96436 70202 96460 70204
rect 96516 70202 96540 70204
rect 96596 70202 96620 70204
rect 96676 70202 96682 70204
rect 96436 70150 96438 70202
rect 96618 70150 96620 70202
rect 96374 70148 96380 70150
rect 96436 70148 96460 70150
rect 96516 70148 96540 70150
rect 96596 70148 96620 70150
rect 96676 70148 96682 70150
rect 96374 70139 96682 70148
rect 97276 70009 97304 70450
rect 97460 70145 97488 70586
rect 97446 70136 97502 70145
rect 97446 70071 97502 70080
rect 97262 70000 97318 70009
rect 97262 69935 97318 69944
rect 97034 69660 97342 69669
rect 97034 69658 97040 69660
rect 97096 69658 97120 69660
rect 97176 69658 97200 69660
rect 97256 69658 97280 69660
rect 97336 69658 97342 69660
rect 97096 69606 97098 69658
rect 97278 69606 97280 69658
rect 97034 69604 97040 69606
rect 97096 69604 97120 69606
rect 97176 69604 97200 69606
rect 97256 69604 97280 69606
rect 97336 69604 97342 69606
rect 97034 69595 97342 69604
rect 96374 69116 96682 69125
rect 96374 69114 96380 69116
rect 96436 69114 96460 69116
rect 96516 69114 96540 69116
rect 96596 69114 96620 69116
rect 96676 69114 96682 69116
rect 96436 69062 96438 69114
rect 96618 69062 96620 69114
rect 96374 69060 96380 69062
rect 96436 69060 96460 69062
rect 96516 69060 96540 69062
rect 96596 69060 96620 69062
rect 96676 69060 96682 69062
rect 96374 69051 96682 69060
rect 97262 68912 97318 68921
rect 97262 68847 97318 68856
rect 97276 68814 97304 68847
rect 97264 68808 97316 68814
rect 97264 68750 97316 68756
rect 97446 68776 97502 68785
rect 97446 68711 97502 68720
rect 97460 68678 97488 68711
rect 97448 68672 97500 68678
rect 97448 68614 97500 68620
rect 97034 68572 97342 68581
rect 97034 68570 97040 68572
rect 97096 68570 97120 68572
rect 97176 68570 97200 68572
rect 97256 68570 97280 68572
rect 97336 68570 97342 68572
rect 97096 68518 97098 68570
rect 97278 68518 97280 68570
rect 97034 68516 97040 68518
rect 97096 68516 97120 68518
rect 97176 68516 97200 68518
rect 97256 68516 97280 68518
rect 97336 68516 97342 68518
rect 97034 68507 97342 68516
rect 97264 68332 97316 68338
rect 97264 68274 97316 68280
rect 96374 68028 96682 68037
rect 96374 68026 96380 68028
rect 96436 68026 96460 68028
rect 96516 68026 96540 68028
rect 96596 68026 96620 68028
rect 96676 68026 96682 68028
rect 96436 67974 96438 68026
rect 96618 67974 96620 68026
rect 96374 67972 96380 67974
rect 96436 67972 96460 67974
rect 96516 67972 96540 67974
rect 96596 67972 96620 67974
rect 96676 67972 96682 67974
rect 96374 67963 96682 67972
rect 97276 67833 97304 68274
rect 97448 68128 97500 68134
rect 97446 68096 97448 68105
rect 97500 68096 97502 68105
rect 97446 68031 97502 68040
rect 97262 67824 97318 67833
rect 97262 67759 97318 67768
rect 97034 67484 97342 67493
rect 97034 67482 97040 67484
rect 97096 67482 97120 67484
rect 97176 67482 97200 67484
rect 97256 67482 97280 67484
rect 97336 67482 97342 67484
rect 97096 67430 97098 67482
rect 97278 67430 97280 67482
rect 97034 67428 97040 67430
rect 97096 67428 97120 67430
rect 97176 67428 97200 67430
rect 97256 67428 97280 67430
rect 97336 67428 97342 67430
rect 97034 67419 97342 67428
rect 97264 67244 97316 67250
rect 97264 67186 97316 67192
rect 96374 66940 96682 66949
rect 96374 66938 96380 66940
rect 96436 66938 96460 66940
rect 96516 66938 96540 66940
rect 96596 66938 96620 66940
rect 96676 66938 96682 66940
rect 96436 66886 96438 66938
rect 96618 66886 96620 66938
rect 96374 66884 96380 66886
rect 96436 66884 96460 66886
rect 96516 66884 96540 66886
rect 96596 66884 96620 66886
rect 96676 66884 96682 66886
rect 96374 66875 96682 66884
rect 97276 66745 97304 67186
rect 97448 67040 97500 67046
rect 97448 66982 97500 66988
rect 97460 66745 97488 66982
rect 97262 66736 97318 66745
rect 97262 66671 97318 66680
rect 97446 66736 97502 66745
rect 97446 66671 97502 66680
rect 97034 66396 97342 66405
rect 97034 66394 97040 66396
rect 97096 66394 97120 66396
rect 97176 66394 97200 66396
rect 97256 66394 97280 66396
rect 97336 66394 97342 66396
rect 97096 66342 97098 66394
rect 97278 66342 97280 66394
rect 97034 66340 97040 66342
rect 97096 66340 97120 66342
rect 97176 66340 97200 66342
rect 97256 66340 97280 66342
rect 97336 66340 97342 66342
rect 97034 66331 97342 66340
rect 96374 65852 96682 65861
rect 96374 65850 96380 65852
rect 96436 65850 96460 65852
rect 96516 65850 96540 65852
rect 96596 65850 96620 65852
rect 96676 65850 96682 65852
rect 96436 65798 96438 65850
rect 96618 65798 96620 65850
rect 96374 65796 96380 65798
rect 96436 65796 96460 65798
rect 96516 65796 96540 65798
rect 96596 65796 96620 65798
rect 96676 65796 96682 65798
rect 96374 65787 96682 65796
rect 97262 65648 97318 65657
rect 97262 65583 97318 65592
rect 97276 65550 97304 65583
rect 97264 65544 97316 65550
rect 97264 65486 97316 65492
rect 97448 65408 97500 65414
rect 97446 65376 97448 65385
rect 97500 65376 97502 65385
rect 97034 65308 97342 65317
rect 97446 65311 97502 65320
rect 97034 65306 97040 65308
rect 97096 65306 97120 65308
rect 97176 65306 97200 65308
rect 97256 65306 97280 65308
rect 97336 65306 97342 65308
rect 97096 65254 97098 65306
rect 97278 65254 97280 65306
rect 97034 65252 97040 65254
rect 97096 65252 97120 65254
rect 97176 65252 97200 65254
rect 97256 65252 97280 65254
rect 97336 65252 97342 65254
rect 97034 65243 97342 65252
rect 97264 65068 97316 65074
rect 97264 65010 97316 65016
rect 96374 64764 96682 64773
rect 96374 64762 96380 64764
rect 96436 64762 96460 64764
rect 96516 64762 96540 64764
rect 96596 64762 96620 64764
rect 96676 64762 96682 64764
rect 96436 64710 96438 64762
rect 96618 64710 96620 64762
rect 96374 64708 96380 64710
rect 96436 64708 96460 64710
rect 96516 64708 96540 64710
rect 96596 64708 96620 64710
rect 96676 64708 96682 64710
rect 96374 64699 96682 64708
rect 97276 64569 97304 65010
rect 97448 64932 97500 64938
rect 97448 64874 97500 64880
rect 97460 64705 97488 64874
rect 97446 64696 97502 64705
rect 97446 64631 97502 64640
rect 97262 64560 97318 64569
rect 97262 64495 97318 64504
rect 97034 64220 97342 64229
rect 97034 64218 97040 64220
rect 97096 64218 97120 64220
rect 97176 64218 97200 64220
rect 97256 64218 97280 64220
rect 97336 64218 97342 64220
rect 97096 64166 97098 64218
rect 97278 64166 97280 64218
rect 97034 64164 97040 64166
rect 97096 64164 97120 64166
rect 97176 64164 97200 64166
rect 97256 64164 97280 64166
rect 97336 64164 97342 64166
rect 97034 64155 97342 64164
rect 96374 63676 96682 63685
rect 96374 63674 96380 63676
rect 96436 63674 96460 63676
rect 96516 63674 96540 63676
rect 96596 63674 96620 63676
rect 96676 63674 96682 63676
rect 96436 63622 96438 63674
rect 96618 63622 96620 63674
rect 96374 63620 96380 63622
rect 96436 63620 96460 63622
rect 96516 63620 96540 63622
rect 96596 63620 96620 63622
rect 96676 63620 96682 63622
rect 96374 63611 96682 63620
rect 97262 63472 97318 63481
rect 97262 63407 97318 63416
rect 97276 63374 97304 63407
rect 97264 63368 97316 63374
rect 97264 63310 97316 63316
rect 97446 63336 97502 63345
rect 97446 63271 97502 63280
rect 97460 63238 97488 63271
rect 97448 63232 97500 63238
rect 97448 63174 97500 63180
rect 97034 63132 97342 63141
rect 97034 63130 97040 63132
rect 97096 63130 97120 63132
rect 97176 63130 97200 63132
rect 97256 63130 97280 63132
rect 97336 63130 97342 63132
rect 97096 63078 97098 63130
rect 97278 63078 97280 63130
rect 97034 63076 97040 63078
rect 97096 63076 97120 63078
rect 97176 63076 97200 63078
rect 97256 63076 97280 63078
rect 97336 63076 97342 63078
rect 97034 63067 97342 63076
rect 97264 62892 97316 62898
rect 97264 62834 97316 62840
rect 96374 62588 96682 62597
rect 96374 62586 96380 62588
rect 96436 62586 96460 62588
rect 96516 62586 96540 62588
rect 96596 62586 96620 62588
rect 96676 62586 96682 62588
rect 96436 62534 96438 62586
rect 96618 62534 96620 62586
rect 96374 62532 96380 62534
rect 96436 62532 96460 62534
rect 96516 62532 96540 62534
rect 96596 62532 96620 62534
rect 96676 62532 96682 62534
rect 96374 62523 96682 62532
rect 97276 62393 97304 62834
rect 97448 62688 97500 62694
rect 97446 62656 97448 62665
rect 97500 62656 97502 62665
rect 97446 62591 97502 62600
rect 97262 62384 97318 62393
rect 97262 62319 97318 62328
rect 97034 62044 97342 62053
rect 97034 62042 97040 62044
rect 97096 62042 97120 62044
rect 97176 62042 97200 62044
rect 97256 62042 97280 62044
rect 97336 62042 97342 62044
rect 97096 61990 97098 62042
rect 97278 61990 97280 62042
rect 97034 61988 97040 61990
rect 97096 61988 97120 61990
rect 97176 61988 97200 61990
rect 97256 61988 97280 61990
rect 97336 61988 97342 61990
rect 97034 61979 97342 61988
rect 97264 61804 97316 61810
rect 97264 61746 97316 61752
rect 96374 61500 96682 61509
rect 96374 61498 96380 61500
rect 96436 61498 96460 61500
rect 96516 61498 96540 61500
rect 96596 61498 96620 61500
rect 96676 61498 96682 61500
rect 96436 61446 96438 61498
rect 96618 61446 96620 61498
rect 96374 61444 96380 61446
rect 96436 61444 96460 61446
rect 96516 61444 96540 61446
rect 96596 61444 96620 61446
rect 96676 61444 96682 61446
rect 96374 61435 96682 61444
rect 97276 61305 97304 61746
rect 97448 61600 97500 61606
rect 97448 61542 97500 61548
rect 97460 61305 97488 61542
rect 97262 61296 97318 61305
rect 97262 61231 97318 61240
rect 97446 61296 97502 61305
rect 97446 61231 97502 61240
rect 97034 60956 97342 60965
rect 97034 60954 97040 60956
rect 97096 60954 97120 60956
rect 97176 60954 97200 60956
rect 97256 60954 97280 60956
rect 97336 60954 97342 60956
rect 97096 60902 97098 60954
rect 97278 60902 97280 60954
rect 97034 60900 97040 60902
rect 97096 60900 97120 60902
rect 97176 60900 97200 60902
rect 97256 60900 97280 60902
rect 97336 60900 97342 60902
rect 97034 60891 97342 60900
rect 96374 60412 96682 60421
rect 96374 60410 96380 60412
rect 96436 60410 96460 60412
rect 96516 60410 96540 60412
rect 96596 60410 96620 60412
rect 96676 60410 96682 60412
rect 96436 60358 96438 60410
rect 96618 60358 96620 60410
rect 96374 60356 96380 60358
rect 96436 60356 96460 60358
rect 96516 60356 96540 60358
rect 96596 60356 96620 60358
rect 96676 60356 96682 60358
rect 96374 60347 96682 60356
rect 97262 60208 97318 60217
rect 97262 60143 97318 60152
rect 97276 60110 97304 60143
rect 97264 60104 97316 60110
rect 97264 60046 97316 60052
rect 97448 59968 97500 59974
rect 97446 59936 97448 59945
rect 97500 59936 97502 59945
rect 97034 59868 97342 59877
rect 97446 59871 97502 59880
rect 97034 59866 97040 59868
rect 97096 59866 97120 59868
rect 97176 59866 97200 59868
rect 97256 59866 97280 59868
rect 97336 59866 97342 59868
rect 97096 59814 97098 59866
rect 97278 59814 97280 59866
rect 97034 59812 97040 59814
rect 97096 59812 97120 59814
rect 97176 59812 97200 59814
rect 97256 59812 97280 59814
rect 97336 59812 97342 59814
rect 97034 59803 97342 59812
rect 97264 59628 97316 59634
rect 97264 59570 97316 59576
rect 96374 59324 96682 59333
rect 96374 59322 96380 59324
rect 96436 59322 96460 59324
rect 96516 59322 96540 59324
rect 96596 59322 96620 59324
rect 96676 59322 96682 59324
rect 96436 59270 96438 59322
rect 96618 59270 96620 59322
rect 96374 59268 96380 59270
rect 96436 59268 96460 59270
rect 96516 59268 96540 59270
rect 96596 59268 96620 59270
rect 96676 59268 96682 59270
rect 96374 59259 96682 59268
rect 97276 59129 97304 59570
rect 97448 59424 97500 59430
rect 97448 59366 97500 59372
rect 97460 59265 97488 59366
rect 97446 59256 97502 59265
rect 97446 59191 97502 59200
rect 97262 59120 97318 59129
rect 97262 59055 97318 59064
rect 97034 58780 97342 58789
rect 97034 58778 97040 58780
rect 97096 58778 97120 58780
rect 97176 58778 97200 58780
rect 97256 58778 97280 58780
rect 97336 58778 97342 58780
rect 97096 58726 97098 58778
rect 97278 58726 97280 58778
rect 97034 58724 97040 58726
rect 97096 58724 97120 58726
rect 97176 58724 97200 58726
rect 97256 58724 97280 58726
rect 97336 58724 97342 58726
rect 97034 58715 97342 58724
rect 96374 58236 96682 58245
rect 96374 58234 96380 58236
rect 96436 58234 96460 58236
rect 96516 58234 96540 58236
rect 96596 58234 96620 58236
rect 96676 58234 96682 58236
rect 96436 58182 96438 58234
rect 96618 58182 96620 58234
rect 96374 58180 96380 58182
rect 96436 58180 96460 58182
rect 96516 58180 96540 58182
rect 96596 58180 96620 58182
rect 96676 58180 96682 58182
rect 96374 58171 96682 58180
rect 97262 58032 97318 58041
rect 97262 57967 97318 57976
rect 97276 57934 97304 57967
rect 97264 57928 97316 57934
rect 97264 57870 97316 57876
rect 97446 57896 97502 57905
rect 97446 57831 97502 57840
rect 97460 57798 97488 57831
rect 97448 57792 97500 57798
rect 97448 57734 97500 57740
rect 97034 57692 97342 57701
rect 97034 57690 97040 57692
rect 97096 57690 97120 57692
rect 97176 57690 97200 57692
rect 97256 57690 97280 57692
rect 97336 57690 97342 57692
rect 97096 57638 97098 57690
rect 97278 57638 97280 57690
rect 97034 57636 97040 57638
rect 97096 57636 97120 57638
rect 97176 57636 97200 57638
rect 97256 57636 97280 57638
rect 97336 57636 97342 57638
rect 97034 57627 97342 57636
rect 97264 57452 97316 57458
rect 97264 57394 97316 57400
rect 96374 57148 96682 57157
rect 96374 57146 96380 57148
rect 96436 57146 96460 57148
rect 96516 57146 96540 57148
rect 96596 57146 96620 57148
rect 96676 57146 96682 57148
rect 96436 57094 96438 57146
rect 96618 57094 96620 57146
rect 96374 57092 96380 57094
rect 96436 57092 96460 57094
rect 96516 57092 96540 57094
rect 96596 57092 96620 57094
rect 96676 57092 96682 57094
rect 96374 57083 96682 57092
rect 97276 56953 97304 57394
rect 97448 57248 97500 57254
rect 97446 57216 97448 57225
rect 97500 57216 97502 57225
rect 97446 57151 97502 57160
rect 97262 56944 97318 56953
rect 97262 56879 97318 56888
rect 97034 56604 97342 56613
rect 97034 56602 97040 56604
rect 97096 56602 97120 56604
rect 97176 56602 97200 56604
rect 97256 56602 97280 56604
rect 97336 56602 97342 56604
rect 97096 56550 97098 56602
rect 97278 56550 97280 56602
rect 97034 56548 97040 56550
rect 97096 56548 97120 56550
rect 97176 56548 97200 56550
rect 97256 56548 97280 56550
rect 97336 56548 97342 56550
rect 97034 56539 97342 56548
rect 97264 56364 97316 56370
rect 97264 56306 97316 56312
rect 96374 56060 96682 56069
rect 96374 56058 96380 56060
rect 96436 56058 96460 56060
rect 96516 56058 96540 56060
rect 96596 56058 96620 56060
rect 96676 56058 96682 56060
rect 96436 56006 96438 56058
rect 96618 56006 96620 56058
rect 96374 56004 96380 56006
rect 96436 56004 96460 56006
rect 96516 56004 96540 56006
rect 96596 56004 96620 56006
rect 96676 56004 96682 56006
rect 96374 55995 96682 56004
rect 97276 55865 97304 56306
rect 97448 56160 97500 56166
rect 97448 56102 97500 56108
rect 97460 55865 97488 56102
rect 97262 55856 97318 55865
rect 97262 55791 97318 55800
rect 97446 55856 97502 55865
rect 97446 55791 97502 55800
rect 97034 55516 97342 55525
rect 97034 55514 97040 55516
rect 97096 55514 97120 55516
rect 97176 55514 97200 55516
rect 97256 55514 97280 55516
rect 97336 55514 97342 55516
rect 97096 55462 97098 55514
rect 97278 55462 97280 55514
rect 97034 55460 97040 55462
rect 97096 55460 97120 55462
rect 97176 55460 97200 55462
rect 97256 55460 97280 55462
rect 97336 55460 97342 55462
rect 97034 55451 97342 55460
rect 96374 54972 96682 54981
rect 96374 54970 96380 54972
rect 96436 54970 96460 54972
rect 96516 54970 96540 54972
rect 96596 54970 96620 54972
rect 96676 54970 96682 54972
rect 96436 54918 96438 54970
rect 96618 54918 96620 54970
rect 96374 54916 96380 54918
rect 96436 54916 96460 54918
rect 96516 54916 96540 54918
rect 96596 54916 96620 54918
rect 96676 54916 96682 54918
rect 96374 54907 96682 54916
rect 97262 54768 97318 54777
rect 97262 54703 97318 54712
rect 97276 54670 97304 54703
rect 97264 54664 97316 54670
rect 97264 54606 97316 54612
rect 97448 54528 97500 54534
rect 97446 54496 97448 54505
rect 97500 54496 97502 54505
rect 97034 54428 97342 54437
rect 97446 54431 97502 54440
rect 97034 54426 97040 54428
rect 97096 54426 97120 54428
rect 97176 54426 97200 54428
rect 97256 54426 97280 54428
rect 97336 54426 97342 54428
rect 97096 54374 97098 54426
rect 97278 54374 97280 54426
rect 97034 54372 97040 54374
rect 97096 54372 97120 54374
rect 97176 54372 97200 54374
rect 97256 54372 97280 54374
rect 97336 54372 97342 54374
rect 97034 54363 97342 54372
rect 97264 54188 97316 54194
rect 97264 54130 97316 54136
rect 96374 53884 96682 53893
rect 96374 53882 96380 53884
rect 96436 53882 96460 53884
rect 96516 53882 96540 53884
rect 96596 53882 96620 53884
rect 96676 53882 96682 53884
rect 96436 53830 96438 53882
rect 96618 53830 96620 53882
rect 96374 53828 96380 53830
rect 96436 53828 96460 53830
rect 96516 53828 96540 53830
rect 96596 53828 96620 53830
rect 96676 53828 96682 53830
rect 96374 53819 96682 53828
rect 97276 53689 97304 54130
rect 97448 53984 97500 53990
rect 97448 53926 97500 53932
rect 97460 53825 97488 53926
rect 97446 53816 97502 53825
rect 97446 53751 97502 53760
rect 97262 53680 97318 53689
rect 97262 53615 97318 53624
rect 97034 53340 97342 53349
rect 97034 53338 97040 53340
rect 97096 53338 97120 53340
rect 97176 53338 97200 53340
rect 97256 53338 97280 53340
rect 97336 53338 97342 53340
rect 97096 53286 97098 53338
rect 97278 53286 97280 53338
rect 97034 53284 97040 53286
rect 97096 53284 97120 53286
rect 97176 53284 97200 53286
rect 97256 53284 97280 53286
rect 97336 53284 97342 53286
rect 97034 53275 97342 53284
rect 96374 52796 96682 52805
rect 96374 52794 96380 52796
rect 96436 52794 96460 52796
rect 96516 52794 96540 52796
rect 96596 52794 96620 52796
rect 96676 52794 96682 52796
rect 96436 52742 96438 52794
rect 96618 52742 96620 52794
rect 96374 52740 96380 52742
rect 96436 52740 96460 52742
rect 96516 52740 96540 52742
rect 96596 52740 96620 52742
rect 96676 52740 96682 52742
rect 96374 52731 96682 52740
rect 97034 52252 97342 52261
rect 97034 52250 97040 52252
rect 97096 52250 97120 52252
rect 97176 52250 97200 52252
rect 97256 52250 97280 52252
rect 97336 52250 97342 52252
rect 97096 52198 97098 52250
rect 97278 52198 97280 52250
rect 97034 52196 97040 52198
rect 97096 52196 97120 52198
rect 97176 52196 97200 52198
rect 97256 52196 97280 52198
rect 97336 52196 97342 52198
rect 97034 52187 97342 52196
rect 96374 51708 96682 51717
rect 96374 51706 96380 51708
rect 96436 51706 96460 51708
rect 96516 51706 96540 51708
rect 96596 51706 96620 51708
rect 96676 51706 96682 51708
rect 96436 51654 96438 51706
rect 96618 51654 96620 51706
rect 96374 51652 96380 51654
rect 96436 51652 96460 51654
rect 96516 51652 96540 51654
rect 96596 51652 96620 51654
rect 96676 51652 96682 51654
rect 96374 51643 96682 51652
rect 97034 51164 97342 51173
rect 97034 51162 97040 51164
rect 97096 51162 97120 51164
rect 97176 51162 97200 51164
rect 97256 51162 97280 51164
rect 97336 51162 97342 51164
rect 97096 51110 97098 51162
rect 97278 51110 97280 51162
rect 97034 51108 97040 51110
rect 97096 51108 97120 51110
rect 97176 51108 97200 51110
rect 97256 51108 97280 51110
rect 97336 51108 97342 51110
rect 97034 51099 97342 51108
rect 92112 50856 92164 50862
rect 92112 50798 92164 50804
rect 92124 50046 92152 50798
rect 96374 50620 96682 50629
rect 96374 50618 96380 50620
rect 96436 50618 96460 50620
rect 96516 50618 96540 50620
rect 96596 50618 96620 50620
rect 96676 50618 96682 50620
rect 96436 50566 96438 50618
rect 96618 50566 96620 50618
rect 96374 50564 96380 50566
rect 96436 50564 96460 50566
rect 96516 50564 96540 50566
rect 96596 50564 96620 50566
rect 96676 50564 96682 50566
rect 96374 50555 96682 50564
rect 97034 50076 97342 50085
rect 97034 50074 97040 50076
rect 97096 50074 97120 50076
rect 97176 50074 97200 50076
rect 97256 50074 97280 50076
rect 97336 50074 97342 50076
rect 91928 50040 91980 50046
rect 91928 49982 91980 49988
rect 92112 50040 92164 50046
rect 97096 50022 97098 50074
rect 97278 50022 97280 50074
rect 97034 50020 97040 50022
rect 97096 50020 97120 50022
rect 97176 50020 97200 50022
rect 97256 50020 97280 50022
rect 97336 50020 97342 50022
rect 97034 50011 97342 50020
rect 92112 49982 92164 49988
rect 91836 48680 91888 48686
rect 91836 48622 91888 48628
rect 55404 48544 55456 48550
rect 53084 48482 53420 48498
rect 55404 48486 55456 48492
rect 91652 48544 91704 48550
rect 91652 48486 91704 48492
rect 53084 48476 53432 48482
rect 53084 48470 53380 48476
rect 53380 48418 53432 48424
rect 50848 8664 50904 8673
rect 50904 8622 51120 8650
rect 50848 8599 50904 8608
rect 51092 5914 51120 8622
rect 90620 8362 90956 8378
rect 90620 8356 90968 8362
rect 90620 8350 90916 8356
rect 90916 8298 90968 8304
rect 91940 8158 91968 49982
rect 96374 49532 96682 49541
rect 96374 49530 96380 49532
rect 96436 49530 96460 49532
rect 96516 49530 96540 49532
rect 96596 49530 96620 49532
rect 96676 49530 96682 49532
rect 96436 49478 96438 49530
rect 96618 49478 96620 49530
rect 96374 49476 96380 49478
rect 96436 49476 96460 49478
rect 96516 49476 96540 49478
rect 96596 49476 96620 49478
rect 96676 49476 96682 49478
rect 96374 49467 96682 49476
rect 97034 48988 97342 48997
rect 97034 48986 97040 48988
rect 97096 48986 97120 48988
rect 97176 48986 97200 48988
rect 97256 48986 97280 48988
rect 97336 48986 97342 48988
rect 97096 48934 97098 48986
rect 97278 48934 97280 48986
rect 97034 48932 97040 48934
rect 97096 48932 97120 48934
rect 97176 48932 97200 48934
rect 97256 48932 97280 48934
rect 97336 48932 97342 48934
rect 97034 48923 97342 48932
rect 96374 48444 96682 48453
rect 96374 48442 96380 48444
rect 96436 48442 96460 48444
rect 96516 48442 96540 48444
rect 96596 48442 96620 48444
rect 96676 48442 96682 48444
rect 96436 48390 96438 48442
rect 96618 48390 96620 48442
rect 96374 48388 96380 48390
rect 96436 48388 96460 48390
rect 96516 48388 96540 48390
rect 96596 48388 96620 48390
rect 96676 48388 96682 48390
rect 96374 48379 96682 48388
rect 97034 47900 97342 47909
rect 97034 47898 97040 47900
rect 97096 47898 97120 47900
rect 97176 47898 97200 47900
rect 97256 47898 97280 47900
rect 97336 47898 97342 47900
rect 97096 47846 97098 47898
rect 97278 47846 97280 47898
rect 97034 47844 97040 47846
rect 97096 47844 97120 47846
rect 97176 47844 97200 47846
rect 97256 47844 97280 47846
rect 97336 47844 97342 47846
rect 97034 47835 97342 47844
rect 96374 47356 96682 47365
rect 96374 47354 96380 47356
rect 96436 47354 96460 47356
rect 96516 47354 96540 47356
rect 96596 47354 96620 47356
rect 96676 47354 96682 47356
rect 96436 47302 96438 47354
rect 96618 47302 96620 47354
rect 96374 47300 96380 47302
rect 96436 47300 96460 47302
rect 96516 47300 96540 47302
rect 96596 47300 96620 47302
rect 96676 47300 96682 47302
rect 96374 47291 96682 47300
rect 97034 46812 97342 46821
rect 97034 46810 97040 46812
rect 97096 46810 97120 46812
rect 97176 46810 97200 46812
rect 97256 46810 97280 46812
rect 97336 46810 97342 46812
rect 97096 46758 97098 46810
rect 97278 46758 97280 46810
rect 97034 46756 97040 46758
rect 97096 46756 97120 46758
rect 97176 46756 97200 46758
rect 97256 46756 97280 46758
rect 97336 46756 97342 46758
rect 97034 46747 97342 46756
rect 96374 46268 96682 46277
rect 96374 46266 96380 46268
rect 96436 46266 96460 46268
rect 96516 46266 96540 46268
rect 96596 46266 96620 46268
rect 96676 46266 96682 46268
rect 96436 46214 96438 46266
rect 96618 46214 96620 46266
rect 96374 46212 96380 46214
rect 96436 46212 96460 46214
rect 96516 46212 96540 46214
rect 96596 46212 96620 46214
rect 96676 46212 96682 46214
rect 96374 46203 96682 46212
rect 97540 45960 97592 45966
rect 97540 45902 97592 45908
rect 97448 45824 97500 45830
rect 97448 45766 97500 45772
rect 97034 45724 97342 45733
rect 97034 45722 97040 45724
rect 97096 45722 97120 45724
rect 97176 45722 97200 45724
rect 97256 45722 97280 45724
rect 97336 45722 97342 45724
rect 97096 45670 97098 45722
rect 97278 45670 97280 45722
rect 97034 45668 97040 45670
rect 97096 45668 97120 45670
rect 97176 45668 97200 45670
rect 97256 45668 97280 45670
rect 97336 45668 97342 45670
rect 97034 45659 97342 45668
rect 97460 45393 97488 45766
rect 97552 45665 97580 45902
rect 97538 45656 97594 45665
rect 97538 45591 97594 45600
rect 97446 45384 97502 45393
rect 97446 45319 97502 45328
rect 96374 45180 96682 45189
rect 96374 45178 96380 45180
rect 96436 45178 96460 45180
rect 96516 45178 96540 45180
rect 96596 45178 96620 45180
rect 96676 45178 96682 45180
rect 96436 45126 96438 45178
rect 96618 45126 96620 45178
rect 96374 45124 96380 45126
rect 96436 45124 96460 45126
rect 96516 45124 96540 45126
rect 96596 45124 96620 45126
rect 96676 45124 96682 45126
rect 96374 45115 96682 45124
rect 97034 44636 97342 44645
rect 97034 44634 97040 44636
rect 97096 44634 97120 44636
rect 97176 44634 97200 44636
rect 97256 44634 97280 44636
rect 97336 44634 97342 44636
rect 97096 44582 97098 44634
rect 97278 44582 97280 44634
rect 97034 44580 97040 44582
rect 97096 44580 97120 44582
rect 97176 44580 97200 44582
rect 97256 44580 97280 44582
rect 97336 44580 97342 44582
rect 97034 44571 97342 44580
rect 97540 44396 97592 44402
rect 97540 44338 97592 44344
rect 97552 44305 97580 44338
rect 97354 44296 97410 44305
rect 97354 44231 97356 44240
rect 97408 44231 97410 44240
rect 97538 44296 97594 44305
rect 97538 44231 97594 44240
rect 97356 44202 97408 44208
rect 96374 44092 96682 44101
rect 96374 44090 96380 44092
rect 96436 44090 96460 44092
rect 96516 44090 96540 44092
rect 96596 44090 96620 44092
rect 96676 44090 96682 44092
rect 96436 44038 96438 44090
rect 96618 44038 96620 44090
rect 96374 44036 96380 44038
rect 96436 44036 96460 44038
rect 96516 44036 96540 44038
rect 96596 44036 96620 44038
rect 96676 44036 96682 44038
rect 96374 44027 96682 44036
rect 97034 43548 97342 43557
rect 97034 43546 97040 43548
rect 97096 43546 97120 43548
rect 97176 43546 97200 43548
rect 97256 43546 97280 43548
rect 97336 43546 97342 43548
rect 97096 43494 97098 43546
rect 97278 43494 97280 43546
rect 97034 43492 97040 43494
rect 97096 43492 97120 43494
rect 97176 43492 97200 43494
rect 97256 43492 97280 43494
rect 97336 43492 97342 43494
rect 97034 43483 97342 43492
rect 97540 43308 97592 43314
rect 97540 43250 97592 43256
rect 97354 43208 97410 43217
rect 97354 43143 97356 43152
rect 97408 43143 97410 43152
rect 97356 43114 97408 43120
rect 96374 43004 96682 43013
rect 96374 43002 96380 43004
rect 96436 43002 96460 43004
rect 96516 43002 96540 43004
rect 96596 43002 96620 43004
rect 96676 43002 96682 43004
rect 96436 42950 96438 43002
rect 96618 42950 96620 43002
rect 96374 42948 96380 42950
rect 96436 42948 96460 42950
rect 96516 42948 96540 42950
rect 96596 42948 96620 42950
rect 96676 42948 96682 42950
rect 96374 42939 96682 42948
rect 97552 42945 97580 43250
rect 97538 42936 97594 42945
rect 97538 42871 97594 42880
rect 97540 42696 97592 42702
rect 97540 42638 97592 42644
rect 97448 42560 97500 42566
rect 97448 42502 97500 42508
rect 97034 42460 97342 42469
rect 97034 42458 97040 42460
rect 97096 42458 97120 42460
rect 97176 42458 97200 42460
rect 97256 42458 97280 42460
rect 97336 42458 97342 42460
rect 97096 42406 97098 42458
rect 97278 42406 97280 42458
rect 97034 42404 97040 42406
rect 97096 42404 97120 42406
rect 97176 42404 97200 42406
rect 97256 42404 97280 42406
rect 97336 42404 97342 42406
rect 97034 42395 97342 42404
rect 97460 42129 97488 42502
rect 97552 42265 97580 42638
rect 97538 42256 97594 42265
rect 97538 42191 97594 42200
rect 97446 42120 97502 42129
rect 97446 42055 97502 42064
rect 96374 41916 96682 41925
rect 96374 41914 96380 41916
rect 96436 41914 96460 41916
rect 96516 41914 96540 41916
rect 96596 41914 96620 41916
rect 96676 41914 96682 41916
rect 96436 41862 96438 41914
rect 96618 41862 96620 41914
rect 96374 41860 96380 41862
rect 96436 41860 96460 41862
rect 96516 41860 96540 41862
rect 96596 41860 96620 41862
rect 96676 41860 96682 41862
rect 96374 41851 96682 41860
rect 97034 41372 97342 41381
rect 97034 41370 97040 41372
rect 97096 41370 97120 41372
rect 97176 41370 97200 41372
rect 97256 41370 97280 41372
rect 97336 41370 97342 41372
rect 97096 41318 97098 41370
rect 97278 41318 97280 41370
rect 97034 41316 97040 41318
rect 97096 41316 97120 41318
rect 97176 41316 97200 41318
rect 97256 41316 97280 41318
rect 97336 41316 97342 41318
rect 97034 41307 97342 41316
rect 97356 41268 97408 41274
rect 97356 41210 97408 41216
rect 97368 41177 97396 41210
rect 97354 41168 97410 41177
rect 97354 41103 97410 41112
rect 97540 41132 97592 41138
rect 97540 41074 97592 41080
rect 97552 40905 97580 41074
rect 97538 40896 97594 40905
rect 96374 40828 96682 40837
rect 97538 40831 97594 40840
rect 96374 40826 96380 40828
rect 96436 40826 96460 40828
rect 96516 40826 96540 40828
rect 96596 40826 96620 40828
rect 96676 40826 96682 40828
rect 96436 40774 96438 40826
rect 96618 40774 96620 40826
rect 96374 40772 96380 40774
rect 96436 40772 96460 40774
rect 96516 40772 96540 40774
rect 96596 40772 96620 40774
rect 96676 40772 96682 40774
rect 96374 40763 96682 40772
rect 97540 40520 97592 40526
rect 97540 40462 97592 40468
rect 97448 40384 97500 40390
rect 97448 40326 97500 40332
rect 97034 40284 97342 40293
rect 97034 40282 97040 40284
rect 97096 40282 97120 40284
rect 97176 40282 97200 40284
rect 97256 40282 97280 40284
rect 97336 40282 97342 40284
rect 97096 40230 97098 40282
rect 97278 40230 97280 40282
rect 97034 40228 97040 40230
rect 97096 40228 97120 40230
rect 97176 40228 97200 40230
rect 97256 40228 97280 40230
rect 97336 40228 97342 40230
rect 97034 40219 97342 40228
rect 97460 39953 97488 40326
rect 97552 40225 97580 40462
rect 97538 40216 97594 40225
rect 97538 40151 97594 40160
rect 97446 39944 97502 39953
rect 97446 39879 97502 39888
rect 96374 39740 96682 39749
rect 96374 39738 96380 39740
rect 96436 39738 96460 39740
rect 96516 39738 96540 39740
rect 96596 39738 96620 39740
rect 96676 39738 96682 39740
rect 96436 39686 96438 39738
rect 96618 39686 96620 39738
rect 96374 39684 96380 39686
rect 96436 39684 96460 39686
rect 96516 39684 96540 39686
rect 96596 39684 96620 39686
rect 96676 39684 96682 39686
rect 96374 39675 96682 39684
rect 97034 39196 97342 39205
rect 97034 39194 97040 39196
rect 97096 39194 97120 39196
rect 97176 39194 97200 39196
rect 97256 39194 97280 39196
rect 97336 39194 97342 39196
rect 97096 39142 97098 39194
rect 97278 39142 97280 39194
rect 97034 39140 97040 39142
rect 97096 39140 97120 39142
rect 97176 39140 97200 39142
rect 97256 39140 97280 39142
rect 97336 39140 97342 39142
rect 97034 39131 97342 39140
rect 97356 39092 97408 39098
rect 97356 39034 97408 39040
rect 97368 39001 97396 39034
rect 97354 38992 97410 39001
rect 97354 38927 97410 38936
rect 97540 38956 97592 38962
rect 97540 38898 97592 38904
rect 97552 38865 97580 38898
rect 97538 38856 97594 38865
rect 97538 38791 97594 38800
rect 96374 38652 96682 38661
rect 96374 38650 96380 38652
rect 96436 38650 96460 38652
rect 96516 38650 96540 38652
rect 96596 38650 96620 38652
rect 96676 38650 96682 38652
rect 96436 38598 96438 38650
rect 96618 38598 96620 38650
rect 96374 38596 96380 38598
rect 96436 38596 96460 38598
rect 96516 38596 96540 38598
rect 96596 38596 96620 38598
rect 96676 38596 96682 38598
rect 96374 38587 96682 38596
rect 97034 38108 97342 38117
rect 97034 38106 97040 38108
rect 97096 38106 97120 38108
rect 97176 38106 97200 38108
rect 97256 38106 97280 38108
rect 97336 38106 97342 38108
rect 97096 38054 97098 38106
rect 97278 38054 97280 38106
rect 97034 38052 97040 38054
rect 97096 38052 97120 38054
rect 97176 38052 97200 38054
rect 97256 38052 97280 38054
rect 97336 38052 97342 38054
rect 97034 38043 97342 38052
rect 97356 38004 97408 38010
rect 97356 37946 97408 37952
rect 97368 37913 97396 37946
rect 97354 37904 97410 37913
rect 97354 37839 97410 37848
rect 97540 37868 97592 37874
rect 97540 37810 97592 37816
rect 96374 37564 96682 37573
rect 96374 37562 96380 37564
rect 96436 37562 96460 37564
rect 96516 37562 96540 37564
rect 96596 37562 96620 37564
rect 96676 37562 96682 37564
rect 96436 37510 96438 37562
rect 96618 37510 96620 37562
rect 96374 37508 96380 37510
rect 96436 37508 96460 37510
rect 96516 37508 96540 37510
rect 96596 37508 96620 37510
rect 96676 37508 96682 37510
rect 96374 37499 96682 37508
rect 97552 37505 97580 37810
rect 97538 37496 97594 37505
rect 97538 37431 97594 37440
rect 96620 37324 96672 37330
rect 96620 37266 96672 37272
rect 96632 36825 96660 37266
rect 97448 37188 97500 37194
rect 97448 37130 97500 37136
rect 97034 37020 97342 37029
rect 97034 37018 97040 37020
rect 97096 37018 97120 37020
rect 97176 37018 97200 37020
rect 97256 37018 97280 37020
rect 97336 37018 97342 37020
rect 97096 36966 97098 37018
rect 97278 36966 97280 37018
rect 97034 36964 97040 36966
rect 97096 36964 97120 36966
rect 97176 36964 97200 36966
rect 97256 36964 97280 36966
rect 97336 36964 97342 36966
rect 97034 36955 97342 36964
rect 97460 36825 97488 37130
rect 96618 36816 96674 36825
rect 96618 36751 96674 36760
rect 97446 36816 97502 36825
rect 97446 36751 97502 36760
rect 96374 36476 96682 36485
rect 96374 36474 96380 36476
rect 96436 36474 96460 36476
rect 96516 36474 96540 36476
rect 96596 36474 96620 36476
rect 96676 36474 96682 36476
rect 96436 36422 96438 36474
rect 96618 36422 96620 36474
rect 96374 36420 96380 36422
rect 96436 36420 96460 36422
rect 96516 36420 96540 36422
rect 96596 36420 96620 36422
rect 96676 36420 96682 36422
rect 96374 36411 96682 36420
rect 97034 35932 97342 35941
rect 97034 35930 97040 35932
rect 97096 35930 97120 35932
rect 97176 35930 97200 35932
rect 97256 35930 97280 35932
rect 97336 35930 97342 35932
rect 97096 35878 97098 35930
rect 97278 35878 97280 35930
rect 97034 35876 97040 35878
rect 97096 35876 97120 35878
rect 97176 35876 97200 35878
rect 97256 35876 97280 35878
rect 97336 35876 97342 35878
rect 97034 35867 97342 35876
rect 97356 35828 97408 35834
rect 97356 35770 97408 35776
rect 97368 35737 97396 35770
rect 97354 35728 97410 35737
rect 97354 35663 97410 35672
rect 97540 35692 97592 35698
rect 97540 35634 97592 35640
rect 97552 35465 97580 35634
rect 97538 35456 97594 35465
rect 96374 35388 96682 35397
rect 97538 35391 97594 35400
rect 96374 35386 96380 35388
rect 96436 35386 96460 35388
rect 96516 35386 96540 35388
rect 96596 35386 96620 35388
rect 96676 35386 96682 35388
rect 96436 35334 96438 35386
rect 96618 35334 96620 35386
rect 96374 35332 96380 35334
rect 96436 35332 96460 35334
rect 96516 35332 96540 35334
rect 96596 35332 96620 35334
rect 96676 35332 96682 35334
rect 96374 35323 96682 35332
rect 97540 35080 97592 35086
rect 97540 35022 97592 35028
rect 97448 34944 97500 34950
rect 97448 34886 97500 34892
rect 97034 34844 97342 34853
rect 97034 34842 97040 34844
rect 97096 34842 97120 34844
rect 97176 34842 97200 34844
rect 97256 34842 97280 34844
rect 97336 34842 97342 34844
rect 97096 34790 97098 34842
rect 97278 34790 97280 34842
rect 97034 34788 97040 34790
rect 97096 34788 97120 34790
rect 97176 34788 97200 34790
rect 97256 34788 97280 34790
rect 97336 34788 97342 34790
rect 97034 34779 97342 34788
rect 97460 34513 97488 34886
rect 97552 34785 97580 35022
rect 97538 34776 97594 34785
rect 97538 34711 97594 34720
rect 97446 34504 97502 34513
rect 97446 34439 97502 34448
rect 96374 34300 96682 34309
rect 96374 34298 96380 34300
rect 96436 34298 96460 34300
rect 96516 34298 96540 34300
rect 96596 34298 96620 34300
rect 96676 34298 96682 34300
rect 96436 34246 96438 34298
rect 96618 34246 96620 34298
rect 96374 34244 96380 34246
rect 96436 34244 96460 34246
rect 96516 34244 96540 34246
rect 96596 34244 96620 34246
rect 96676 34244 96682 34246
rect 96374 34235 96682 34244
rect 97034 33756 97342 33765
rect 97034 33754 97040 33756
rect 97096 33754 97120 33756
rect 97176 33754 97200 33756
rect 97256 33754 97280 33756
rect 97336 33754 97342 33756
rect 97096 33702 97098 33754
rect 97278 33702 97280 33754
rect 97034 33700 97040 33702
rect 97096 33700 97120 33702
rect 97176 33700 97200 33702
rect 97256 33700 97280 33702
rect 97336 33700 97342 33702
rect 97034 33691 97342 33700
rect 97356 33652 97408 33658
rect 97356 33594 97408 33600
rect 97368 33561 97396 33594
rect 97354 33552 97410 33561
rect 97354 33487 97410 33496
rect 97540 33516 97592 33522
rect 97540 33458 97592 33464
rect 97552 33425 97580 33458
rect 97538 33416 97594 33425
rect 97538 33351 97594 33360
rect 96374 33212 96682 33221
rect 96374 33210 96380 33212
rect 96436 33210 96460 33212
rect 96516 33210 96540 33212
rect 96596 33210 96620 33212
rect 96676 33210 96682 33212
rect 96436 33158 96438 33210
rect 96618 33158 96620 33210
rect 96374 33156 96380 33158
rect 96436 33156 96460 33158
rect 96516 33156 96540 33158
rect 96596 33156 96620 33158
rect 96676 33156 96682 33158
rect 96374 33147 96682 33156
rect 97034 32668 97342 32677
rect 97034 32666 97040 32668
rect 97096 32666 97120 32668
rect 97176 32666 97200 32668
rect 97256 32666 97280 32668
rect 97336 32666 97342 32668
rect 97096 32614 97098 32666
rect 97278 32614 97280 32666
rect 97034 32612 97040 32614
rect 97096 32612 97120 32614
rect 97176 32612 97200 32614
rect 97256 32612 97280 32614
rect 97336 32612 97342 32614
rect 97034 32603 97342 32612
rect 97264 32496 97316 32502
rect 97262 32464 97264 32473
rect 97316 32464 97318 32473
rect 97262 32399 97318 32408
rect 97448 32428 97500 32434
rect 97448 32370 97500 32376
rect 96374 32124 96682 32133
rect 96374 32122 96380 32124
rect 96436 32122 96460 32124
rect 96516 32122 96540 32124
rect 96596 32122 96620 32124
rect 96676 32122 96682 32124
rect 96436 32070 96438 32122
rect 96618 32070 96620 32122
rect 96374 32068 96380 32070
rect 96436 32068 96460 32070
rect 96516 32068 96540 32070
rect 96596 32068 96620 32070
rect 96676 32068 96682 32070
rect 96374 32059 96682 32068
rect 97460 32065 97488 32370
rect 97446 32056 97502 32065
rect 97446 31991 97502 32000
rect 96620 31952 96672 31958
rect 96620 31894 96672 31900
rect 96632 31385 96660 31894
rect 97540 31816 97592 31822
rect 97540 31758 97592 31764
rect 97034 31580 97342 31589
rect 97034 31578 97040 31580
rect 97096 31578 97120 31580
rect 97176 31578 97200 31580
rect 97256 31578 97280 31580
rect 97336 31578 97342 31580
rect 97096 31526 97098 31578
rect 97278 31526 97280 31578
rect 97034 31524 97040 31526
rect 97096 31524 97120 31526
rect 97176 31524 97200 31526
rect 97256 31524 97280 31526
rect 97336 31524 97342 31526
rect 97034 31515 97342 31524
rect 97552 31385 97580 31758
rect 96618 31376 96674 31385
rect 96618 31311 96674 31320
rect 97538 31376 97594 31385
rect 97538 31311 97594 31320
rect 96374 31036 96682 31045
rect 96374 31034 96380 31036
rect 96436 31034 96460 31036
rect 96516 31034 96540 31036
rect 96596 31034 96620 31036
rect 96676 31034 96682 31036
rect 96436 30982 96438 31034
rect 96618 30982 96620 31034
rect 96374 30980 96380 30982
rect 96436 30980 96460 30982
rect 96516 30980 96540 30982
rect 96596 30980 96620 30982
rect 96676 30980 96682 30982
rect 96374 30971 96682 30980
rect 97540 30592 97592 30598
rect 97540 30534 97592 30540
rect 97034 30492 97342 30501
rect 97034 30490 97040 30492
rect 97096 30490 97120 30492
rect 97176 30490 97200 30492
rect 97256 30490 97280 30492
rect 97336 30490 97342 30492
rect 97096 30438 97098 30490
rect 97278 30438 97280 30490
rect 97034 30436 97040 30438
rect 97096 30436 97120 30438
rect 97176 30436 97200 30438
rect 97256 30436 97280 30438
rect 97336 30436 97342 30438
rect 97034 30427 97342 30436
rect 97262 30288 97318 30297
rect 97262 30223 97264 30232
rect 97316 30223 97318 30232
rect 97264 30194 97316 30200
rect 97552 30190 97580 30534
rect 97540 30184 97592 30190
rect 97540 30126 97592 30132
rect 97552 30025 97580 30126
rect 97538 30016 97594 30025
rect 96374 29948 96682 29957
rect 97538 29951 97594 29960
rect 96374 29946 96380 29948
rect 96436 29946 96460 29948
rect 96516 29946 96540 29948
rect 96596 29946 96620 29948
rect 96676 29946 96682 29948
rect 96436 29894 96438 29946
rect 96618 29894 96620 29946
rect 96374 29892 96380 29894
rect 96436 29892 96460 29894
rect 96516 29892 96540 29894
rect 96596 29892 96620 29894
rect 96676 29892 96682 29894
rect 96374 29883 96682 29892
rect 97540 29640 97592 29646
rect 97540 29582 97592 29588
rect 97448 29504 97500 29510
rect 97448 29446 97500 29452
rect 97034 29404 97342 29413
rect 97034 29402 97040 29404
rect 97096 29402 97120 29404
rect 97176 29402 97200 29404
rect 97256 29402 97280 29404
rect 97336 29402 97342 29404
rect 97096 29350 97098 29402
rect 97278 29350 97280 29402
rect 97034 29348 97040 29350
rect 97096 29348 97120 29350
rect 97176 29348 97200 29350
rect 97256 29348 97280 29350
rect 97336 29348 97342 29350
rect 97034 29339 97342 29348
rect 97460 29209 97488 29446
rect 97552 29345 97580 29582
rect 97538 29336 97594 29345
rect 97538 29271 97594 29280
rect 97446 29200 97502 29209
rect 97446 29135 97502 29144
rect 96374 28860 96682 28869
rect 96374 28858 96380 28860
rect 96436 28858 96460 28860
rect 96516 28858 96540 28860
rect 96596 28858 96620 28860
rect 96676 28858 96682 28860
rect 96436 28806 96438 28858
rect 96618 28806 96620 28858
rect 96374 28804 96380 28806
rect 96436 28804 96460 28806
rect 96516 28804 96540 28806
rect 96596 28804 96620 28806
rect 96676 28804 96682 28806
rect 96374 28795 96682 28804
rect 97034 28316 97342 28325
rect 97034 28314 97040 28316
rect 97096 28314 97120 28316
rect 97176 28314 97200 28316
rect 97256 28314 97280 28316
rect 97336 28314 97342 28316
rect 97096 28262 97098 28314
rect 97278 28262 97280 28314
rect 97034 28260 97040 28262
rect 97096 28260 97120 28262
rect 97176 28260 97200 28262
rect 97256 28260 97280 28262
rect 97336 28260 97342 28262
rect 97034 28251 97342 28260
rect 97262 28112 97318 28121
rect 97262 28047 97264 28056
rect 97316 28047 97318 28056
rect 97264 28018 97316 28024
rect 97446 27976 97502 27985
rect 97446 27911 97448 27920
rect 97500 27911 97502 27920
rect 97448 27882 97500 27888
rect 96374 27772 96682 27781
rect 96374 27770 96380 27772
rect 96436 27770 96460 27772
rect 96516 27770 96540 27772
rect 96596 27770 96620 27772
rect 96676 27770 96682 27772
rect 96436 27718 96438 27770
rect 96618 27718 96620 27770
rect 96374 27716 96380 27718
rect 96436 27716 96460 27718
rect 96516 27716 96540 27718
rect 96596 27716 96620 27718
rect 96676 27716 96682 27718
rect 96374 27707 96682 27716
rect 97034 27228 97342 27237
rect 97034 27226 97040 27228
rect 97096 27226 97120 27228
rect 97176 27226 97200 27228
rect 97256 27226 97280 27228
rect 97336 27226 97342 27228
rect 97096 27174 97098 27226
rect 97278 27174 97280 27226
rect 97034 27172 97040 27174
rect 97096 27172 97120 27174
rect 97176 27172 97200 27174
rect 97256 27172 97280 27174
rect 97336 27172 97342 27174
rect 97034 27163 97342 27172
rect 97262 27024 97318 27033
rect 97262 26959 97264 26968
rect 97316 26959 97318 26968
rect 97264 26930 97316 26936
rect 97448 26784 97500 26790
rect 97448 26726 97500 26732
rect 96374 26684 96682 26693
rect 96374 26682 96380 26684
rect 96436 26682 96460 26684
rect 96516 26682 96540 26684
rect 96596 26682 96620 26684
rect 96676 26682 96682 26684
rect 96436 26630 96438 26682
rect 96618 26630 96620 26682
rect 96374 26628 96380 26630
rect 96436 26628 96460 26630
rect 96516 26628 96540 26630
rect 96596 26628 96620 26630
rect 96676 26628 96682 26630
rect 96374 26619 96682 26628
rect 97460 26625 97488 26726
rect 97446 26616 97502 26625
rect 97446 26551 97502 26560
rect 97448 26512 97500 26518
rect 97448 26454 97500 26460
rect 96896 26376 96948 26382
rect 96896 26318 96948 26324
rect 96908 25945 96936 26318
rect 97034 26140 97342 26149
rect 97034 26138 97040 26140
rect 97096 26138 97120 26140
rect 97176 26138 97200 26140
rect 97256 26138 97280 26140
rect 97336 26138 97342 26140
rect 97096 26086 97098 26138
rect 97278 26086 97280 26138
rect 97034 26084 97040 26086
rect 97096 26084 97120 26086
rect 97176 26084 97200 26086
rect 97256 26084 97280 26086
rect 97336 26084 97342 26086
rect 97034 26075 97342 26084
rect 97460 25945 97488 26454
rect 96894 25936 96950 25945
rect 96894 25871 96950 25880
rect 97446 25936 97502 25945
rect 97446 25871 97502 25880
rect 96374 25596 96682 25605
rect 96374 25594 96380 25596
rect 96436 25594 96460 25596
rect 96516 25594 96540 25596
rect 96596 25594 96620 25596
rect 96676 25594 96682 25596
rect 96436 25542 96438 25594
rect 96618 25542 96620 25594
rect 96374 25540 96380 25542
rect 96436 25540 96460 25542
rect 96516 25540 96540 25542
rect 96596 25540 96620 25542
rect 96676 25540 96682 25542
rect 96374 25531 96682 25540
rect 97034 25052 97342 25061
rect 97034 25050 97040 25052
rect 97096 25050 97120 25052
rect 97176 25050 97200 25052
rect 97256 25050 97280 25052
rect 97336 25050 97342 25052
rect 97096 24998 97098 25050
rect 97278 24998 97280 25050
rect 97034 24996 97040 24998
rect 97096 24996 97120 24998
rect 97176 24996 97200 24998
rect 97256 24996 97280 24998
rect 97336 24996 97342 24998
rect 97034 24987 97342 24996
rect 97262 24848 97318 24857
rect 97262 24783 97264 24792
rect 97316 24783 97318 24792
rect 97264 24754 97316 24760
rect 97448 24608 97500 24614
rect 97446 24576 97448 24585
rect 97500 24576 97502 24585
rect 96374 24508 96682 24517
rect 97446 24511 97502 24520
rect 96374 24506 96380 24508
rect 96436 24506 96460 24508
rect 96516 24506 96540 24508
rect 96596 24506 96620 24508
rect 96676 24506 96682 24508
rect 96436 24454 96438 24506
rect 96618 24454 96620 24506
rect 96374 24452 96380 24454
rect 96436 24452 96460 24454
rect 96516 24452 96540 24454
rect 96596 24452 96620 24454
rect 96676 24452 96682 24454
rect 96374 24443 96682 24452
rect 96620 24200 96672 24206
rect 96620 24142 96672 24148
rect 96632 23769 96660 24142
rect 97448 24064 97500 24070
rect 97448 24006 97500 24012
rect 97034 23964 97342 23973
rect 97034 23962 97040 23964
rect 97096 23962 97120 23964
rect 97176 23962 97200 23964
rect 97256 23962 97280 23964
rect 97336 23962 97342 23964
rect 97096 23910 97098 23962
rect 97278 23910 97280 23962
rect 97034 23908 97040 23910
rect 97096 23908 97120 23910
rect 97176 23908 97200 23910
rect 97256 23908 97280 23910
rect 97336 23908 97342 23910
rect 97034 23899 97342 23908
rect 97460 23905 97488 24006
rect 97446 23896 97502 23905
rect 97446 23831 97502 23840
rect 96618 23760 96674 23769
rect 96618 23695 96674 23704
rect 96374 23420 96682 23429
rect 96374 23418 96380 23420
rect 96436 23418 96460 23420
rect 96516 23418 96540 23420
rect 96596 23418 96620 23420
rect 96676 23418 96682 23420
rect 96436 23366 96438 23418
rect 96618 23366 96620 23418
rect 96374 23364 96380 23366
rect 96436 23364 96460 23366
rect 96516 23364 96540 23366
rect 96596 23364 96620 23366
rect 96676 23364 96682 23366
rect 96374 23355 96682 23364
rect 97034 22876 97342 22885
rect 97034 22874 97040 22876
rect 97096 22874 97120 22876
rect 97176 22874 97200 22876
rect 97256 22874 97280 22876
rect 97336 22874 97342 22876
rect 97096 22822 97098 22874
rect 97278 22822 97280 22874
rect 97034 22820 97040 22822
rect 97096 22820 97120 22822
rect 97176 22820 97200 22822
rect 97256 22820 97280 22822
rect 97336 22820 97342 22822
rect 97034 22811 97342 22820
rect 97262 22672 97318 22681
rect 97262 22607 97264 22616
rect 97316 22607 97318 22616
rect 97264 22578 97316 22584
rect 97446 22536 97502 22545
rect 97446 22471 97448 22480
rect 97500 22471 97502 22480
rect 97448 22442 97500 22448
rect 96374 22332 96682 22341
rect 96374 22330 96380 22332
rect 96436 22330 96460 22332
rect 96516 22330 96540 22332
rect 96596 22330 96620 22332
rect 96676 22330 96682 22332
rect 96436 22278 96438 22330
rect 96618 22278 96620 22330
rect 96374 22276 96380 22278
rect 96436 22276 96460 22278
rect 96516 22276 96540 22278
rect 96596 22276 96620 22278
rect 96676 22276 96682 22278
rect 96374 22267 96682 22276
rect 97034 21788 97342 21797
rect 97034 21786 97040 21788
rect 97096 21786 97120 21788
rect 97176 21786 97200 21788
rect 97256 21786 97280 21788
rect 97336 21786 97342 21788
rect 97096 21734 97098 21786
rect 97278 21734 97280 21786
rect 97034 21732 97040 21734
rect 97096 21732 97120 21734
rect 97176 21732 97200 21734
rect 97256 21732 97280 21734
rect 97336 21732 97342 21734
rect 97034 21723 97342 21732
rect 97262 21584 97318 21593
rect 97262 21519 97264 21528
rect 97316 21519 97318 21528
rect 97264 21490 97316 21496
rect 97448 21344 97500 21350
rect 97448 21286 97500 21292
rect 96374 21244 96682 21253
rect 96374 21242 96380 21244
rect 96436 21242 96460 21244
rect 96516 21242 96540 21244
rect 96596 21242 96620 21244
rect 96676 21242 96682 21244
rect 96436 21190 96438 21242
rect 96618 21190 96620 21242
rect 96374 21188 96380 21190
rect 96436 21188 96460 21190
rect 96516 21188 96540 21190
rect 96596 21188 96620 21190
rect 96676 21188 96682 21190
rect 96374 21179 96682 21188
rect 97460 21185 97488 21286
rect 97446 21176 97502 21185
rect 97446 21111 97502 21120
rect 96620 20936 96672 20942
rect 96620 20878 96672 20884
rect 96632 20505 96660 20878
rect 97448 20800 97500 20806
rect 97448 20742 97500 20748
rect 97034 20700 97342 20709
rect 97034 20698 97040 20700
rect 97096 20698 97120 20700
rect 97176 20698 97200 20700
rect 97256 20698 97280 20700
rect 97336 20698 97342 20700
rect 97096 20646 97098 20698
rect 97278 20646 97280 20698
rect 97034 20644 97040 20646
rect 97096 20644 97120 20646
rect 97176 20644 97200 20646
rect 97256 20644 97280 20646
rect 97336 20644 97342 20646
rect 97034 20635 97342 20644
rect 97460 20505 97488 20742
rect 96618 20496 96674 20505
rect 96618 20431 96674 20440
rect 97446 20496 97502 20505
rect 97446 20431 97502 20440
rect 96374 20156 96682 20165
rect 96374 20154 96380 20156
rect 96436 20154 96460 20156
rect 96516 20154 96540 20156
rect 96596 20154 96620 20156
rect 96676 20154 96682 20156
rect 96436 20102 96438 20154
rect 96618 20102 96620 20154
rect 96374 20100 96380 20102
rect 96436 20100 96460 20102
rect 96516 20100 96540 20102
rect 96596 20100 96620 20102
rect 96676 20100 96682 20102
rect 96374 20091 96682 20100
rect 97034 19612 97342 19621
rect 97034 19610 97040 19612
rect 97096 19610 97120 19612
rect 97176 19610 97200 19612
rect 97256 19610 97280 19612
rect 97336 19610 97342 19612
rect 97096 19558 97098 19610
rect 97278 19558 97280 19610
rect 97034 19556 97040 19558
rect 97096 19556 97120 19558
rect 97176 19556 97200 19558
rect 97256 19556 97280 19558
rect 97336 19556 97342 19558
rect 97034 19547 97342 19556
rect 97448 19508 97500 19514
rect 97448 19450 97500 19456
rect 97264 19372 97316 19378
rect 97264 19314 97316 19320
rect 97276 19281 97304 19314
rect 97262 19272 97318 19281
rect 97262 19207 97318 19216
rect 97460 19145 97488 19450
rect 97446 19136 97502 19145
rect 96374 19068 96682 19077
rect 97446 19071 97502 19080
rect 96374 19066 96380 19068
rect 96436 19066 96460 19068
rect 96516 19066 96540 19068
rect 96596 19066 96620 19068
rect 96676 19066 96682 19068
rect 96436 19014 96438 19066
rect 96618 19014 96620 19066
rect 96374 19012 96380 19014
rect 96436 19012 96460 19014
rect 96516 19012 96540 19014
rect 96596 19012 96620 19014
rect 96676 19012 96682 19014
rect 96374 19003 96682 19012
rect 96620 18760 96672 18766
rect 96620 18702 96672 18708
rect 96632 18329 96660 18702
rect 97448 18624 97500 18630
rect 97448 18566 97500 18572
rect 97034 18524 97342 18533
rect 97034 18522 97040 18524
rect 97096 18522 97120 18524
rect 97176 18522 97200 18524
rect 97256 18522 97280 18524
rect 97336 18522 97342 18524
rect 97096 18470 97098 18522
rect 97278 18470 97280 18522
rect 97034 18468 97040 18470
rect 97096 18468 97120 18470
rect 97176 18468 97200 18470
rect 97256 18468 97280 18470
rect 97336 18468 97342 18470
rect 97034 18459 97342 18468
rect 97460 18465 97488 18566
rect 97446 18456 97502 18465
rect 97446 18391 97502 18400
rect 96618 18320 96674 18329
rect 96618 18255 96674 18264
rect 96374 17980 96682 17989
rect 96374 17978 96380 17980
rect 96436 17978 96460 17980
rect 96516 17978 96540 17980
rect 96596 17978 96620 17980
rect 96676 17978 96682 17980
rect 96436 17926 96438 17978
rect 96618 17926 96620 17978
rect 96374 17924 96380 17926
rect 96436 17924 96460 17926
rect 96516 17924 96540 17926
rect 96596 17924 96620 17926
rect 96676 17924 96682 17926
rect 96374 17915 96682 17924
rect 97034 17436 97342 17445
rect 97034 17434 97040 17436
rect 97096 17434 97120 17436
rect 97176 17434 97200 17436
rect 97256 17434 97280 17436
rect 97336 17434 97342 17436
rect 97096 17382 97098 17434
rect 97278 17382 97280 17434
rect 97034 17380 97040 17382
rect 97096 17380 97120 17382
rect 97176 17380 97200 17382
rect 97256 17380 97280 17382
rect 97336 17380 97342 17382
rect 97034 17371 97342 17380
rect 97262 17232 97318 17241
rect 97262 17167 97264 17176
rect 97316 17167 97318 17176
rect 97264 17138 97316 17144
rect 97446 17096 97502 17105
rect 97446 17031 97448 17040
rect 97500 17031 97502 17040
rect 97448 17002 97500 17008
rect 96374 16892 96682 16901
rect 96374 16890 96380 16892
rect 96436 16890 96460 16892
rect 96516 16890 96540 16892
rect 96596 16890 96620 16892
rect 96676 16890 96682 16892
rect 96436 16838 96438 16890
rect 96618 16838 96620 16890
rect 96374 16836 96380 16838
rect 96436 16836 96460 16838
rect 96516 16836 96540 16838
rect 96596 16836 96620 16838
rect 96676 16836 96682 16838
rect 96374 16827 96682 16836
rect 97034 16348 97342 16357
rect 97034 16346 97040 16348
rect 97096 16346 97120 16348
rect 97176 16346 97200 16348
rect 97256 16346 97280 16348
rect 97336 16346 97342 16348
rect 97096 16294 97098 16346
rect 97278 16294 97280 16346
rect 97034 16292 97040 16294
rect 97096 16292 97120 16294
rect 97176 16292 97200 16294
rect 97256 16292 97280 16294
rect 97336 16292 97342 16294
rect 97034 16283 97342 16292
rect 97262 16144 97318 16153
rect 97262 16079 97264 16088
rect 97316 16079 97318 16088
rect 97264 16050 97316 16056
rect 97448 15904 97500 15910
rect 97448 15846 97500 15852
rect 96374 15804 96682 15813
rect 96374 15802 96380 15804
rect 96436 15802 96460 15804
rect 96516 15802 96540 15804
rect 96596 15802 96620 15804
rect 96676 15802 96682 15804
rect 96436 15750 96438 15802
rect 96618 15750 96620 15802
rect 96374 15748 96380 15750
rect 96436 15748 96460 15750
rect 96516 15748 96540 15750
rect 96596 15748 96620 15750
rect 96676 15748 96682 15750
rect 96374 15739 96682 15748
rect 97460 15745 97488 15846
rect 97446 15736 97502 15745
rect 97446 15671 97502 15680
rect 96620 15496 96672 15502
rect 96620 15438 96672 15444
rect 96632 15065 96660 15438
rect 97448 15360 97500 15366
rect 97448 15302 97500 15308
rect 97034 15260 97342 15269
rect 97034 15258 97040 15260
rect 97096 15258 97120 15260
rect 97176 15258 97200 15260
rect 97256 15258 97280 15260
rect 97336 15258 97342 15260
rect 97096 15206 97098 15258
rect 97278 15206 97280 15258
rect 97034 15204 97040 15206
rect 97096 15204 97120 15206
rect 97176 15204 97200 15206
rect 97256 15204 97280 15206
rect 97336 15204 97342 15206
rect 97034 15195 97342 15204
rect 97460 15065 97488 15302
rect 96618 15056 96674 15065
rect 96618 14991 96674 15000
rect 97446 15056 97502 15065
rect 97446 14991 97502 15000
rect 96374 14716 96682 14725
rect 96374 14714 96380 14716
rect 96436 14714 96460 14716
rect 96516 14714 96540 14716
rect 96596 14714 96620 14716
rect 96676 14714 96682 14716
rect 96436 14662 96438 14714
rect 96618 14662 96620 14714
rect 96374 14660 96380 14662
rect 96436 14660 96460 14662
rect 96516 14660 96540 14662
rect 96596 14660 96620 14662
rect 96676 14660 96682 14662
rect 96374 14651 96682 14660
rect 97034 14172 97342 14181
rect 97034 14170 97040 14172
rect 97096 14170 97120 14172
rect 97176 14170 97200 14172
rect 97256 14170 97280 14172
rect 97336 14170 97342 14172
rect 97096 14118 97098 14170
rect 97278 14118 97280 14170
rect 97034 14116 97040 14118
rect 97096 14116 97120 14118
rect 97176 14116 97200 14118
rect 97256 14116 97280 14118
rect 97336 14116 97342 14118
rect 97034 14107 97342 14116
rect 97448 14068 97500 14074
rect 97448 14010 97500 14016
rect 97262 13968 97318 13977
rect 97262 13903 97264 13912
rect 97316 13903 97318 13912
rect 97264 13874 97316 13880
rect 97460 13705 97488 14010
rect 97446 13696 97502 13705
rect 96374 13628 96682 13637
rect 97446 13631 97502 13640
rect 96374 13626 96380 13628
rect 96436 13626 96460 13628
rect 96516 13626 96540 13628
rect 96596 13626 96620 13628
rect 96676 13626 96682 13628
rect 96436 13574 96438 13626
rect 96618 13574 96620 13626
rect 96374 13572 96380 13574
rect 96436 13572 96460 13574
rect 96516 13572 96540 13574
rect 96596 13572 96620 13574
rect 96676 13572 96682 13574
rect 96374 13563 96682 13572
rect 96620 13320 96672 13326
rect 96620 13262 96672 13268
rect 96632 12889 96660 13262
rect 97448 13184 97500 13190
rect 97448 13126 97500 13132
rect 97034 13084 97342 13093
rect 97034 13082 97040 13084
rect 97096 13082 97120 13084
rect 97176 13082 97200 13084
rect 97256 13082 97280 13084
rect 97336 13082 97342 13084
rect 97096 13030 97098 13082
rect 97278 13030 97280 13082
rect 97034 13028 97040 13030
rect 97096 13028 97120 13030
rect 97176 13028 97200 13030
rect 97256 13028 97280 13030
rect 97336 13028 97342 13030
rect 97034 13019 97342 13028
rect 97460 13025 97488 13126
rect 97446 13016 97502 13025
rect 97446 12951 97502 12960
rect 96618 12880 96674 12889
rect 96618 12815 96674 12824
rect 96374 12540 96682 12549
rect 96374 12538 96380 12540
rect 96436 12538 96460 12540
rect 96516 12538 96540 12540
rect 96596 12538 96620 12540
rect 96676 12538 96682 12540
rect 96436 12486 96438 12538
rect 96618 12486 96620 12538
rect 96374 12484 96380 12486
rect 96436 12484 96460 12486
rect 96516 12484 96540 12486
rect 96596 12484 96620 12486
rect 96676 12484 96682 12486
rect 96374 12475 96682 12484
rect 97034 11996 97342 12005
rect 97034 11994 97040 11996
rect 97096 11994 97120 11996
rect 97176 11994 97200 11996
rect 97256 11994 97280 11996
rect 97336 11994 97342 11996
rect 97096 11942 97098 11994
rect 97278 11942 97280 11994
rect 97034 11940 97040 11942
rect 97096 11940 97120 11942
rect 97176 11940 97200 11942
rect 97256 11940 97280 11942
rect 97336 11940 97342 11942
rect 97034 11931 97342 11940
rect 97262 11792 97318 11801
rect 97262 11727 97264 11736
rect 97316 11727 97318 11736
rect 97264 11698 97316 11704
rect 97446 11656 97502 11665
rect 97446 11591 97448 11600
rect 97500 11591 97502 11600
rect 97448 11562 97500 11568
rect 96374 11452 96682 11461
rect 96374 11450 96380 11452
rect 96436 11450 96460 11452
rect 96516 11450 96540 11452
rect 96596 11450 96620 11452
rect 96676 11450 96682 11452
rect 96436 11398 96438 11450
rect 96618 11398 96620 11450
rect 96374 11396 96380 11398
rect 96436 11396 96460 11398
rect 96516 11396 96540 11398
rect 96596 11396 96620 11398
rect 96676 11396 96682 11398
rect 96374 11387 96682 11396
rect 97034 10908 97342 10917
rect 97034 10906 97040 10908
rect 97096 10906 97120 10908
rect 97176 10906 97200 10908
rect 97256 10906 97280 10908
rect 97336 10906 97342 10908
rect 97096 10854 97098 10906
rect 97278 10854 97280 10906
rect 97034 10852 97040 10854
rect 97096 10852 97120 10854
rect 97176 10852 97200 10854
rect 97256 10852 97280 10854
rect 97336 10852 97342 10854
rect 97034 10843 97342 10852
rect 96374 10364 96682 10373
rect 96374 10362 96380 10364
rect 96436 10362 96460 10364
rect 96516 10362 96540 10364
rect 96596 10362 96620 10364
rect 96676 10362 96682 10364
rect 96436 10310 96438 10362
rect 96618 10310 96620 10362
rect 96374 10308 96380 10310
rect 96436 10308 96460 10310
rect 96516 10308 96540 10310
rect 96596 10308 96620 10310
rect 96676 10308 96682 10310
rect 96374 10299 96682 10308
rect 97034 9820 97342 9829
rect 97034 9818 97040 9820
rect 97096 9818 97120 9820
rect 97176 9818 97200 9820
rect 97256 9818 97280 9820
rect 97336 9818 97342 9820
rect 97096 9766 97098 9818
rect 97278 9766 97280 9818
rect 97034 9764 97040 9766
rect 97096 9764 97120 9766
rect 97176 9764 97200 9766
rect 97256 9764 97280 9766
rect 97336 9764 97342 9766
rect 97034 9755 97342 9764
rect 96374 9276 96682 9285
rect 96374 9274 96380 9276
rect 96436 9274 96460 9276
rect 96516 9274 96540 9276
rect 96596 9274 96620 9276
rect 96676 9274 96682 9276
rect 96436 9222 96438 9274
rect 96618 9222 96620 9274
rect 96374 9220 96380 9222
rect 96436 9220 96460 9222
rect 96516 9220 96540 9222
rect 96596 9220 96620 9222
rect 96676 9220 96682 9222
rect 96374 9211 96682 9220
rect 97034 8732 97342 8741
rect 97034 8730 97040 8732
rect 97096 8730 97120 8732
rect 97176 8730 97200 8732
rect 97256 8730 97280 8732
rect 97336 8730 97342 8732
rect 97096 8678 97098 8730
rect 97278 8678 97280 8730
rect 97034 8676 97040 8678
rect 97096 8676 97120 8678
rect 97176 8676 97200 8678
rect 97256 8676 97280 8678
rect 97336 8676 97342 8678
rect 97034 8667 97342 8676
rect 97540 8492 97592 8498
rect 97540 8434 97592 8440
rect 97552 8265 97580 8434
rect 97538 8256 97594 8265
rect 96374 8188 96682 8197
rect 97538 8191 97594 8200
rect 96374 8186 96380 8188
rect 96436 8186 96460 8188
rect 96516 8186 96540 8188
rect 96596 8186 96620 8188
rect 96676 8186 96682 8188
rect 54484 8152 54536 8158
rect 54188 8100 54484 8106
rect 91928 8152 91980 8158
rect 54188 8094 54536 8100
rect 54188 8092 54524 8094
rect 51966 7834 51994 8092
rect 53070 7834 53098 8092
rect 54174 8078 54524 8092
rect 54174 7834 54202 8078
rect 51966 7806 52040 7834
rect 53070 7806 53144 7834
rect 50620 5908 50672 5914
rect 50620 5850 50672 5856
rect 51080 5908 51132 5914
rect 51080 5850 51132 5856
rect 52012 5778 52040 7806
rect 52000 5772 52052 5778
rect 52000 5714 52052 5720
rect 53116 5710 53144 7806
rect 54128 7806 54202 7834
rect 56382 7834 56410 8092
rect 57486 7834 57514 8092
rect 58604 8078 58756 8106
rect 59708 8078 60044 8106
rect 60812 8078 60964 8106
rect 56382 7806 56456 7834
rect 53104 5704 53156 5710
rect 53104 5646 53156 5652
rect 54128 5642 54156 7806
rect 54116 5636 54168 5642
rect 54116 5578 54168 5584
rect 48780 2644 48832 2650
rect 48780 2586 48832 2592
rect 45468 2508 45520 2514
rect 45468 2450 45520 2456
rect 46388 2508 46440 2514
rect 46388 2450 46440 2456
rect 47492 2508 47544 2514
rect 47492 2450 47544 2456
rect 56428 2446 56456 7806
rect 57440 7806 57514 7834
rect 57440 2446 57468 7806
rect 58728 2446 58756 8078
rect 60016 2446 60044 8078
rect 60936 2446 60964 8078
rect 61902 7834 61930 8092
rect 63020 8078 63264 8106
rect 61902 7806 61976 7834
rect 61948 2446 61976 7806
rect 63236 2446 63264 8078
rect 64110 7834 64138 8092
rect 65214 7834 65242 8092
rect 66332 8078 66760 8106
rect 67436 8078 67772 8106
rect 68540 8078 68692 8106
rect 64110 7806 64184 7834
rect 64156 2446 64184 7806
rect 65168 7806 65242 7834
rect 65168 2446 65196 7806
rect 65654 6012 65962 6021
rect 65654 6010 65660 6012
rect 65716 6010 65740 6012
rect 65796 6010 65820 6012
rect 65876 6010 65900 6012
rect 65956 6010 65962 6012
rect 65716 5958 65718 6010
rect 65898 5958 65900 6010
rect 65654 5956 65660 5958
rect 65716 5956 65740 5958
rect 65796 5956 65820 5958
rect 65876 5956 65900 5958
rect 65956 5956 65962 5958
rect 65654 5947 65962 5956
rect 66314 5468 66622 5477
rect 66314 5466 66320 5468
rect 66376 5466 66400 5468
rect 66456 5466 66480 5468
rect 66536 5466 66560 5468
rect 66616 5466 66622 5468
rect 66376 5414 66378 5466
rect 66558 5414 66560 5466
rect 66314 5412 66320 5414
rect 66376 5412 66400 5414
rect 66456 5412 66480 5414
rect 66536 5412 66560 5414
rect 66616 5412 66622 5414
rect 66314 5403 66622 5412
rect 65654 4924 65962 4933
rect 65654 4922 65660 4924
rect 65716 4922 65740 4924
rect 65796 4922 65820 4924
rect 65876 4922 65900 4924
rect 65956 4922 65962 4924
rect 65716 4870 65718 4922
rect 65898 4870 65900 4922
rect 65654 4868 65660 4870
rect 65716 4868 65740 4870
rect 65796 4868 65820 4870
rect 65876 4868 65900 4870
rect 65956 4868 65962 4870
rect 65654 4859 65962 4868
rect 66314 4380 66622 4389
rect 66314 4378 66320 4380
rect 66376 4378 66400 4380
rect 66456 4378 66480 4380
rect 66536 4378 66560 4380
rect 66616 4378 66622 4380
rect 66376 4326 66378 4378
rect 66558 4326 66560 4378
rect 66314 4324 66320 4326
rect 66376 4324 66400 4326
rect 66456 4324 66480 4326
rect 66536 4324 66560 4326
rect 66616 4324 66622 4326
rect 66314 4315 66622 4324
rect 65654 3836 65962 3845
rect 65654 3834 65660 3836
rect 65716 3834 65740 3836
rect 65796 3834 65820 3836
rect 65876 3834 65900 3836
rect 65956 3834 65962 3836
rect 65716 3782 65718 3834
rect 65898 3782 65900 3834
rect 65654 3780 65660 3782
rect 65716 3780 65740 3782
rect 65796 3780 65820 3782
rect 65876 3780 65900 3782
rect 65956 3780 65962 3782
rect 65654 3771 65962 3780
rect 66314 3292 66622 3301
rect 66314 3290 66320 3292
rect 66376 3290 66400 3292
rect 66456 3290 66480 3292
rect 66536 3290 66560 3292
rect 66616 3290 66622 3292
rect 66376 3238 66378 3290
rect 66558 3238 66560 3290
rect 66314 3236 66320 3238
rect 66376 3236 66400 3238
rect 66456 3236 66480 3238
rect 66536 3236 66560 3238
rect 66616 3236 66622 3238
rect 66314 3227 66622 3236
rect 65654 2748 65962 2757
rect 65654 2746 65660 2748
rect 65716 2746 65740 2748
rect 65796 2746 65820 2748
rect 65876 2746 65900 2748
rect 65956 2746 65962 2748
rect 65716 2694 65718 2746
rect 65898 2694 65900 2746
rect 65654 2692 65660 2694
rect 65716 2692 65740 2694
rect 65796 2692 65820 2694
rect 65876 2692 65900 2694
rect 65956 2692 65962 2694
rect 65654 2683 65962 2692
rect 66732 2446 66760 8078
rect 67744 2446 67772 8078
rect 68664 2446 68692 8078
rect 69630 7834 69658 8092
rect 70748 8078 70992 8106
rect 69630 7806 69704 7834
rect 69676 2446 69704 7806
rect 70964 2446 70992 8078
rect 71838 7834 71866 8092
rect 72942 7834 72970 8092
rect 74060 8078 74212 8106
rect 75164 8078 75500 8106
rect 71838 7806 71912 7834
rect 71884 2446 71912 7806
rect 72896 7806 72970 7834
rect 72896 2446 72924 7806
rect 74184 2650 74212 8078
rect 75472 2650 75500 8078
rect 76254 7834 76282 8092
rect 77358 7834 77386 8092
rect 78476 8078 78720 8106
rect 76254 7806 76328 7834
rect 77358 7806 77432 7834
rect 76300 2650 76328 7806
rect 77404 2650 77432 7806
rect 78692 2650 78720 8078
rect 79566 7834 79594 8092
rect 80684 8078 80836 8106
rect 81788 8078 81940 8106
rect 82892 8078 83228 8106
rect 79520 7806 79594 7834
rect 79520 2650 79548 7806
rect 80808 2650 80836 8078
rect 81912 2650 81940 8078
rect 83200 2650 83228 8078
rect 83982 7834 84010 8092
rect 85086 7834 85114 8092
rect 86204 8078 86448 8106
rect 83982 7806 84056 7834
rect 85086 7806 85160 7834
rect 84028 2650 84056 7806
rect 85132 2650 85160 7806
rect 74172 2644 74224 2650
rect 74172 2586 74224 2592
rect 75460 2644 75512 2650
rect 75460 2586 75512 2592
rect 76288 2644 76340 2650
rect 76288 2586 76340 2592
rect 77392 2644 77444 2650
rect 77392 2586 77444 2592
rect 78680 2644 78732 2650
rect 78680 2586 78732 2592
rect 79508 2644 79560 2650
rect 79508 2586 79560 2592
rect 80796 2644 80848 2650
rect 80796 2586 80848 2592
rect 81900 2644 81952 2650
rect 81900 2586 81952 2592
rect 83188 2644 83240 2650
rect 83188 2586 83240 2592
rect 84016 2644 84068 2650
rect 84016 2586 84068 2592
rect 85120 2644 85172 2650
rect 85120 2586 85172 2592
rect 86420 2582 86448 8078
rect 87294 7834 87322 8092
rect 88412 8078 88748 8106
rect 89516 8078 89852 8106
rect 96436 8134 96438 8186
rect 96618 8134 96620 8186
rect 96374 8132 96380 8134
rect 96436 8132 96460 8134
rect 96516 8132 96540 8134
rect 96596 8132 96620 8134
rect 96676 8132 96682 8134
rect 96374 8123 96682 8132
rect 91928 8094 91980 8100
rect 87294 7806 87368 7834
rect 86408 2576 86460 2582
rect 86408 2518 86460 2524
rect 87340 2514 87368 7806
rect 88720 2514 88748 8078
rect 89536 2848 89588 2854
rect 89536 2790 89588 2796
rect 87328 2508 87380 2514
rect 87328 2450 87380 2456
rect 88708 2508 88760 2514
rect 88708 2450 88760 2456
rect 89548 2446 89576 2790
rect 89824 2514 89852 8078
rect 97034 7644 97342 7653
rect 97034 7642 97040 7644
rect 97096 7642 97120 7644
rect 97176 7642 97200 7644
rect 97256 7642 97280 7644
rect 97336 7642 97342 7644
rect 97096 7590 97098 7642
rect 97278 7590 97280 7642
rect 97034 7588 97040 7590
rect 97096 7588 97120 7590
rect 97176 7588 97200 7590
rect 97256 7588 97280 7590
rect 97336 7588 97342 7590
rect 97034 7579 97342 7588
rect 96374 7100 96682 7109
rect 96374 7098 96380 7100
rect 96436 7098 96460 7100
rect 96516 7098 96540 7100
rect 96596 7098 96620 7100
rect 96676 7098 96682 7100
rect 96436 7046 96438 7098
rect 96618 7046 96620 7098
rect 96374 7044 96380 7046
rect 96436 7044 96460 7046
rect 96516 7044 96540 7046
rect 96596 7044 96620 7046
rect 96676 7044 96682 7046
rect 96374 7035 96682 7044
rect 97034 6556 97342 6565
rect 97034 6554 97040 6556
rect 97096 6554 97120 6556
rect 97176 6554 97200 6556
rect 97256 6554 97280 6556
rect 97336 6554 97342 6556
rect 97096 6502 97098 6554
rect 97278 6502 97280 6554
rect 97034 6500 97040 6502
rect 97096 6500 97120 6502
rect 97176 6500 97200 6502
rect 97256 6500 97280 6502
rect 97336 6500 97342 6502
rect 97034 6491 97342 6500
rect 96374 6012 96682 6021
rect 96374 6010 96380 6012
rect 96436 6010 96460 6012
rect 96516 6010 96540 6012
rect 96596 6010 96620 6012
rect 96676 6010 96682 6012
rect 96436 5958 96438 6010
rect 96618 5958 96620 6010
rect 96374 5956 96380 5958
rect 96436 5956 96460 5958
rect 96516 5956 96540 5958
rect 96596 5956 96620 5958
rect 96676 5956 96682 5958
rect 96374 5947 96682 5956
rect 97034 5468 97342 5477
rect 97034 5466 97040 5468
rect 97096 5466 97120 5468
rect 97176 5466 97200 5468
rect 97256 5466 97280 5468
rect 97336 5466 97342 5468
rect 97096 5414 97098 5466
rect 97278 5414 97280 5466
rect 97034 5412 97040 5414
rect 97096 5412 97120 5414
rect 97176 5412 97200 5414
rect 97256 5412 97280 5414
rect 97336 5412 97342 5414
rect 97034 5403 97342 5412
rect 96374 4924 96682 4933
rect 96374 4922 96380 4924
rect 96436 4922 96460 4924
rect 96516 4922 96540 4924
rect 96596 4922 96620 4924
rect 96676 4922 96682 4924
rect 96436 4870 96438 4922
rect 96618 4870 96620 4922
rect 96374 4868 96380 4870
rect 96436 4868 96460 4870
rect 96516 4868 96540 4870
rect 96596 4868 96620 4870
rect 96676 4868 96682 4870
rect 96374 4859 96682 4868
rect 97034 4380 97342 4389
rect 97034 4378 97040 4380
rect 97096 4378 97120 4380
rect 97176 4378 97200 4380
rect 97256 4378 97280 4380
rect 97336 4378 97342 4380
rect 97096 4326 97098 4378
rect 97278 4326 97280 4378
rect 97034 4324 97040 4326
rect 97096 4324 97120 4326
rect 97176 4324 97200 4326
rect 97256 4324 97280 4326
rect 97336 4324 97342 4326
rect 97034 4315 97342 4324
rect 96374 3836 96682 3845
rect 96374 3834 96380 3836
rect 96436 3834 96460 3836
rect 96516 3834 96540 3836
rect 96596 3834 96620 3836
rect 96676 3834 96682 3836
rect 96436 3782 96438 3834
rect 96618 3782 96620 3834
rect 96374 3780 96380 3782
rect 96436 3780 96460 3782
rect 96516 3780 96540 3782
rect 96596 3780 96620 3782
rect 96676 3780 96682 3782
rect 96374 3771 96682 3780
rect 97034 3292 97342 3301
rect 97034 3290 97040 3292
rect 97096 3290 97120 3292
rect 97176 3290 97200 3292
rect 97256 3290 97280 3292
rect 97336 3290 97342 3292
rect 97096 3238 97098 3290
rect 97278 3238 97280 3290
rect 97034 3236 97040 3238
rect 97096 3236 97120 3238
rect 97176 3236 97200 3238
rect 97256 3236 97280 3238
rect 97336 3236 97342 3238
rect 97034 3227 97342 3236
rect 96374 2748 96682 2757
rect 96374 2746 96380 2748
rect 96436 2746 96460 2748
rect 96516 2746 96540 2748
rect 96596 2746 96620 2748
rect 96676 2746 96682 2748
rect 96436 2694 96438 2746
rect 96618 2694 96620 2746
rect 96374 2692 96380 2694
rect 96436 2692 96460 2694
rect 96516 2692 96540 2694
rect 96596 2692 96620 2694
rect 96676 2692 96682 2694
rect 96374 2683 96682 2692
rect 89812 2508 89864 2514
rect 89812 2450 89864 2456
rect 14556 2440 14608 2446
rect 14556 2382 14608 2388
rect 15568 2440 15620 2446
rect 15568 2382 15620 2388
rect 16856 2440 16908 2446
rect 16856 2382 16908 2388
rect 17776 2440 17828 2446
rect 17776 2382 17828 2388
rect 18788 2440 18840 2446
rect 18788 2382 18840 2388
rect 20076 2440 20128 2446
rect 20076 2382 20128 2388
rect 20996 2440 21048 2446
rect 20996 2382 21048 2388
rect 22284 2440 22336 2446
rect 22284 2382 22336 2388
rect 23296 2440 23348 2446
rect 23296 2382 23348 2388
rect 24584 2440 24636 2446
rect 24584 2382 24636 2388
rect 25504 2440 25556 2446
rect 25504 2382 25556 2388
rect 26516 2440 26568 2446
rect 26516 2382 26568 2388
rect 27804 2440 27856 2446
rect 27804 2382 27856 2388
rect 29092 2440 29144 2446
rect 29092 2382 29144 2388
rect 30012 2440 30064 2446
rect 30012 2382 30064 2388
rect 31024 2440 31076 2446
rect 31024 2382 31076 2388
rect 56416 2440 56468 2446
rect 56416 2382 56468 2388
rect 57428 2440 57480 2446
rect 57428 2382 57480 2388
rect 58716 2440 58768 2446
rect 58716 2382 58768 2388
rect 60004 2440 60056 2446
rect 60004 2382 60056 2388
rect 60924 2440 60976 2446
rect 60924 2382 60976 2388
rect 61936 2440 61988 2446
rect 61936 2382 61988 2388
rect 63224 2440 63276 2446
rect 63224 2382 63276 2388
rect 64144 2440 64196 2446
rect 64144 2382 64196 2388
rect 65156 2440 65208 2446
rect 65156 2382 65208 2388
rect 66720 2440 66772 2446
rect 66720 2382 66772 2388
rect 67732 2440 67784 2446
rect 67732 2382 67784 2388
rect 68652 2440 68704 2446
rect 68652 2382 68704 2388
rect 69664 2440 69716 2446
rect 69664 2382 69716 2388
rect 70952 2440 71004 2446
rect 70952 2382 71004 2388
rect 71872 2440 71924 2446
rect 71872 2382 71924 2388
rect 72884 2440 72936 2446
rect 72884 2382 72936 2388
rect 89536 2440 89588 2446
rect 89536 2382 89588 2388
rect 12256 2304 12308 2310
rect 12256 2246 12308 2252
rect 14188 2304 14240 2310
rect 14188 2246 14240 2252
rect 15476 2304 15528 2310
rect 15476 2246 15528 2252
rect 16764 2304 16816 2310
rect 16764 2246 16816 2252
rect 17408 2304 17460 2310
rect 17408 2246 17460 2252
rect 18696 2304 18748 2310
rect 18696 2246 18748 2252
rect 19984 2304 20036 2310
rect 19984 2246 20036 2252
rect 21272 2304 21324 2310
rect 21272 2246 21324 2252
rect 21916 2304 21968 2310
rect 21916 2246 21968 2252
rect 23204 2304 23256 2310
rect 23204 2246 23256 2252
rect 24492 2304 24544 2310
rect 24492 2246 24544 2252
rect 25136 2304 25188 2310
rect 25136 2246 25188 2252
rect 26424 2304 26476 2310
rect 26424 2246 26476 2252
rect 27712 2304 27764 2310
rect 27712 2246 27764 2252
rect 29000 2304 29052 2310
rect 29000 2246 29052 2252
rect 29644 2304 29696 2310
rect 29644 2246 29696 2252
rect 30932 2304 30984 2310
rect 30932 2246 30984 2252
rect 32220 2304 32272 2310
rect 32220 2246 32272 2252
rect 32864 2304 32916 2310
rect 32864 2246 32916 2252
rect 34152 2304 34204 2310
rect 34152 2246 34204 2252
rect 35440 2304 35492 2310
rect 35440 2246 35492 2252
rect 36728 2304 36780 2310
rect 36728 2246 36780 2252
rect 37372 2304 37424 2310
rect 37372 2246 37424 2252
rect 38660 2304 38712 2310
rect 38660 2246 38712 2252
rect 39948 2304 40000 2310
rect 39948 2246 40000 2252
rect 40592 2304 40644 2310
rect 40592 2246 40644 2252
rect 41880 2304 41932 2310
rect 41880 2246 41932 2252
rect 43168 2304 43220 2310
rect 43168 2246 43220 2252
rect 44456 2304 44508 2310
rect 44456 2246 44508 2252
rect 45100 2304 45152 2310
rect 45100 2246 45152 2252
rect 46388 2304 46440 2310
rect 46388 2246 46440 2252
rect 47676 2304 47728 2310
rect 47676 2246 47728 2252
rect 48320 2304 48372 2310
rect 48320 2246 48372 2252
rect 56048 2304 56100 2310
rect 56048 2246 56100 2252
rect 57336 2304 57388 2310
rect 57336 2246 57388 2252
rect 58624 2304 58676 2310
rect 58624 2246 58676 2252
rect 59912 2304 59964 2310
rect 59912 2246 59964 2252
rect 60556 2304 60608 2310
rect 60556 2246 60608 2252
rect 61844 2304 61896 2310
rect 61844 2246 61896 2252
rect 63132 2304 63184 2310
rect 63132 2246 63184 2252
rect 63776 2304 63828 2310
rect 63776 2246 63828 2252
rect 65064 2304 65116 2310
rect 65064 2246 65116 2252
rect 66720 2304 66772 2310
rect 66720 2246 66772 2252
rect 67640 2304 67692 2310
rect 67640 2246 67692 2252
rect 68284 2304 68336 2310
rect 68284 2246 68336 2252
rect 69572 2304 69624 2310
rect 69572 2246 69624 2252
rect 70860 2304 70912 2310
rect 70860 2246 70912 2252
rect 71504 2304 71556 2310
rect 71504 2246 71556 2252
rect 72792 2304 72844 2310
rect 72792 2246 72844 2252
rect 74080 2304 74132 2310
rect 74080 2246 74132 2252
rect 75368 2304 75420 2310
rect 75368 2246 75420 2252
rect 76012 2304 76064 2310
rect 76012 2246 76064 2252
rect 77300 2304 77352 2310
rect 77300 2246 77352 2252
rect 78588 2304 78640 2310
rect 78588 2246 78640 2252
rect 79232 2304 79284 2310
rect 79232 2246 79284 2252
rect 80520 2304 80572 2310
rect 80520 2246 80572 2252
rect 81808 2304 81860 2310
rect 81808 2246 81860 2252
rect 83096 2304 83148 2310
rect 83096 2246 83148 2252
rect 83740 2304 83792 2310
rect 83740 2246 83792 2252
rect 85028 2304 85080 2310
rect 85028 2246 85080 2252
rect 86316 2304 86368 2310
rect 86316 2246 86368 2252
rect 86960 2304 87012 2310
rect 86960 2246 87012 2252
rect 88248 2304 88300 2310
rect 88248 2246 88300 2252
rect 12268 800 12296 2246
rect 14200 800 14228 2246
rect 15488 800 15516 2246
rect 16776 800 16804 2246
rect 17420 800 17448 2246
rect 18708 800 18736 2246
rect 19996 800 20024 2246
rect 21284 800 21312 2246
rect 21928 800 21956 2246
rect 23216 800 23244 2246
rect 24504 800 24532 2246
rect 25148 800 25176 2246
rect 26436 800 26464 2246
rect 27724 800 27752 2246
rect 29012 800 29040 2246
rect 29656 800 29684 2246
rect 30944 800 30972 2246
rect 32232 800 32260 2246
rect 32876 800 32904 2246
rect 34164 800 34192 2246
rect 35452 800 35480 2246
rect 35594 2204 35902 2213
rect 35594 2202 35600 2204
rect 35656 2202 35680 2204
rect 35736 2202 35760 2204
rect 35816 2202 35840 2204
rect 35896 2202 35902 2204
rect 35656 2150 35658 2202
rect 35838 2150 35840 2202
rect 35594 2148 35600 2150
rect 35656 2148 35680 2150
rect 35736 2148 35760 2150
rect 35816 2148 35840 2150
rect 35896 2148 35902 2150
rect 35594 2139 35902 2148
rect 36740 800 36768 2246
rect 37384 800 37412 2246
rect 38672 800 38700 2246
rect 39960 800 39988 2246
rect 40604 800 40632 2246
rect 41892 800 41920 2246
rect 43180 800 43208 2246
rect 44468 800 44496 2246
rect 45112 800 45140 2246
rect 46400 800 46428 2246
rect 47688 800 47716 2246
rect 48332 800 48360 2246
rect 56060 800 56088 2246
rect 57348 800 57376 2246
rect 58636 800 58664 2246
rect 59924 800 59952 2246
rect 60568 800 60596 2246
rect 61856 800 61884 2246
rect 63144 800 63172 2246
rect 63788 800 63816 2246
rect 65076 800 65104 2246
rect 66314 2204 66622 2213
rect 66314 2202 66320 2204
rect 66376 2202 66400 2204
rect 66456 2202 66480 2204
rect 66536 2202 66560 2204
rect 66616 2202 66622 2204
rect 66376 2150 66378 2202
rect 66558 2150 66560 2202
rect 66314 2148 66320 2150
rect 66376 2148 66400 2150
rect 66456 2148 66480 2150
rect 66536 2148 66560 2150
rect 66616 2148 66622 2150
rect 66314 2139 66622 2148
rect 66364 870 66484 898
rect 66364 800 66392 870
rect 10322 0 10378 800
rect 11610 0 11666 800
rect 12254 0 12310 800
rect 14186 0 14242 800
rect 15474 0 15530 800
rect 16762 0 16818 800
rect 17406 0 17462 800
rect 18694 0 18750 800
rect 19982 0 20038 800
rect 21270 0 21326 800
rect 21914 0 21970 800
rect 23202 0 23258 800
rect 24490 0 24546 800
rect 25134 0 25190 800
rect 26422 0 26478 800
rect 27710 0 27766 800
rect 28998 0 29054 800
rect 29642 0 29698 800
rect 30930 0 30986 800
rect 32218 0 32274 800
rect 32862 0 32918 800
rect 34150 0 34206 800
rect 35438 0 35494 800
rect 36726 0 36782 800
rect 37370 0 37426 800
rect 38658 0 38714 800
rect 39946 0 40002 800
rect 40590 0 40646 800
rect 41878 0 41934 800
rect 43166 0 43222 800
rect 44454 0 44510 800
rect 45098 0 45154 800
rect 46386 0 46442 800
rect 47674 0 47730 800
rect 48318 0 48374 800
rect 56046 0 56102 800
rect 57334 0 57390 800
rect 58622 0 58678 800
rect 59910 0 59966 800
rect 60554 0 60610 800
rect 61842 0 61898 800
rect 63130 0 63186 800
rect 63774 0 63830 800
rect 65062 0 65118 800
rect 66350 0 66406 800
rect 66456 762 66484 870
rect 66732 762 66760 2246
rect 67652 800 67680 2246
rect 68296 800 68324 2246
rect 69584 800 69612 2246
rect 70872 800 70900 2246
rect 71516 800 71544 2246
rect 72804 800 72832 2246
rect 74092 800 74120 2246
rect 75380 800 75408 2246
rect 76024 800 76052 2246
rect 77312 800 77340 2246
rect 78600 800 78628 2246
rect 79244 800 79272 2246
rect 80532 800 80560 2246
rect 81820 800 81848 2246
rect 83108 800 83136 2246
rect 83752 800 83780 2246
rect 85040 800 85068 2246
rect 86328 800 86356 2246
rect 86972 800 87000 2246
rect 88260 800 88288 2246
rect 89548 800 89576 2382
rect 97034 2204 97342 2213
rect 97034 2202 97040 2204
rect 97096 2202 97120 2204
rect 97176 2202 97200 2204
rect 97256 2202 97280 2204
rect 97336 2202 97342 2204
rect 97096 2150 97098 2202
rect 97278 2150 97280 2202
rect 97034 2148 97040 2150
rect 97096 2148 97120 2150
rect 97176 2148 97200 2150
rect 97256 2148 97280 2150
rect 97336 2148 97342 2150
rect 97034 2139 97342 2148
rect 66456 734 66760 762
rect 67638 0 67694 800
rect 68282 0 68338 800
rect 69570 0 69626 800
rect 70858 0 70914 800
rect 71502 0 71558 800
rect 72790 0 72846 800
rect 74078 0 74134 800
rect 75366 0 75422 800
rect 76010 0 76066 800
rect 77298 0 77354 800
rect 78586 0 78642 800
rect 79230 0 79286 800
rect 80518 0 80574 800
rect 81806 0 81862 800
rect 83094 0 83150 800
rect 83738 0 83794 800
rect 85026 0 85082 800
rect 86314 0 86370 800
rect 86958 0 87014 800
rect 88246 0 88302 800
rect 89534 0 89590 800
<< via2 >>
rect 4880 95770 4936 95772
rect 4960 95770 5016 95772
rect 5040 95770 5096 95772
rect 5120 95770 5176 95772
rect 4880 95718 4926 95770
rect 4926 95718 4936 95770
rect 4960 95718 4990 95770
rect 4990 95718 5002 95770
rect 5002 95718 5016 95770
rect 5040 95718 5054 95770
rect 5054 95718 5066 95770
rect 5066 95718 5096 95770
rect 5120 95718 5130 95770
rect 5130 95718 5176 95770
rect 4880 95716 4936 95718
rect 4960 95716 5016 95718
rect 5040 95716 5096 95718
rect 5120 95716 5176 95718
rect 4220 95226 4276 95228
rect 4300 95226 4356 95228
rect 4380 95226 4436 95228
rect 4460 95226 4516 95228
rect 4220 95174 4266 95226
rect 4266 95174 4276 95226
rect 4300 95174 4330 95226
rect 4330 95174 4342 95226
rect 4342 95174 4356 95226
rect 4380 95174 4394 95226
rect 4394 95174 4406 95226
rect 4406 95174 4436 95226
rect 4460 95174 4470 95226
rect 4470 95174 4516 95226
rect 4220 95172 4276 95174
rect 4300 95172 4356 95174
rect 4380 95172 4436 95174
rect 4460 95172 4516 95174
rect 4880 94682 4936 94684
rect 4960 94682 5016 94684
rect 5040 94682 5096 94684
rect 5120 94682 5176 94684
rect 4880 94630 4926 94682
rect 4926 94630 4936 94682
rect 4960 94630 4990 94682
rect 4990 94630 5002 94682
rect 5002 94630 5016 94682
rect 5040 94630 5054 94682
rect 5054 94630 5066 94682
rect 5066 94630 5096 94682
rect 5120 94630 5130 94682
rect 5130 94630 5176 94682
rect 4880 94628 4936 94630
rect 4960 94628 5016 94630
rect 5040 94628 5096 94630
rect 5120 94628 5176 94630
rect 4220 94138 4276 94140
rect 4300 94138 4356 94140
rect 4380 94138 4436 94140
rect 4460 94138 4516 94140
rect 4220 94086 4266 94138
rect 4266 94086 4276 94138
rect 4300 94086 4330 94138
rect 4330 94086 4342 94138
rect 4342 94086 4356 94138
rect 4380 94086 4394 94138
rect 4394 94086 4406 94138
rect 4406 94086 4436 94138
rect 4460 94086 4470 94138
rect 4470 94086 4516 94138
rect 4220 94084 4276 94086
rect 4300 94084 4356 94086
rect 4380 94084 4436 94086
rect 4460 94084 4516 94086
rect 4880 93594 4936 93596
rect 4960 93594 5016 93596
rect 5040 93594 5096 93596
rect 5120 93594 5176 93596
rect 4880 93542 4926 93594
rect 4926 93542 4936 93594
rect 4960 93542 4990 93594
rect 4990 93542 5002 93594
rect 5002 93542 5016 93594
rect 5040 93542 5054 93594
rect 5054 93542 5066 93594
rect 5066 93542 5096 93594
rect 5120 93542 5130 93594
rect 5130 93542 5176 93594
rect 4880 93540 4936 93542
rect 4960 93540 5016 93542
rect 5040 93540 5096 93542
rect 5120 93540 5176 93542
rect 4220 93050 4276 93052
rect 4300 93050 4356 93052
rect 4380 93050 4436 93052
rect 4460 93050 4516 93052
rect 4220 92998 4266 93050
rect 4266 92998 4276 93050
rect 4300 92998 4330 93050
rect 4330 92998 4342 93050
rect 4342 92998 4356 93050
rect 4380 92998 4394 93050
rect 4394 92998 4406 93050
rect 4406 92998 4436 93050
rect 4460 92998 4470 93050
rect 4470 92998 4516 93050
rect 4220 92996 4276 92998
rect 4300 92996 4356 92998
rect 4380 92996 4436 92998
rect 4460 92996 4516 92998
rect 4880 92506 4936 92508
rect 4960 92506 5016 92508
rect 5040 92506 5096 92508
rect 5120 92506 5176 92508
rect 4880 92454 4926 92506
rect 4926 92454 4936 92506
rect 4960 92454 4990 92506
rect 4990 92454 5002 92506
rect 5002 92454 5016 92506
rect 5040 92454 5054 92506
rect 5054 92454 5066 92506
rect 5066 92454 5096 92506
rect 5120 92454 5130 92506
rect 5130 92454 5176 92506
rect 4880 92452 4936 92454
rect 4960 92452 5016 92454
rect 5040 92452 5096 92454
rect 5120 92452 5176 92454
rect 4220 91962 4276 91964
rect 4300 91962 4356 91964
rect 4380 91962 4436 91964
rect 4460 91962 4516 91964
rect 4220 91910 4266 91962
rect 4266 91910 4276 91962
rect 4300 91910 4330 91962
rect 4330 91910 4342 91962
rect 4342 91910 4356 91962
rect 4380 91910 4394 91962
rect 4394 91910 4406 91962
rect 4406 91910 4436 91962
rect 4460 91910 4470 91962
rect 4470 91910 4516 91962
rect 4220 91908 4276 91910
rect 4300 91908 4356 91910
rect 4380 91908 4436 91910
rect 4460 91908 4516 91910
rect 4880 91418 4936 91420
rect 4960 91418 5016 91420
rect 5040 91418 5096 91420
rect 5120 91418 5176 91420
rect 4880 91366 4926 91418
rect 4926 91366 4936 91418
rect 4960 91366 4990 91418
rect 4990 91366 5002 91418
rect 5002 91366 5016 91418
rect 5040 91366 5054 91418
rect 5054 91366 5066 91418
rect 5066 91366 5096 91418
rect 5120 91366 5130 91418
rect 5130 91366 5176 91418
rect 4880 91364 4936 91366
rect 4960 91364 5016 91366
rect 5040 91364 5096 91366
rect 5120 91364 5176 91366
rect 4220 90874 4276 90876
rect 4300 90874 4356 90876
rect 4380 90874 4436 90876
rect 4460 90874 4516 90876
rect 4220 90822 4266 90874
rect 4266 90822 4276 90874
rect 4300 90822 4330 90874
rect 4330 90822 4342 90874
rect 4342 90822 4356 90874
rect 4380 90822 4394 90874
rect 4394 90822 4406 90874
rect 4406 90822 4436 90874
rect 4460 90822 4470 90874
rect 4470 90822 4516 90874
rect 4220 90820 4276 90822
rect 4300 90820 4356 90822
rect 4380 90820 4436 90822
rect 4460 90820 4516 90822
rect 4880 90330 4936 90332
rect 4960 90330 5016 90332
rect 5040 90330 5096 90332
rect 5120 90330 5176 90332
rect 4880 90278 4926 90330
rect 4926 90278 4936 90330
rect 4960 90278 4990 90330
rect 4990 90278 5002 90330
rect 5002 90278 5016 90330
rect 5040 90278 5054 90330
rect 5054 90278 5066 90330
rect 5066 90278 5096 90330
rect 5120 90278 5130 90330
rect 5130 90278 5176 90330
rect 4880 90276 4936 90278
rect 4960 90276 5016 90278
rect 5040 90276 5096 90278
rect 5120 90276 5176 90278
rect 4220 89786 4276 89788
rect 4300 89786 4356 89788
rect 4380 89786 4436 89788
rect 4460 89786 4516 89788
rect 4220 89734 4266 89786
rect 4266 89734 4276 89786
rect 4300 89734 4330 89786
rect 4330 89734 4342 89786
rect 4342 89734 4356 89786
rect 4380 89734 4394 89786
rect 4394 89734 4406 89786
rect 4406 89734 4436 89786
rect 4460 89734 4470 89786
rect 4470 89734 4516 89786
rect 4220 89732 4276 89734
rect 4300 89732 4356 89734
rect 4380 89732 4436 89734
rect 4460 89732 4516 89734
rect 4880 89242 4936 89244
rect 4960 89242 5016 89244
rect 5040 89242 5096 89244
rect 5120 89242 5176 89244
rect 4880 89190 4926 89242
rect 4926 89190 4936 89242
rect 4960 89190 4990 89242
rect 4990 89190 5002 89242
rect 5002 89190 5016 89242
rect 5040 89190 5054 89242
rect 5054 89190 5066 89242
rect 5066 89190 5096 89242
rect 5120 89190 5130 89242
rect 5130 89190 5176 89242
rect 4880 89188 4936 89190
rect 4960 89188 5016 89190
rect 5040 89188 5096 89190
rect 5120 89188 5176 89190
rect 4220 88698 4276 88700
rect 4300 88698 4356 88700
rect 4380 88698 4436 88700
rect 4460 88698 4516 88700
rect 4220 88646 4266 88698
rect 4266 88646 4276 88698
rect 4300 88646 4330 88698
rect 4330 88646 4342 88698
rect 4342 88646 4356 88698
rect 4380 88646 4394 88698
rect 4394 88646 4406 88698
rect 4406 88646 4436 88698
rect 4460 88646 4470 88698
rect 4470 88646 4516 88698
rect 4220 88644 4276 88646
rect 4300 88644 4356 88646
rect 4380 88644 4436 88646
rect 4460 88644 4516 88646
rect 4880 88154 4936 88156
rect 4960 88154 5016 88156
rect 5040 88154 5096 88156
rect 5120 88154 5176 88156
rect 4880 88102 4926 88154
rect 4926 88102 4936 88154
rect 4960 88102 4990 88154
rect 4990 88102 5002 88154
rect 5002 88102 5016 88154
rect 5040 88102 5054 88154
rect 5054 88102 5066 88154
rect 5066 88102 5096 88154
rect 5120 88102 5130 88154
rect 5130 88102 5176 88154
rect 4880 88100 4936 88102
rect 4960 88100 5016 88102
rect 5040 88100 5096 88102
rect 5120 88100 5176 88102
rect 4220 87610 4276 87612
rect 4300 87610 4356 87612
rect 4380 87610 4436 87612
rect 4460 87610 4516 87612
rect 4220 87558 4266 87610
rect 4266 87558 4276 87610
rect 4300 87558 4330 87610
rect 4330 87558 4342 87610
rect 4342 87558 4356 87610
rect 4380 87558 4394 87610
rect 4394 87558 4406 87610
rect 4406 87558 4436 87610
rect 4460 87558 4470 87610
rect 4470 87558 4516 87610
rect 4220 87556 4276 87558
rect 4300 87556 4356 87558
rect 4380 87556 4436 87558
rect 4460 87556 4516 87558
rect 846 87216 902 87272
rect 4880 87066 4936 87068
rect 4960 87066 5016 87068
rect 5040 87066 5096 87068
rect 5120 87066 5176 87068
rect 4880 87014 4926 87066
rect 4926 87014 4936 87066
rect 4960 87014 4990 87066
rect 4990 87014 5002 87066
rect 5002 87014 5016 87066
rect 5040 87014 5054 87066
rect 5054 87014 5066 87066
rect 5066 87014 5096 87066
rect 5120 87014 5130 87066
rect 5130 87014 5176 87066
rect 4880 87012 4936 87014
rect 4960 87012 5016 87014
rect 5040 87012 5096 87014
rect 5120 87012 5176 87014
rect 846 86572 848 86592
rect 848 86572 900 86592
rect 900 86572 902 86592
rect 846 86536 902 86572
rect 4220 86522 4276 86524
rect 4300 86522 4356 86524
rect 4380 86522 4436 86524
rect 4460 86522 4516 86524
rect 4220 86470 4266 86522
rect 4266 86470 4276 86522
rect 4300 86470 4330 86522
rect 4330 86470 4342 86522
rect 4342 86470 4356 86522
rect 4380 86470 4394 86522
rect 4394 86470 4406 86522
rect 4406 86470 4436 86522
rect 4460 86470 4470 86522
rect 4470 86470 4516 86522
rect 4220 86468 4276 86470
rect 4300 86468 4356 86470
rect 4380 86468 4436 86470
rect 4460 86468 4516 86470
rect 4880 85978 4936 85980
rect 4960 85978 5016 85980
rect 5040 85978 5096 85980
rect 5120 85978 5176 85980
rect 4880 85926 4926 85978
rect 4926 85926 4936 85978
rect 4960 85926 4990 85978
rect 4990 85926 5002 85978
rect 5002 85926 5016 85978
rect 5040 85926 5054 85978
rect 5054 85926 5066 85978
rect 5066 85926 5096 85978
rect 5120 85926 5130 85978
rect 5130 85926 5176 85978
rect 4880 85924 4936 85926
rect 4960 85924 5016 85926
rect 5040 85924 5096 85926
rect 5120 85924 5176 85926
rect 4220 85434 4276 85436
rect 4300 85434 4356 85436
rect 4380 85434 4436 85436
rect 4460 85434 4516 85436
rect 4220 85382 4266 85434
rect 4266 85382 4276 85434
rect 4300 85382 4330 85434
rect 4330 85382 4342 85434
rect 4342 85382 4356 85434
rect 4380 85382 4394 85434
rect 4394 85382 4406 85434
rect 4406 85382 4436 85434
rect 4460 85382 4470 85434
rect 4470 85382 4516 85434
rect 4220 85380 4276 85382
rect 4300 85380 4356 85382
rect 4380 85380 4436 85382
rect 4460 85380 4516 85382
rect 846 84940 848 84960
rect 848 84940 900 84960
rect 900 84940 902 84960
rect 846 84904 902 84940
rect 4880 84890 4936 84892
rect 4960 84890 5016 84892
rect 5040 84890 5096 84892
rect 5120 84890 5176 84892
rect 4880 84838 4926 84890
rect 4926 84838 4936 84890
rect 4960 84838 4990 84890
rect 4990 84838 5002 84890
rect 5002 84838 5016 84890
rect 5040 84838 5054 84890
rect 5054 84838 5066 84890
rect 5066 84838 5096 84890
rect 5120 84838 5130 84890
rect 5130 84838 5176 84890
rect 4880 84836 4936 84838
rect 4960 84836 5016 84838
rect 5040 84836 5096 84838
rect 5120 84836 5176 84838
rect 846 84516 902 84552
rect 846 84496 848 84516
rect 848 84496 900 84516
rect 900 84496 902 84516
rect 4220 84346 4276 84348
rect 4300 84346 4356 84348
rect 4380 84346 4436 84348
rect 4460 84346 4516 84348
rect 4220 84294 4266 84346
rect 4266 84294 4276 84346
rect 4300 84294 4330 84346
rect 4330 84294 4342 84346
rect 4342 84294 4356 84346
rect 4380 84294 4394 84346
rect 4394 84294 4406 84346
rect 4406 84294 4436 84346
rect 4460 84294 4470 84346
rect 4470 84294 4516 84346
rect 4220 84292 4276 84294
rect 4300 84292 4356 84294
rect 4380 84292 4436 84294
rect 4460 84292 4516 84294
rect 1674 84088 1730 84144
rect 4880 83802 4936 83804
rect 4960 83802 5016 83804
rect 5040 83802 5096 83804
rect 5120 83802 5176 83804
rect 4880 83750 4926 83802
rect 4926 83750 4936 83802
rect 4960 83750 4990 83802
rect 4990 83750 5002 83802
rect 5002 83750 5016 83802
rect 5040 83750 5054 83802
rect 5054 83750 5066 83802
rect 5066 83750 5096 83802
rect 5120 83750 5130 83802
rect 5130 83750 5176 83802
rect 4880 83748 4936 83750
rect 4960 83748 5016 83750
rect 5040 83748 5096 83750
rect 5120 83748 5176 83750
rect 4220 83258 4276 83260
rect 4300 83258 4356 83260
rect 4380 83258 4436 83260
rect 4460 83258 4516 83260
rect 4220 83206 4266 83258
rect 4266 83206 4276 83258
rect 4300 83206 4330 83258
rect 4330 83206 4342 83258
rect 4342 83206 4356 83258
rect 4380 83206 4394 83258
rect 4394 83206 4406 83258
rect 4406 83206 4436 83258
rect 4460 83206 4470 83258
rect 4470 83206 4516 83258
rect 4220 83204 4276 83206
rect 4300 83204 4356 83206
rect 4380 83204 4436 83206
rect 4460 83204 4516 83206
rect 846 83136 902 83192
rect 4880 82714 4936 82716
rect 4960 82714 5016 82716
rect 5040 82714 5096 82716
rect 5120 82714 5176 82716
rect 4880 82662 4926 82714
rect 4926 82662 4936 82714
rect 4960 82662 4990 82714
rect 4990 82662 5002 82714
rect 5002 82662 5016 82714
rect 5040 82662 5054 82714
rect 5054 82662 5066 82714
rect 5066 82662 5096 82714
rect 5120 82662 5130 82714
rect 5130 82662 5176 82714
rect 4880 82660 4936 82662
rect 4960 82660 5016 82662
rect 5040 82660 5096 82662
rect 5120 82660 5176 82662
rect 4220 82170 4276 82172
rect 4300 82170 4356 82172
rect 4380 82170 4436 82172
rect 4460 82170 4516 82172
rect 4220 82118 4266 82170
rect 4266 82118 4276 82170
rect 4300 82118 4330 82170
rect 4330 82118 4342 82170
rect 4342 82118 4356 82170
rect 4380 82118 4394 82170
rect 4394 82118 4406 82170
rect 4406 82118 4436 82170
rect 4460 82118 4470 82170
rect 4470 82118 4516 82170
rect 4220 82116 4276 82118
rect 4300 82116 4356 82118
rect 4380 82116 4436 82118
rect 4460 82116 4516 82118
rect 846 81776 902 81832
rect 4880 81626 4936 81628
rect 4960 81626 5016 81628
rect 5040 81626 5096 81628
rect 5120 81626 5176 81628
rect 4880 81574 4926 81626
rect 4926 81574 4936 81626
rect 4960 81574 4990 81626
rect 4990 81574 5002 81626
rect 5002 81574 5016 81626
rect 5040 81574 5054 81626
rect 5054 81574 5066 81626
rect 5066 81574 5096 81626
rect 5120 81574 5130 81626
rect 5130 81574 5176 81626
rect 4880 81572 4936 81574
rect 4960 81572 5016 81574
rect 5040 81572 5096 81574
rect 5120 81572 5176 81574
rect 846 81132 848 81152
rect 848 81132 900 81152
rect 900 81132 902 81152
rect 846 81096 902 81132
rect 4220 81082 4276 81084
rect 4300 81082 4356 81084
rect 4380 81082 4436 81084
rect 4460 81082 4516 81084
rect 4220 81030 4266 81082
rect 4266 81030 4276 81082
rect 4300 81030 4330 81082
rect 4330 81030 4342 81082
rect 4342 81030 4356 81082
rect 4380 81030 4394 81082
rect 4394 81030 4406 81082
rect 4406 81030 4436 81082
rect 4460 81030 4470 81082
rect 4470 81030 4516 81082
rect 4220 81028 4276 81030
rect 4300 81028 4356 81030
rect 4380 81028 4436 81030
rect 4460 81028 4516 81030
rect 4880 80538 4936 80540
rect 4960 80538 5016 80540
rect 5040 80538 5096 80540
rect 5120 80538 5176 80540
rect 4880 80486 4926 80538
rect 4926 80486 4936 80538
rect 4960 80486 4990 80538
rect 4990 80486 5002 80538
rect 5002 80486 5016 80538
rect 5040 80486 5054 80538
rect 5054 80486 5066 80538
rect 5066 80486 5096 80538
rect 5120 80486 5130 80538
rect 5130 80486 5176 80538
rect 4880 80484 4936 80486
rect 4960 80484 5016 80486
rect 5040 80484 5096 80486
rect 5120 80484 5176 80486
rect 4220 79994 4276 79996
rect 4300 79994 4356 79996
rect 4380 79994 4436 79996
rect 4460 79994 4516 79996
rect 4220 79942 4266 79994
rect 4266 79942 4276 79994
rect 4300 79942 4330 79994
rect 4330 79942 4342 79994
rect 4342 79942 4356 79994
rect 4380 79942 4394 79994
rect 4394 79942 4406 79994
rect 4406 79942 4436 79994
rect 4460 79942 4470 79994
rect 4470 79942 4516 79994
rect 4220 79940 4276 79942
rect 4300 79940 4356 79942
rect 4380 79940 4436 79942
rect 4460 79940 4516 79942
rect 846 79500 848 79520
rect 848 79500 900 79520
rect 900 79500 902 79520
rect 846 79464 902 79500
rect 4880 79450 4936 79452
rect 4960 79450 5016 79452
rect 5040 79450 5096 79452
rect 5120 79450 5176 79452
rect 4880 79398 4926 79450
rect 4926 79398 4936 79450
rect 4960 79398 4990 79450
rect 4990 79398 5002 79450
rect 5002 79398 5016 79450
rect 5040 79398 5054 79450
rect 5054 79398 5066 79450
rect 5066 79398 5096 79450
rect 5120 79398 5130 79450
rect 5130 79398 5176 79450
rect 4880 79396 4936 79398
rect 4960 79396 5016 79398
rect 5040 79396 5096 79398
rect 5120 79396 5176 79398
rect 846 79076 902 79112
rect 846 79056 848 79076
rect 848 79056 900 79076
rect 900 79056 902 79076
rect 4220 78906 4276 78908
rect 4300 78906 4356 78908
rect 4380 78906 4436 78908
rect 4460 78906 4516 78908
rect 4220 78854 4266 78906
rect 4266 78854 4276 78906
rect 4300 78854 4330 78906
rect 4330 78854 4342 78906
rect 4342 78854 4356 78906
rect 4380 78854 4394 78906
rect 4394 78854 4406 78906
rect 4406 78854 4436 78906
rect 4460 78854 4470 78906
rect 4470 78854 4516 78906
rect 4220 78852 4276 78854
rect 4300 78852 4356 78854
rect 4380 78852 4436 78854
rect 4460 78852 4516 78854
rect 4880 78362 4936 78364
rect 4960 78362 5016 78364
rect 5040 78362 5096 78364
rect 5120 78362 5176 78364
rect 4880 78310 4926 78362
rect 4926 78310 4936 78362
rect 4960 78310 4990 78362
rect 4990 78310 5002 78362
rect 5002 78310 5016 78362
rect 5040 78310 5054 78362
rect 5054 78310 5066 78362
rect 5066 78310 5096 78362
rect 5120 78310 5130 78362
rect 5130 78310 5176 78362
rect 4880 78308 4936 78310
rect 4960 78308 5016 78310
rect 5040 78308 5096 78310
rect 5120 78308 5176 78310
rect 4220 77818 4276 77820
rect 4300 77818 4356 77820
rect 4380 77818 4436 77820
rect 4460 77818 4516 77820
rect 4220 77766 4266 77818
rect 4266 77766 4276 77818
rect 4300 77766 4330 77818
rect 4330 77766 4342 77818
rect 4342 77766 4356 77818
rect 4380 77766 4394 77818
rect 4394 77766 4406 77818
rect 4406 77766 4436 77818
rect 4460 77766 4470 77818
rect 4470 77766 4516 77818
rect 4220 77764 4276 77766
rect 4300 77764 4356 77766
rect 4380 77764 4436 77766
rect 4460 77764 4516 77766
rect 846 77696 902 77752
rect 4880 77274 4936 77276
rect 4960 77274 5016 77276
rect 5040 77274 5096 77276
rect 5120 77274 5176 77276
rect 4880 77222 4926 77274
rect 4926 77222 4936 77274
rect 4960 77222 4990 77274
rect 4990 77222 5002 77274
rect 5002 77222 5016 77274
rect 5040 77222 5054 77274
rect 5054 77222 5066 77274
rect 5066 77222 5096 77274
rect 5120 77222 5130 77274
rect 5130 77222 5176 77274
rect 4880 77220 4936 77222
rect 4960 77220 5016 77222
rect 5040 77220 5096 77222
rect 5120 77220 5176 77222
rect 4220 76730 4276 76732
rect 4300 76730 4356 76732
rect 4380 76730 4436 76732
rect 4460 76730 4516 76732
rect 4220 76678 4266 76730
rect 4266 76678 4276 76730
rect 4300 76678 4330 76730
rect 4330 76678 4342 76730
rect 4342 76678 4356 76730
rect 4380 76678 4394 76730
rect 4394 76678 4406 76730
rect 4406 76678 4436 76730
rect 4460 76678 4470 76730
rect 4470 76678 4516 76730
rect 4220 76676 4276 76678
rect 4300 76676 4356 76678
rect 4380 76676 4436 76678
rect 4460 76676 4516 76678
rect 846 76336 902 76392
rect 4880 76186 4936 76188
rect 4960 76186 5016 76188
rect 5040 76186 5096 76188
rect 5120 76186 5176 76188
rect 4880 76134 4926 76186
rect 4926 76134 4936 76186
rect 4960 76134 4990 76186
rect 4990 76134 5002 76186
rect 5002 76134 5016 76186
rect 5040 76134 5054 76186
rect 5054 76134 5066 76186
rect 5066 76134 5096 76186
rect 5120 76134 5130 76186
rect 5130 76134 5176 76186
rect 4880 76132 4936 76134
rect 4960 76132 5016 76134
rect 5040 76132 5096 76134
rect 5120 76132 5176 76134
rect 846 75656 902 75712
rect 4220 75642 4276 75644
rect 4300 75642 4356 75644
rect 4380 75642 4436 75644
rect 4460 75642 4516 75644
rect 4220 75590 4266 75642
rect 4266 75590 4276 75642
rect 4300 75590 4330 75642
rect 4330 75590 4342 75642
rect 4342 75590 4356 75642
rect 4380 75590 4394 75642
rect 4394 75590 4406 75642
rect 4406 75590 4436 75642
rect 4460 75590 4470 75642
rect 4470 75590 4516 75642
rect 4220 75588 4276 75590
rect 4300 75588 4356 75590
rect 4380 75588 4436 75590
rect 4460 75588 4516 75590
rect 1674 75384 1730 75440
rect 4880 75098 4936 75100
rect 4960 75098 5016 75100
rect 5040 75098 5096 75100
rect 5120 75098 5176 75100
rect 4880 75046 4926 75098
rect 4926 75046 4936 75098
rect 4960 75046 4990 75098
rect 4990 75046 5002 75098
rect 5002 75046 5016 75098
rect 5040 75046 5054 75098
rect 5054 75046 5066 75098
rect 5066 75046 5096 75098
rect 5120 75046 5130 75098
rect 5130 75046 5176 75098
rect 4880 75044 4936 75046
rect 4960 75044 5016 75046
rect 5040 75044 5096 75046
rect 5120 75044 5176 75046
rect 4220 74554 4276 74556
rect 4300 74554 4356 74556
rect 4380 74554 4436 74556
rect 4460 74554 4516 74556
rect 4220 74502 4266 74554
rect 4266 74502 4276 74554
rect 4300 74502 4330 74554
rect 4330 74502 4342 74554
rect 4342 74502 4356 74554
rect 4380 74502 4394 74554
rect 4394 74502 4406 74554
rect 4406 74502 4436 74554
rect 4460 74502 4470 74554
rect 4470 74502 4516 74554
rect 4220 74500 4276 74502
rect 4300 74500 4356 74502
rect 4380 74500 4436 74502
rect 4460 74500 4516 74502
rect 846 74060 848 74080
rect 848 74060 900 74080
rect 900 74060 902 74080
rect 846 74024 902 74060
rect 4880 74010 4936 74012
rect 4960 74010 5016 74012
rect 5040 74010 5096 74012
rect 5120 74010 5176 74012
rect 4880 73958 4926 74010
rect 4926 73958 4936 74010
rect 4960 73958 4990 74010
rect 4990 73958 5002 74010
rect 5002 73958 5016 74010
rect 5040 73958 5054 74010
rect 5054 73958 5066 74010
rect 5066 73958 5096 74010
rect 5120 73958 5130 74010
rect 5130 73958 5176 74010
rect 4880 73956 4936 73958
rect 4960 73956 5016 73958
rect 5040 73956 5096 73958
rect 5120 73956 5176 73958
rect 846 73636 902 73672
rect 846 73616 848 73636
rect 848 73616 900 73636
rect 900 73616 902 73636
rect 4220 73466 4276 73468
rect 4300 73466 4356 73468
rect 4380 73466 4436 73468
rect 4460 73466 4516 73468
rect 4220 73414 4266 73466
rect 4266 73414 4276 73466
rect 4300 73414 4330 73466
rect 4330 73414 4342 73466
rect 4342 73414 4356 73466
rect 4380 73414 4394 73466
rect 4394 73414 4406 73466
rect 4406 73414 4436 73466
rect 4460 73414 4470 73466
rect 4470 73414 4516 73466
rect 4220 73412 4276 73414
rect 4300 73412 4356 73414
rect 4380 73412 4436 73414
rect 4460 73412 4516 73414
rect 4880 72922 4936 72924
rect 4960 72922 5016 72924
rect 5040 72922 5096 72924
rect 5120 72922 5176 72924
rect 4880 72870 4926 72922
rect 4926 72870 4936 72922
rect 4960 72870 4990 72922
rect 4990 72870 5002 72922
rect 5002 72870 5016 72922
rect 5040 72870 5054 72922
rect 5054 72870 5066 72922
rect 5066 72870 5096 72922
rect 5120 72870 5130 72922
rect 5130 72870 5176 72922
rect 4880 72868 4936 72870
rect 4960 72868 5016 72870
rect 5040 72868 5096 72870
rect 5120 72868 5176 72870
rect 4220 72378 4276 72380
rect 4300 72378 4356 72380
rect 4380 72378 4436 72380
rect 4460 72378 4516 72380
rect 4220 72326 4266 72378
rect 4266 72326 4276 72378
rect 4300 72326 4330 72378
rect 4330 72326 4342 72378
rect 4342 72326 4356 72378
rect 4380 72326 4394 72378
rect 4394 72326 4406 72378
rect 4406 72326 4436 72378
rect 4460 72326 4470 72378
rect 4470 72326 4516 72378
rect 4220 72324 4276 72326
rect 4300 72324 4356 72326
rect 4380 72324 4436 72326
rect 4460 72324 4516 72326
rect 846 72256 902 72312
rect 4880 71834 4936 71836
rect 4960 71834 5016 71836
rect 5040 71834 5096 71836
rect 5120 71834 5176 71836
rect 4880 71782 4926 71834
rect 4926 71782 4936 71834
rect 4960 71782 4990 71834
rect 4990 71782 5002 71834
rect 5002 71782 5016 71834
rect 5040 71782 5054 71834
rect 5054 71782 5066 71834
rect 5066 71782 5096 71834
rect 5120 71782 5130 71834
rect 5130 71782 5176 71834
rect 4880 71780 4936 71782
rect 4960 71780 5016 71782
rect 5040 71780 5096 71782
rect 5120 71780 5176 71782
rect 4220 71290 4276 71292
rect 4300 71290 4356 71292
rect 4380 71290 4436 71292
rect 4460 71290 4516 71292
rect 4220 71238 4266 71290
rect 4266 71238 4276 71290
rect 4300 71238 4330 71290
rect 4330 71238 4342 71290
rect 4342 71238 4356 71290
rect 4380 71238 4394 71290
rect 4394 71238 4406 71290
rect 4406 71238 4436 71290
rect 4460 71238 4470 71290
rect 4470 71238 4516 71290
rect 4220 71236 4276 71238
rect 4300 71236 4356 71238
rect 4380 71236 4436 71238
rect 4460 71236 4516 71238
rect 846 70896 902 70952
rect 4880 70746 4936 70748
rect 4960 70746 5016 70748
rect 5040 70746 5096 70748
rect 5120 70746 5176 70748
rect 4880 70694 4926 70746
rect 4926 70694 4936 70746
rect 4960 70694 4990 70746
rect 4990 70694 5002 70746
rect 5002 70694 5016 70746
rect 5040 70694 5054 70746
rect 5054 70694 5066 70746
rect 5066 70694 5096 70746
rect 5120 70694 5130 70746
rect 5130 70694 5176 70746
rect 4880 70692 4936 70694
rect 4960 70692 5016 70694
rect 5040 70692 5096 70694
rect 5120 70692 5176 70694
rect 1306 70080 1362 70136
rect 4220 70202 4276 70204
rect 4300 70202 4356 70204
rect 4380 70202 4436 70204
rect 4460 70202 4516 70204
rect 4220 70150 4266 70202
rect 4266 70150 4276 70202
rect 4300 70150 4330 70202
rect 4330 70150 4342 70202
rect 4342 70150 4356 70202
rect 4380 70150 4394 70202
rect 4394 70150 4406 70202
rect 4406 70150 4436 70202
rect 4460 70150 4470 70202
rect 4470 70150 4516 70202
rect 4220 70148 4276 70150
rect 4300 70148 4356 70150
rect 4380 70148 4436 70150
rect 4460 70148 4516 70150
rect 1582 69944 1638 70000
rect 4880 69658 4936 69660
rect 4960 69658 5016 69660
rect 5040 69658 5096 69660
rect 5120 69658 5176 69660
rect 4880 69606 4926 69658
rect 4926 69606 4936 69658
rect 4960 69606 4990 69658
rect 4990 69606 5002 69658
rect 5002 69606 5016 69658
rect 5040 69606 5054 69658
rect 5054 69606 5066 69658
rect 5066 69606 5096 69658
rect 5120 69606 5130 69658
rect 5130 69606 5176 69658
rect 4880 69604 4936 69606
rect 4960 69604 5016 69606
rect 5040 69604 5096 69606
rect 5120 69604 5176 69606
rect 4220 69114 4276 69116
rect 4300 69114 4356 69116
rect 4380 69114 4436 69116
rect 4460 69114 4516 69116
rect 4220 69062 4266 69114
rect 4266 69062 4276 69114
rect 4300 69062 4330 69114
rect 4330 69062 4342 69114
rect 4342 69062 4356 69114
rect 4380 69062 4394 69114
rect 4394 69062 4406 69114
rect 4406 69062 4436 69114
rect 4460 69062 4470 69114
rect 4470 69062 4516 69114
rect 4220 69060 4276 69062
rect 4300 69060 4356 69062
rect 4380 69060 4436 69062
rect 4460 69060 4516 69062
rect 1122 68740 1178 68776
rect 1122 68720 1124 68740
rect 1124 68720 1176 68740
rect 1176 68720 1178 68740
rect 4880 68570 4936 68572
rect 4960 68570 5016 68572
rect 5040 68570 5096 68572
rect 5120 68570 5176 68572
rect 4880 68518 4926 68570
rect 4926 68518 4936 68570
rect 4960 68518 4990 68570
rect 4990 68518 5002 68570
rect 5002 68518 5016 68570
rect 5040 68518 5054 68570
rect 5054 68518 5066 68570
rect 5066 68518 5096 68570
rect 5120 68518 5130 68570
rect 5130 68518 5176 68570
rect 4880 68516 4936 68518
rect 4960 68516 5016 68518
rect 5040 68516 5096 68518
rect 5120 68516 5176 68518
rect 1306 68040 1362 68096
rect 4220 68026 4276 68028
rect 4300 68026 4356 68028
rect 4380 68026 4436 68028
rect 4460 68026 4516 68028
rect 4220 67974 4266 68026
rect 4266 67974 4276 68026
rect 4300 67974 4330 68026
rect 4330 67974 4342 68026
rect 4342 67974 4356 68026
rect 4380 67974 4394 68026
rect 4394 67974 4406 68026
rect 4406 67974 4436 68026
rect 4460 67974 4470 68026
rect 4470 67974 4516 68026
rect 4220 67972 4276 67974
rect 4300 67972 4356 67974
rect 4380 67972 4436 67974
rect 4460 67972 4516 67974
rect 4880 67482 4936 67484
rect 4960 67482 5016 67484
rect 5040 67482 5096 67484
rect 5120 67482 5176 67484
rect 4880 67430 4926 67482
rect 4926 67430 4936 67482
rect 4960 67430 4990 67482
rect 4990 67430 5002 67482
rect 5002 67430 5016 67482
rect 5040 67430 5054 67482
rect 5054 67430 5066 67482
rect 5066 67430 5096 67482
rect 5120 67430 5130 67482
rect 5130 67430 5176 67482
rect 4880 67428 4936 67430
rect 4960 67428 5016 67430
rect 5040 67428 5096 67430
rect 5120 67428 5176 67430
rect 4220 66938 4276 66940
rect 4300 66938 4356 66940
rect 4380 66938 4436 66940
rect 4460 66938 4516 66940
rect 4220 66886 4266 66938
rect 4266 66886 4276 66938
rect 4300 66886 4330 66938
rect 4330 66886 4342 66938
rect 4342 66886 4356 66938
rect 4380 66886 4394 66938
rect 4394 66886 4406 66938
rect 4406 66886 4436 66938
rect 4460 66886 4470 66938
rect 4470 66886 4516 66938
rect 4220 66884 4276 66886
rect 4300 66884 4356 66886
rect 4380 66884 4436 66886
rect 4460 66884 4516 66886
rect 1306 66680 1362 66736
rect 4880 66394 4936 66396
rect 4960 66394 5016 66396
rect 5040 66394 5096 66396
rect 5120 66394 5176 66396
rect 4880 66342 4926 66394
rect 4926 66342 4936 66394
rect 4960 66342 4990 66394
rect 4990 66342 5002 66394
rect 5002 66342 5016 66394
rect 5040 66342 5054 66394
rect 5054 66342 5066 66394
rect 5066 66342 5096 66394
rect 5120 66342 5130 66394
rect 5130 66342 5176 66394
rect 4880 66340 4936 66342
rect 4960 66340 5016 66342
rect 5040 66340 5096 66342
rect 5120 66340 5176 66342
rect 4220 65850 4276 65852
rect 4300 65850 4356 65852
rect 4380 65850 4436 65852
rect 4460 65850 4516 65852
rect 4220 65798 4266 65850
rect 4266 65798 4276 65850
rect 4300 65798 4330 65850
rect 4330 65798 4342 65850
rect 4342 65798 4356 65850
rect 4380 65798 4394 65850
rect 4394 65798 4406 65850
rect 4406 65798 4436 65850
rect 4460 65798 4470 65850
rect 4470 65798 4516 65850
rect 4220 65796 4276 65798
rect 4300 65796 4356 65798
rect 4380 65796 4436 65798
rect 4460 65796 4516 65798
rect 1122 65320 1178 65376
rect 4880 65306 4936 65308
rect 4960 65306 5016 65308
rect 5040 65306 5096 65308
rect 5120 65306 5176 65308
rect 4880 65254 4926 65306
rect 4926 65254 4936 65306
rect 4960 65254 4990 65306
rect 4990 65254 5002 65306
rect 5002 65254 5016 65306
rect 5040 65254 5054 65306
rect 5054 65254 5066 65306
rect 5066 65254 5096 65306
rect 5120 65254 5130 65306
rect 5130 65254 5176 65306
rect 4880 65252 4936 65254
rect 4960 65252 5016 65254
rect 5040 65252 5096 65254
rect 5120 65252 5176 65254
rect 1306 64640 1362 64696
rect 4220 64762 4276 64764
rect 4300 64762 4356 64764
rect 4380 64762 4436 64764
rect 4460 64762 4516 64764
rect 4220 64710 4266 64762
rect 4266 64710 4276 64762
rect 4300 64710 4330 64762
rect 4330 64710 4342 64762
rect 4342 64710 4356 64762
rect 4380 64710 4394 64762
rect 4394 64710 4406 64762
rect 4406 64710 4436 64762
rect 4460 64710 4470 64762
rect 4470 64710 4516 64762
rect 4220 64708 4276 64710
rect 4300 64708 4356 64710
rect 4380 64708 4436 64710
rect 4460 64708 4516 64710
rect 1674 64504 1730 64560
rect 4880 64218 4936 64220
rect 4960 64218 5016 64220
rect 5040 64218 5096 64220
rect 5120 64218 5176 64220
rect 4880 64166 4926 64218
rect 4926 64166 4936 64218
rect 4960 64166 4990 64218
rect 4990 64166 5002 64218
rect 5002 64166 5016 64218
rect 5040 64166 5054 64218
rect 5054 64166 5066 64218
rect 5066 64166 5096 64218
rect 5120 64166 5130 64218
rect 5130 64166 5176 64218
rect 4880 64164 4936 64166
rect 4960 64164 5016 64166
rect 5040 64164 5096 64166
rect 5120 64164 5176 64166
rect 4220 63674 4276 63676
rect 4300 63674 4356 63676
rect 4380 63674 4436 63676
rect 4460 63674 4516 63676
rect 4220 63622 4266 63674
rect 4266 63622 4276 63674
rect 4300 63622 4330 63674
rect 4330 63622 4342 63674
rect 4342 63622 4356 63674
rect 4380 63622 4394 63674
rect 4394 63622 4406 63674
rect 4406 63622 4436 63674
rect 4460 63622 4470 63674
rect 4470 63622 4516 63674
rect 4220 63620 4276 63622
rect 4300 63620 4356 63622
rect 4380 63620 4436 63622
rect 4460 63620 4516 63622
rect 1122 63300 1178 63336
rect 1122 63280 1124 63300
rect 1124 63280 1176 63300
rect 1176 63280 1178 63300
rect 4880 63130 4936 63132
rect 4960 63130 5016 63132
rect 5040 63130 5096 63132
rect 5120 63130 5176 63132
rect 4880 63078 4926 63130
rect 4926 63078 4936 63130
rect 4960 63078 4990 63130
rect 4990 63078 5002 63130
rect 5002 63078 5016 63130
rect 5040 63078 5054 63130
rect 5054 63078 5066 63130
rect 5066 63078 5096 63130
rect 5120 63078 5130 63130
rect 5130 63078 5176 63130
rect 4880 63076 4936 63078
rect 4960 63076 5016 63078
rect 5040 63076 5096 63078
rect 5120 63076 5176 63078
rect 1306 62600 1362 62656
rect 4220 62586 4276 62588
rect 4300 62586 4356 62588
rect 4380 62586 4436 62588
rect 4460 62586 4516 62588
rect 4220 62534 4266 62586
rect 4266 62534 4276 62586
rect 4300 62534 4330 62586
rect 4330 62534 4342 62586
rect 4342 62534 4356 62586
rect 4380 62534 4394 62586
rect 4394 62534 4406 62586
rect 4406 62534 4436 62586
rect 4460 62534 4470 62586
rect 4470 62534 4516 62586
rect 4220 62532 4276 62534
rect 4300 62532 4356 62534
rect 4380 62532 4436 62534
rect 4460 62532 4516 62534
rect 4880 62042 4936 62044
rect 4960 62042 5016 62044
rect 5040 62042 5096 62044
rect 5120 62042 5176 62044
rect 4880 61990 4926 62042
rect 4926 61990 4936 62042
rect 4960 61990 4990 62042
rect 4990 61990 5002 62042
rect 5002 61990 5016 62042
rect 5040 61990 5054 62042
rect 5054 61990 5066 62042
rect 5066 61990 5096 62042
rect 5120 61990 5130 62042
rect 5130 61990 5176 62042
rect 4880 61988 4936 61990
rect 4960 61988 5016 61990
rect 5040 61988 5096 61990
rect 5120 61988 5176 61990
rect 4220 61498 4276 61500
rect 4300 61498 4356 61500
rect 4380 61498 4436 61500
rect 4460 61498 4516 61500
rect 4220 61446 4266 61498
rect 4266 61446 4276 61498
rect 4300 61446 4330 61498
rect 4330 61446 4342 61498
rect 4342 61446 4356 61498
rect 4380 61446 4394 61498
rect 4394 61446 4406 61498
rect 4406 61446 4436 61498
rect 4460 61446 4470 61498
rect 4470 61446 4516 61498
rect 4220 61444 4276 61446
rect 4300 61444 4356 61446
rect 4380 61444 4436 61446
rect 4460 61444 4516 61446
rect 1306 61240 1362 61296
rect 4880 60954 4936 60956
rect 4960 60954 5016 60956
rect 5040 60954 5096 60956
rect 5120 60954 5176 60956
rect 4880 60902 4926 60954
rect 4926 60902 4936 60954
rect 4960 60902 4990 60954
rect 4990 60902 5002 60954
rect 5002 60902 5016 60954
rect 5040 60902 5054 60954
rect 5054 60902 5066 60954
rect 5066 60902 5096 60954
rect 5120 60902 5130 60954
rect 5130 60902 5176 60954
rect 4880 60900 4936 60902
rect 4960 60900 5016 60902
rect 5040 60900 5096 60902
rect 5120 60900 5176 60902
rect 4220 60410 4276 60412
rect 4300 60410 4356 60412
rect 4380 60410 4436 60412
rect 4460 60410 4516 60412
rect 4220 60358 4266 60410
rect 4266 60358 4276 60410
rect 4300 60358 4330 60410
rect 4330 60358 4342 60410
rect 4342 60358 4356 60410
rect 4380 60358 4394 60410
rect 4394 60358 4406 60410
rect 4406 60358 4436 60410
rect 4460 60358 4470 60410
rect 4470 60358 4516 60410
rect 4220 60356 4276 60358
rect 4300 60356 4356 60358
rect 4380 60356 4436 60358
rect 4460 60356 4516 60358
rect 1214 59880 1270 59936
rect 4880 59866 4936 59868
rect 4960 59866 5016 59868
rect 5040 59866 5096 59868
rect 5120 59866 5176 59868
rect 4880 59814 4926 59866
rect 4926 59814 4936 59866
rect 4960 59814 4990 59866
rect 4990 59814 5002 59866
rect 5002 59814 5016 59866
rect 5040 59814 5054 59866
rect 5054 59814 5066 59866
rect 5066 59814 5096 59866
rect 5120 59814 5130 59866
rect 5130 59814 5176 59866
rect 4880 59812 4936 59814
rect 4960 59812 5016 59814
rect 5040 59812 5096 59814
rect 5120 59812 5176 59814
rect 1214 59200 1270 59256
rect 4220 59322 4276 59324
rect 4300 59322 4356 59324
rect 4380 59322 4436 59324
rect 4460 59322 4516 59324
rect 4220 59270 4266 59322
rect 4266 59270 4276 59322
rect 4300 59270 4330 59322
rect 4330 59270 4342 59322
rect 4342 59270 4356 59322
rect 4380 59270 4394 59322
rect 4394 59270 4406 59322
rect 4406 59270 4436 59322
rect 4460 59270 4470 59322
rect 4470 59270 4516 59322
rect 4220 59268 4276 59270
rect 4300 59268 4356 59270
rect 4380 59268 4436 59270
rect 4460 59268 4516 59270
rect 1582 59064 1638 59120
rect 4880 58778 4936 58780
rect 4960 58778 5016 58780
rect 5040 58778 5096 58780
rect 5120 58778 5176 58780
rect 4880 58726 4926 58778
rect 4926 58726 4936 58778
rect 4960 58726 4990 58778
rect 4990 58726 5002 58778
rect 5002 58726 5016 58778
rect 5040 58726 5054 58778
rect 5054 58726 5066 58778
rect 5066 58726 5096 58778
rect 5120 58726 5130 58778
rect 5130 58726 5176 58778
rect 4880 58724 4936 58726
rect 4960 58724 5016 58726
rect 5040 58724 5096 58726
rect 5120 58724 5176 58726
rect 4220 58234 4276 58236
rect 4300 58234 4356 58236
rect 4380 58234 4436 58236
rect 4460 58234 4516 58236
rect 4220 58182 4266 58234
rect 4266 58182 4276 58234
rect 4300 58182 4330 58234
rect 4330 58182 4342 58234
rect 4342 58182 4356 58234
rect 4380 58182 4394 58234
rect 4394 58182 4406 58234
rect 4406 58182 4436 58234
rect 4460 58182 4470 58234
rect 4470 58182 4516 58234
rect 4220 58180 4276 58182
rect 4300 58180 4356 58182
rect 4380 58180 4436 58182
rect 4460 58180 4516 58182
rect 1582 57976 1638 58032
rect 1306 57876 1308 57896
rect 1308 57876 1360 57896
rect 1360 57876 1362 57896
rect 1306 57840 1362 57876
rect 4880 57690 4936 57692
rect 4960 57690 5016 57692
rect 5040 57690 5096 57692
rect 5120 57690 5176 57692
rect 4880 57638 4926 57690
rect 4926 57638 4936 57690
rect 4960 57638 4990 57690
rect 4990 57638 5002 57690
rect 5002 57638 5016 57690
rect 5040 57638 5054 57690
rect 5054 57638 5066 57690
rect 5066 57638 5096 57690
rect 5120 57638 5130 57690
rect 5130 57638 5176 57690
rect 4880 57636 4936 57638
rect 4960 57636 5016 57638
rect 5040 57636 5096 57638
rect 5120 57636 5176 57638
rect 1306 57160 1362 57216
rect 4220 57146 4276 57148
rect 4300 57146 4356 57148
rect 4380 57146 4436 57148
rect 4460 57146 4516 57148
rect 4220 57094 4266 57146
rect 4266 57094 4276 57146
rect 4300 57094 4330 57146
rect 4330 57094 4342 57146
rect 4342 57094 4356 57146
rect 4380 57094 4394 57146
rect 4394 57094 4406 57146
rect 4406 57094 4436 57146
rect 4460 57094 4470 57146
rect 4470 57094 4516 57146
rect 4220 57092 4276 57094
rect 4300 57092 4356 57094
rect 4380 57092 4436 57094
rect 4460 57092 4516 57094
rect 4880 56602 4936 56604
rect 4960 56602 5016 56604
rect 5040 56602 5096 56604
rect 5120 56602 5176 56604
rect 4880 56550 4926 56602
rect 4926 56550 4936 56602
rect 4960 56550 4990 56602
rect 4990 56550 5002 56602
rect 5002 56550 5016 56602
rect 5040 56550 5054 56602
rect 5054 56550 5066 56602
rect 5066 56550 5096 56602
rect 5120 56550 5130 56602
rect 5130 56550 5176 56602
rect 4880 56548 4936 56550
rect 4960 56548 5016 56550
rect 5040 56548 5096 56550
rect 5120 56548 5176 56550
rect 4220 56058 4276 56060
rect 4300 56058 4356 56060
rect 4380 56058 4436 56060
rect 4460 56058 4516 56060
rect 4220 56006 4266 56058
rect 4266 56006 4276 56058
rect 4300 56006 4330 56058
rect 4330 56006 4342 56058
rect 4342 56006 4356 56058
rect 4380 56006 4394 56058
rect 4394 56006 4406 56058
rect 4406 56006 4436 56058
rect 4460 56006 4470 56058
rect 4470 56006 4516 56058
rect 4220 56004 4276 56006
rect 4300 56004 4356 56006
rect 4380 56004 4436 56006
rect 4460 56004 4516 56006
rect 1306 55800 1362 55856
rect 4880 55514 4936 55516
rect 4960 55514 5016 55516
rect 5040 55514 5096 55516
rect 5120 55514 5176 55516
rect 4880 55462 4926 55514
rect 4926 55462 4936 55514
rect 4960 55462 4990 55514
rect 4990 55462 5002 55514
rect 5002 55462 5016 55514
rect 5040 55462 5054 55514
rect 5054 55462 5066 55514
rect 5066 55462 5096 55514
rect 5120 55462 5130 55514
rect 5130 55462 5176 55514
rect 4880 55460 4936 55462
rect 4960 55460 5016 55462
rect 5040 55460 5096 55462
rect 5120 55460 5176 55462
rect 4220 54970 4276 54972
rect 4300 54970 4356 54972
rect 4380 54970 4436 54972
rect 4460 54970 4516 54972
rect 4220 54918 4266 54970
rect 4266 54918 4276 54970
rect 4300 54918 4330 54970
rect 4330 54918 4342 54970
rect 4342 54918 4356 54970
rect 4380 54918 4394 54970
rect 4394 54918 4406 54970
rect 4406 54918 4436 54970
rect 4460 54918 4470 54970
rect 4470 54918 4516 54970
rect 4220 54916 4276 54918
rect 4300 54916 4356 54918
rect 4380 54916 4436 54918
rect 4460 54916 4516 54918
rect 1306 54440 1362 54496
rect 4880 54426 4936 54428
rect 4960 54426 5016 54428
rect 5040 54426 5096 54428
rect 5120 54426 5176 54428
rect 4880 54374 4926 54426
rect 4926 54374 4936 54426
rect 4960 54374 4990 54426
rect 4990 54374 5002 54426
rect 5002 54374 5016 54426
rect 5040 54374 5054 54426
rect 5054 54374 5066 54426
rect 5066 54374 5096 54426
rect 5120 54374 5130 54426
rect 5130 54374 5176 54426
rect 4880 54372 4936 54374
rect 4960 54372 5016 54374
rect 5040 54372 5096 54374
rect 5120 54372 5176 54374
rect 1214 53760 1270 53816
rect 4220 53882 4276 53884
rect 4300 53882 4356 53884
rect 4380 53882 4436 53884
rect 4460 53882 4516 53884
rect 4220 53830 4266 53882
rect 4266 53830 4276 53882
rect 4300 53830 4330 53882
rect 4330 53830 4342 53882
rect 4342 53830 4356 53882
rect 4380 53830 4394 53882
rect 4394 53830 4406 53882
rect 4406 53830 4436 53882
rect 4460 53830 4470 53882
rect 4470 53830 4516 53882
rect 4220 53828 4276 53830
rect 4300 53828 4356 53830
rect 4380 53828 4436 53830
rect 4460 53828 4516 53830
rect 1582 53624 1638 53680
rect 4880 53338 4936 53340
rect 4960 53338 5016 53340
rect 5040 53338 5096 53340
rect 5120 53338 5176 53340
rect 4880 53286 4926 53338
rect 4926 53286 4936 53338
rect 4960 53286 4990 53338
rect 4990 53286 5002 53338
rect 5002 53286 5016 53338
rect 5040 53286 5054 53338
rect 5054 53286 5066 53338
rect 5066 53286 5096 53338
rect 5120 53286 5130 53338
rect 5130 53286 5176 53338
rect 4880 53284 4936 53286
rect 4960 53284 5016 53286
rect 5040 53284 5096 53286
rect 5120 53284 5176 53286
rect 4220 52794 4276 52796
rect 4300 52794 4356 52796
rect 4380 52794 4436 52796
rect 4460 52794 4516 52796
rect 4220 52742 4266 52794
rect 4266 52742 4276 52794
rect 4300 52742 4330 52794
rect 4330 52742 4342 52794
rect 4342 52742 4356 52794
rect 4380 52742 4394 52794
rect 4394 52742 4406 52794
rect 4406 52742 4436 52794
rect 4460 52742 4470 52794
rect 4470 52742 4516 52794
rect 4220 52740 4276 52742
rect 4300 52740 4356 52742
rect 4380 52740 4436 52742
rect 4460 52740 4516 52742
rect 4880 52250 4936 52252
rect 4960 52250 5016 52252
rect 5040 52250 5096 52252
rect 5120 52250 5176 52252
rect 4880 52198 4926 52250
rect 4926 52198 4936 52250
rect 4960 52198 4990 52250
rect 4990 52198 5002 52250
rect 5002 52198 5016 52250
rect 5040 52198 5054 52250
rect 5054 52198 5066 52250
rect 5066 52198 5096 52250
rect 5120 52198 5130 52250
rect 5130 52198 5176 52250
rect 4880 52196 4936 52198
rect 4960 52196 5016 52198
rect 5040 52196 5096 52198
rect 5120 52196 5176 52198
rect 4220 51706 4276 51708
rect 4300 51706 4356 51708
rect 4380 51706 4436 51708
rect 4460 51706 4516 51708
rect 4220 51654 4266 51706
rect 4266 51654 4276 51706
rect 4300 51654 4330 51706
rect 4330 51654 4342 51706
rect 4342 51654 4356 51706
rect 4380 51654 4394 51706
rect 4394 51654 4406 51706
rect 4406 51654 4436 51706
rect 4460 51654 4470 51706
rect 4470 51654 4516 51706
rect 4220 51652 4276 51654
rect 4300 51652 4356 51654
rect 4380 51652 4436 51654
rect 4460 51652 4516 51654
rect 4880 51162 4936 51164
rect 4960 51162 5016 51164
rect 5040 51162 5096 51164
rect 5120 51162 5176 51164
rect 4880 51110 4926 51162
rect 4926 51110 4936 51162
rect 4960 51110 4990 51162
rect 4990 51110 5002 51162
rect 5002 51110 5016 51162
rect 5040 51110 5054 51162
rect 5054 51110 5066 51162
rect 5066 51110 5096 51162
rect 5120 51110 5130 51162
rect 5130 51110 5176 51162
rect 4880 51108 4936 51110
rect 4960 51108 5016 51110
rect 5040 51108 5096 51110
rect 5120 51108 5176 51110
rect 4220 50618 4276 50620
rect 4300 50618 4356 50620
rect 4380 50618 4436 50620
rect 4460 50618 4516 50620
rect 4220 50566 4266 50618
rect 4266 50566 4276 50618
rect 4300 50566 4330 50618
rect 4330 50566 4342 50618
rect 4342 50566 4356 50618
rect 4380 50566 4394 50618
rect 4394 50566 4406 50618
rect 4406 50566 4436 50618
rect 4460 50566 4470 50618
rect 4470 50566 4516 50618
rect 4220 50564 4276 50566
rect 4300 50564 4356 50566
rect 4380 50564 4436 50566
rect 4460 50564 4516 50566
rect 4880 50074 4936 50076
rect 4960 50074 5016 50076
rect 5040 50074 5096 50076
rect 5120 50074 5176 50076
rect 4880 50022 4926 50074
rect 4926 50022 4936 50074
rect 4960 50022 4990 50074
rect 4990 50022 5002 50074
rect 5002 50022 5016 50074
rect 5040 50022 5054 50074
rect 5054 50022 5066 50074
rect 5066 50022 5096 50074
rect 5120 50022 5130 50074
rect 5130 50022 5176 50074
rect 4880 50020 4936 50022
rect 4960 50020 5016 50022
rect 5040 50020 5096 50022
rect 5120 50020 5176 50022
rect 4220 49530 4276 49532
rect 4300 49530 4356 49532
rect 4380 49530 4436 49532
rect 4460 49530 4516 49532
rect 4220 49478 4266 49530
rect 4266 49478 4276 49530
rect 4300 49478 4330 49530
rect 4330 49478 4342 49530
rect 4342 49478 4356 49530
rect 4380 49478 4394 49530
rect 4394 49478 4406 49530
rect 4406 49478 4436 49530
rect 4460 49478 4470 49530
rect 4470 49478 4516 49530
rect 4220 49476 4276 49478
rect 4300 49476 4356 49478
rect 4380 49476 4436 49478
rect 4460 49476 4516 49478
rect 4880 48986 4936 48988
rect 4960 48986 5016 48988
rect 5040 48986 5096 48988
rect 5120 48986 5176 48988
rect 4880 48934 4926 48986
rect 4926 48934 4936 48986
rect 4960 48934 4990 48986
rect 4990 48934 5002 48986
rect 5002 48934 5016 48986
rect 5040 48934 5054 48986
rect 5054 48934 5066 48986
rect 5066 48934 5096 48986
rect 5120 48934 5130 48986
rect 5130 48934 5176 48986
rect 4880 48932 4936 48934
rect 4960 48932 5016 48934
rect 5040 48932 5096 48934
rect 5120 48932 5176 48934
rect 35600 95770 35656 95772
rect 35680 95770 35736 95772
rect 35760 95770 35816 95772
rect 35840 95770 35896 95772
rect 35600 95718 35646 95770
rect 35646 95718 35656 95770
rect 35680 95718 35710 95770
rect 35710 95718 35722 95770
rect 35722 95718 35736 95770
rect 35760 95718 35774 95770
rect 35774 95718 35786 95770
rect 35786 95718 35816 95770
rect 35840 95718 35850 95770
rect 35850 95718 35896 95770
rect 35600 95716 35656 95718
rect 35680 95716 35736 95718
rect 35760 95716 35816 95718
rect 35840 95716 35896 95718
rect 34940 95226 34996 95228
rect 35020 95226 35076 95228
rect 35100 95226 35156 95228
rect 35180 95226 35236 95228
rect 34940 95174 34986 95226
rect 34986 95174 34996 95226
rect 35020 95174 35050 95226
rect 35050 95174 35062 95226
rect 35062 95174 35076 95226
rect 35100 95174 35114 95226
rect 35114 95174 35126 95226
rect 35126 95174 35156 95226
rect 35180 95174 35190 95226
rect 35190 95174 35236 95226
rect 34940 95172 34996 95174
rect 35020 95172 35076 95174
rect 35100 95172 35156 95174
rect 35180 95172 35236 95174
rect 34940 94138 34996 94140
rect 35020 94138 35076 94140
rect 35100 94138 35156 94140
rect 35180 94138 35236 94140
rect 34940 94086 34986 94138
rect 34986 94086 34996 94138
rect 35020 94086 35050 94138
rect 35050 94086 35062 94138
rect 35062 94086 35076 94138
rect 35100 94086 35114 94138
rect 35114 94086 35126 94138
rect 35126 94086 35156 94138
rect 35180 94086 35190 94138
rect 35190 94086 35236 94138
rect 34940 94084 34996 94086
rect 35020 94084 35076 94086
rect 35100 94084 35156 94086
rect 35180 94084 35236 94086
rect 34940 93050 34996 93052
rect 35020 93050 35076 93052
rect 35100 93050 35156 93052
rect 35180 93050 35236 93052
rect 34940 92998 34986 93050
rect 34986 92998 34996 93050
rect 35020 92998 35050 93050
rect 35050 92998 35062 93050
rect 35062 92998 35076 93050
rect 35100 92998 35114 93050
rect 35114 92998 35126 93050
rect 35126 92998 35156 93050
rect 35180 92998 35190 93050
rect 35190 92998 35236 93050
rect 34940 92996 34996 92998
rect 35020 92996 35076 92998
rect 35100 92996 35156 92998
rect 35180 92996 35236 92998
rect 35600 94682 35656 94684
rect 35680 94682 35736 94684
rect 35760 94682 35816 94684
rect 35840 94682 35896 94684
rect 35600 94630 35646 94682
rect 35646 94630 35656 94682
rect 35680 94630 35710 94682
rect 35710 94630 35722 94682
rect 35722 94630 35736 94682
rect 35760 94630 35774 94682
rect 35774 94630 35786 94682
rect 35786 94630 35816 94682
rect 35840 94630 35850 94682
rect 35850 94630 35896 94682
rect 35600 94628 35656 94630
rect 35680 94628 35736 94630
rect 35760 94628 35816 94630
rect 35840 94628 35896 94630
rect 35600 93594 35656 93596
rect 35680 93594 35736 93596
rect 35760 93594 35816 93596
rect 35840 93594 35896 93596
rect 35600 93542 35646 93594
rect 35646 93542 35656 93594
rect 35680 93542 35710 93594
rect 35710 93542 35722 93594
rect 35722 93542 35736 93594
rect 35760 93542 35774 93594
rect 35774 93542 35786 93594
rect 35786 93542 35816 93594
rect 35840 93542 35850 93594
rect 35850 93542 35896 93594
rect 35600 93540 35656 93542
rect 35680 93540 35736 93542
rect 35760 93540 35816 93542
rect 35840 93540 35896 93542
rect 66320 95770 66376 95772
rect 66400 95770 66456 95772
rect 66480 95770 66536 95772
rect 66560 95770 66616 95772
rect 66320 95718 66366 95770
rect 66366 95718 66376 95770
rect 66400 95718 66430 95770
rect 66430 95718 66442 95770
rect 66442 95718 66456 95770
rect 66480 95718 66494 95770
rect 66494 95718 66506 95770
rect 66506 95718 66536 95770
rect 66560 95718 66570 95770
rect 66570 95718 66616 95770
rect 66320 95716 66376 95718
rect 66400 95716 66456 95718
rect 66480 95716 66536 95718
rect 66560 95716 66616 95718
rect 97040 95770 97096 95772
rect 97120 95770 97176 95772
rect 97200 95770 97256 95772
rect 97280 95770 97336 95772
rect 97040 95718 97086 95770
rect 97086 95718 97096 95770
rect 97120 95718 97150 95770
rect 97150 95718 97162 95770
rect 97162 95718 97176 95770
rect 97200 95718 97214 95770
rect 97214 95718 97226 95770
rect 97226 95718 97256 95770
rect 97280 95718 97290 95770
rect 97290 95718 97336 95770
rect 97040 95716 97096 95718
rect 97120 95716 97176 95718
rect 97200 95716 97256 95718
rect 97280 95716 97336 95718
rect 13266 90480 13322 90536
rect 8298 87488 8354 87544
rect 8298 86672 8354 86728
rect 8298 85312 8354 85368
rect 8298 83408 8354 83464
rect 8298 82048 8354 82104
rect 8298 81232 8354 81288
rect 8298 79872 8354 79928
rect 8298 79056 8354 79112
rect 8298 77968 8354 78024
rect 8298 76608 8354 76664
rect 8298 74432 8354 74488
rect 8298 73616 8354 73672
rect 8298 72528 8354 72584
rect 8298 71168 8354 71224
rect 8298 68584 8354 68640
rect 8298 68040 8354 68096
rect 8298 66952 8354 67008
rect 8298 65728 8354 65784
rect 8298 63144 8354 63200
rect 8298 62600 8354 62656
rect 8298 61512 8354 61568
rect 8298 60308 8354 60344
rect 8298 60288 8300 60308
rect 8300 60288 8352 60308
rect 8352 60288 8354 60308
rect 8298 57160 8354 57216
rect 8298 56072 8354 56128
rect 8298 54868 8354 54904
rect 8298 54848 8300 54868
rect 8300 54848 8352 54868
rect 8352 54848 8354 54868
rect 4220 48442 4276 48444
rect 4300 48442 4356 48444
rect 4380 48442 4436 48444
rect 4460 48442 4516 48444
rect 4220 48390 4266 48442
rect 4266 48390 4276 48442
rect 4300 48390 4330 48442
rect 4330 48390 4342 48442
rect 4342 48390 4356 48442
rect 4380 48390 4394 48442
rect 4394 48390 4406 48442
rect 4406 48390 4436 48442
rect 4460 48390 4470 48442
rect 4470 48390 4516 48442
rect 4220 48388 4276 48390
rect 4300 48388 4356 48390
rect 4380 48388 4436 48390
rect 4460 48388 4516 48390
rect 1214 48320 1270 48376
rect 4880 47898 4936 47900
rect 4960 47898 5016 47900
rect 5040 47898 5096 47900
rect 5120 47898 5176 47900
rect 4880 47846 4926 47898
rect 4926 47846 4936 47898
rect 4960 47846 4990 47898
rect 4990 47846 5002 47898
rect 5002 47846 5016 47898
rect 5040 47846 5054 47898
rect 5054 47846 5066 47898
rect 5066 47846 5096 47898
rect 5120 47846 5130 47898
rect 5130 47846 5176 47898
rect 4880 47844 4936 47846
rect 4960 47844 5016 47846
rect 5040 47844 5096 47846
rect 5120 47844 5176 47846
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 4880 46810 4936 46812
rect 4960 46810 5016 46812
rect 5040 46810 5096 46812
rect 5120 46810 5176 46812
rect 4880 46758 4926 46810
rect 4926 46758 4936 46810
rect 4960 46758 4990 46810
rect 4990 46758 5002 46810
rect 5002 46758 5016 46810
rect 5040 46758 5054 46810
rect 5054 46758 5066 46810
rect 5066 46758 5096 46810
rect 5120 46758 5130 46810
rect 5130 46758 5176 46810
rect 4880 46756 4936 46758
rect 4960 46756 5016 46758
rect 5040 46756 5096 46758
rect 5120 46756 5176 46758
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 846 45772 848 45792
rect 848 45772 900 45792
rect 900 45772 902 45792
rect 846 45736 902 45772
rect 4880 45722 4936 45724
rect 4960 45722 5016 45724
rect 5040 45722 5096 45724
rect 5120 45722 5176 45724
rect 4880 45670 4926 45722
rect 4926 45670 4936 45722
rect 4960 45670 4990 45722
rect 4990 45670 5002 45722
rect 5002 45670 5016 45722
rect 5040 45670 5054 45722
rect 5054 45670 5066 45722
rect 5066 45670 5096 45722
rect 5120 45670 5130 45722
rect 5130 45670 5176 45722
rect 4880 45668 4936 45670
rect 4960 45668 5016 45670
rect 5040 45668 5096 45670
rect 5120 45668 5176 45670
rect 1674 45328 1730 45384
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4880 44634 4936 44636
rect 4960 44634 5016 44636
rect 5040 44634 5096 44636
rect 5120 44634 5176 44636
rect 4880 44582 4926 44634
rect 4926 44582 4936 44634
rect 4960 44582 4990 44634
rect 4990 44582 5002 44634
rect 5002 44582 5016 44634
rect 5040 44582 5054 44634
rect 5054 44582 5066 44634
rect 5066 44582 5096 44634
rect 5120 44582 5130 44634
rect 5130 44582 5176 44634
rect 4880 44580 4936 44582
rect 4960 44580 5016 44582
rect 5040 44580 5096 44582
rect 5120 44580 5176 44582
rect 846 44376 902 44432
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4880 43546 4936 43548
rect 4960 43546 5016 43548
rect 5040 43546 5096 43548
rect 5120 43546 5176 43548
rect 4880 43494 4926 43546
rect 4926 43494 4936 43546
rect 4960 43494 4990 43546
rect 4990 43494 5002 43546
rect 5002 43494 5016 43546
rect 5040 43494 5054 43546
rect 5054 43494 5066 43546
rect 5066 43494 5096 43546
rect 5120 43494 5130 43546
rect 5130 43494 5176 43546
rect 4880 43492 4936 43494
rect 4960 43492 5016 43494
rect 5040 43492 5096 43494
rect 5120 43492 5176 43494
rect 846 43052 848 43072
rect 848 43052 900 43072
rect 900 43052 902 43072
rect 846 43016 902 43052
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4880 42458 4936 42460
rect 4960 42458 5016 42460
rect 5040 42458 5096 42460
rect 5120 42458 5176 42460
rect 4880 42406 4926 42458
rect 4926 42406 4936 42458
rect 4960 42406 4990 42458
rect 4990 42406 5002 42458
rect 5002 42406 5016 42458
rect 5040 42406 5054 42458
rect 5054 42406 5066 42458
rect 5066 42406 5096 42458
rect 5120 42406 5130 42458
rect 5130 42406 5176 42458
rect 4880 42404 4936 42406
rect 4960 42404 5016 42406
rect 5040 42404 5096 42406
rect 5120 42404 5176 42406
rect 846 42336 902 42392
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4880 41370 4936 41372
rect 4960 41370 5016 41372
rect 5040 41370 5096 41372
rect 5120 41370 5176 41372
rect 4880 41318 4926 41370
rect 4926 41318 4936 41370
rect 4960 41318 4990 41370
rect 4990 41318 5002 41370
rect 5002 41318 5016 41370
rect 5040 41318 5054 41370
rect 5054 41318 5066 41370
rect 5066 41318 5096 41370
rect 5120 41318 5130 41370
rect 5130 41318 5176 41370
rect 4880 41316 4936 41318
rect 4960 41316 5016 41318
rect 5040 41316 5096 41318
rect 5120 41316 5176 41318
rect 846 40996 902 41032
rect 846 40976 848 40996
rect 848 40976 900 40996
rect 900 40976 902 40996
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 846 40332 848 40352
rect 848 40332 900 40352
rect 900 40332 902 40352
rect 846 40296 902 40332
rect 4880 40282 4936 40284
rect 4960 40282 5016 40284
rect 5040 40282 5096 40284
rect 5120 40282 5176 40284
rect 4880 40230 4926 40282
rect 4926 40230 4936 40282
rect 4960 40230 4990 40282
rect 4990 40230 5002 40282
rect 5002 40230 5016 40282
rect 5040 40230 5054 40282
rect 5054 40230 5066 40282
rect 5066 40230 5096 40282
rect 5120 40230 5130 40282
rect 5130 40230 5176 40282
rect 4880 40228 4936 40230
rect 4960 40228 5016 40230
rect 5040 40228 5096 40230
rect 5120 40228 5176 40230
rect 1674 39888 1730 39944
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4880 39194 4936 39196
rect 4960 39194 5016 39196
rect 5040 39194 5096 39196
rect 5120 39194 5176 39196
rect 4880 39142 4926 39194
rect 4926 39142 4936 39194
rect 4960 39142 4990 39194
rect 4990 39142 5002 39194
rect 5002 39142 5016 39194
rect 5040 39142 5054 39194
rect 5054 39142 5066 39194
rect 5066 39142 5096 39194
rect 5120 39142 5130 39194
rect 5130 39142 5176 39194
rect 4880 39140 4936 39142
rect 4960 39140 5016 39142
rect 5040 39140 5096 39142
rect 5120 39140 5176 39142
rect 846 38700 848 38720
rect 848 38700 900 38720
rect 900 38700 902 38720
rect 846 38664 902 38700
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4880 38106 4936 38108
rect 4960 38106 5016 38108
rect 5040 38106 5096 38108
rect 5120 38106 5176 38108
rect 4880 38054 4926 38106
rect 4926 38054 4936 38106
rect 4960 38054 4990 38106
rect 4990 38054 5002 38106
rect 5002 38054 5016 38106
rect 5040 38054 5054 38106
rect 5054 38054 5066 38106
rect 5066 38054 5096 38106
rect 5120 38054 5130 38106
rect 5130 38054 5176 38106
rect 4880 38052 4936 38054
rect 4960 38052 5016 38054
rect 5040 38052 5096 38054
rect 5120 38052 5176 38054
rect 846 37612 848 37632
rect 848 37612 900 37632
rect 900 37612 902 37632
rect 846 37576 902 37612
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4880 37018 4936 37020
rect 4960 37018 5016 37020
rect 5040 37018 5096 37020
rect 5120 37018 5176 37020
rect 4880 36966 4926 37018
rect 4926 36966 4936 37018
rect 4960 36966 4990 37018
rect 4990 36966 5002 37018
rect 5002 36966 5016 37018
rect 5040 36966 5054 37018
rect 5054 36966 5066 37018
rect 5066 36966 5096 37018
rect 5120 36966 5130 37018
rect 5130 36966 5176 37018
rect 4880 36964 4936 36966
rect 4960 36964 5016 36966
rect 5040 36964 5096 36966
rect 5120 36964 5176 36966
rect 846 36896 902 36952
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4880 35930 4936 35932
rect 4960 35930 5016 35932
rect 5040 35930 5096 35932
rect 5120 35930 5176 35932
rect 4880 35878 4926 35930
rect 4926 35878 4936 35930
rect 4960 35878 4990 35930
rect 4990 35878 5002 35930
rect 5002 35878 5016 35930
rect 5040 35878 5054 35930
rect 5054 35878 5066 35930
rect 5066 35878 5096 35930
rect 5120 35878 5130 35930
rect 5130 35878 5176 35930
rect 4880 35876 4936 35878
rect 4960 35876 5016 35878
rect 5040 35876 5096 35878
rect 5120 35876 5176 35878
rect 846 35556 902 35592
rect 846 35536 848 35556
rect 848 35536 900 35556
rect 900 35536 902 35556
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 846 34892 848 34912
rect 848 34892 900 34912
rect 900 34892 902 34912
rect 846 34856 902 34892
rect 4880 34842 4936 34844
rect 4960 34842 5016 34844
rect 5040 34842 5096 34844
rect 5120 34842 5176 34844
rect 4880 34790 4926 34842
rect 4926 34790 4936 34842
rect 4960 34790 4990 34842
rect 4990 34790 5002 34842
rect 5002 34790 5016 34842
rect 5040 34790 5054 34842
rect 5054 34790 5066 34842
rect 5066 34790 5096 34842
rect 5120 34790 5130 34842
rect 5130 34790 5176 34842
rect 4880 34788 4936 34790
rect 4960 34788 5016 34790
rect 5040 34788 5096 34790
rect 5120 34788 5176 34790
rect 1674 34448 1730 34504
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4880 33754 4936 33756
rect 4960 33754 5016 33756
rect 5040 33754 5096 33756
rect 5120 33754 5176 33756
rect 4880 33702 4926 33754
rect 4926 33702 4936 33754
rect 4960 33702 4990 33754
rect 4990 33702 5002 33754
rect 5002 33702 5016 33754
rect 5040 33702 5054 33754
rect 5054 33702 5066 33754
rect 5066 33702 5096 33754
rect 5120 33702 5130 33754
rect 5130 33702 5176 33754
rect 4880 33700 4936 33702
rect 4960 33700 5016 33702
rect 5040 33700 5096 33702
rect 5120 33700 5176 33702
rect 846 33260 848 33280
rect 848 33260 900 33280
rect 900 33260 902 33280
rect 846 33224 902 33260
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4880 32666 4936 32668
rect 4960 32666 5016 32668
rect 5040 32666 5096 32668
rect 5120 32666 5176 32668
rect 4880 32614 4926 32666
rect 4926 32614 4936 32666
rect 4960 32614 4990 32666
rect 4990 32614 5002 32666
rect 5002 32614 5016 32666
rect 5040 32614 5054 32666
rect 5054 32614 5066 32666
rect 5066 32614 5096 32666
rect 5120 32614 5130 32666
rect 5130 32614 5176 32666
rect 4880 32612 4936 32614
rect 4960 32612 5016 32614
rect 5040 32612 5096 32614
rect 5120 32612 5176 32614
rect 846 32172 848 32192
rect 848 32172 900 32192
rect 900 32172 902 32192
rect 846 32136 902 32172
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 846 31456 902 31512
rect 4880 31578 4936 31580
rect 4960 31578 5016 31580
rect 5040 31578 5096 31580
rect 5120 31578 5176 31580
rect 4880 31526 4926 31578
rect 4926 31526 4936 31578
rect 4960 31526 4990 31578
rect 4990 31526 5002 31578
rect 5002 31526 5016 31578
rect 5040 31526 5054 31578
rect 5054 31526 5066 31578
rect 5066 31526 5096 31578
rect 5120 31526 5130 31578
rect 5130 31526 5176 31578
rect 4880 31524 4936 31526
rect 4960 31524 5016 31526
rect 5040 31524 5096 31526
rect 5120 31524 5176 31526
rect 1674 31184 1730 31240
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4880 30490 4936 30492
rect 4960 30490 5016 30492
rect 5040 30490 5096 30492
rect 5120 30490 5176 30492
rect 4880 30438 4926 30490
rect 4926 30438 4936 30490
rect 4960 30438 4990 30490
rect 4990 30438 5002 30490
rect 5002 30438 5016 30490
rect 5040 30438 5054 30490
rect 5054 30438 5066 30490
rect 5066 30438 5096 30490
rect 5120 30438 5130 30490
rect 5130 30438 5176 30490
rect 4880 30436 4936 30438
rect 4960 30436 5016 30438
rect 5040 30436 5096 30438
rect 5120 30436 5176 30438
rect 846 30116 902 30152
rect 846 30096 848 30116
rect 848 30096 900 30116
rect 900 30096 902 30116
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 846 29452 848 29472
rect 848 29452 900 29472
rect 900 29452 902 29472
rect 846 29416 902 29452
rect 4880 29402 4936 29404
rect 4960 29402 5016 29404
rect 5040 29402 5096 29404
rect 5120 29402 5176 29404
rect 4880 29350 4926 29402
rect 4926 29350 4936 29402
rect 4960 29350 4990 29402
rect 4990 29350 5002 29402
rect 5002 29350 5016 29402
rect 5040 29350 5054 29402
rect 5054 29350 5066 29402
rect 5066 29350 5096 29402
rect 5120 29350 5130 29402
rect 5130 29350 5176 29402
rect 4880 29348 4936 29350
rect 4960 29348 5016 29350
rect 5040 29348 5096 29350
rect 5120 29348 5176 29350
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4880 28314 4936 28316
rect 4960 28314 5016 28316
rect 5040 28314 5096 28316
rect 5120 28314 5176 28316
rect 4880 28262 4926 28314
rect 4926 28262 4936 28314
rect 4960 28262 4990 28314
rect 4990 28262 5002 28314
rect 5002 28262 5016 28314
rect 5040 28262 5054 28314
rect 5054 28262 5066 28314
rect 5066 28262 5096 28314
rect 5120 28262 5130 28314
rect 5130 28262 5176 28314
rect 4880 28260 4936 28262
rect 4960 28260 5016 28262
rect 5040 28260 5096 28262
rect 5120 28260 5176 28262
rect 1306 27920 1362 27976
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4880 27226 4936 27228
rect 4960 27226 5016 27228
rect 5040 27226 5096 27228
rect 5120 27226 5176 27228
rect 4880 27174 4926 27226
rect 4926 27174 4936 27226
rect 4960 27174 4990 27226
rect 4990 27174 5002 27226
rect 5002 27174 5016 27226
rect 5040 27174 5054 27226
rect 5054 27174 5066 27226
rect 5066 27174 5096 27226
rect 5120 27174 5130 27226
rect 5130 27174 5176 27226
rect 4880 27172 4936 27174
rect 4960 27172 5016 27174
rect 5040 27172 5096 27174
rect 5120 27172 5176 27174
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 1306 26560 1362 26616
rect 1306 25880 1362 25936
rect 4880 26138 4936 26140
rect 4960 26138 5016 26140
rect 5040 26138 5096 26140
rect 5120 26138 5176 26140
rect 4880 26086 4926 26138
rect 4926 26086 4936 26138
rect 4960 26086 4990 26138
rect 4990 26086 5002 26138
rect 5002 26086 5016 26138
rect 5040 26086 5054 26138
rect 5054 26086 5066 26138
rect 5066 26086 5096 26138
rect 5120 26086 5130 26138
rect 5130 26086 5176 26138
rect 4880 26084 4936 26086
rect 4960 26084 5016 26086
rect 5040 26084 5096 26086
rect 5120 26084 5176 26086
rect 1674 25744 1730 25800
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4880 25050 4936 25052
rect 4960 25050 5016 25052
rect 5040 25050 5096 25052
rect 5120 25050 5176 25052
rect 4880 24998 4926 25050
rect 4926 24998 4936 25050
rect 4960 24998 4990 25050
rect 4990 24998 5002 25050
rect 5002 24998 5016 25050
rect 5040 24998 5054 25050
rect 5054 24998 5066 25050
rect 5066 24998 5096 25050
rect 5120 24998 5130 25050
rect 5130 24998 5176 25050
rect 4880 24996 4936 24998
rect 4960 24996 5016 24998
rect 5040 24996 5096 24998
rect 5120 24996 5176 24998
rect 1306 24520 1362 24576
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4880 23962 4936 23964
rect 4960 23962 5016 23964
rect 5040 23962 5096 23964
rect 5120 23962 5176 23964
rect 4880 23910 4926 23962
rect 4926 23910 4936 23962
rect 4960 23910 4990 23962
rect 4990 23910 5002 23962
rect 5002 23910 5016 23962
rect 5040 23910 5054 23962
rect 5054 23910 5066 23962
rect 5066 23910 5096 23962
rect 5120 23910 5130 23962
rect 5130 23910 5176 23962
rect 4880 23908 4936 23910
rect 4960 23908 5016 23910
rect 5040 23908 5096 23910
rect 5120 23908 5176 23910
rect 1306 23840 1362 23896
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4880 22874 4936 22876
rect 4960 22874 5016 22876
rect 5040 22874 5096 22876
rect 5120 22874 5176 22876
rect 4880 22822 4926 22874
rect 4926 22822 4936 22874
rect 4960 22822 4990 22874
rect 4990 22822 5002 22874
rect 5002 22822 5016 22874
rect 5040 22822 5054 22874
rect 5054 22822 5066 22874
rect 5066 22822 5096 22874
rect 5120 22822 5130 22874
rect 5130 22822 5176 22874
rect 4880 22820 4936 22822
rect 4960 22820 5016 22822
rect 5040 22820 5096 22822
rect 5120 22820 5176 22822
rect 1122 22480 1178 22536
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4880 21786 4936 21788
rect 4960 21786 5016 21788
rect 5040 21786 5096 21788
rect 5120 21786 5176 21788
rect 4880 21734 4926 21786
rect 4926 21734 4936 21786
rect 4960 21734 4990 21786
rect 4990 21734 5002 21786
rect 5002 21734 5016 21786
rect 5040 21734 5054 21786
rect 5054 21734 5066 21786
rect 5066 21734 5096 21786
rect 5120 21734 5130 21786
rect 5130 21734 5176 21786
rect 4880 21732 4936 21734
rect 4960 21732 5016 21734
rect 5040 21732 5096 21734
rect 5120 21732 5176 21734
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 1306 21120 1362 21176
rect 1306 20440 1362 20496
rect 4880 20698 4936 20700
rect 4960 20698 5016 20700
rect 5040 20698 5096 20700
rect 5120 20698 5176 20700
rect 4880 20646 4926 20698
rect 4926 20646 4936 20698
rect 4960 20646 4990 20698
rect 4990 20646 5002 20698
rect 5002 20646 5016 20698
rect 5040 20646 5054 20698
rect 5054 20646 5066 20698
rect 5066 20646 5096 20698
rect 5120 20646 5130 20698
rect 5130 20646 5176 20698
rect 4880 20644 4936 20646
rect 4960 20644 5016 20646
rect 5040 20644 5096 20646
rect 5120 20644 5176 20646
rect 1858 20304 1914 20360
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4880 19610 4936 19612
rect 4960 19610 5016 19612
rect 5040 19610 5096 19612
rect 5120 19610 5176 19612
rect 4880 19558 4926 19610
rect 4926 19558 4936 19610
rect 4960 19558 4990 19610
rect 4990 19558 5002 19610
rect 5002 19558 5016 19610
rect 5040 19558 5054 19610
rect 5054 19558 5066 19610
rect 5066 19558 5096 19610
rect 5120 19558 5130 19610
rect 5130 19558 5176 19610
rect 4880 19556 4936 19558
rect 4960 19556 5016 19558
rect 5040 19556 5096 19558
rect 5120 19556 5176 19558
rect 1490 19080 1546 19136
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4880 18522 4936 18524
rect 4960 18522 5016 18524
rect 5040 18522 5096 18524
rect 5120 18522 5176 18524
rect 4880 18470 4926 18522
rect 4926 18470 4936 18522
rect 4960 18470 4990 18522
rect 4990 18470 5002 18522
rect 5002 18470 5016 18522
rect 5040 18470 5054 18522
rect 5054 18470 5066 18522
rect 5066 18470 5096 18522
rect 5120 18470 5130 18522
rect 5130 18470 5176 18522
rect 4880 18468 4936 18470
rect 4960 18468 5016 18470
rect 5040 18468 5096 18470
rect 5120 18468 5176 18470
rect 1306 18400 1362 18456
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4880 17434 4936 17436
rect 4960 17434 5016 17436
rect 5040 17434 5096 17436
rect 5120 17434 5176 17436
rect 4880 17382 4926 17434
rect 4926 17382 4936 17434
rect 4960 17382 4990 17434
rect 4990 17382 5002 17434
rect 5002 17382 5016 17434
rect 5040 17382 5054 17434
rect 5054 17382 5066 17434
rect 5066 17382 5096 17434
rect 5120 17382 5130 17434
rect 5130 17382 5176 17434
rect 4880 17380 4936 17382
rect 4960 17380 5016 17382
rect 5040 17380 5096 17382
rect 5120 17380 5176 17382
rect 1122 17040 1178 17096
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4880 16346 4936 16348
rect 4960 16346 5016 16348
rect 5040 16346 5096 16348
rect 5120 16346 5176 16348
rect 4880 16294 4926 16346
rect 4926 16294 4936 16346
rect 4960 16294 4990 16346
rect 4990 16294 5002 16346
rect 5002 16294 5016 16346
rect 5040 16294 5054 16346
rect 5054 16294 5066 16346
rect 5066 16294 5096 16346
rect 5120 16294 5130 16346
rect 5130 16294 5176 16346
rect 4880 16292 4936 16294
rect 4960 16292 5016 16294
rect 5040 16292 5096 16294
rect 5120 16292 5176 16294
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 1214 15680 1270 15736
rect 1306 15000 1362 15056
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 1858 14864 1914 14920
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 1306 13640 1362 13696
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 1306 12960 1362 13016
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 1122 11600 1178 11656
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 65660 95226 65716 95228
rect 65740 95226 65796 95228
rect 65820 95226 65876 95228
rect 65900 95226 65956 95228
rect 65660 95174 65706 95226
rect 65706 95174 65716 95226
rect 65740 95174 65770 95226
rect 65770 95174 65782 95226
rect 65782 95174 65796 95226
rect 65820 95174 65834 95226
rect 65834 95174 65846 95226
rect 65846 95174 65876 95226
rect 65900 95174 65910 95226
rect 65910 95174 65956 95226
rect 65660 95172 65716 95174
rect 65740 95172 65796 95174
rect 65820 95172 65876 95174
rect 65900 95172 65956 95174
rect 66320 94682 66376 94684
rect 66400 94682 66456 94684
rect 66480 94682 66536 94684
rect 66560 94682 66616 94684
rect 66320 94630 66366 94682
rect 66366 94630 66376 94682
rect 66400 94630 66430 94682
rect 66430 94630 66442 94682
rect 66442 94630 66456 94682
rect 66480 94630 66494 94682
rect 66494 94630 66506 94682
rect 66506 94630 66536 94682
rect 66560 94630 66570 94682
rect 66570 94630 66616 94682
rect 66320 94628 66376 94630
rect 66400 94628 66456 94630
rect 66480 94628 66536 94630
rect 66560 94628 66616 94630
rect 65660 94138 65716 94140
rect 65740 94138 65796 94140
rect 65820 94138 65876 94140
rect 65900 94138 65956 94140
rect 65660 94086 65706 94138
rect 65706 94086 65716 94138
rect 65740 94086 65770 94138
rect 65770 94086 65782 94138
rect 65782 94086 65796 94138
rect 65820 94086 65834 94138
rect 65834 94086 65846 94138
rect 65846 94086 65876 94138
rect 65900 94086 65910 94138
rect 65910 94086 65956 94138
rect 65660 94084 65716 94086
rect 65740 94084 65796 94086
rect 65820 94084 65876 94086
rect 65900 94084 65956 94086
rect 66320 93594 66376 93596
rect 66400 93594 66456 93596
rect 66480 93594 66536 93596
rect 66560 93594 66616 93596
rect 66320 93542 66366 93594
rect 66366 93542 66376 93594
rect 66400 93542 66430 93594
rect 66430 93542 66442 93594
rect 66442 93542 66456 93594
rect 66480 93542 66494 93594
rect 66494 93542 66506 93594
rect 66506 93542 66536 93594
rect 66560 93542 66570 93594
rect 66570 93542 66616 93594
rect 66320 93540 66376 93542
rect 66400 93540 66456 93542
rect 66480 93540 66536 93542
rect 66560 93540 66616 93542
rect 65660 93050 65716 93052
rect 65740 93050 65796 93052
rect 65820 93050 65876 93052
rect 65900 93050 65956 93052
rect 65660 92998 65706 93050
rect 65706 92998 65716 93050
rect 65740 92998 65770 93050
rect 65770 92998 65782 93050
rect 65782 92998 65796 93050
rect 65820 92998 65834 93050
rect 65834 92998 65846 93050
rect 65846 92998 65876 93050
rect 65900 92998 65910 93050
rect 65910 92998 65956 93050
rect 65660 92996 65716 92998
rect 65740 92996 65796 92998
rect 65820 92996 65876 92998
rect 65900 92996 65956 92998
rect 96380 95226 96436 95228
rect 96460 95226 96516 95228
rect 96540 95226 96596 95228
rect 96620 95226 96676 95228
rect 96380 95174 96426 95226
rect 96426 95174 96436 95226
rect 96460 95174 96490 95226
rect 96490 95174 96502 95226
rect 96502 95174 96516 95226
rect 96540 95174 96554 95226
rect 96554 95174 96566 95226
rect 96566 95174 96596 95226
rect 96620 95174 96630 95226
rect 96630 95174 96676 95226
rect 96380 95172 96436 95174
rect 96460 95172 96516 95174
rect 96540 95172 96596 95174
rect 96620 95172 96676 95174
rect 97040 94682 97096 94684
rect 97120 94682 97176 94684
rect 97200 94682 97256 94684
rect 97280 94682 97336 94684
rect 97040 94630 97086 94682
rect 97086 94630 97096 94682
rect 97120 94630 97150 94682
rect 97150 94630 97162 94682
rect 97162 94630 97176 94682
rect 97200 94630 97214 94682
rect 97214 94630 97226 94682
rect 97226 94630 97256 94682
rect 97280 94630 97290 94682
rect 97290 94630 97336 94682
rect 97040 94628 97096 94630
rect 97120 94628 97176 94630
rect 97200 94628 97256 94630
rect 97280 94628 97336 94630
rect 96380 94138 96436 94140
rect 96460 94138 96516 94140
rect 96540 94138 96596 94140
rect 96620 94138 96676 94140
rect 96380 94086 96426 94138
rect 96426 94086 96436 94138
rect 96460 94086 96490 94138
rect 96490 94086 96502 94138
rect 96502 94086 96516 94138
rect 96540 94086 96554 94138
rect 96554 94086 96566 94138
rect 96566 94086 96596 94138
rect 96620 94086 96630 94138
rect 96630 94086 96676 94138
rect 96380 94084 96436 94086
rect 96460 94084 96516 94086
rect 96540 94084 96596 94086
rect 96620 94084 96676 94086
rect 8298 44396 8354 44432
rect 8298 44376 8300 44396
rect 8300 44376 8352 44396
rect 8352 44376 8354 44396
rect 8298 43308 8354 43344
rect 8298 43288 8300 43308
rect 8300 43288 8352 43308
rect 8352 43288 8354 43308
rect 8298 42644 8300 42664
rect 8300 42644 8352 42664
rect 8352 42644 8354 42664
rect 8298 42608 8354 42644
rect 8298 41132 8354 41168
rect 8298 41112 8300 41132
rect 8300 41112 8352 41132
rect 8352 41112 8354 41132
rect 8298 38956 8354 38992
rect 8298 38936 8300 38956
rect 8300 38936 8352 38956
rect 8352 38936 8354 38956
rect 8298 37868 8354 37904
rect 8298 37848 8300 37868
rect 8300 37848 8352 37868
rect 8352 37848 8354 37868
rect 8298 37204 8300 37224
rect 8300 37204 8352 37224
rect 8352 37204 8354 37224
rect 8298 37168 8354 37204
rect 8298 35692 8354 35728
rect 8298 35672 8300 35692
rect 8300 35672 8352 35692
rect 8352 35672 8354 35692
rect 8298 33516 8354 33552
rect 8298 33496 8300 33516
rect 8300 33496 8352 33516
rect 8352 33496 8354 33516
rect 8298 32428 8354 32464
rect 8298 32408 8300 32428
rect 8300 32408 8352 32428
rect 8352 32408 8354 32428
rect 8298 30252 8354 30288
rect 8298 30232 8300 30252
rect 8300 30232 8352 30252
rect 8352 30232 8354 30252
rect 8298 29588 8300 29608
rect 8300 29588 8352 29608
rect 8352 29588 8354 29608
rect 8298 29552 8354 29588
rect 8298 28056 8354 28112
rect 8298 26988 8354 27024
rect 8298 26968 8300 26988
rect 8300 26968 8352 26988
rect 8352 26968 8354 26988
rect 8298 24812 8354 24848
rect 8298 24792 8300 24812
rect 8300 24792 8352 24812
rect 8352 24792 8354 24812
rect 8298 23976 8354 24032
rect 8298 22636 8354 22672
rect 8298 22616 8300 22636
rect 8300 22616 8352 22636
rect 8352 22616 8354 22636
rect 8298 21548 8354 21584
rect 8298 21528 8300 21548
rect 8300 21528 8352 21548
rect 8352 21528 8354 21548
rect 8298 18944 8354 19000
rect 8298 18536 8354 18592
rect 8298 17176 8354 17232
rect 8298 16088 8354 16144
rect 8298 13932 8354 13968
rect 8298 13912 8300 13932
rect 8300 13912 8352 13932
rect 8352 13912 8354 13932
rect 8298 13232 8354 13288
rect 8298 11736 8354 11792
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 35600 5466 35656 5468
rect 35680 5466 35736 5468
rect 35760 5466 35816 5468
rect 35840 5466 35896 5468
rect 35600 5414 35646 5466
rect 35646 5414 35656 5466
rect 35680 5414 35710 5466
rect 35710 5414 35722 5466
rect 35722 5414 35736 5466
rect 35760 5414 35774 5466
rect 35774 5414 35786 5466
rect 35786 5414 35816 5466
rect 35840 5414 35850 5466
rect 35850 5414 35896 5466
rect 35600 5412 35656 5414
rect 35680 5412 35736 5414
rect 35760 5412 35816 5414
rect 35840 5412 35896 5414
rect 35600 4378 35656 4380
rect 35680 4378 35736 4380
rect 35760 4378 35816 4380
rect 35840 4378 35896 4380
rect 35600 4326 35646 4378
rect 35646 4326 35656 4378
rect 35680 4326 35710 4378
rect 35710 4326 35722 4378
rect 35722 4326 35736 4378
rect 35760 4326 35774 4378
rect 35774 4326 35786 4378
rect 35786 4326 35816 4378
rect 35840 4326 35850 4378
rect 35850 4326 35896 4378
rect 35600 4324 35656 4326
rect 35680 4324 35736 4326
rect 35760 4324 35816 4326
rect 35840 4324 35896 4326
rect 35600 3290 35656 3292
rect 35680 3290 35736 3292
rect 35760 3290 35816 3292
rect 35840 3290 35896 3292
rect 35600 3238 35646 3290
rect 35646 3238 35656 3290
rect 35680 3238 35710 3290
rect 35710 3238 35722 3290
rect 35722 3238 35736 3290
rect 35760 3238 35774 3290
rect 35774 3238 35786 3290
rect 35786 3238 35816 3290
rect 35840 3238 35850 3290
rect 35850 3238 35896 3290
rect 35600 3236 35656 3238
rect 35680 3236 35736 3238
rect 35760 3236 35816 3238
rect 35840 3236 35896 3238
rect 97040 93594 97096 93596
rect 97120 93594 97176 93596
rect 97200 93594 97256 93596
rect 97280 93594 97336 93596
rect 97040 93542 97086 93594
rect 97086 93542 97096 93594
rect 97120 93542 97150 93594
rect 97150 93542 97162 93594
rect 97162 93542 97176 93594
rect 97200 93542 97214 93594
rect 97214 93542 97226 93594
rect 97226 93542 97256 93594
rect 97280 93542 97290 93594
rect 97290 93542 97336 93594
rect 97040 93540 97096 93542
rect 97120 93540 97176 93542
rect 97200 93540 97256 93542
rect 97280 93540 97336 93542
rect 96380 93050 96436 93052
rect 96460 93050 96516 93052
rect 96540 93050 96596 93052
rect 96620 93050 96676 93052
rect 96380 92998 96426 93050
rect 96426 92998 96436 93050
rect 96460 92998 96490 93050
rect 96490 92998 96502 93050
rect 96502 92998 96516 93050
rect 96540 92998 96554 93050
rect 96554 92998 96566 93050
rect 96566 92998 96596 93050
rect 96620 92998 96630 93050
rect 96630 92998 96676 93050
rect 96380 92996 96436 92998
rect 96460 92996 96516 92998
rect 96540 92996 96596 92998
rect 96620 92996 96676 92998
rect 97040 92506 97096 92508
rect 97120 92506 97176 92508
rect 97200 92506 97256 92508
rect 97280 92506 97336 92508
rect 97040 92454 97086 92506
rect 97086 92454 97096 92506
rect 97120 92454 97150 92506
rect 97150 92454 97162 92506
rect 97162 92454 97176 92506
rect 97200 92454 97214 92506
rect 97214 92454 97226 92506
rect 97226 92454 97256 92506
rect 97280 92454 97290 92506
rect 97290 92454 97336 92506
rect 97040 92452 97096 92454
rect 97120 92452 97176 92454
rect 97200 92452 97256 92454
rect 97280 92452 97336 92454
rect 96380 91962 96436 91964
rect 96460 91962 96516 91964
rect 96540 91962 96596 91964
rect 96620 91962 96676 91964
rect 96380 91910 96426 91962
rect 96426 91910 96436 91962
rect 96460 91910 96490 91962
rect 96490 91910 96502 91962
rect 96502 91910 96516 91962
rect 96540 91910 96554 91962
rect 96554 91910 96566 91962
rect 96566 91910 96596 91962
rect 96620 91910 96630 91962
rect 96630 91910 96676 91962
rect 96380 91908 96436 91910
rect 96460 91908 96516 91910
rect 96540 91908 96596 91910
rect 96620 91908 96676 91910
rect 97040 91418 97096 91420
rect 97120 91418 97176 91420
rect 97200 91418 97256 91420
rect 97280 91418 97336 91420
rect 97040 91366 97086 91418
rect 97086 91366 97096 91418
rect 97120 91366 97150 91418
rect 97150 91366 97162 91418
rect 97162 91366 97176 91418
rect 97200 91366 97214 91418
rect 97214 91366 97226 91418
rect 97226 91366 97256 91418
rect 97280 91366 97290 91418
rect 97290 91366 97336 91418
rect 97040 91364 97096 91366
rect 97120 91364 97176 91366
rect 97200 91364 97256 91366
rect 97280 91364 97336 91366
rect 96380 90874 96436 90876
rect 96460 90874 96516 90876
rect 96540 90874 96596 90876
rect 96620 90874 96676 90876
rect 96380 90822 96426 90874
rect 96426 90822 96436 90874
rect 96460 90822 96490 90874
rect 96490 90822 96502 90874
rect 96502 90822 96516 90874
rect 96540 90822 96554 90874
rect 96554 90822 96566 90874
rect 96566 90822 96596 90874
rect 96620 90822 96630 90874
rect 96630 90822 96676 90874
rect 96380 90820 96436 90822
rect 96460 90820 96516 90822
rect 96540 90820 96596 90822
rect 96620 90820 96676 90822
rect 97040 90330 97096 90332
rect 97120 90330 97176 90332
rect 97200 90330 97256 90332
rect 97280 90330 97336 90332
rect 97040 90278 97086 90330
rect 97086 90278 97096 90330
rect 97120 90278 97150 90330
rect 97150 90278 97162 90330
rect 97162 90278 97176 90330
rect 97200 90278 97214 90330
rect 97214 90278 97226 90330
rect 97226 90278 97256 90330
rect 97280 90278 97290 90330
rect 97290 90278 97336 90330
rect 97040 90276 97096 90278
rect 97120 90276 97176 90278
rect 97200 90276 97256 90278
rect 97280 90276 97336 90278
rect 96380 89786 96436 89788
rect 96460 89786 96516 89788
rect 96540 89786 96596 89788
rect 96620 89786 96676 89788
rect 96380 89734 96426 89786
rect 96426 89734 96436 89786
rect 96460 89734 96490 89786
rect 96490 89734 96502 89786
rect 96502 89734 96516 89786
rect 96540 89734 96554 89786
rect 96554 89734 96566 89786
rect 96566 89734 96596 89786
rect 96620 89734 96630 89786
rect 96630 89734 96676 89786
rect 96380 89732 96436 89734
rect 96460 89732 96516 89734
rect 96540 89732 96596 89734
rect 96620 89732 96676 89734
rect 97040 89242 97096 89244
rect 97120 89242 97176 89244
rect 97200 89242 97256 89244
rect 97280 89242 97336 89244
rect 97040 89190 97086 89242
rect 97086 89190 97096 89242
rect 97120 89190 97150 89242
rect 97150 89190 97162 89242
rect 97162 89190 97176 89242
rect 97200 89190 97214 89242
rect 97214 89190 97226 89242
rect 97226 89190 97256 89242
rect 97280 89190 97290 89242
rect 97290 89190 97336 89242
rect 97040 89188 97096 89190
rect 97120 89188 97176 89190
rect 97200 89188 97256 89190
rect 97280 89188 97336 89190
rect 96380 88698 96436 88700
rect 96460 88698 96516 88700
rect 96540 88698 96596 88700
rect 96620 88698 96676 88700
rect 96380 88646 96426 88698
rect 96426 88646 96436 88698
rect 96460 88646 96490 88698
rect 96490 88646 96502 88698
rect 96502 88646 96516 88698
rect 96540 88646 96554 88698
rect 96554 88646 96566 88698
rect 96566 88646 96596 88698
rect 96620 88646 96630 88698
rect 96630 88646 96676 88698
rect 96380 88644 96436 88646
rect 96460 88644 96516 88646
rect 96540 88644 96596 88646
rect 96620 88644 96676 88646
rect 97040 88154 97096 88156
rect 97120 88154 97176 88156
rect 97200 88154 97256 88156
rect 97280 88154 97336 88156
rect 97040 88102 97086 88154
rect 97086 88102 97096 88154
rect 97120 88102 97150 88154
rect 97150 88102 97162 88154
rect 97162 88102 97176 88154
rect 97200 88102 97214 88154
rect 97214 88102 97226 88154
rect 97226 88102 97256 88154
rect 97280 88102 97290 88154
rect 97290 88102 97336 88154
rect 97040 88100 97096 88102
rect 97120 88100 97176 88102
rect 97200 88100 97256 88102
rect 97280 88100 97336 88102
rect 96380 87610 96436 87612
rect 96460 87610 96516 87612
rect 96540 87610 96596 87612
rect 96620 87610 96676 87612
rect 96380 87558 96426 87610
rect 96426 87558 96436 87610
rect 96460 87558 96490 87610
rect 96490 87558 96502 87610
rect 96502 87558 96516 87610
rect 96540 87558 96554 87610
rect 96554 87558 96566 87610
rect 96566 87558 96596 87610
rect 96620 87558 96630 87610
rect 96630 87558 96676 87610
rect 96380 87556 96436 87558
rect 96460 87556 96516 87558
rect 96540 87556 96596 87558
rect 96620 87556 96676 87558
rect 97354 87388 97356 87408
rect 97356 87388 97408 87408
rect 97408 87388 97410 87408
rect 97354 87352 97410 87388
rect 97538 87080 97594 87136
rect 97040 87066 97096 87068
rect 97120 87066 97176 87068
rect 97200 87066 97256 87068
rect 97280 87066 97336 87068
rect 97040 87014 97086 87066
rect 97086 87014 97096 87066
rect 97120 87014 97150 87066
rect 97150 87014 97162 87066
rect 97162 87014 97176 87066
rect 97200 87014 97214 87066
rect 97214 87014 97226 87066
rect 97226 87014 97256 87066
rect 97280 87014 97290 87066
rect 97290 87014 97336 87066
rect 97040 87012 97096 87014
rect 97120 87012 97176 87014
rect 97200 87012 97256 87014
rect 97280 87012 97336 87014
rect 96380 86522 96436 86524
rect 96460 86522 96516 86524
rect 96540 86522 96596 86524
rect 96620 86522 96676 86524
rect 96380 86470 96426 86522
rect 96426 86470 96436 86522
rect 96460 86470 96490 86522
rect 96490 86470 96502 86522
rect 96502 86470 96516 86522
rect 96540 86470 96554 86522
rect 96554 86470 96566 86522
rect 96566 86470 96596 86522
rect 96620 86470 96630 86522
rect 96630 86470 96676 86522
rect 96380 86468 96436 86470
rect 96460 86468 96516 86470
rect 96540 86468 96596 86470
rect 96620 86468 96676 86470
rect 97538 86400 97594 86456
rect 97354 86264 97410 86320
rect 97040 85978 97096 85980
rect 97120 85978 97176 85980
rect 97200 85978 97256 85980
rect 97280 85978 97336 85980
rect 97040 85926 97086 85978
rect 97086 85926 97096 85978
rect 97120 85926 97150 85978
rect 97150 85926 97162 85978
rect 97162 85926 97176 85978
rect 97200 85926 97214 85978
rect 97214 85926 97226 85978
rect 97226 85926 97256 85978
rect 97280 85926 97290 85978
rect 97290 85926 97336 85978
rect 97040 85924 97096 85926
rect 97120 85924 97176 85926
rect 97200 85924 97256 85926
rect 97280 85924 97336 85926
rect 96380 85434 96436 85436
rect 96460 85434 96516 85436
rect 96540 85434 96596 85436
rect 96620 85434 96676 85436
rect 96380 85382 96426 85434
rect 96426 85382 96436 85434
rect 96460 85382 96490 85434
rect 96490 85382 96502 85434
rect 96502 85382 96516 85434
rect 96540 85382 96554 85434
rect 96554 85382 96566 85434
rect 96566 85382 96596 85434
rect 96620 85382 96630 85434
rect 96630 85382 96676 85434
rect 96380 85380 96436 85382
rect 96460 85380 96516 85382
rect 96540 85380 96596 85382
rect 96620 85380 96676 85382
rect 97354 85212 97356 85232
rect 97356 85212 97408 85232
rect 97408 85212 97410 85232
rect 97354 85176 97410 85212
rect 97538 85076 97540 85096
rect 97540 85076 97592 85096
rect 97592 85076 97594 85096
rect 97538 85040 97594 85076
rect 97040 84890 97096 84892
rect 97120 84890 97176 84892
rect 97200 84890 97256 84892
rect 97280 84890 97336 84892
rect 97040 84838 97086 84890
rect 97086 84838 97096 84890
rect 97120 84838 97150 84890
rect 97150 84838 97162 84890
rect 97162 84838 97176 84890
rect 97200 84838 97214 84890
rect 97214 84838 97226 84890
rect 97226 84838 97256 84890
rect 97280 84838 97290 84890
rect 97290 84838 97336 84890
rect 97040 84836 97096 84838
rect 97120 84836 97176 84838
rect 97200 84836 97256 84838
rect 97280 84836 97336 84838
rect 96380 84346 96436 84348
rect 96460 84346 96516 84348
rect 96540 84346 96596 84348
rect 96620 84346 96676 84348
rect 96380 84294 96426 84346
rect 96426 84294 96436 84346
rect 96460 84294 96490 84346
rect 96490 84294 96502 84346
rect 96502 84294 96516 84346
rect 96540 84294 96554 84346
rect 96554 84294 96566 84346
rect 96566 84294 96596 84346
rect 96620 84294 96630 84346
rect 96630 84294 96676 84346
rect 96380 84292 96436 84294
rect 96460 84292 96516 84294
rect 96540 84292 96596 84294
rect 96620 84292 96676 84294
rect 97538 84360 97594 84416
rect 97354 84088 97410 84144
rect 97040 83802 97096 83804
rect 97120 83802 97176 83804
rect 97200 83802 97256 83804
rect 97280 83802 97336 83804
rect 97040 83750 97086 83802
rect 97086 83750 97096 83802
rect 97120 83750 97150 83802
rect 97150 83750 97162 83802
rect 97162 83750 97176 83802
rect 97200 83750 97214 83802
rect 97214 83750 97226 83802
rect 97226 83750 97256 83802
rect 97280 83750 97290 83802
rect 97290 83750 97336 83802
rect 97040 83748 97096 83750
rect 97120 83748 97176 83750
rect 97200 83748 97256 83750
rect 97280 83748 97336 83750
rect 96380 83258 96436 83260
rect 96460 83258 96516 83260
rect 96540 83258 96596 83260
rect 96620 83258 96676 83260
rect 96380 83206 96426 83258
rect 96426 83206 96436 83258
rect 96460 83206 96490 83258
rect 96490 83206 96502 83258
rect 96502 83206 96516 83258
rect 96540 83206 96554 83258
rect 96554 83206 96566 83258
rect 96566 83206 96596 83258
rect 96620 83206 96630 83258
rect 96630 83206 96676 83258
rect 96380 83204 96436 83206
rect 96460 83204 96516 83206
rect 96540 83204 96596 83206
rect 96620 83204 96676 83206
rect 97354 83000 97410 83056
rect 97538 83000 97594 83056
rect 97040 82714 97096 82716
rect 97120 82714 97176 82716
rect 97200 82714 97256 82716
rect 97280 82714 97336 82716
rect 97040 82662 97086 82714
rect 97086 82662 97096 82714
rect 97120 82662 97150 82714
rect 97150 82662 97162 82714
rect 97162 82662 97176 82714
rect 97200 82662 97214 82714
rect 97214 82662 97226 82714
rect 97226 82662 97256 82714
rect 97280 82662 97290 82714
rect 97290 82662 97336 82714
rect 97040 82660 97096 82662
rect 97120 82660 97176 82662
rect 97200 82660 97256 82662
rect 97280 82660 97336 82662
rect 96380 82170 96436 82172
rect 96460 82170 96516 82172
rect 96540 82170 96596 82172
rect 96620 82170 96676 82172
rect 96380 82118 96426 82170
rect 96426 82118 96436 82170
rect 96460 82118 96490 82170
rect 96490 82118 96502 82170
rect 96502 82118 96516 82170
rect 96540 82118 96554 82170
rect 96554 82118 96566 82170
rect 96566 82118 96596 82170
rect 96620 82118 96630 82170
rect 96630 82118 96676 82170
rect 96380 82116 96436 82118
rect 96460 82116 96516 82118
rect 96540 82116 96596 82118
rect 96620 82116 96676 82118
rect 97354 81948 97356 81968
rect 97356 81948 97408 81968
rect 97408 81948 97410 81968
rect 97354 81912 97410 81948
rect 97538 81640 97594 81696
rect 97040 81626 97096 81628
rect 97120 81626 97176 81628
rect 97200 81626 97256 81628
rect 97280 81626 97336 81628
rect 97040 81574 97086 81626
rect 97086 81574 97096 81626
rect 97120 81574 97150 81626
rect 97150 81574 97162 81626
rect 97162 81574 97176 81626
rect 97200 81574 97214 81626
rect 97214 81574 97226 81626
rect 97226 81574 97256 81626
rect 97280 81574 97290 81626
rect 97290 81574 97336 81626
rect 97040 81572 97096 81574
rect 97120 81572 97176 81574
rect 97200 81572 97256 81574
rect 97280 81572 97336 81574
rect 96380 81082 96436 81084
rect 96460 81082 96516 81084
rect 96540 81082 96596 81084
rect 96620 81082 96676 81084
rect 96380 81030 96426 81082
rect 96426 81030 96436 81082
rect 96460 81030 96490 81082
rect 96490 81030 96502 81082
rect 96502 81030 96516 81082
rect 96540 81030 96554 81082
rect 96554 81030 96566 81082
rect 96566 81030 96596 81082
rect 96620 81030 96630 81082
rect 96630 81030 96676 81082
rect 96380 81028 96436 81030
rect 96460 81028 96516 81030
rect 96540 81028 96596 81030
rect 96620 81028 96676 81030
rect 97538 80960 97594 81016
rect 97354 80824 97410 80880
rect 97040 80538 97096 80540
rect 97120 80538 97176 80540
rect 97200 80538 97256 80540
rect 97280 80538 97336 80540
rect 97040 80486 97086 80538
rect 97086 80486 97096 80538
rect 97120 80486 97150 80538
rect 97150 80486 97162 80538
rect 97162 80486 97176 80538
rect 97200 80486 97214 80538
rect 97214 80486 97226 80538
rect 97226 80486 97256 80538
rect 97280 80486 97290 80538
rect 97290 80486 97336 80538
rect 97040 80484 97096 80486
rect 97120 80484 97176 80486
rect 97200 80484 97256 80486
rect 97280 80484 97336 80486
rect 96380 79994 96436 79996
rect 96460 79994 96516 79996
rect 96540 79994 96596 79996
rect 96620 79994 96676 79996
rect 96380 79942 96426 79994
rect 96426 79942 96436 79994
rect 96460 79942 96490 79994
rect 96490 79942 96502 79994
rect 96502 79942 96516 79994
rect 96540 79942 96554 79994
rect 96554 79942 96566 79994
rect 96566 79942 96596 79994
rect 96620 79942 96630 79994
rect 96630 79942 96676 79994
rect 96380 79940 96436 79942
rect 96460 79940 96516 79942
rect 96540 79940 96596 79942
rect 96620 79940 96676 79942
rect 97354 79772 97356 79792
rect 97356 79772 97408 79792
rect 97408 79772 97410 79792
rect 97354 79736 97410 79772
rect 97538 79636 97540 79656
rect 97540 79636 97592 79656
rect 97592 79636 97594 79656
rect 97538 79600 97594 79636
rect 97040 79450 97096 79452
rect 97120 79450 97176 79452
rect 97200 79450 97256 79452
rect 97280 79450 97336 79452
rect 97040 79398 97086 79450
rect 97086 79398 97096 79450
rect 97120 79398 97150 79450
rect 97150 79398 97162 79450
rect 97162 79398 97176 79450
rect 97200 79398 97214 79450
rect 97214 79398 97226 79450
rect 97226 79398 97256 79450
rect 97280 79398 97290 79450
rect 97290 79398 97336 79450
rect 97040 79396 97096 79398
rect 97120 79396 97176 79398
rect 97200 79396 97256 79398
rect 97280 79396 97336 79398
rect 96380 78906 96436 78908
rect 96460 78906 96516 78908
rect 96540 78906 96596 78908
rect 96620 78906 96676 78908
rect 96380 78854 96426 78906
rect 96426 78854 96436 78906
rect 96460 78854 96490 78906
rect 96490 78854 96502 78906
rect 96502 78854 96516 78906
rect 96540 78854 96554 78906
rect 96554 78854 96566 78906
rect 96566 78854 96596 78906
rect 96620 78854 96630 78906
rect 96630 78854 96676 78906
rect 96380 78852 96436 78854
rect 96460 78852 96516 78854
rect 96540 78852 96596 78854
rect 96620 78852 96676 78854
rect 97446 78920 97502 78976
rect 97262 78648 97318 78704
rect 97040 78362 97096 78364
rect 97120 78362 97176 78364
rect 97200 78362 97256 78364
rect 97280 78362 97336 78364
rect 97040 78310 97086 78362
rect 97086 78310 97096 78362
rect 97120 78310 97150 78362
rect 97150 78310 97162 78362
rect 97162 78310 97176 78362
rect 97200 78310 97214 78362
rect 97214 78310 97226 78362
rect 97226 78310 97256 78362
rect 97280 78310 97290 78362
rect 97290 78310 97336 78362
rect 97040 78308 97096 78310
rect 97120 78308 97176 78310
rect 97200 78308 97256 78310
rect 97280 78308 97336 78310
rect 96380 77818 96436 77820
rect 96460 77818 96516 77820
rect 96540 77818 96596 77820
rect 96620 77818 96676 77820
rect 96380 77766 96426 77818
rect 96426 77766 96436 77818
rect 96460 77766 96490 77818
rect 96490 77766 96502 77818
rect 96502 77766 96516 77818
rect 96540 77766 96554 77818
rect 96554 77766 96566 77818
rect 96566 77766 96596 77818
rect 96620 77766 96630 77818
rect 96630 77766 96676 77818
rect 96380 77764 96436 77766
rect 96460 77764 96516 77766
rect 96540 77764 96596 77766
rect 96620 77764 96676 77766
rect 97354 77560 97410 77616
rect 97538 77560 97594 77616
rect 97040 77274 97096 77276
rect 97120 77274 97176 77276
rect 97200 77274 97256 77276
rect 97280 77274 97336 77276
rect 97040 77222 97086 77274
rect 97086 77222 97096 77274
rect 97120 77222 97150 77274
rect 97150 77222 97162 77274
rect 97162 77222 97176 77274
rect 97200 77222 97214 77274
rect 97214 77222 97226 77274
rect 97226 77222 97256 77274
rect 97280 77222 97290 77274
rect 97290 77222 97336 77274
rect 97040 77220 97096 77222
rect 97120 77220 97176 77222
rect 97200 77220 97256 77222
rect 97280 77220 97336 77222
rect 96380 76730 96436 76732
rect 96460 76730 96516 76732
rect 96540 76730 96596 76732
rect 96620 76730 96676 76732
rect 96380 76678 96426 76730
rect 96426 76678 96436 76730
rect 96460 76678 96490 76730
rect 96490 76678 96502 76730
rect 96502 76678 96516 76730
rect 96540 76678 96554 76730
rect 96554 76678 96566 76730
rect 96566 76678 96596 76730
rect 96620 76678 96630 76730
rect 96630 76678 96676 76730
rect 96380 76676 96436 76678
rect 96460 76676 96516 76678
rect 96540 76676 96596 76678
rect 96620 76676 96676 76678
rect 97354 76508 97356 76528
rect 97356 76508 97408 76528
rect 97408 76508 97410 76528
rect 97354 76472 97410 76508
rect 97538 76200 97594 76256
rect 97040 76186 97096 76188
rect 97120 76186 97176 76188
rect 97200 76186 97256 76188
rect 97280 76186 97336 76188
rect 97040 76134 97086 76186
rect 97086 76134 97096 76186
rect 97120 76134 97150 76186
rect 97150 76134 97162 76186
rect 97162 76134 97176 76186
rect 97200 76134 97214 76186
rect 97214 76134 97226 76186
rect 97226 76134 97256 76186
rect 97280 76134 97290 76186
rect 97290 76134 97336 76186
rect 97040 76132 97096 76134
rect 97120 76132 97176 76134
rect 97200 76132 97256 76134
rect 97280 76132 97336 76134
rect 96380 75642 96436 75644
rect 96460 75642 96516 75644
rect 96540 75642 96596 75644
rect 96620 75642 96676 75644
rect 96380 75590 96426 75642
rect 96426 75590 96436 75642
rect 96460 75590 96490 75642
rect 96490 75590 96502 75642
rect 96502 75590 96516 75642
rect 96540 75590 96554 75642
rect 96554 75590 96566 75642
rect 96566 75590 96596 75642
rect 96620 75590 96630 75642
rect 96630 75590 96676 75642
rect 96380 75588 96436 75590
rect 96460 75588 96516 75590
rect 96540 75588 96596 75590
rect 96620 75588 96676 75590
rect 97538 75520 97594 75576
rect 97354 75384 97410 75440
rect 97040 75098 97096 75100
rect 97120 75098 97176 75100
rect 97200 75098 97256 75100
rect 97280 75098 97336 75100
rect 97040 75046 97086 75098
rect 97086 75046 97096 75098
rect 97120 75046 97150 75098
rect 97150 75046 97162 75098
rect 97162 75046 97176 75098
rect 97200 75046 97214 75098
rect 97214 75046 97226 75098
rect 97226 75046 97256 75098
rect 97280 75046 97290 75098
rect 97290 75046 97336 75098
rect 97040 75044 97096 75046
rect 97120 75044 97176 75046
rect 97200 75044 97256 75046
rect 97280 75044 97336 75046
rect 96380 74554 96436 74556
rect 96460 74554 96516 74556
rect 96540 74554 96596 74556
rect 96620 74554 96676 74556
rect 96380 74502 96426 74554
rect 96426 74502 96436 74554
rect 96460 74502 96490 74554
rect 96490 74502 96502 74554
rect 96502 74502 96516 74554
rect 96540 74502 96554 74554
rect 96554 74502 96566 74554
rect 96566 74502 96596 74554
rect 96620 74502 96630 74554
rect 96630 74502 96676 74554
rect 96380 74500 96436 74502
rect 96460 74500 96516 74502
rect 96540 74500 96596 74502
rect 96620 74500 96676 74502
rect 97262 74332 97264 74352
rect 97264 74332 97316 74352
rect 97316 74332 97318 74352
rect 97262 74296 97318 74332
rect 97446 74180 97502 74216
rect 97446 74160 97448 74180
rect 97448 74160 97500 74180
rect 97500 74160 97502 74180
rect 97040 74010 97096 74012
rect 97120 74010 97176 74012
rect 97200 74010 97256 74012
rect 97280 74010 97336 74012
rect 97040 73958 97086 74010
rect 97086 73958 97096 74010
rect 97120 73958 97150 74010
rect 97150 73958 97162 74010
rect 97162 73958 97176 74010
rect 97200 73958 97214 74010
rect 97214 73958 97226 74010
rect 97226 73958 97256 74010
rect 97280 73958 97290 74010
rect 97290 73958 97336 74010
rect 97040 73956 97096 73958
rect 97120 73956 97176 73958
rect 97200 73956 97256 73958
rect 97280 73956 97336 73958
rect 96380 73466 96436 73468
rect 96460 73466 96516 73468
rect 96540 73466 96596 73468
rect 96620 73466 96676 73468
rect 96380 73414 96426 73466
rect 96426 73414 96436 73466
rect 96460 73414 96490 73466
rect 96490 73414 96502 73466
rect 96502 73414 96516 73466
rect 96540 73414 96554 73466
rect 96554 73414 96566 73466
rect 96566 73414 96596 73466
rect 96620 73414 96630 73466
rect 96630 73414 96676 73466
rect 96380 73412 96436 73414
rect 96460 73412 96516 73414
rect 96540 73412 96596 73414
rect 96620 73412 96676 73414
rect 97538 73480 97594 73536
rect 97354 73208 97410 73264
rect 97040 72922 97096 72924
rect 97120 72922 97176 72924
rect 97200 72922 97256 72924
rect 97280 72922 97336 72924
rect 97040 72870 97086 72922
rect 97086 72870 97096 72922
rect 97120 72870 97150 72922
rect 97150 72870 97162 72922
rect 97162 72870 97176 72922
rect 97200 72870 97214 72922
rect 97214 72870 97226 72922
rect 97226 72870 97256 72922
rect 97280 72870 97290 72922
rect 97290 72870 97336 72922
rect 97040 72868 97096 72870
rect 97120 72868 97176 72870
rect 97200 72868 97256 72870
rect 97280 72868 97336 72870
rect 96380 72378 96436 72380
rect 96460 72378 96516 72380
rect 96540 72378 96596 72380
rect 96620 72378 96676 72380
rect 96380 72326 96426 72378
rect 96426 72326 96436 72378
rect 96460 72326 96490 72378
rect 96490 72326 96502 72378
rect 96502 72326 96516 72378
rect 96540 72326 96554 72378
rect 96554 72326 96566 72378
rect 96566 72326 96596 72378
rect 96620 72326 96630 72378
rect 96630 72326 96676 72378
rect 96380 72324 96436 72326
rect 96460 72324 96516 72326
rect 96540 72324 96596 72326
rect 96620 72324 96676 72326
rect 97262 72120 97318 72176
rect 97538 72156 97540 72176
rect 97540 72156 97592 72176
rect 97592 72156 97594 72176
rect 97538 72120 97594 72156
rect 97040 71834 97096 71836
rect 97120 71834 97176 71836
rect 97200 71834 97256 71836
rect 97280 71834 97336 71836
rect 97040 71782 97086 71834
rect 97086 71782 97096 71834
rect 97120 71782 97150 71834
rect 97150 71782 97162 71834
rect 97162 71782 97176 71834
rect 97200 71782 97214 71834
rect 97214 71782 97226 71834
rect 97226 71782 97256 71834
rect 97280 71782 97290 71834
rect 97290 71782 97336 71834
rect 97040 71780 97096 71782
rect 97120 71780 97176 71782
rect 97200 71780 97256 71782
rect 97280 71780 97336 71782
rect 96380 71290 96436 71292
rect 96460 71290 96516 71292
rect 96540 71290 96596 71292
rect 96620 71290 96676 71292
rect 96380 71238 96426 71290
rect 96426 71238 96436 71290
rect 96460 71238 96490 71290
rect 96490 71238 96502 71290
rect 96502 71238 96516 71290
rect 96540 71238 96554 71290
rect 96554 71238 96566 71290
rect 96566 71238 96596 71290
rect 96620 71238 96630 71290
rect 96630 71238 96676 71290
rect 96380 71236 96436 71238
rect 96460 71236 96516 71238
rect 96540 71236 96596 71238
rect 96620 71236 96676 71238
rect 97354 71068 97356 71088
rect 97356 71068 97408 71088
rect 97408 71068 97410 71088
rect 97354 71032 97410 71068
rect 97538 70760 97594 70816
rect 97040 70746 97096 70748
rect 97120 70746 97176 70748
rect 97200 70746 97256 70748
rect 97280 70746 97336 70748
rect 97040 70694 97086 70746
rect 97086 70694 97096 70746
rect 97120 70694 97150 70746
rect 97150 70694 97162 70746
rect 97162 70694 97176 70746
rect 97200 70694 97214 70746
rect 97214 70694 97226 70746
rect 97226 70694 97256 70746
rect 97280 70694 97290 70746
rect 97290 70694 97336 70746
rect 97040 70692 97096 70694
rect 97120 70692 97176 70694
rect 97200 70692 97256 70694
rect 97280 70692 97336 70694
rect 96380 70202 96436 70204
rect 96460 70202 96516 70204
rect 96540 70202 96596 70204
rect 96620 70202 96676 70204
rect 96380 70150 96426 70202
rect 96426 70150 96436 70202
rect 96460 70150 96490 70202
rect 96490 70150 96502 70202
rect 96502 70150 96516 70202
rect 96540 70150 96554 70202
rect 96554 70150 96566 70202
rect 96566 70150 96596 70202
rect 96620 70150 96630 70202
rect 96630 70150 96676 70202
rect 96380 70148 96436 70150
rect 96460 70148 96516 70150
rect 96540 70148 96596 70150
rect 96620 70148 96676 70150
rect 97446 70080 97502 70136
rect 97262 69944 97318 70000
rect 97040 69658 97096 69660
rect 97120 69658 97176 69660
rect 97200 69658 97256 69660
rect 97280 69658 97336 69660
rect 97040 69606 97086 69658
rect 97086 69606 97096 69658
rect 97120 69606 97150 69658
rect 97150 69606 97162 69658
rect 97162 69606 97176 69658
rect 97200 69606 97214 69658
rect 97214 69606 97226 69658
rect 97226 69606 97256 69658
rect 97280 69606 97290 69658
rect 97290 69606 97336 69658
rect 97040 69604 97096 69606
rect 97120 69604 97176 69606
rect 97200 69604 97256 69606
rect 97280 69604 97336 69606
rect 96380 69114 96436 69116
rect 96460 69114 96516 69116
rect 96540 69114 96596 69116
rect 96620 69114 96676 69116
rect 96380 69062 96426 69114
rect 96426 69062 96436 69114
rect 96460 69062 96490 69114
rect 96490 69062 96502 69114
rect 96502 69062 96516 69114
rect 96540 69062 96554 69114
rect 96554 69062 96566 69114
rect 96566 69062 96596 69114
rect 96620 69062 96630 69114
rect 96630 69062 96676 69114
rect 96380 69060 96436 69062
rect 96460 69060 96516 69062
rect 96540 69060 96596 69062
rect 96620 69060 96676 69062
rect 97262 68856 97318 68912
rect 97446 68720 97502 68776
rect 97040 68570 97096 68572
rect 97120 68570 97176 68572
rect 97200 68570 97256 68572
rect 97280 68570 97336 68572
rect 97040 68518 97086 68570
rect 97086 68518 97096 68570
rect 97120 68518 97150 68570
rect 97150 68518 97162 68570
rect 97162 68518 97176 68570
rect 97200 68518 97214 68570
rect 97214 68518 97226 68570
rect 97226 68518 97256 68570
rect 97280 68518 97290 68570
rect 97290 68518 97336 68570
rect 97040 68516 97096 68518
rect 97120 68516 97176 68518
rect 97200 68516 97256 68518
rect 97280 68516 97336 68518
rect 96380 68026 96436 68028
rect 96460 68026 96516 68028
rect 96540 68026 96596 68028
rect 96620 68026 96676 68028
rect 96380 67974 96426 68026
rect 96426 67974 96436 68026
rect 96460 67974 96490 68026
rect 96490 67974 96502 68026
rect 96502 67974 96516 68026
rect 96540 67974 96554 68026
rect 96554 67974 96566 68026
rect 96566 67974 96596 68026
rect 96620 67974 96630 68026
rect 96630 67974 96676 68026
rect 96380 67972 96436 67974
rect 96460 67972 96516 67974
rect 96540 67972 96596 67974
rect 96620 67972 96676 67974
rect 97446 68076 97448 68096
rect 97448 68076 97500 68096
rect 97500 68076 97502 68096
rect 97446 68040 97502 68076
rect 97262 67768 97318 67824
rect 97040 67482 97096 67484
rect 97120 67482 97176 67484
rect 97200 67482 97256 67484
rect 97280 67482 97336 67484
rect 97040 67430 97086 67482
rect 97086 67430 97096 67482
rect 97120 67430 97150 67482
rect 97150 67430 97162 67482
rect 97162 67430 97176 67482
rect 97200 67430 97214 67482
rect 97214 67430 97226 67482
rect 97226 67430 97256 67482
rect 97280 67430 97290 67482
rect 97290 67430 97336 67482
rect 97040 67428 97096 67430
rect 97120 67428 97176 67430
rect 97200 67428 97256 67430
rect 97280 67428 97336 67430
rect 96380 66938 96436 66940
rect 96460 66938 96516 66940
rect 96540 66938 96596 66940
rect 96620 66938 96676 66940
rect 96380 66886 96426 66938
rect 96426 66886 96436 66938
rect 96460 66886 96490 66938
rect 96490 66886 96502 66938
rect 96502 66886 96516 66938
rect 96540 66886 96554 66938
rect 96554 66886 96566 66938
rect 96566 66886 96596 66938
rect 96620 66886 96630 66938
rect 96630 66886 96676 66938
rect 96380 66884 96436 66886
rect 96460 66884 96516 66886
rect 96540 66884 96596 66886
rect 96620 66884 96676 66886
rect 97262 66680 97318 66736
rect 97446 66680 97502 66736
rect 97040 66394 97096 66396
rect 97120 66394 97176 66396
rect 97200 66394 97256 66396
rect 97280 66394 97336 66396
rect 97040 66342 97086 66394
rect 97086 66342 97096 66394
rect 97120 66342 97150 66394
rect 97150 66342 97162 66394
rect 97162 66342 97176 66394
rect 97200 66342 97214 66394
rect 97214 66342 97226 66394
rect 97226 66342 97256 66394
rect 97280 66342 97290 66394
rect 97290 66342 97336 66394
rect 97040 66340 97096 66342
rect 97120 66340 97176 66342
rect 97200 66340 97256 66342
rect 97280 66340 97336 66342
rect 96380 65850 96436 65852
rect 96460 65850 96516 65852
rect 96540 65850 96596 65852
rect 96620 65850 96676 65852
rect 96380 65798 96426 65850
rect 96426 65798 96436 65850
rect 96460 65798 96490 65850
rect 96490 65798 96502 65850
rect 96502 65798 96516 65850
rect 96540 65798 96554 65850
rect 96554 65798 96566 65850
rect 96566 65798 96596 65850
rect 96620 65798 96630 65850
rect 96630 65798 96676 65850
rect 96380 65796 96436 65798
rect 96460 65796 96516 65798
rect 96540 65796 96596 65798
rect 96620 65796 96676 65798
rect 97262 65592 97318 65648
rect 97446 65356 97448 65376
rect 97448 65356 97500 65376
rect 97500 65356 97502 65376
rect 97446 65320 97502 65356
rect 97040 65306 97096 65308
rect 97120 65306 97176 65308
rect 97200 65306 97256 65308
rect 97280 65306 97336 65308
rect 97040 65254 97086 65306
rect 97086 65254 97096 65306
rect 97120 65254 97150 65306
rect 97150 65254 97162 65306
rect 97162 65254 97176 65306
rect 97200 65254 97214 65306
rect 97214 65254 97226 65306
rect 97226 65254 97256 65306
rect 97280 65254 97290 65306
rect 97290 65254 97336 65306
rect 97040 65252 97096 65254
rect 97120 65252 97176 65254
rect 97200 65252 97256 65254
rect 97280 65252 97336 65254
rect 96380 64762 96436 64764
rect 96460 64762 96516 64764
rect 96540 64762 96596 64764
rect 96620 64762 96676 64764
rect 96380 64710 96426 64762
rect 96426 64710 96436 64762
rect 96460 64710 96490 64762
rect 96490 64710 96502 64762
rect 96502 64710 96516 64762
rect 96540 64710 96554 64762
rect 96554 64710 96566 64762
rect 96566 64710 96596 64762
rect 96620 64710 96630 64762
rect 96630 64710 96676 64762
rect 96380 64708 96436 64710
rect 96460 64708 96516 64710
rect 96540 64708 96596 64710
rect 96620 64708 96676 64710
rect 97446 64640 97502 64696
rect 97262 64504 97318 64560
rect 97040 64218 97096 64220
rect 97120 64218 97176 64220
rect 97200 64218 97256 64220
rect 97280 64218 97336 64220
rect 97040 64166 97086 64218
rect 97086 64166 97096 64218
rect 97120 64166 97150 64218
rect 97150 64166 97162 64218
rect 97162 64166 97176 64218
rect 97200 64166 97214 64218
rect 97214 64166 97226 64218
rect 97226 64166 97256 64218
rect 97280 64166 97290 64218
rect 97290 64166 97336 64218
rect 97040 64164 97096 64166
rect 97120 64164 97176 64166
rect 97200 64164 97256 64166
rect 97280 64164 97336 64166
rect 96380 63674 96436 63676
rect 96460 63674 96516 63676
rect 96540 63674 96596 63676
rect 96620 63674 96676 63676
rect 96380 63622 96426 63674
rect 96426 63622 96436 63674
rect 96460 63622 96490 63674
rect 96490 63622 96502 63674
rect 96502 63622 96516 63674
rect 96540 63622 96554 63674
rect 96554 63622 96566 63674
rect 96566 63622 96596 63674
rect 96620 63622 96630 63674
rect 96630 63622 96676 63674
rect 96380 63620 96436 63622
rect 96460 63620 96516 63622
rect 96540 63620 96596 63622
rect 96620 63620 96676 63622
rect 97262 63416 97318 63472
rect 97446 63280 97502 63336
rect 97040 63130 97096 63132
rect 97120 63130 97176 63132
rect 97200 63130 97256 63132
rect 97280 63130 97336 63132
rect 97040 63078 97086 63130
rect 97086 63078 97096 63130
rect 97120 63078 97150 63130
rect 97150 63078 97162 63130
rect 97162 63078 97176 63130
rect 97200 63078 97214 63130
rect 97214 63078 97226 63130
rect 97226 63078 97256 63130
rect 97280 63078 97290 63130
rect 97290 63078 97336 63130
rect 97040 63076 97096 63078
rect 97120 63076 97176 63078
rect 97200 63076 97256 63078
rect 97280 63076 97336 63078
rect 96380 62586 96436 62588
rect 96460 62586 96516 62588
rect 96540 62586 96596 62588
rect 96620 62586 96676 62588
rect 96380 62534 96426 62586
rect 96426 62534 96436 62586
rect 96460 62534 96490 62586
rect 96490 62534 96502 62586
rect 96502 62534 96516 62586
rect 96540 62534 96554 62586
rect 96554 62534 96566 62586
rect 96566 62534 96596 62586
rect 96620 62534 96630 62586
rect 96630 62534 96676 62586
rect 96380 62532 96436 62534
rect 96460 62532 96516 62534
rect 96540 62532 96596 62534
rect 96620 62532 96676 62534
rect 97446 62636 97448 62656
rect 97448 62636 97500 62656
rect 97500 62636 97502 62656
rect 97446 62600 97502 62636
rect 97262 62328 97318 62384
rect 97040 62042 97096 62044
rect 97120 62042 97176 62044
rect 97200 62042 97256 62044
rect 97280 62042 97336 62044
rect 97040 61990 97086 62042
rect 97086 61990 97096 62042
rect 97120 61990 97150 62042
rect 97150 61990 97162 62042
rect 97162 61990 97176 62042
rect 97200 61990 97214 62042
rect 97214 61990 97226 62042
rect 97226 61990 97256 62042
rect 97280 61990 97290 62042
rect 97290 61990 97336 62042
rect 97040 61988 97096 61990
rect 97120 61988 97176 61990
rect 97200 61988 97256 61990
rect 97280 61988 97336 61990
rect 96380 61498 96436 61500
rect 96460 61498 96516 61500
rect 96540 61498 96596 61500
rect 96620 61498 96676 61500
rect 96380 61446 96426 61498
rect 96426 61446 96436 61498
rect 96460 61446 96490 61498
rect 96490 61446 96502 61498
rect 96502 61446 96516 61498
rect 96540 61446 96554 61498
rect 96554 61446 96566 61498
rect 96566 61446 96596 61498
rect 96620 61446 96630 61498
rect 96630 61446 96676 61498
rect 96380 61444 96436 61446
rect 96460 61444 96516 61446
rect 96540 61444 96596 61446
rect 96620 61444 96676 61446
rect 97262 61240 97318 61296
rect 97446 61240 97502 61296
rect 97040 60954 97096 60956
rect 97120 60954 97176 60956
rect 97200 60954 97256 60956
rect 97280 60954 97336 60956
rect 97040 60902 97086 60954
rect 97086 60902 97096 60954
rect 97120 60902 97150 60954
rect 97150 60902 97162 60954
rect 97162 60902 97176 60954
rect 97200 60902 97214 60954
rect 97214 60902 97226 60954
rect 97226 60902 97256 60954
rect 97280 60902 97290 60954
rect 97290 60902 97336 60954
rect 97040 60900 97096 60902
rect 97120 60900 97176 60902
rect 97200 60900 97256 60902
rect 97280 60900 97336 60902
rect 96380 60410 96436 60412
rect 96460 60410 96516 60412
rect 96540 60410 96596 60412
rect 96620 60410 96676 60412
rect 96380 60358 96426 60410
rect 96426 60358 96436 60410
rect 96460 60358 96490 60410
rect 96490 60358 96502 60410
rect 96502 60358 96516 60410
rect 96540 60358 96554 60410
rect 96554 60358 96566 60410
rect 96566 60358 96596 60410
rect 96620 60358 96630 60410
rect 96630 60358 96676 60410
rect 96380 60356 96436 60358
rect 96460 60356 96516 60358
rect 96540 60356 96596 60358
rect 96620 60356 96676 60358
rect 97262 60152 97318 60208
rect 97446 59916 97448 59936
rect 97448 59916 97500 59936
rect 97500 59916 97502 59936
rect 97446 59880 97502 59916
rect 97040 59866 97096 59868
rect 97120 59866 97176 59868
rect 97200 59866 97256 59868
rect 97280 59866 97336 59868
rect 97040 59814 97086 59866
rect 97086 59814 97096 59866
rect 97120 59814 97150 59866
rect 97150 59814 97162 59866
rect 97162 59814 97176 59866
rect 97200 59814 97214 59866
rect 97214 59814 97226 59866
rect 97226 59814 97256 59866
rect 97280 59814 97290 59866
rect 97290 59814 97336 59866
rect 97040 59812 97096 59814
rect 97120 59812 97176 59814
rect 97200 59812 97256 59814
rect 97280 59812 97336 59814
rect 96380 59322 96436 59324
rect 96460 59322 96516 59324
rect 96540 59322 96596 59324
rect 96620 59322 96676 59324
rect 96380 59270 96426 59322
rect 96426 59270 96436 59322
rect 96460 59270 96490 59322
rect 96490 59270 96502 59322
rect 96502 59270 96516 59322
rect 96540 59270 96554 59322
rect 96554 59270 96566 59322
rect 96566 59270 96596 59322
rect 96620 59270 96630 59322
rect 96630 59270 96676 59322
rect 96380 59268 96436 59270
rect 96460 59268 96516 59270
rect 96540 59268 96596 59270
rect 96620 59268 96676 59270
rect 97446 59200 97502 59256
rect 97262 59064 97318 59120
rect 97040 58778 97096 58780
rect 97120 58778 97176 58780
rect 97200 58778 97256 58780
rect 97280 58778 97336 58780
rect 97040 58726 97086 58778
rect 97086 58726 97096 58778
rect 97120 58726 97150 58778
rect 97150 58726 97162 58778
rect 97162 58726 97176 58778
rect 97200 58726 97214 58778
rect 97214 58726 97226 58778
rect 97226 58726 97256 58778
rect 97280 58726 97290 58778
rect 97290 58726 97336 58778
rect 97040 58724 97096 58726
rect 97120 58724 97176 58726
rect 97200 58724 97256 58726
rect 97280 58724 97336 58726
rect 96380 58234 96436 58236
rect 96460 58234 96516 58236
rect 96540 58234 96596 58236
rect 96620 58234 96676 58236
rect 96380 58182 96426 58234
rect 96426 58182 96436 58234
rect 96460 58182 96490 58234
rect 96490 58182 96502 58234
rect 96502 58182 96516 58234
rect 96540 58182 96554 58234
rect 96554 58182 96566 58234
rect 96566 58182 96596 58234
rect 96620 58182 96630 58234
rect 96630 58182 96676 58234
rect 96380 58180 96436 58182
rect 96460 58180 96516 58182
rect 96540 58180 96596 58182
rect 96620 58180 96676 58182
rect 97262 57976 97318 58032
rect 97446 57840 97502 57896
rect 97040 57690 97096 57692
rect 97120 57690 97176 57692
rect 97200 57690 97256 57692
rect 97280 57690 97336 57692
rect 97040 57638 97086 57690
rect 97086 57638 97096 57690
rect 97120 57638 97150 57690
rect 97150 57638 97162 57690
rect 97162 57638 97176 57690
rect 97200 57638 97214 57690
rect 97214 57638 97226 57690
rect 97226 57638 97256 57690
rect 97280 57638 97290 57690
rect 97290 57638 97336 57690
rect 97040 57636 97096 57638
rect 97120 57636 97176 57638
rect 97200 57636 97256 57638
rect 97280 57636 97336 57638
rect 96380 57146 96436 57148
rect 96460 57146 96516 57148
rect 96540 57146 96596 57148
rect 96620 57146 96676 57148
rect 96380 57094 96426 57146
rect 96426 57094 96436 57146
rect 96460 57094 96490 57146
rect 96490 57094 96502 57146
rect 96502 57094 96516 57146
rect 96540 57094 96554 57146
rect 96554 57094 96566 57146
rect 96566 57094 96596 57146
rect 96620 57094 96630 57146
rect 96630 57094 96676 57146
rect 96380 57092 96436 57094
rect 96460 57092 96516 57094
rect 96540 57092 96596 57094
rect 96620 57092 96676 57094
rect 97446 57196 97448 57216
rect 97448 57196 97500 57216
rect 97500 57196 97502 57216
rect 97446 57160 97502 57196
rect 97262 56888 97318 56944
rect 97040 56602 97096 56604
rect 97120 56602 97176 56604
rect 97200 56602 97256 56604
rect 97280 56602 97336 56604
rect 97040 56550 97086 56602
rect 97086 56550 97096 56602
rect 97120 56550 97150 56602
rect 97150 56550 97162 56602
rect 97162 56550 97176 56602
rect 97200 56550 97214 56602
rect 97214 56550 97226 56602
rect 97226 56550 97256 56602
rect 97280 56550 97290 56602
rect 97290 56550 97336 56602
rect 97040 56548 97096 56550
rect 97120 56548 97176 56550
rect 97200 56548 97256 56550
rect 97280 56548 97336 56550
rect 96380 56058 96436 56060
rect 96460 56058 96516 56060
rect 96540 56058 96596 56060
rect 96620 56058 96676 56060
rect 96380 56006 96426 56058
rect 96426 56006 96436 56058
rect 96460 56006 96490 56058
rect 96490 56006 96502 56058
rect 96502 56006 96516 56058
rect 96540 56006 96554 56058
rect 96554 56006 96566 56058
rect 96566 56006 96596 56058
rect 96620 56006 96630 56058
rect 96630 56006 96676 56058
rect 96380 56004 96436 56006
rect 96460 56004 96516 56006
rect 96540 56004 96596 56006
rect 96620 56004 96676 56006
rect 97262 55800 97318 55856
rect 97446 55800 97502 55856
rect 97040 55514 97096 55516
rect 97120 55514 97176 55516
rect 97200 55514 97256 55516
rect 97280 55514 97336 55516
rect 97040 55462 97086 55514
rect 97086 55462 97096 55514
rect 97120 55462 97150 55514
rect 97150 55462 97162 55514
rect 97162 55462 97176 55514
rect 97200 55462 97214 55514
rect 97214 55462 97226 55514
rect 97226 55462 97256 55514
rect 97280 55462 97290 55514
rect 97290 55462 97336 55514
rect 97040 55460 97096 55462
rect 97120 55460 97176 55462
rect 97200 55460 97256 55462
rect 97280 55460 97336 55462
rect 96380 54970 96436 54972
rect 96460 54970 96516 54972
rect 96540 54970 96596 54972
rect 96620 54970 96676 54972
rect 96380 54918 96426 54970
rect 96426 54918 96436 54970
rect 96460 54918 96490 54970
rect 96490 54918 96502 54970
rect 96502 54918 96516 54970
rect 96540 54918 96554 54970
rect 96554 54918 96566 54970
rect 96566 54918 96596 54970
rect 96620 54918 96630 54970
rect 96630 54918 96676 54970
rect 96380 54916 96436 54918
rect 96460 54916 96516 54918
rect 96540 54916 96596 54918
rect 96620 54916 96676 54918
rect 97262 54712 97318 54768
rect 97446 54476 97448 54496
rect 97448 54476 97500 54496
rect 97500 54476 97502 54496
rect 97446 54440 97502 54476
rect 97040 54426 97096 54428
rect 97120 54426 97176 54428
rect 97200 54426 97256 54428
rect 97280 54426 97336 54428
rect 97040 54374 97086 54426
rect 97086 54374 97096 54426
rect 97120 54374 97150 54426
rect 97150 54374 97162 54426
rect 97162 54374 97176 54426
rect 97200 54374 97214 54426
rect 97214 54374 97226 54426
rect 97226 54374 97256 54426
rect 97280 54374 97290 54426
rect 97290 54374 97336 54426
rect 97040 54372 97096 54374
rect 97120 54372 97176 54374
rect 97200 54372 97256 54374
rect 97280 54372 97336 54374
rect 96380 53882 96436 53884
rect 96460 53882 96516 53884
rect 96540 53882 96596 53884
rect 96620 53882 96676 53884
rect 96380 53830 96426 53882
rect 96426 53830 96436 53882
rect 96460 53830 96490 53882
rect 96490 53830 96502 53882
rect 96502 53830 96516 53882
rect 96540 53830 96554 53882
rect 96554 53830 96566 53882
rect 96566 53830 96596 53882
rect 96620 53830 96630 53882
rect 96630 53830 96676 53882
rect 96380 53828 96436 53830
rect 96460 53828 96516 53830
rect 96540 53828 96596 53830
rect 96620 53828 96676 53830
rect 97446 53760 97502 53816
rect 97262 53624 97318 53680
rect 97040 53338 97096 53340
rect 97120 53338 97176 53340
rect 97200 53338 97256 53340
rect 97280 53338 97336 53340
rect 97040 53286 97086 53338
rect 97086 53286 97096 53338
rect 97120 53286 97150 53338
rect 97150 53286 97162 53338
rect 97162 53286 97176 53338
rect 97200 53286 97214 53338
rect 97214 53286 97226 53338
rect 97226 53286 97256 53338
rect 97280 53286 97290 53338
rect 97290 53286 97336 53338
rect 97040 53284 97096 53286
rect 97120 53284 97176 53286
rect 97200 53284 97256 53286
rect 97280 53284 97336 53286
rect 96380 52794 96436 52796
rect 96460 52794 96516 52796
rect 96540 52794 96596 52796
rect 96620 52794 96676 52796
rect 96380 52742 96426 52794
rect 96426 52742 96436 52794
rect 96460 52742 96490 52794
rect 96490 52742 96502 52794
rect 96502 52742 96516 52794
rect 96540 52742 96554 52794
rect 96554 52742 96566 52794
rect 96566 52742 96596 52794
rect 96620 52742 96630 52794
rect 96630 52742 96676 52794
rect 96380 52740 96436 52742
rect 96460 52740 96516 52742
rect 96540 52740 96596 52742
rect 96620 52740 96676 52742
rect 97040 52250 97096 52252
rect 97120 52250 97176 52252
rect 97200 52250 97256 52252
rect 97280 52250 97336 52252
rect 97040 52198 97086 52250
rect 97086 52198 97096 52250
rect 97120 52198 97150 52250
rect 97150 52198 97162 52250
rect 97162 52198 97176 52250
rect 97200 52198 97214 52250
rect 97214 52198 97226 52250
rect 97226 52198 97256 52250
rect 97280 52198 97290 52250
rect 97290 52198 97336 52250
rect 97040 52196 97096 52198
rect 97120 52196 97176 52198
rect 97200 52196 97256 52198
rect 97280 52196 97336 52198
rect 96380 51706 96436 51708
rect 96460 51706 96516 51708
rect 96540 51706 96596 51708
rect 96620 51706 96676 51708
rect 96380 51654 96426 51706
rect 96426 51654 96436 51706
rect 96460 51654 96490 51706
rect 96490 51654 96502 51706
rect 96502 51654 96516 51706
rect 96540 51654 96554 51706
rect 96554 51654 96566 51706
rect 96566 51654 96596 51706
rect 96620 51654 96630 51706
rect 96630 51654 96676 51706
rect 96380 51652 96436 51654
rect 96460 51652 96516 51654
rect 96540 51652 96596 51654
rect 96620 51652 96676 51654
rect 97040 51162 97096 51164
rect 97120 51162 97176 51164
rect 97200 51162 97256 51164
rect 97280 51162 97336 51164
rect 97040 51110 97086 51162
rect 97086 51110 97096 51162
rect 97120 51110 97150 51162
rect 97150 51110 97162 51162
rect 97162 51110 97176 51162
rect 97200 51110 97214 51162
rect 97214 51110 97226 51162
rect 97226 51110 97256 51162
rect 97280 51110 97290 51162
rect 97290 51110 97336 51162
rect 97040 51108 97096 51110
rect 97120 51108 97176 51110
rect 97200 51108 97256 51110
rect 97280 51108 97336 51110
rect 96380 50618 96436 50620
rect 96460 50618 96516 50620
rect 96540 50618 96596 50620
rect 96620 50618 96676 50620
rect 96380 50566 96426 50618
rect 96426 50566 96436 50618
rect 96460 50566 96490 50618
rect 96490 50566 96502 50618
rect 96502 50566 96516 50618
rect 96540 50566 96554 50618
rect 96554 50566 96566 50618
rect 96566 50566 96596 50618
rect 96620 50566 96630 50618
rect 96630 50566 96676 50618
rect 96380 50564 96436 50566
rect 96460 50564 96516 50566
rect 96540 50564 96596 50566
rect 96620 50564 96676 50566
rect 97040 50074 97096 50076
rect 97120 50074 97176 50076
rect 97200 50074 97256 50076
rect 97280 50074 97336 50076
rect 97040 50022 97086 50074
rect 97086 50022 97096 50074
rect 97120 50022 97150 50074
rect 97150 50022 97162 50074
rect 97162 50022 97176 50074
rect 97200 50022 97214 50074
rect 97214 50022 97226 50074
rect 97226 50022 97256 50074
rect 97280 50022 97290 50074
rect 97290 50022 97336 50074
rect 97040 50020 97096 50022
rect 97120 50020 97176 50022
rect 97200 50020 97256 50022
rect 97280 50020 97336 50022
rect 50848 8608 50904 8664
rect 96380 49530 96436 49532
rect 96460 49530 96516 49532
rect 96540 49530 96596 49532
rect 96620 49530 96676 49532
rect 96380 49478 96426 49530
rect 96426 49478 96436 49530
rect 96460 49478 96490 49530
rect 96490 49478 96502 49530
rect 96502 49478 96516 49530
rect 96540 49478 96554 49530
rect 96554 49478 96566 49530
rect 96566 49478 96596 49530
rect 96620 49478 96630 49530
rect 96630 49478 96676 49530
rect 96380 49476 96436 49478
rect 96460 49476 96516 49478
rect 96540 49476 96596 49478
rect 96620 49476 96676 49478
rect 97040 48986 97096 48988
rect 97120 48986 97176 48988
rect 97200 48986 97256 48988
rect 97280 48986 97336 48988
rect 97040 48934 97086 48986
rect 97086 48934 97096 48986
rect 97120 48934 97150 48986
rect 97150 48934 97162 48986
rect 97162 48934 97176 48986
rect 97200 48934 97214 48986
rect 97214 48934 97226 48986
rect 97226 48934 97256 48986
rect 97280 48934 97290 48986
rect 97290 48934 97336 48986
rect 97040 48932 97096 48934
rect 97120 48932 97176 48934
rect 97200 48932 97256 48934
rect 97280 48932 97336 48934
rect 96380 48442 96436 48444
rect 96460 48442 96516 48444
rect 96540 48442 96596 48444
rect 96620 48442 96676 48444
rect 96380 48390 96426 48442
rect 96426 48390 96436 48442
rect 96460 48390 96490 48442
rect 96490 48390 96502 48442
rect 96502 48390 96516 48442
rect 96540 48390 96554 48442
rect 96554 48390 96566 48442
rect 96566 48390 96596 48442
rect 96620 48390 96630 48442
rect 96630 48390 96676 48442
rect 96380 48388 96436 48390
rect 96460 48388 96516 48390
rect 96540 48388 96596 48390
rect 96620 48388 96676 48390
rect 97040 47898 97096 47900
rect 97120 47898 97176 47900
rect 97200 47898 97256 47900
rect 97280 47898 97336 47900
rect 97040 47846 97086 47898
rect 97086 47846 97096 47898
rect 97120 47846 97150 47898
rect 97150 47846 97162 47898
rect 97162 47846 97176 47898
rect 97200 47846 97214 47898
rect 97214 47846 97226 47898
rect 97226 47846 97256 47898
rect 97280 47846 97290 47898
rect 97290 47846 97336 47898
rect 97040 47844 97096 47846
rect 97120 47844 97176 47846
rect 97200 47844 97256 47846
rect 97280 47844 97336 47846
rect 96380 47354 96436 47356
rect 96460 47354 96516 47356
rect 96540 47354 96596 47356
rect 96620 47354 96676 47356
rect 96380 47302 96426 47354
rect 96426 47302 96436 47354
rect 96460 47302 96490 47354
rect 96490 47302 96502 47354
rect 96502 47302 96516 47354
rect 96540 47302 96554 47354
rect 96554 47302 96566 47354
rect 96566 47302 96596 47354
rect 96620 47302 96630 47354
rect 96630 47302 96676 47354
rect 96380 47300 96436 47302
rect 96460 47300 96516 47302
rect 96540 47300 96596 47302
rect 96620 47300 96676 47302
rect 97040 46810 97096 46812
rect 97120 46810 97176 46812
rect 97200 46810 97256 46812
rect 97280 46810 97336 46812
rect 97040 46758 97086 46810
rect 97086 46758 97096 46810
rect 97120 46758 97150 46810
rect 97150 46758 97162 46810
rect 97162 46758 97176 46810
rect 97200 46758 97214 46810
rect 97214 46758 97226 46810
rect 97226 46758 97256 46810
rect 97280 46758 97290 46810
rect 97290 46758 97336 46810
rect 97040 46756 97096 46758
rect 97120 46756 97176 46758
rect 97200 46756 97256 46758
rect 97280 46756 97336 46758
rect 96380 46266 96436 46268
rect 96460 46266 96516 46268
rect 96540 46266 96596 46268
rect 96620 46266 96676 46268
rect 96380 46214 96426 46266
rect 96426 46214 96436 46266
rect 96460 46214 96490 46266
rect 96490 46214 96502 46266
rect 96502 46214 96516 46266
rect 96540 46214 96554 46266
rect 96554 46214 96566 46266
rect 96566 46214 96596 46266
rect 96620 46214 96630 46266
rect 96630 46214 96676 46266
rect 96380 46212 96436 46214
rect 96460 46212 96516 46214
rect 96540 46212 96596 46214
rect 96620 46212 96676 46214
rect 97040 45722 97096 45724
rect 97120 45722 97176 45724
rect 97200 45722 97256 45724
rect 97280 45722 97336 45724
rect 97040 45670 97086 45722
rect 97086 45670 97096 45722
rect 97120 45670 97150 45722
rect 97150 45670 97162 45722
rect 97162 45670 97176 45722
rect 97200 45670 97214 45722
rect 97214 45670 97226 45722
rect 97226 45670 97256 45722
rect 97280 45670 97290 45722
rect 97290 45670 97336 45722
rect 97040 45668 97096 45670
rect 97120 45668 97176 45670
rect 97200 45668 97256 45670
rect 97280 45668 97336 45670
rect 97538 45600 97594 45656
rect 97446 45328 97502 45384
rect 96380 45178 96436 45180
rect 96460 45178 96516 45180
rect 96540 45178 96596 45180
rect 96620 45178 96676 45180
rect 96380 45126 96426 45178
rect 96426 45126 96436 45178
rect 96460 45126 96490 45178
rect 96490 45126 96502 45178
rect 96502 45126 96516 45178
rect 96540 45126 96554 45178
rect 96554 45126 96566 45178
rect 96566 45126 96596 45178
rect 96620 45126 96630 45178
rect 96630 45126 96676 45178
rect 96380 45124 96436 45126
rect 96460 45124 96516 45126
rect 96540 45124 96596 45126
rect 96620 45124 96676 45126
rect 97040 44634 97096 44636
rect 97120 44634 97176 44636
rect 97200 44634 97256 44636
rect 97280 44634 97336 44636
rect 97040 44582 97086 44634
rect 97086 44582 97096 44634
rect 97120 44582 97150 44634
rect 97150 44582 97162 44634
rect 97162 44582 97176 44634
rect 97200 44582 97214 44634
rect 97214 44582 97226 44634
rect 97226 44582 97256 44634
rect 97280 44582 97290 44634
rect 97290 44582 97336 44634
rect 97040 44580 97096 44582
rect 97120 44580 97176 44582
rect 97200 44580 97256 44582
rect 97280 44580 97336 44582
rect 97354 44260 97410 44296
rect 97354 44240 97356 44260
rect 97356 44240 97408 44260
rect 97408 44240 97410 44260
rect 97538 44240 97594 44296
rect 96380 44090 96436 44092
rect 96460 44090 96516 44092
rect 96540 44090 96596 44092
rect 96620 44090 96676 44092
rect 96380 44038 96426 44090
rect 96426 44038 96436 44090
rect 96460 44038 96490 44090
rect 96490 44038 96502 44090
rect 96502 44038 96516 44090
rect 96540 44038 96554 44090
rect 96554 44038 96566 44090
rect 96566 44038 96596 44090
rect 96620 44038 96630 44090
rect 96630 44038 96676 44090
rect 96380 44036 96436 44038
rect 96460 44036 96516 44038
rect 96540 44036 96596 44038
rect 96620 44036 96676 44038
rect 97040 43546 97096 43548
rect 97120 43546 97176 43548
rect 97200 43546 97256 43548
rect 97280 43546 97336 43548
rect 97040 43494 97086 43546
rect 97086 43494 97096 43546
rect 97120 43494 97150 43546
rect 97150 43494 97162 43546
rect 97162 43494 97176 43546
rect 97200 43494 97214 43546
rect 97214 43494 97226 43546
rect 97226 43494 97256 43546
rect 97280 43494 97290 43546
rect 97290 43494 97336 43546
rect 97040 43492 97096 43494
rect 97120 43492 97176 43494
rect 97200 43492 97256 43494
rect 97280 43492 97336 43494
rect 97354 43172 97410 43208
rect 97354 43152 97356 43172
rect 97356 43152 97408 43172
rect 97408 43152 97410 43172
rect 96380 43002 96436 43004
rect 96460 43002 96516 43004
rect 96540 43002 96596 43004
rect 96620 43002 96676 43004
rect 96380 42950 96426 43002
rect 96426 42950 96436 43002
rect 96460 42950 96490 43002
rect 96490 42950 96502 43002
rect 96502 42950 96516 43002
rect 96540 42950 96554 43002
rect 96554 42950 96566 43002
rect 96566 42950 96596 43002
rect 96620 42950 96630 43002
rect 96630 42950 96676 43002
rect 96380 42948 96436 42950
rect 96460 42948 96516 42950
rect 96540 42948 96596 42950
rect 96620 42948 96676 42950
rect 97538 42880 97594 42936
rect 97040 42458 97096 42460
rect 97120 42458 97176 42460
rect 97200 42458 97256 42460
rect 97280 42458 97336 42460
rect 97040 42406 97086 42458
rect 97086 42406 97096 42458
rect 97120 42406 97150 42458
rect 97150 42406 97162 42458
rect 97162 42406 97176 42458
rect 97200 42406 97214 42458
rect 97214 42406 97226 42458
rect 97226 42406 97256 42458
rect 97280 42406 97290 42458
rect 97290 42406 97336 42458
rect 97040 42404 97096 42406
rect 97120 42404 97176 42406
rect 97200 42404 97256 42406
rect 97280 42404 97336 42406
rect 97538 42200 97594 42256
rect 97446 42064 97502 42120
rect 96380 41914 96436 41916
rect 96460 41914 96516 41916
rect 96540 41914 96596 41916
rect 96620 41914 96676 41916
rect 96380 41862 96426 41914
rect 96426 41862 96436 41914
rect 96460 41862 96490 41914
rect 96490 41862 96502 41914
rect 96502 41862 96516 41914
rect 96540 41862 96554 41914
rect 96554 41862 96566 41914
rect 96566 41862 96596 41914
rect 96620 41862 96630 41914
rect 96630 41862 96676 41914
rect 96380 41860 96436 41862
rect 96460 41860 96516 41862
rect 96540 41860 96596 41862
rect 96620 41860 96676 41862
rect 97040 41370 97096 41372
rect 97120 41370 97176 41372
rect 97200 41370 97256 41372
rect 97280 41370 97336 41372
rect 97040 41318 97086 41370
rect 97086 41318 97096 41370
rect 97120 41318 97150 41370
rect 97150 41318 97162 41370
rect 97162 41318 97176 41370
rect 97200 41318 97214 41370
rect 97214 41318 97226 41370
rect 97226 41318 97256 41370
rect 97280 41318 97290 41370
rect 97290 41318 97336 41370
rect 97040 41316 97096 41318
rect 97120 41316 97176 41318
rect 97200 41316 97256 41318
rect 97280 41316 97336 41318
rect 97354 41112 97410 41168
rect 97538 40840 97594 40896
rect 96380 40826 96436 40828
rect 96460 40826 96516 40828
rect 96540 40826 96596 40828
rect 96620 40826 96676 40828
rect 96380 40774 96426 40826
rect 96426 40774 96436 40826
rect 96460 40774 96490 40826
rect 96490 40774 96502 40826
rect 96502 40774 96516 40826
rect 96540 40774 96554 40826
rect 96554 40774 96566 40826
rect 96566 40774 96596 40826
rect 96620 40774 96630 40826
rect 96630 40774 96676 40826
rect 96380 40772 96436 40774
rect 96460 40772 96516 40774
rect 96540 40772 96596 40774
rect 96620 40772 96676 40774
rect 97040 40282 97096 40284
rect 97120 40282 97176 40284
rect 97200 40282 97256 40284
rect 97280 40282 97336 40284
rect 97040 40230 97086 40282
rect 97086 40230 97096 40282
rect 97120 40230 97150 40282
rect 97150 40230 97162 40282
rect 97162 40230 97176 40282
rect 97200 40230 97214 40282
rect 97214 40230 97226 40282
rect 97226 40230 97256 40282
rect 97280 40230 97290 40282
rect 97290 40230 97336 40282
rect 97040 40228 97096 40230
rect 97120 40228 97176 40230
rect 97200 40228 97256 40230
rect 97280 40228 97336 40230
rect 97538 40160 97594 40216
rect 97446 39888 97502 39944
rect 96380 39738 96436 39740
rect 96460 39738 96516 39740
rect 96540 39738 96596 39740
rect 96620 39738 96676 39740
rect 96380 39686 96426 39738
rect 96426 39686 96436 39738
rect 96460 39686 96490 39738
rect 96490 39686 96502 39738
rect 96502 39686 96516 39738
rect 96540 39686 96554 39738
rect 96554 39686 96566 39738
rect 96566 39686 96596 39738
rect 96620 39686 96630 39738
rect 96630 39686 96676 39738
rect 96380 39684 96436 39686
rect 96460 39684 96516 39686
rect 96540 39684 96596 39686
rect 96620 39684 96676 39686
rect 97040 39194 97096 39196
rect 97120 39194 97176 39196
rect 97200 39194 97256 39196
rect 97280 39194 97336 39196
rect 97040 39142 97086 39194
rect 97086 39142 97096 39194
rect 97120 39142 97150 39194
rect 97150 39142 97162 39194
rect 97162 39142 97176 39194
rect 97200 39142 97214 39194
rect 97214 39142 97226 39194
rect 97226 39142 97256 39194
rect 97280 39142 97290 39194
rect 97290 39142 97336 39194
rect 97040 39140 97096 39142
rect 97120 39140 97176 39142
rect 97200 39140 97256 39142
rect 97280 39140 97336 39142
rect 97354 38936 97410 38992
rect 97538 38800 97594 38856
rect 96380 38650 96436 38652
rect 96460 38650 96516 38652
rect 96540 38650 96596 38652
rect 96620 38650 96676 38652
rect 96380 38598 96426 38650
rect 96426 38598 96436 38650
rect 96460 38598 96490 38650
rect 96490 38598 96502 38650
rect 96502 38598 96516 38650
rect 96540 38598 96554 38650
rect 96554 38598 96566 38650
rect 96566 38598 96596 38650
rect 96620 38598 96630 38650
rect 96630 38598 96676 38650
rect 96380 38596 96436 38598
rect 96460 38596 96516 38598
rect 96540 38596 96596 38598
rect 96620 38596 96676 38598
rect 97040 38106 97096 38108
rect 97120 38106 97176 38108
rect 97200 38106 97256 38108
rect 97280 38106 97336 38108
rect 97040 38054 97086 38106
rect 97086 38054 97096 38106
rect 97120 38054 97150 38106
rect 97150 38054 97162 38106
rect 97162 38054 97176 38106
rect 97200 38054 97214 38106
rect 97214 38054 97226 38106
rect 97226 38054 97256 38106
rect 97280 38054 97290 38106
rect 97290 38054 97336 38106
rect 97040 38052 97096 38054
rect 97120 38052 97176 38054
rect 97200 38052 97256 38054
rect 97280 38052 97336 38054
rect 97354 37848 97410 37904
rect 96380 37562 96436 37564
rect 96460 37562 96516 37564
rect 96540 37562 96596 37564
rect 96620 37562 96676 37564
rect 96380 37510 96426 37562
rect 96426 37510 96436 37562
rect 96460 37510 96490 37562
rect 96490 37510 96502 37562
rect 96502 37510 96516 37562
rect 96540 37510 96554 37562
rect 96554 37510 96566 37562
rect 96566 37510 96596 37562
rect 96620 37510 96630 37562
rect 96630 37510 96676 37562
rect 96380 37508 96436 37510
rect 96460 37508 96516 37510
rect 96540 37508 96596 37510
rect 96620 37508 96676 37510
rect 97538 37440 97594 37496
rect 97040 37018 97096 37020
rect 97120 37018 97176 37020
rect 97200 37018 97256 37020
rect 97280 37018 97336 37020
rect 97040 36966 97086 37018
rect 97086 36966 97096 37018
rect 97120 36966 97150 37018
rect 97150 36966 97162 37018
rect 97162 36966 97176 37018
rect 97200 36966 97214 37018
rect 97214 36966 97226 37018
rect 97226 36966 97256 37018
rect 97280 36966 97290 37018
rect 97290 36966 97336 37018
rect 97040 36964 97096 36966
rect 97120 36964 97176 36966
rect 97200 36964 97256 36966
rect 97280 36964 97336 36966
rect 96618 36760 96674 36816
rect 97446 36760 97502 36816
rect 96380 36474 96436 36476
rect 96460 36474 96516 36476
rect 96540 36474 96596 36476
rect 96620 36474 96676 36476
rect 96380 36422 96426 36474
rect 96426 36422 96436 36474
rect 96460 36422 96490 36474
rect 96490 36422 96502 36474
rect 96502 36422 96516 36474
rect 96540 36422 96554 36474
rect 96554 36422 96566 36474
rect 96566 36422 96596 36474
rect 96620 36422 96630 36474
rect 96630 36422 96676 36474
rect 96380 36420 96436 36422
rect 96460 36420 96516 36422
rect 96540 36420 96596 36422
rect 96620 36420 96676 36422
rect 97040 35930 97096 35932
rect 97120 35930 97176 35932
rect 97200 35930 97256 35932
rect 97280 35930 97336 35932
rect 97040 35878 97086 35930
rect 97086 35878 97096 35930
rect 97120 35878 97150 35930
rect 97150 35878 97162 35930
rect 97162 35878 97176 35930
rect 97200 35878 97214 35930
rect 97214 35878 97226 35930
rect 97226 35878 97256 35930
rect 97280 35878 97290 35930
rect 97290 35878 97336 35930
rect 97040 35876 97096 35878
rect 97120 35876 97176 35878
rect 97200 35876 97256 35878
rect 97280 35876 97336 35878
rect 97354 35672 97410 35728
rect 97538 35400 97594 35456
rect 96380 35386 96436 35388
rect 96460 35386 96516 35388
rect 96540 35386 96596 35388
rect 96620 35386 96676 35388
rect 96380 35334 96426 35386
rect 96426 35334 96436 35386
rect 96460 35334 96490 35386
rect 96490 35334 96502 35386
rect 96502 35334 96516 35386
rect 96540 35334 96554 35386
rect 96554 35334 96566 35386
rect 96566 35334 96596 35386
rect 96620 35334 96630 35386
rect 96630 35334 96676 35386
rect 96380 35332 96436 35334
rect 96460 35332 96516 35334
rect 96540 35332 96596 35334
rect 96620 35332 96676 35334
rect 97040 34842 97096 34844
rect 97120 34842 97176 34844
rect 97200 34842 97256 34844
rect 97280 34842 97336 34844
rect 97040 34790 97086 34842
rect 97086 34790 97096 34842
rect 97120 34790 97150 34842
rect 97150 34790 97162 34842
rect 97162 34790 97176 34842
rect 97200 34790 97214 34842
rect 97214 34790 97226 34842
rect 97226 34790 97256 34842
rect 97280 34790 97290 34842
rect 97290 34790 97336 34842
rect 97040 34788 97096 34790
rect 97120 34788 97176 34790
rect 97200 34788 97256 34790
rect 97280 34788 97336 34790
rect 97538 34720 97594 34776
rect 97446 34448 97502 34504
rect 96380 34298 96436 34300
rect 96460 34298 96516 34300
rect 96540 34298 96596 34300
rect 96620 34298 96676 34300
rect 96380 34246 96426 34298
rect 96426 34246 96436 34298
rect 96460 34246 96490 34298
rect 96490 34246 96502 34298
rect 96502 34246 96516 34298
rect 96540 34246 96554 34298
rect 96554 34246 96566 34298
rect 96566 34246 96596 34298
rect 96620 34246 96630 34298
rect 96630 34246 96676 34298
rect 96380 34244 96436 34246
rect 96460 34244 96516 34246
rect 96540 34244 96596 34246
rect 96620 34244 96676 34246
rect 97040 33754 97096 33756
rect 97120 33754 97176 33756
rect 97200 33754 97256 33756
rect 97280 33754 97336 33756
rect 97040 33702 97086 33754
rect 97086 33702 97096 33754
rect 97120 33702 97150 33754
rect 97150 33702 97162 33754
rect 97162 33702 97176 33754
rect 97200 33702 97214 33754
rect 97214 33702 97226 33754
rect 97226 33702 97256 33754
rect 97280 33702 97290 33754
rect 97290 33702 97336 33754
rect 97040 33700 97096 33702
rect 97120 33700 97176 33702
rect 97200 33700 97256 33702
rect 97280 33700 97336 33702
rect 97354 33496 97410 33552
rect 97538 33360 97594 33416
rect 96380 33210 96436 33212
rect 96460 33210 96516 33212
rect 96540 33210 96596 33212
rect 96620 33210 96676 33212
rect 96380 33158 96426 33210
rect 96426 33158 96436 33210
rect 96460 33158 96490 33210
rect 96490 33158 96502 33210
rect 96502 33158 96516 33210
rect 96540 33158 96554 33210
rect 96554 33158 96566 33210
rect 96566 33158 96596 33210
rect 96620 33158 96630 33210
rect 96630 33158 96676 33210
rect 96380 33156 96436 33158
rect 96460 33156 96516 33158
rect 96540 33156 96596 33158
rect 96620 33156 96676 33158
rect 97040 32666 97096 32668
rect 97120 32666 97176 32668
rect 97200 32666 97256 32668
rect 97280 32666 97336 32668
rect 97040 32614 97086 32666
rect 97086 32614 97096 32666
rect 97120 32614 97150 32666
rect 97150 32614 97162 32666
rect 97162 32614 97176 32666
rect 97200 32614 97214 32666
rect 97214 32614 97226 32666
rect 97226 32614 97256 32666
rect 97280 32614 97290 32666
rect 97290 32614 97336 32666
rect 97040 32612 97096 32614
rect 97120 32612 97176 32614
rect 97200 32612 97256 32614
rect 97280 32612 97336 32614
rect 97262 32444 97264 32464
rect 97264 32444 97316 32464
rect 97316 32444 97318 32464
rect 97262 32408 97318 32444
rect 96380 32122 96436 32124
rect 96460 32122 96516 32124
rect 96540 32122 96596 32124
rect 96620 32122 96676 32124
rect 96380 32070 96426 32122
rect 96426 32070 96436 32122
rect 96460 32070 96490 32122
rect 96490 32070 96502 32122
rect 96502 32070 96516 32122
rect 96540 32070 96554 32122
rect 96554 32070 96566 32122
rect 96566 32070 96596 32122
rect 96620 32070 96630 32122
rect 96630 32070 96676 32122
rect 96380 32068 96436 32070
rect 96460 32068 96516 32070
rect 96540 32068 96596 32070
rect 96620 32068 96676 32070
rect 97446 32000 97502 32056
rect 97040 31578 97096 31580
rect 97120 31578 97176 31580
rect 97200 31578 97256 31580
rect 97280 31578 97336 31580
rect 97040 31526 97086 31578
rect 97086 31526 97096 31578
rect 97120 31526 97150 31578
rect 97150 31526 97162 31578
rect 97162 31526 97176 31578
rect 97200 31526 97214 31578
rect 97214 31526 97226 31578
rect 97226 31526 97256 31578
rect 97280 31526 97290 31578
rect 97290 31526 97336 31578
rect 97040 31524 97096 31526
rect 97120 31524 97176 31526
rect 97200 31524 97256 31526
rect 97280 31524 97336 31526
rect 96618 31320 96674 31376
rect 97538 31320 97594 31376
rect 96380 31034 96436 31036
rect 96460 31034 96516 31036
rect 96540 31034 96596 31036
rect 96620 31034 96676 31036
rect 96380 30982 96426 31034
rect 96426 30982 96436 31034
rect 96460 30982 96490 31034
rect 96490 30982 96502 31034
rect 96502 30982 96516 31034
rect 96540 30982 96554 31034
rect 96554 30982 96566 31034
rect 96566 30982 96596 31034
rect 96620 30982 96630 31034
rect 96630 30982 96676 31034
rect 96380 30980 96436 30982
rect 96460 30980 96516 30982
rect 96540 30980 96596 30982
rect 96620 30980 96676 30982
rect 97040 30490 97096 30492
rect 97120 30490 97176 30492
rect 97200 30490 97256 30492
rect 97280 30490 97336 30492
rect 97040 30438 97086 30490
rect 97086 30438 97096 30490
rect 97120 30438 97150 30490
rect 97150 30438 97162 30490
rect 97162 30438 97176 30490
rect 97200 30438 97214 30490
rect 97214 30438 97226 30490
rect 97226 30438 97256 30490
rect 97280 30438 97290 30490
rect 97290 30438 97336 30490
rect 97040 30436 97096 30438
rect 97120 30436 97176 30438
rect 97200 30436 97256 30438
rect 97280 30436 97336 30438
rect 97262 30252 97318 30288
rect 97262 30232 97264 30252
rect 97264 30232 97316 30252
rect 97316 30232 97318 30252
rect 97538 29960 97594 30016
rect 96380 29946 96436 29948
rect 96460 29946 96516 29948
rect 96540 29946 96596 29948
rect 96620 29946 96676 29948
rect 96380 29894 96426 29946
rect 96426 29894 96436 29946
rect 96460 29894 96490 29946
rect 96490 29894 96502 29946
rect 96502 29894 96516 29946
rect 96540 29894 96554 29946
rect 96554 29894 96566 29946
rect 96566 29894 96596 29946
rect 96620 29894 96630 29946
rect 96630 29894 96676 29946
rect 96380 29892 96436 29894
rect 96460 29892 96516 29894
rect 96540 29892 96596 29894
rect 96620 29892 96676 29894
rect 97040 29402 97096 29404
rect 97120 29402 97176 29404
rect 97200 29402 97256 29404
rect 97280 29402 97336 29404
rect 97040 29350 97086 29402
rect 97086 29350 97096 29402
rect 97120 29350 97150 29402
rect 97150 29350 97162 29402
rect 97162 29350 97176 29402
rect 97200 29350 97214 29402
rect 97214 29350 97226 29402
rect 97226 29350 97256 29402
rect 97280 29350 97290 29402
rect 97290 29350 97336 29402
rect 97040 29348 97096 29350
rect 97120 29348 97176 29350
rect 97200 29348 97256 29350
rect 97280 29348 97336 29350
rect 97538 29280 97594 29336
rect 97446 29144 97502 29200
rect 96380 28858 96436 28860
rect 96460 28858 96516 28860
rect 96540 28858 96596 28860
rect 96620 28858 96676 28860
rect 96380 28806 96426 28858
rect 96426 28806 96436 28858
rect 96460 28806 96490 28858
rect 96490 28806 96502 28858
rect 96502 28806 96516 28858
rect 96540 28806 96554 28858
rect 96554 28806 96566 28858
rect 96566 28806 96596 28858
rect 96620 28806 96630 28858
rect 96630 28806 96676 28858
rect 96380 28804 96436 28806
rect 96460 28804 96516 28806
rect 96540 28804 96596 28806
rect 96620 28804 96676 28806
rect 97040 28314 97096 28316
rect 97120 28314 97176 28316
rect 97200 28314 97256 28316
rect 97280 28314 97336 28316
rect 97040 28262 97086 28314
rect 97086 28262 97096 28314
rect 97120 28262 97150 28314
rect 97150 28262 97162 28314
rect 97162 28262 97176 28314
rect 97200 28262 97214 28314
rect 97214 28262 97226 28314
rect 97226 28262 97256 28314
rect 97280 28262 97290 28314
rect 97290 28262 97336 28314
rect 97040 28260 97096 28262
rect 97120 28260 97176 28262
rect 97200 28260 97256 28262
rect 97280 28260 97336 28262
rect 97262 28076 97318 28112
rect 97262 28056 97264 28076
rect 97264 28056 97316 28076
rect 97316 28056 97318 28076
rect 97446 27940 97502 27976
rect 97446 27920 97448 27940
rect 97448 27920 97500 27940
rect 97500 27920 97502 27940
rect 96380 27770 96436 27772
rect 96460 27770 96516 27772
rect 96540 27770 96596 27772
rect 96620 27770 96676 27772
rect 96380 27718 96426 27770
rect 96426 27718 96436 27770
rect 96460 27718 96490 27770
rect 96490 27718 96502 27770
rect 96502 27718 96516 27770
rect 96540 27718 96554 27770
rect 96554 27718 96566 27770
rect 96566 27718 96596 27770
rect 96620 27718 96630 27770
rect 96630 27718 96676 27770
rect 96380 27716 96436 27718
rect 96460 27716 96516 27718
rect 96540 27716 96596 27718
rect 96620 27716 96676 27718
rect 97040 27226 97096 27228
rect 97120 27226 97176 27228
rect 97200 27226 97256 27228
rect 97280 27226 97336 27228
rect 97040 27174 97086 27226
rect 97086 27174 97096 27226
rect 97120 27174 97150 27226
rect 97150 27174 97162 27226
rect 97162 27174 97176 27226
rect 97200 27174 97214 27226
rect 97214 27174 97226 27226
rect 97226 27174 97256 27226
rect 97280 27174 97290 27226
rect 97290 27174 97336 27226
rect 97040 27172 97096 27174
rect 97120 27172 97176 27174
rect 97200 27172 97256 27174
rect 97280 27172 97336 27174
rect 97262 26988 97318 27024
rect 97262 26968 97264 26988
rect 97264 26968 97316 26988
rect 97316 26968 97318 26988
rect 96380 26682 96436 26684
rect 96460 26682 96516 26684
rect 96540 26682 96596 26684
rect 96620 26682 96676 26684
rect 96380 26630 96426 26682
rect 96426 26630 96436 26682
rect 96460 26630 96490 26682
rect 96490 26630 96502 26682
rect 96502 26630 96516 26682
rect 96540 26630 96554 26682
rect 96554 26630 96566 26682
rect 96566 26630 96596 26682
rect 96620 26630 96630 26682
rect 96630 26630 96676 26682
rect 96380 26628 96436 26630
rect 96460 26628 96516 26630
rect 96540 26628 96596 26630
rect 96620 26628 96676 26630
rect 97446 26560 97502 26616
rect 97040 26138 97096 26140
rect 97120 26138 97176 26140
rect 97200 26138 97256 26140
rect 97280 26138 97336 26140
rect 97040 26086 97086 26138
rect 97086 26086 97096 26138
rect 97120 26086 97150 26138
rect 97150 26086 97162 26138
rect 97162 26086 97176 26138
rect 97200 26086 97214 26138
rect 97214 26086 97226 26138
rect 97226 26086 97256 26138
rect 97280 26086 97290 26138
rect 97290 26086 97336 26138
rect 97040 26084 97096 26086
rect 97120 26084 97176 26086
rect 97200 26084 97256 26086
rect 97280 26084 97336 26086
rect 96894 25880 96950 25936
rect 97446 25880 97502 25936
rect 96380 25594 96436 25596
rect 96460 25594 96516 25596
rect 96540 25594 96596 25596
rect 96620 25594 96676 25596
rect 96380 25542 96426 25594
rect 96426 25542 96436 25594
rect 96460 25542 96490 25594
rect 96490 25542 96502 25594
rect 96502 25542 96516 25594
rect 96540 25542 96554 25594
rect 96554 25542 96566 25594
rect 96566 25542 96596 25594
rect 96620 25542 96630 25594
rect 96630 25542 96676 25594
rect 96380 25540 96436 25542
rect 96460 25540 96516 25542
rect 96540 25540 96596 25542
rect 96620 25540 96676 25542
rect 97040 25050 97096 25052
rect 97120 25050 97176 25052
rect 97200 25050 97256 25052
rect 97280 25050 97336 25052
rect 97040 24998 97086 25050
rect 97086 24998 97096 25050
rect 97120 24998 97150 25050
rect 97150 24998 97162 25050
rect 97162 24998 97176 25050
rect 97200 24998 97214 25050
rect 97214 24998 97226 25050
rect 97226 24998 97256 25050
rect 97280 24998 97290 25050
rect 97290 24998 97336 25050
rect 97040 24996 97096 24998
rect 97120 24996 97176 24998
rect 97200 24996 97256 24998
rect 97280 24996 97336 24998
rect 97262 24812 97318 24848
rect 97262 24792 97264 24812
rect 97264 24792 97316 24812
rect 97316 24792 97318 24812
rect 97446 24556 97448 24576
rect 97448 24556 97500 24576
rect 97500 24556 97502 24576
rect 97446 24520 97502 24556
rect 96380 24506 96436 24508
rect 96460 24506 96516 24508
rect 96540 24506 96596 24508
rect 96620 24506 96676 24508
rect 96380 24454 96426 24506
rect 96426 24454 96436 24506
rect 96460 24454 96490 24506
rect 96490 24454 96502 24506
rect 96502 24454 96516 24506
rect 96540 24454 96554 24506
rect 96554 24454 96566 24506
rect 96566 24454 96596 24506
rect 96620 24454 96630 24506
rect 96630 24454 96676 24506
rect 96380 24452 96436 24454
rect 96460 24452 96516 24454
rect 96540 24452 96596 24454
rect 96620 24452 96676 24454
rect 97040 23962 97096 23964
rect 97120 23962 97176 23964
rect 97200 23962 97256 23964
rect 97280 23962 97336 23964
rect 97040 23910 97086 23962
rect 97086 23910 97096 23962
rect 97120 23910 97150 23962
rect 97150 23910 97162 23962
rect 97162 23910 97176 23962
rect 97200 23910 97214 23962
rect 97214 23910 97226 23962
rect 97226 23910 97256 23962
rect 97280 23910 97290 23962
rect 97290 23910 97336 23962
rect 97040 23908 97096 23910
rect 97120 23908 97176 23910
rect 97200 23908 97256 23910
rect 97280 23908 97336 23910
rect 97446 23840 97502 23896
rect 96618 23704 96674 23760
rect 96380 23418 96436 23420
rect 96460 23418 96516 23420
rect 96540 23418 96596 23420
rect 96620 23418 96676 23420
rect 96380 23366 96426 23418
rect 96426 23366 96436 23418
rect 96460 23366 96490 23418
rect 96490 23366 96502 23418
rect 96502 23366 96516 23418
rect 96540 23366 96554 23418
rect 96554 23366 96566 23418
rect 96566 23366 96596 23418
rect 96620 23366 96630 23418
rect 96630 23366 96676 23418
rect 96380 23364 96436 23366
rect 96460 23364 96516 23366
rect 96540 23364 96596 23366
rect 96620 23364 96676 23366
rect 97040 22874 97096 22876
rect 97120 22874 97176 22876
rect 97200 22874 97256 22876
rect 97280 22874 97336 22876
rect 97040 22822 97086 22874
rect 97086 22822 97096 22874
rect 97120 22822 97150 22874
rect 97150 22822 97162 22874
rect 97162 22822 97176 22874
rect 97200 22822 97214 22874
rect 97214 22822 97226 22874
rect 97226 22822 97256 22874
rect 97280 22822 97290 22874
rect 97290 22822 97336 22874
rect 97040 22820 97096 22822
rect 97120 22820 97176 22822
rect 97200 22820 97256 22822
rect 97280 22820 97336 22822
rect 97262 22636 97318 22672
rect 97262 22616 97264 22636
rect 97264 22616 97316 22636
rect 97316 22616 97318 22636
rect 97446 22500 97502 22536
rect 97446 22480 97448 22500
rect 97448 22480 97500 22500
rect 97500 22480 97502 22500
rect 96380 22330 96436 22332
rect 96460 22330 96516 22332
rect 96540 22330 96596 22332
rect 96620 22330 96676 22332
rect 96380 22278 96426 22330
rect 96426 22278 96436 22330
rect 96460 22278 96490 22330
rect 96490 22278 96502 22330
rect 96502 22278 96516 22330
rect 96540 22278 96554 22330
rect 96554 22278 96566 22330
rect 96566 22278 96596 22330
rect 96620 22278 96630 22330
rect 96630 22278 96676 22330
rect 96380 22276 96436 22278
rect 96460 22276 96516 22278
rect 96540 22276 96596 22278
rect 96620 22276 96676 22278
rect 97040 21786 97096 21788
rect 97120 21786 97176 21788
rect 97200 21786 97256 21788
rect 97280 21786 97336 21788
rect 97040 21734 97086 21786
rect 97086 21734 97096 21786
rect 97120 21734 97150 21786
rect 97150 21734 97162 21786
rect 97162 21734 97176 21786
rect 97200 21734 97214 21786
rect 97214 21734 97226 21786
rect 97226 21734 97256 21786
rect 97280 21734 97290 21786
rect 97290 21734 97336 21786
rect 97040 21732 97096 21734
rect 97120 21732 97176 21734
rect 97200 21732 97256 21734
rect 97280 21732 97336 21734
rect 97262 21548 97318 21584
rect 97262 21528 97264 21548
rect 97264 21528 97316 21548
rect 97316 21528 97318 21548
rect 96380 21242 96436 21244
rect 96460 21242 96516 21244
rect 96540 21242 96596 21244
rect 96620 21242 96676 21244
rect 96380 21190 96426 21242
rect 96426 21190 96436 21242
rect 96460 21190 96490 21242
rect 96490 21190 96502 21242
rect 96502 21190 96516 21242
rect 96540 21190 96554 21242
rect 96554 21190 96566 21242
rect 96566 21190 96596 21242
rect 96620 21190 96630 21242
rect 96630 21190 96676 21242
rect 96380 21188 96436 21190
rect 96460 21188 96516 21190
rect 96540 21188 96596 21190
rect 96620 21188 96676 21190
rect 97446 21120 97502 21176
rect 97040 20698 97096 20700
rect 97120 20698 97176 20700
rect 97200 20698 97256 20700
rect 97280 20698 97336 20700
rect 97040 20646 97086 20698
rect 97086 20646 97096 20698
rect 97120 20646 97150 20698
rect 97150 20646 97162 20698
rect 97162 20646 97176 20698
rect 97200 20646 97214 20698
rect 97214 20646 97226 20698
rect 97226 20646 97256 20698
rect 97280 20646 97290 20698
rect 97290 20646 97336 20698
rect 97040 20644 97096 20646
rect 97120 20644 97176 20646
rect 97200 20644 97256 20646
rect 97280 20644 97336 20646
rect 96618 20440 96674 20496
rect 97446 20440 97502 20496
rect 96380 20154 96436 20156
rect 96460 20154 96516 20156
rect 96540 20154 96596 20156
rect 96620 20154 96676 20156
rect 96380 20102 96426 20154
rect 96426 20102 96436 20154
rect 96460 20102 96490 20154
rect 96490 20102 96502 20154
rect 96502 20102 96516 20154
rect 96540 20102 96554 20154
rect 96554 20102 96566 20154
rect 96566 20102 96596 20154
rect 96620 20102 96630 20154
rect 96630 20102 96676 20154
rect 96380 20100 96436 20102
rect 96460 20100 96516 20102
rect 96540 20100 96596 20102
rect 96620 20100 96676 20102
rect 97040 19610 97096 19612
rect 97120 19610 97176 19612
rect 97200 19610 97256 19612
rect 97280 19610 97336 19612
rect 97040 19558 97086 19610
rect 97086 19558 97096 19610
rect 97120 19558 97150 19610
rect 97150 19558 97162 19610
rect 97162 19558 97176 19610
rect 97200 19558 97214 19610
rect 97214 19558 97226 19610
rect 97226 19558 97256 19610
rect 97280 19558 97290 19610
rect 97290 19558 97336 19610
rect 97040 19556 97096 19558
rect 97120 19556 97176 19558
rect 97200 19556 97256 19558
rect 97280 19556 97336 19558
rect 97262 19216 97318 19272
rect 97446 19080 97502 19136
rect 96380 19066 96436 19068
rect 96460 19066 96516 19068
rect 96540 19066 96596 19068
rect 96620 19066 96676 19068
rect 96380 19014 96426 19066
rect 96426 19014 96436 19066
rect 96460 19014 96490 19066
rect 96490 19014 96502 19066
rect 96502 19014 96516 19066
rect 96540 19014 96554 19066
rect 96554 19014 96566 19066
rect 96566 19014 96596 19066
rect 96620 19014 96630 19066
rect 96630 19014 96676 19066
rect 96380 19012 96436 19014
rect 96460 19012 96516 19014
rect 96540 19012 96596 19014
rect 96620 19012 96676 19014
rect 97040 18522 97096 18524
rect 97120 18522 97176 18524
rect 97200 18522 97256 18524
rect 97280 18522 97336 18524
rect 97040 18470 97086 18522
rect 97086 18470 97096 18522
rect 97120 18470 97150 18522
rect 97150 18470 97162 18522
rect 97162 18470 97176 18522
rect 97200 18470 97214 18522
rect 97214 18470 97226 18522
rect 97226 18470 97256 18522
rect 97280 18470 97290 18522
rect 97290 18470 97336 18522
rect 97040 18468 97096 18470
rect 97120 18468 97176 18470
rect 97200 18468 97256 18470
rect 97280 18468 97336 18470
rect 97446 18400 97502 18456
rect 96618 18264 96674 18320
rect 96380 17978 96436 17980
rect 96460 17978 96516 17980
rect 96540 17978 96596 17980
rect 96620 17978 96676 17980
rect 96380 17926 96426 17978
rect 96426 17926 96436 17978
rect 96460 17926 96490 17978
rect 96490 17926 96502 17978
rect 96502 17926 96516 17978
rect 96540 17926 96554 17978
rect 96554 17926 96566 17978
rect 96566 17926 96596 17978
rect 96620 17926 96630 17978
rect 96630 17926 96676 17978
rect 96380 17924 96436 17926
rect 96460 17924 96516 17926
rect 96540 17924 96596 17926
rect 96620 17924 96676 17926
rect 97040 17434 97096 17436
rect 97120 17434 97176 17436
rect 97200 17434 97256 17436
rect 97280 17434 97336 17436
rect 97040 17382 97086 17434
rect 97086 17382 97096 17434
rect 97120 17382 97150 17434
rect 97150 17382 97162 17434
rect 97162 17382 97176 17434
rect 97200 17382 97214 17434
rect 97214 17382 97226 17434
rect 97226 17382 97256 17434
rect 97280 17382 97290 17434
rect 97290 17382 97336 17434
rect 97040 17380 97096 17382
rect 97120 17380 97176 17382
rect 97200 17380 97256 17382
rect 97280 17380 97336 17382
rect 97262 17196 97318 17232
rect 97262 17176 97264 17196
rect 97264 17176 97316 17196
rect 97316 17176 97318 17196
rect 97446 17060 97502 17096
rect 97446 17040 97448 17060
rect 97448 17040 97500 17060
rect 97500 17040 97502 17060
rect 96380 16890 96436 16892
rect 96460 16890 96516 16892
rect 96540 16890 96596 16892
rect 96620 16890 96676 16892
rect 96380 16838 96426 16890
rect 96426 16838 96436 16890
rect 96460 16838 96490 16890
rect 96490 16838 96502 16890
rect 96502 16838 96516 16890
rect 96540 16838 96554 16890
rect 96554 16838 96566 16890
rect 96566 16838 96596 16890
rect 96620 16838 96630 16890
rect 96630 16838 96676 16890
rect 96380 16836 96436 16838
rect 96460 16836 96516 16838
rect 96540 16836 96596 16838
rect 96620 16836 96676 16838
rect 97040 16346 97096 16348
rect 97120 16346 97176 16348
rect 97200 16346 97256 16348
rect 97280 16346 97336 16348
rect 97040 16294 97086 16346
rect 97086 16294 97096 16346
rect 97120 16294 97150 16346
rect 97150 16294 97162 16346
rect 97162 16294 97176 16346
rect 97200 16294 97214 16346
rect 97214 16294 97226 16346
rect 97226 16294 97256 16346
rect 97280 16294 97290 16346
rect 97290 16294 97336 16346
rect 97040 16292 97096 16294
rect 97120 16292 97176 16294
rect 97200 16292 97256 16294
rect 97280 16292 97336 16294
rect 97262 16108 97318 16144
rect 97262 16088 97264 16108
rect 97264 16088 97316 16108
rect 97316 16088 97318 16108
rect 96380 15802 96436 15804
rect 96460 15802 96516 15804
rect 96540 15802 96596 15804
rect 96620 15802 96676 15804
rect 96380 15750 96426 15802
rect 96426 15750 96436 15802
rect 96460 15750 96490 15802
rect 96490 15750 96502 15802
rect 96502 15750 96516 15802
rect 96540 15750 96554 15802
rect 96554 15750 96566 15802
rect 96566 15750 96596 15802
rect 96620 15750 96630 15802
rect 96630 15750 96676 15802
rect 96380 15748 96436 15750
rect 96460 15748 96516 15750
rect 96540 15748 96596 15750
rect 96620 15748 96676 15750
rect 97446 15680 97502 15736
rect 97040 15258 97096 15260
rect 97120 15258 97176 15260
rect 97200 15258 97256 15260
rect 97280 15258 97336 15260
rect 97040 15206 97086 15258
rect 97086 15206 97096 15258
rect 97120 15206 97150 15258
rect 97150 15206 97162 15258
rect 97162 15206 97176 15258
rect 97200 15206 97214 15258
rect 97214 15206 97226 15258
rect 97226 15206 97256 15258
rect 97280 15206 97290 15258
rect 97290 15206 97336 15258
rect 97040 15204 97096 15206
rect 97120 15204 97176 15206
rect 97200 15204 97256 15206
rect 97280 15204 97336 15206
rect 96618 15000 96674 15056
rect 97446 15000 97502 15056
rect 96380 14714 96436 14716
rect 96460 14714 96516 14716
rect 96540 14714 96596 14716
rect 96620 14714 96676 14716
rect 96380 14662 96426 14714
rect 96426 14662 96436 14714
rect 96460 14662 96490 14714
rect 96490 14662 96502 14714
rect 96502 14662 96516 14714
rect 96540 14662 96554 14714
rect 96554 14662 96566 14714
rect 96566 14662 96596 14714
rect 96620 14662 96630 14714
rect 96630 14662 96676 14714
rect 96380 14660 96436 14662
rect 96460 14660 96516 14662
rect 96540 14660 96596 14662
rect 96620 14660 96676 14662
rect 97040 14170 97096 14172
rect 97120 14170 97176 14172
rect 97200 14170 97256 14172
rect 97280 14170 97336 14172
rect 97040 14118 97086 14170
rect 97086 14118 97096 14170
rect 97120 14118 97150 14170
rect 97150 14118 97162 14170
rect 97162 14118 97176 14170
rect 97200 14118 97214 14170
rect 97214 14118 97226 14170
rect 97226 14118 97256 14170
rect 97280 14118 97290 14170
rect 97290 14118 97336 14170
rect 97040 14116 97096 14118
rect 97120 14116 97176 14118
rect 97200 14116 97256 14118
rect 97280 14116 97336 14118
rect 97262 13932 97318 13968
rect 97262 13912 97264 13932
rect 97264 13912 97316 13932
rect 97316 13912 97318 13932
rect 97446 13640 97502 13696
rect 96380 13626 96436 13628
rect 96460 13626 96516 13628
rect 96540 13626 96596 13628
rect 96620 13626 96676 13628
rect 96380 13574 96426 13626
rect 96426 13574 96436 13626
rect 96460 13574 96490 13626
rect 96490 13574 96502 13626
rect 96502 13574 96516 13626
rect 96540 13574 96554 13626
rect 96554 13574 96566 13626
rect 96566 13574 96596 13626
rect 96620 13574 96630 13626
rect 96630 13574 96676 13626
rect 96380 13572 96436 13574
rect 96460 13572 96516 13574
rect 96540 13572 96596 13574
rect 96620 13572 96676 13574
rect 97040 13082 97096 13084
rect 97120 13082 97176 13084
rect 97200 13082 97256 13084
rect 97280 13082 97336 13084
rect 97040 13030 97086 13082
rect 97086 13030 97096 13082
rect 97120 13030 97150 13082
rect 97150 13030 97162 13082
rect 97162 13030 97176 13082
rect 97200 13030 97214 13082
rect 97214 13030 97226 13082
rect 97226 13030 97256 13082
rect 97280 13030 97290 13082
rect 97290 13030 97336 13082
rect 97040 13028 97096 13030
rect 97120 13028 97176 13030
rect 97200 13028 97256 13030
rect 97280 13028 97336 13030
rect 97446 12960 97502 13016
rect 96618 12824 96674 12880
rect 96380 12538 96436 12540
rect 96460 12538 96516 12540
rect 96540 12538 96596 12540
rect 96620 12538 96676 12540
rect 96380 12486 96426 12538
rect 96426 12486 96436 12538
rect 96460 12486 96490 12538
rect 96490 12486 96502 12538
rect 96502 12486 96516 12538
rect 96540 12486 96554 12538
rect 96554 12486 96566 12538
rect 96566 12486 96596 12538
rect 96620 12486 96630 12538
rect 96630 12486 96676 12538
rect 96380 12484 96436 12486
rect 96460 12484 96516 12486
rect 96540 12484 96596 12486
rect 96620 12484 96676 12486
rect 97040 11994 97096 11996
rect 97120 11994 97176 11996
rect 97200 11994 97256 11996
rect 97280 11994 97336 11996
rect 97040 11942 97086 11994
rect 97086 11942 97096 11994
rect 97120 11942 97150 11994
rect 97150 11942 97162 11994
rect 97162 11942 97176 11994
rect 97200 11942 97214 11994
rect 97214 11942 97226 11994
rect 97226 11942 97256 11994
rect 97280 11942 97290 11994
rect 97290 11942 97336 11994
rect 97040 11940 97096 11942
rect 97120 11940 97176 11942
rect 97200 11940 97256 11942
rect 97280 11940 97336 11942
rect 97262 11756 97318 11792
rect 97262 11736 97264 11756
rect 97264 11736 97316 11756
rect 97316 11736 97318 11756
rect 97446 11620 97502 11656
rect 97446 11600 97448 11620
rect 97448 11600 97500 11620
rect 97500 11600 97502 11620
rect 96380 11450 96436 11452
rect 96460 11450 96516 11452
rect 96540 11450 96596 11452
rect 96620 11450 96676 11452
rect 96380 11398 96426 11450
rect 96426 11398 96436 11450
rect 96460 11398 96490 11450
rect 96490 11398 96502 11450
rect 96502 11398 96516 11450
rect 96540 11398 96554 11450
rect 96554 11398 96566 11450
rect 96566 11398 96596 11450
rect 96620 11398 96630 11450
rect 96630 11398 96676 11450
rect 96380 11396 96436 11398
rect 96460 11396 96516 11398
rect 96540 11396 96596 11398
rect 96620 11396 96676 11398
rect 97040 10906 97096 10908
rect 97120 10906 97176 10908
rect 97200 10906 97256 10908
rect 97280 10906 97336 10908
rect 97040 10854 97086 10906
rect 97086 10854 97096 10906
rect 97120 10854 97150 10906
rect 97150 10854 97162 10906
rect 97162 10854 97176 10906
rect 97200 10854 97214 10906
rect 97214 10854 97226 10906
rect 97226 10854 97256 10906
rect 97280 10854 97290 10906
rect 97290 10854 97336 10906
rect 97040 10852 97096 10854
rect 97120 10852 97176 10854
rect 97200 10852 97256 10854
rect 97280 10852 97336 10854
rect 96380 10362 96436 10364
rect 96460 10362 96516 10364
rect 96540 10362 96596 10364
rect 96620 10362 96676 10364
rect 96380 10310 96426 10362
rect 96426 10310 96436 10362
rect 96460 10310 96490 10362
rect 96490 10310 96502 10362
rect 96502 10310 96516 10362
rect 96540 10310 96554 10362
rect 96554 10310 96566 10362
rect 96566 10310 96596 10362
rect 96620 10310 96630 10362
rect 96630 10310 96676 10362
rect 96380 10308 96436 10310
rect 96460 10308 96516 10310
rect 96540 10308 96596 10310
rect 96620 10308 96676 10310
rect 97040 9818 97096 9820
rect 97120 9818 97176 9820
rect 97200 9818 97256 9820
rect 97280 9818 97336 9820
rect 97040 9766 97086 9818
rect 97086 9766 97096 9818
rect 97120 9766 97150 9818
rect 97150 9766 97162 9818
rect 97162 9766 97176 9818
rect 97200 9766 97214 9818
rect 97214 9766 97226 9818
rect 97226 9766 97256 9818
rect 97280 9766 97290 9818
rect 97290 9766 97336 9818
rect 97040 9764 97096 9766
rect 97120 9764 97176 9766
rect 97200 9764 97256 9766
rect 97280 9764 97336 9766
rect 96380 9274 96436 9276
rect 96460 9274 96516 9276
rect 96540 9274 96596 9276
rect 96620 9274 96676 9276
rect 96380 9222 96426 9274
rect 96426 9222 96436 9274
rect 96460 9222 96490 9274
rect 96490 9222 96502 9274
rect 96502 9222 96516 9274
rect 96540 9222 96554 9274
rect 96554 9222 96566 9274
rect 96566 9222 96596 9274
rect 96620 9222 96630 9274
rect 96630 9222 96676 9274
rect 96380 9220 96436 9222
rect 96460 9220 96516 9222
rect 96540 9220 96596 9222
rect 96620 9220 96676 9222
rect 97040 8730 97096 8732
rect 97120 8730 97176 8732
rect 97200 8730 97256 8732
rect 97280 8730 97336 8732
rect 97040 8678 97086 8730
rect 97086 8678 97096 8730
rect 97120 8678 97150 8730
rect 97150 8678 97162 8730
rect 97162 8678 97176 8730
rect 97200 8678 97214 8730
rect 97214 8678 97226 8730
rect 97226 8678 97256 8730
rect 97280 8678 97290 8730
rect 97290 8678 97336 8730
rect 97040 8676 97096 8678
rect 97120 8676 97176 8678
rect 97200 8676 97256 8678
rect 97280 8676 97336 8678
rect 97538 8200 97594 8256
rect 96380 8186 96436 8188
rect 96460 8186 96516 8188
rect 96540 8186 96596 8188
rect 96620 8186 96676 8188
rect 65660 6010 65716 6012
rect 65740 6010 65796 6012
rect 65820 6010 65876 6012
rect 65900 6010 65956 6012
rect 65660 5958 65706 6010
rect 65706 5958 65716 6010
rect 65740 5958 65770 6010
rect 65770 5958 65782 6010
rect 65782 5958 65796 6010
rect 65820 5958 65834 6010
rect 65834 5958 65846 6010
rect 65846 5958 65876 6010
rect 65900 5958 65910 6010
rect 65910 5958 65956 6010
rect 65660 5956 65716 5958
rect 65740 5956 65796 5958
rect 65820 5956 65876 5958
rect 65900 5956 65956 5958
rect 66320 5466 66376 5468
rect 66400 5466 66456 5468
rect 66480 5466 66536 5468
rect 66560 5466 66616 5468
rect 66320 5414 66366 5466
rect 66366 5414 66376 5466
rect 66400 5414 66430 5466
rect 66430 5414 66442 5466
rect 66442 5414 66456 5466
rect 66480 5414 66494 5466
rect 66494 5414 66506 5466
rect 66506 5414 66536 5466
rect 66560 5414 66570 5466
rect 66570 5414 66616 5466
rect 66320 5412 66376 5414
rect 66400 5412 66456 5414
rect 66480 5412 66536 5414
rect 66560 5412 66616 5414
rect 65660 4922 65716 4924
rect 65740 4922 65796 4924
rect 65820 4922 65876 4924
rect 65900 4922 65956 4924
rect 65660 4870 65706 4922
rect 65706 4870 65716 4922
rect 65740 4870 65770 4922
rect 65770 4870 65782 4922
rect 65782 4870 65796 4922
rect 65820 4870 65834 4922
rect 65834 4870 65846 4922
rect 65846 4870 65876 4922
rect 65900 4870 65910 4922
rect 65910 4870 65956 4922
rect 65660 4868 65716 4870
rect 65740 4868 65796 4870
rect 65820 4868 65876 4870
rect 65900 4868 65956 4870
rect 66320 4378 66376 4380
rect 66400 4378 66456 4380
rect 66480 4378 66536 4380
rect 66560 4378 66616 4380
rect 66320 4326 66366 4378
rect 66366 4326 66376 4378
rect 66400 4326 66430 4378
rect 66430 4326 66442 4378
rect 66442 4326 66456 4378
rect 66480 4326 66494 4378
rect 66494 4326 66506 4378
rect 66506 4326 66536 4378
rect 66560 4326 66570 4378
rect 66570 4326 66616 4378
rect 66320 4324 66376 4326
rect 66400 4324 66456 4326
rect 66480 4324 66536 4326
rect 66560 4324 66616 4326
rect 65660 3834 65716 3836
rect 65740 3834 65796 3836
rect 65820 3834 65876 3836
rect 65900 3834 65956 3836
rect 65660 3782 65706 3834
rect 65706 3782 65716 3834
rect 65740 3782 65770 3834
rect 65770 3782 65782 3834
rect 65782 3782 65796 3834
rect 65820 3782 65834 3834
rect 65834 3782 65846 3834
rect 65846 3782 65876 3834
rect 65900 3782 65910 3834
rect 65910 3782 65956 3834
rect 65660 3780 65716 3782
rect 65740 3780 65796 3782
rect 65820 3780 65876 3782
rect 65900 3780 65956 3782
rect 66320 3290 66376 3292
rect 66400 3290 66456 3292
rect 66480 3290 66536 3292
rect 66560 3290 66616 3292
rect 66320 3238 66366 3290
rect 66366 3238 66376 3290
rect 66400 3238 66430 3290
rect 66430 3238 66442 3290
rect 66442 3238 66456 3290
rect 66480 3238 66494 3290
rect 66494 3238 66506 3290
rect 66506 3238 66536 3290
rect 66560 3238 66570 3290
rect 66570 3238 66616 3290
rect 66320 3236 66376 3238
rect 66400 3236 66456 3238
rect 66480 3236 66536 3238
rect 66560 3236 66616 3238
rect 65660 2746 65716 2748
rect 65740 2746 65796 2748
rect 65820 2746 65876 2748
rect 65900 2746 65956 2748
rect 65660 2694 65706 2746
rect 65706 2694 65716 2746
rect 65740 2694 65770 2746
rect 65770 2694 65782 2746
rect 65782 2694 65796 2746
rect 65820 2694 65834 2746
rect 65834 2694 65846 2746
rect 65846 2694 65876 2746
rect 65900 2694 65910 2746
rect 65910 2694 65956 2746
rect 65660 2692 65716 2694
rect 65740 2692 65796 2694
rect 65820 2692 65876 2694
rect 65900 2692 65956 2694
rect 96380 8134 96426 8186
rect 96426 8134 96436 8186
rect 96460 8134 96490 8186
rect 96490 8134 96502 8186
rect 96502 8134 96516 8186
rect 96540 8134 96554 8186
rect 96554 8134 96566 8186
rect 96566 8134 96596 8186
rect 96620 8134 96630 8186
rect 96630 8134 96676 8186
rect 96380 8132 96436 8134
rect 96460 8132 96516 8134
rect 96540 8132 96596 8134
rect 96620 8132 96676 8134
rect 97040 7642 97096 7644
rect 97120 7642 97176 7644
rect 97200 7642 97256 7644
rect 97280 7642 97336 7644
rect 97040 7590 97086 7642
rect 97086 7590 97096 7642
rect 97120 7590 97150 7642
rect 97150 7590 97162 7642
rect 97162 7590 97176 7642
rect 97200 7590 97214 7642
rect 97214 7590 97226 7642
rect 97226 7590 97256 7642
rect 97280 7590 97290 7642
rect 97290 7590 97336 7642
rect 97040 7588 97096 7590
rect 97120 7588 97176 7590
rect 97200 7588 97256 7590
rect 97280 7588 97336 7590
rect 96380 7098 96436 7100
rect 96460 7098 96516 7100
rect 96540 7098 96596 7100
rect 96620 7098 96676 7100
rect 96380 7046 96426 7098
rect 96426 7046 96436 7098
rect 96460 7046 96490 7098
rect 96490 7046 96502 7098
rect 96502 7046 96516 7098
rect 96540 7046 96554 7098
rect 96554 7046 96566 7098
rect 96566 7046 96596 7098
rect 96620 7046 96630 7098
rect 96630 7046 96676 7098
rect 96380 7044 96436 7046
rect 96460 7044 96516 7046
rect 96540 7044 96596 7046
rect 96620 7044 96676 7046
rect 97040 6554 97096 6556
rect 97120 6554 97176 6556
rect 97200 6554 97256 6556
rect 97280 6554 97336 6556
rect 97040 6502 97086 6554
rect 97086 6502 97096 6554
rect 97120 6502 97150 6554
rect 97150 6502 97162 6554
rect 97162 6502 97176 6554
rect 97200 6502 97214 6554
rect 97214 6502 97226 6554
rect 97226 6502 97256 6554
rect 97280 6502 97290 6554
rect 97290 6502 97336 6554
rect 97040 6500 97096 6502
rect 97120 6500 97176 6502
rect 97200 6500 97256 6502
rect 97280 6500 97336 6502
rect 96380 6010 96436 6012
rect 96460 6010 96516 6012
rect 96540 6010 96596 6012
rect 96620 6010 96676 6012
rect 96380 5958 96426 6010
rect 96426 5958 96436 6010
rect 96460 5958 96490 6010
rect 96490 5958 96502 6010
rect 96502 5958 96516 6010
rect 96540 5958 96554 6010
rect 96554 5958 96566 6010
rect 96566 5958 96596 6010
rect 96620 5958 96630 6010
rect 96630 5958 96676 6010
rect 96380 5956 96436 5958
rect 96460 5956 96516 5958
rect 96540 5956 96596 5958
rect 96620 5956 96676 5958
rect 97040 5466 97096 5468
rect 97120 5466 97176 5468
rect 97200 5466 97256 5468
rect 97280 5466 97336 5468
rect 97040 5414 97086 5466
rect 97086 5414 97096 5466
rect 97120 5414 97150 5466
rect 97150 5414 97162 5466
rect 97162 5414 97176 5466
rect 97200 5414 97214 5466
rect 97214 5414 97226 5466
rect 97226 5414 97256 5466
rect 97280 5414 97290 5466
rect 97290 5414 97336 5466
rect 97040 5412 97096 5414
rect 97120 5412 97176 5414
rect 97200 5412 97256 5414
rect 97280 5412 97336 5414
rect 96380 4922 96436 4924
rect 96460 4922 96516 4924
rect 96540 4922 96596 4924
rect 96620 4922 96676 4924
rect 96380 4870 96426 4922
rect 96426 4870 96436 4922
rect 96460 4870 96490 4922
rect 96490 4870 96502 4922
rect 96502 4870 96516 4922
rect 96540 4870 96554 4922
rect 96554 4870 96566 4922
rect 96566 4870 96596 4922
rect 96620 4870 96630 4922
rect 96630 4870 96676 4922
rect 96380 4868 96436 4870
rect 96460 4868 96516 4870
rect 96540 4868 96596 4870
rect 96620 4868 96676 4870
rect 97040 4378 97096 4380
rect 97120 4378 97176 4380
rect 97200 4378 97256 4380
rect 97280 4378 97336 4380
rect 97040 4326 97086 4378
rect 97086 4326 97096 4378
rect 97120 4326 97150 4378
rect 97150 4326 97162 4378
rect 97162 4326 97176 4378
rect 97200 4326 97214 4378
rect 97214 4326 97226 4378
rect 97226 4326 97256 4378
rect 97280 4326 97290 4378
rect 97290 4326 97336 4378
rect 97040 4324 97096 4326
rect 97120 4324 97176 4326
rect 97200 4324 97256 4326
rect 97280 4324 97336 4326
rect 96380 3834 96436 3836
rect 96460 3834 96516 3836
rect 96540 3834 96596 3836
rect 96620 3834 96676 3836
rect 96380 3782 96426 3834
rect 96426 3782 96436 3834
rect 96460 3782 96490 3834
rect 96490 3782 96502 3834
rect 96502 3782 96516 3834
rect 96540 3782 96554 3834
rect 96554 3782 96566 3834
rect 96566 3782 96596 3834
rect 96620 3782 96630 3834
rect 96630 3782 96676 3834
rect 96380 3780 96436 3782
rect 96460 3780 96516 3782
rect 96540 3780 96596 3782
rect 96620 3780 96676 3782
rect 97040 3290 97096 3292
rect 97120 3290 97176 3292
rect 97200 3290 97256 3292
rect 97280 3290 97336 3292
rect 97040 3238 97086 3290
rect 97086 3238 97096 3290
rect 97120 3238 97150 3290
rect 97150 3238 97162 3290
rect 97162 3238 97176 3290
rect 97200 3238 97214 3290
rect 97214 3238 97226 3290
rect 97226 3238 97256 3290
rect 97280 3238 97290 3290
rect 97290 3238 97336 3290
rect 97040 3236 97096 3238
rect 97120 3236 97176 3238
rect 97200 3236 97256 3238
rect 97280 3236 97336 3238
rect 96380 2746 96436 2748
rect 96460 2746 96516 2748
rect 96540 2746 96596 2748
rect 96620 2746 96676 2748
rect 96380 2694 96426 2746
rect 96426 2694 96436 2746
rect 96460 2694 96490 2746
rect 96490 2694 96502 2746
rect 96502 2694 96516 2746
rect 96540 2694 96554 2746
rect 96554 2694 96566 2746
rect 96566 2694 96596 2746
rect 96620 2694 96630 2746
rect 96630 2694 96676 2746
rect 96380 2692 96436 2694
rect 96460 2692 96516 2694
rect 96540 2692 96596 2694
rect 96620 2692 96676 2694
rect 35600 2202 35656 2204
rect 35680 2202 35736 2204
rect 35760 2202 35816 2204
rect 35840 2202 35896 2204
rect 35600 2150 35646 2202
rect 35646 2150 35656 2202
rect 35680 2150 35710 2202
rect 35710 2150 35722 2202
rect 35722 2150 35736 2202
rect 35760 2150 35774 2202
rect 35774 2150 35786 2202
rect 35786 2150 35816 2202
rect 35840 2150 35850 2202
rect 35850 2150 35896 2202
rect 35600 2148 35656 2150
rect 35680 2148 35736 2150
rect 35760 2148 35816 2150
rect 35840 2148 35896 2150
rect 66320 2202 66376 2204
rect 66400 2202 66456 2204
rect 66480 2202 66536 2204
rect 66560 2202 66616 2204
rect 66320 2150 66366 2202
rect 66366 2150 66376 2202
rect 66400 2150 66430 2202
rect 66430 2150 66442 2202
rect 66442 2150 66456 2202
rect 66480 2150 66494 2202
rect 66494 2150 66506 2202
rect 66506 2150 66536 2202
rect 66560 2150 66570 2202
rect 66570 2150 66616 2202
rect 66320 2148 66376 2150
rect 66400 2148 66456 2150
rect 66480 2148 66536 2150
rect 66560 2148 66616 2150
rect 97040 2202 97096 2204
rect 97120 2202 97176 2204
rect 97200 2202 97256 2204
rect 97280 2202 97336 2204
rect 97040 2150 97086 2202
rect 97086 2150 97096 2202
rect 97120 2150 97150 2202
rect 97150 2150 97162 2202
rect 97162 2150 97176 2202
rect 97200 2150 97214 2202
rect 97214 2150 97226 2202
rect 97226 2150 97256 2202
rect 97280 2150 97290 2202
rect 97290 2150 97336 2202
rect 97040 2148 97096 2150
rect 97120 2148 97176 2150
rect 97200 2148 97256 2150
rect 97280 2148 97336 2150
<< metal3 >>
rect 4870 95776 5186 95777
rect 4870 95712 4876 95776
rect 4940 95712 4956 95776
rect 5020 95712 5036 95776
rect 5100 95712 5116 95776
rect 5180 95712 5186 95776
rect 4870 95711 5186 95712
rect 35590 95776 35906 95777
rect 35590 95712 35596 95776
rect 35660 95712 35676 95776
rect 35740 95712 35756 95776
rect 35820 95712 35836 95776
rect 35900 95712 35906 95776
rect 35590 95711 35906 95712
rect 66310 95776 66626 95777
rect 66310 95712 66316 95776
rect 66380 95712 66396 95776
rect 66460 95712 66476 95776
rect 66540 95712 66556 95776
rect 66620 95712 66626 95776
rect 66310 95711 66626 95712
rect 97030 95776 97346 95777
rect 97030 95712 97036 95776
rect 97100 95712 97116 95776
rect 97180 95712 97196 95776
rect 97260 95712 97276 95776
rect 97340 95712 97346 95776
rect 97030 95711 97346 95712
rect 4210 95232 4526 95233
rect 4210 95168 4216 95232
rect 4280 95168 4296 95232
rect 4360 95168 4376 95232
rect 4440 95168 4456 95232
rect 4520 95168 4526 95232
rect 4210 95167 4526 95168
rect 34930 95232 35246 95233
rect 34930 95168 34936 95232
rect 35000 95168 35016 95232
rect 35080 95168 35096 95232
rect 35160 95168 35176 95232
rect 35240 95168 35246 95232
rect 34930 95167 35246 95168
rect 65650 95232 65966 95233
rect 65650 95168 65656 95232
rect 65720 95168 65736 95232
rect 65800 95168 65816 95232
rect 65880 95168 65896 95232
rect 65960 95168 65966 95232
rect 65650 95167 65966 95168
rect 96370 95232 96686 95233
rect 96370 95168 96376 95232
rect 96440 95168 96456 95232
rect 96520 95168 96536 95232
rect 96600 95168 96616 95232
rect 96680 95168 96686 95232
rect 96370 95167 96686 95168
rect 4870 94688 5186 94689
rect 4870 94624 4876 94688
rect 4940 94624 4956 94688
rect 5020 94624 5036 94688
rect 5100 94624 5116 94688
rect 5180 94624 5186 94688
rect 4870 94623 5186 94624
rect 35590 94688 35906 94689
rect 35590 94624 35596 94688
rect 35660 94624 35676 94688
rect 35740 94624 35756 94688
rect 35820 94624 35836 94688
rect 35900 94624 35906 94688
rect 35590 94623 35906 94624
rect 66310 94688 66626 94689
rect 66310 94624 66316 94688
rect 66380 94624 66396 94688
rect 66460 94624 66476 94688
rect 66540 94624 66556 94688
rect 66620 94624 66626 94688
rect 66310 94623 66626 94624
rect 97030 94688 97346 94689
rect 97030 94624 97036 94688
rect 97100 94624 97116 94688
rect 97180 94624 97196 94688
rect 97260 94624 97276 94688
rect 97340 94624 97346 94688
rect 97030 94623 97346 94624
rect 4210 94144 4526 94145
rect 4210 94080 4216 94144
rect 4280 94080 4296 94144
rect 4360 94080 4376 94144
rect 4440 94080 4456 94144
rect 4520 94080 4526 94144
rect 4210 94079 4526 94080
rect 34930 94144 35246 94145
rect 34930 94080 34936 94144
rect 35000 94080 35016 94144
rect 35080 94080 35096 94144
rect 35160 94080 35176 94144
rect 35240 94080 35246 94144
rect 34930 94079 35246 94080
rect 65650 94144 65966 94145
rect 65650 94080 65656 94144
rect 65720 94080 65736 94144
rect 65800 94080 65816 94144
rect 65880 94080 65896 94144
rect 65960 94080 65966 94144
rect 65650 94079 65966 94080
rect 96370 94144 96686 94145
rect 96370 94080 96376 94144
rect 96440 94080 96456 94144
rect 96520 94080 96536 94144
rect 96600 94080 96616 94144
rect 96680 94080 96686 94144
rect 96370 94079 96686 94080
rect 4870 93600 5186 93601
rect 4870 93536 4876 93600
rect 4940 93536 4956 93600
rect 5020 93536 5036 93600
rect 5100 93536 5116 93600
rect 5180 93536 5186 93600
rect 4870 93535 5186 93536
rect 35590 93600 35906 93601
rect 35590 93536 35596 93600
rect 35660 93536 35676 93600
rect 35740 93536 35756 93600
rect 35820 93536 35836 93600
rect 35900 93536 35906 93600
rect 35590 93535 35906 93536
rect 66310 93600 66626 93601
rect 66310 93536 66316 93600
rect 66380 93536 66396 93600
rect 66460 93536 66476 93600
rect 66540 93536 66556 93600
rect 66620 93536 66626 93600
rect 66310 93535 66626 93536
rect 97030 93600 97346 93601
rect 97030 93536 97036 93600
rect 97100 93536 97116 93600
rect 97180 93536 97196 93600
rect 97260 93536 97276 93600
rect 97340 93536 97346 93600
rect 97030 93535 97346 93536
rect 4210 93056 4526 93057
rect 4210 92992 4216 93056
rect 4280 92992 4296 93056
rect 4360 92992 4376 93056
rect 4440 92992 4456 93056
rect 4520 92992 4526 93056
rect 4210 92991 4526 92992
rect 34930 93056 35246 93057
rect 34930 92992 34936 93056
rect 35000 92992 35016 93056
rect 35080 92992 35096 93056
rect 35160 92992 35176 93056
rect 35240 92992 35246 93056
rect 34930 92991 35246 92992
rect 65650 93056 65966 93057
rect 65650 92992 65656 93056
rect 65720 92992 65736 93056
rect 65800 92992 65816 93056
rect 65880 92992 65896 93056
rect 65960 92992 65966 93056
rect 65650 92991 65966 92992
rect 96370 93056 96686 93057
rect 96370 92992 96376 93056
rect 96440 92992 96456 93056
rect 96520 92992 96536 93056
rect 96600 92992 96616 93056
rect 96680 92992 96686 93056
rect 96370 92991 96686 92992
rect 4870 92512 5186 92513
rect 4870 92448 4876 92512
rect 4940 92448 4956 92512
rect 5020 92448 5036 92512
rect 5100 92448 5116 92512
rect 5180 92448 5186 92512
rect 4870 92447 5186 92448
rect 97030 92512 97346 92513
rect 97030 92448 97036 92512
rect 97100 92448 97116 92512
rect 97180 92448 97196 92512
rect 97260 92448 97276 92512
rect 97340 92448 97346 92512
rect 97030 92447 97346 92448
rect 4210 91968 4526 91969
rect 4210 91904 4216 91968
rect 4280 91904 4296 91968
rect 4360 91904 4376 91968
rect 4440 91904 4456 91968
rect 4520 91904 4526 91968
rect 4210 91903 4526 91904
rect 96370 91968 96686 91969
rect 96370 91904 96376 91968
rect 96440 91904 96456 91968
rect 96520 91904 96536 91968
rect 96600 91904 96616 91968
rect 96680 91904 96686 91968
rect 96370 91903 96686 91904
rect 4870 91424 5186 91425
rect 4870 91360 4876 91424
rect 4940 91360 4956 91424
rect 5020 91360 5036 91424
rect 5100 91360 5116 91424
rect 5180 91360 5186 91424
rect 4870 91359 5186 91360
rect 97030 91424 97346 91425
rect 97030 91360 97036 91424
rect 97100 91360 97116 91424
rect 97180 91360 97196 91424
rect 97260 91360 97276 91424
rect 97340 91360 97346 91424
rect 97030 91359 97346 91360
rect 4210 90880 4526 90881
rect 4210 90816 4216 90880
rect 4280 90816 4296 90880
rect 4360 90816 4376 90880
rect 4440 90816 4456 90880
rect 4520 90816 4526 90880
rect 4210 90815 4526 90816
rect 96370 90880 96686 90881
rect 96370 90816 96376 90880
rect 96440 90816 96456 90880
rect 96520 90816 96536 90880
rect 96600 90816 96616 90880
rect 96680 90816 96686 90880
rect 96370 90815 96686 90816
rect 13261 90538 13327 90541
rect 50838 90538 50844 90540
rect 13261 90536 50844 90538
rect 13261 90480 13266 90536
rect 13322 90480 50844 90536
rect 13261 90478 50844 90480
rect 13261 90475 13327 90478
rect 50838 90476 50844 90478
rect 50908 90476 50914 90540
rect 4870 90336 5186 90337
rect 4870 90272 4876 90336
rect 4940 90272 4956 90336
rect 5020 90272 5036 90336
rect 5100 90272 5116 90336
rect 5180 90272 5186 90336
rect 4870 90271 5186 90272
rect 97030 90336 97346 90337
rect 97030 90272 97036 90336
rect 97100 90272 97116 90336
rect 97180 90272 97196 90336
rect 97260 90272 97276 90336
rect 97340 90272 97346 90336
rect 97030 90271 97346 90272
rect 4210 89792 4526 89793
rect 4210 89728 4216 89792
rect 4280 89728 4296 89792
rect 4360 89728 4376 89792
rect 4440 89728 4456 89792
rect 4520 89728 4526 89792
rect 4210 89727 4526 89728
rect 96370 89792 96686 89793
rect 96370 89728 96376 89792
rect 96440 89728 96456 89792
rect 96520 89728 96536 89792
rect 96600 89728 96616 89792
rect 96680 89728 96686 89792
rect 96370 89727 96686 89728
rect 4870 89248 5186 89249
rect 4870 89184 4876 89248
rect 4940 89184 4956 89248
rect 5020 89184 5036 89248
rect 5100 89184 5116 89248
rect 5180 89184 5186 89248
rect 4870 89183 5186 89184
rect 97030 89248 97346 89249
rect 97030 89184 97036 89248
rect 97100 89184 97116 89248
rect 97180 89184 97196 89248
rect 97260 89184 97276 89248
rect 97340 89184 97346 89248
rect 97030 89183 97346 89184
rect 4210 88704 4526 88705
rect 4210 88640 4216 88704
rect 4280 88640 4296 88704
rect 4360 88640 4376 88704
rect 4440 88640 4456 88704
rect 4520 88640 4526 88704
rect 4210 88639 4526 88640
rect 96370 88704 96686 88705
rect 96370 88640 96376 88704
rect 96440 88640 96456 88704
rect 96520 88640 96536 88704
rect 96600 88640 96616 88704
rect 96680 88640 96686 88704
rect 96370 88639 96686 88640
rect 4870 88160 5186 88161
rect 4870 88096 4876 88160
rect 4940 88096 4956 88160
rect 5020 88096 5036 88160
rect 5100 88096 5116 88160
rect 5180 88096 5186 88160
rect 4870 88095 5186 88096
rect 97030 88160 97346 88161
rect 97030 88096 97036 88160
rect 97100 88096 97116 88160
rect 97180 88096 97196 88160
rect 97260 88096 97276 88160
rect 97340 88096 97346 88160
rect 97030 88095 97346 88096
rect 4210 87616 4526 87617
rect 4210 87552 4216 87616
rect 4280 87552 4296 87616
rect 4360 87552 4376 87616
rect 4440 87552 4456 87616
rect 4520 87552 4526 87616
rect 4210 87551 4526 87552
rect 96370 87616 96686 87617
rect 96370 87552 96376 87616
rect 96440 87552 96456 87616
rect 96520 87552 96536 87616
rect 96600 87552 96616 87616
rect 96680 87552 96686 87616
rect 96370 87551 96686 87552
rect 8293 87546 8359 87549
rect 8293 87544 8402 87546
rect 8293 87488 8298 87544
rect 8354 87488 8402 87544
rect 8293 87483 8402 87488
rect 8342 87380 8402 87483
rect 97349 87410 97415 87413
rect 91908 87408 97415 87410
rect 91908 87352 97354 87408
rect 97410 87352 97415 87408
rect 91908 87350 97415 87352
rect 97349 87347 97415 87350
rect 841 87274 907 87277
rect 798 87272 907 87274
rect 798 87216 846 87272
rect 902 87216 907 87272
rect 798 87211 907 87216
rect 798 87168 858 87211
rect 0 87078 858 87168
rect 97533 87138 97599 87141
rect 98200 87138 99000 87168
rect 97533 87136 99000 87138
rect 97533 87080 97538 87136
rect 97594 87080 99000 87136
rect 97533 87078 99000 87080
rect 0 87048 800 87078
rect 97533 87075 97599 87078
rect 4870 87072 5186 87073
rect 4870 87008 4876 87072
rect 4940 87008 4956 87072
rect 5020 87008 5036 87072
rect 5100 87008 5116 87072
rect 5180 87008 5186 87072
rect 4870 87007 5186 87008
rect 97030 87072 97346 87073
rect 97030 87008 97036 87072
rect 97100 87008 97116 87072
rect 97180 87008 97196 87072
rect 97260 87008 97276 87072
rect 97340 87008 97346 87072
rect 98200 87048 99000 87078
rect 97030 87007 97346 87008
rect 8293 86730 8359 86733
rect 8293 86728 8402 86730
rect 8293 86672 8298 86728
rect 8354 86672 8402 86728
rect 8293 86667 8402 86672
rect 841 86594 907 86597
rect 798 86592 907 86594
rect 798 86536 846 86592
rect 902 86536 907 86592
rect 798 86531 907 86536
rect 798 86488 858 86531
rect 0 86398 858 86488
rect 4210 86528 4526 86529
rect 4210 86464 4216 86528
rect 4280 86464 4296 86528
rect 4360 86464 4376 86528
rect 4440 86464 4456 86528
rect 4520 86464 4526 86528
rect 4210 86463 4526 86464
rect 0 86368 800 86398
rect 8342 86292 8402 86667
rect 96370 86528 96686 86529
rect 96370 86464 96376 86528
rect 96440 86464 96456 86528
rect 96520 86464 96536 86528
rect 96600 86464 96616 86528
rect 96680 86464 96686 86528
rect 96370 86463 96686 86464
rect 97533 86458 97599 86461
rect 98200 86458 99000 86488
rect 97533 86456 99000 86458
rect 97533 86400 97538 86456
rect 97594 86400 99000 86456
rect 97533 86398 99000 86400
rect 97533 86395 97599 86398
rect 98200 86368 99000 86398
rect 97349 86322 97415 86325
rect 91908 86320 97415 86322
rect 91908 86264 97354 86320
rect 97410 86264 97415 86320
rect 91908 86262 97415 86264
rect 97349 86259 97415 86262
rect 4870 85984 5186 85985
rect 4870 85920 4876 85984
rect 4940 85920 4956 85984
rect 5020 85920 5036 85984
rect 5100 85920 5116 85984
rect 5180 85920 5186 85984
rect 4870 85919 5186 85920
rect 97030 85984 97346 85985
rect 97030 85920 97036 85984
rect 97100 85920 97116 85984
rect 97180 85920 97196 85984
rect 97260 85920 97276 85984
rect 97340 85920 97346 85984
rect 97030 85919 97346 85920
rect 4210 85440 4526 85441
rect 4210 85376 4216 85440
rect 4280 85376 4296 85440
rect 4360 85376 4376 85440
rect 4440 85376 4456 85440
rect 4520 85376 4526 85440
rect 4210 85375 4526 85376
rect 96370 85440 96686 85441
rect 96370 85376 96376 85440
rect 96440 85376 96456 85440
rect 96520 85376 96536 85440
rect 96600 85376 96616 85440
rect 96680 85376 96686 85440
rect 96370 85375 96686 85376
rect 8293 85370 8359 85373
rect 8293 85368 8402 85370
rect 8293 85312 8298 85368
rect 8354 85312 8402 85368
rect 8293 85307 8402 85312
rect 8342 85204 8402 85307
rect 97349 85234 97415 85237
rect 91908 85232 97415 85234
rect 91908 85176 97354 85232
rect 97410 85176 97415 85232
rect 91908 85174 97415 85176
rect 97349 85171 97415 85174
rect 0 85098 800 85128
rect 97533 85098 97599 85101
rect 98200 85098 99000 85128
rect 0 85008 858 85098
rect 97533 85096 99000 85098
rect 97533 85040 97538 85096
rect 97594 85040 99000 85096
rect 97533 85038 99000 85040
rect 97533 85035 97599 85038
rect 98200 85008 99000 85038
rect 798 84965 858 85008
rect 798 84960 907 84965
rect 798 84904 846 84960
rect 902 84904 907 84960
rect 798 84902 907 84904
rect 841 84899 907 84902
rect 4870 84896 5186 84897
rect 4870 84832 4876 84896
rect 4940 84832 4956 84896
rect 5020 84832 5036 84896
rect 5100 84832 5116 84896
rect 5180 84832 5186 84896
rect 4870 84831 5186 84832
rect 97030 84896 97346 84897
rect 97030 84832 97036 84896
rect 97100 84832 97116 84896
rect 97180 84832 97196 84896
rect 97260 84832 97276 84896
rect 97340 84832 97346 84896
rect 97030 84831 97346 84832
rect 841 84554 907 84557
rect 798 84552 907 84554
rect 798 84496 846 84552
rect 902 84496 907 84552
rect 798 84491 907 84496
rect 798 84448 858 84491
rect 0 84358 858 84448
rect 97533 84418 97599 84421
rect 98200 84418 99000 84448
rect 97533 84416 99000 84418
rect 97533 84360 97538 84416
rect 97594 84360 99000 84416
rect 97533 84358 99000 84360
rect 0 84328 800 84358
rect 97533 84355 97599 84358
rect 4210 84352 4526 84353
rect 4210 84288 4216 84352
rect 4280 84288 4296 84352
rect 4360 84288 4376 84352
rect 4440 84288 4456 84352
rect 4520 84288 4526 84352
rect 4210 84287 4526 84288
rect 96370 84352 96686 84353
rect 96370 84288 96376 84352
rect 96440 84288 96456 84352
rect 96520 84288 96536 84352
rect 96600 84288 96616 84352
rect 96680 84288 96686 84352
rect 98200 84328 99000 84358
rect 96370 84287 96686 84288
rect 1669 84146 1735 84149
rect 97349 84146 97415 84149
rect 1669 84144 8188 84146
rect 1669 84088 1674 84144
rect 1730 84088 8188 84144
rect 1669 84086 8188 84088
rect 91908 84144 97415 84146
rect 91908 84088 97354 84144
rect 97410 84088 97415 84144
rect 91908 84086 97415 84088
rect 1669 84083 1735 84086
rect 97349 84083 97415 84086
rect 4870 83808 5186 83809
rect 4870 83744 4876 83808
rect 4940 83744 4956 83808
rect 5020 83744 5036 83808
rect 5100 83744 5116 83808
rect 5180 83744 5186 83808
rect 4870 83743 5186 83744
rect 97030 83808 97346 83809
rect 97030 83744 97036 83808
rect 97100 83744 97116 83808
rect 97180 83744 97196 83808
rect 97260 83744 97276 83808
rect 97340 83744 97346 83808
rect 97030 83743 97346 83744
rect 8293 83466 8359 83469
rect 8293 83464 8402 83466
rect 8293 83408 8298 83464
rect 8354 83408 8402 83464
rect 8293 83403 8402 83408
rect 4210 83264 4526 83265
rect 4210 83200 4216 83264
rect 4280 83200 4296 83264
rect 4360 83200 4376 83264
rect 4440 83200 4456 83264
rect 4520 83200 4526 83264
rect 4210 83199 4526 83200
rect 841 83194 907 83197
rect 798 83192 907 83194
rect 798 83136 846 83192
rect 902 83136 907 83192
rect 798 83131 907 83136
rect 798 83088 858 83131
rect 0 82998 858 83088
rect 8342 83028 8402 83403
rect 96370 83264 96686 83265
rect 96370 83200 96376 83264
rect 96440 83200 96456 83264
rect 96520 83200 96536 83264
rect 96600 83200 96616 83264
rect 96680 83200 96686 83264
rect 96370 83199 96686 83200
rect 97349 83058 97415 83061
rect 91908 83056 97415 83058
rect 91908 83000 97354 83056
rect 97410 83000 97415 83056
rect 91908 82998 97415 83000
rect 0 82968 800 82998
rect 97349 82995 97415 82998
rect 97533 83058 97599 83061
rect 98200 83058 99000 83088
rect 97533 83056 99000 83058
rect 97533 83000 97538 83056
rect 97594 83000 99000 83056
rect 97533 82998 99000 83000
rect 97533 82995 97599 82998
rect 98200 82968 99000 82998
rect 4870 82720 5186 82721
rect 4870 82656 4876 82720
rect 4940 82656 4956 82720
rect 5020 82656 5036 82720
rect 5100 82656 5116 82720
rect 5180 82656 5186 82720
rect 4870 82655 5186 82656
rect 97030 82720 97346 82721
rect 97030 82656 97036 82720
rect 97100 82656 97116 82720
rect 97180 82656 97196 82720
rect 97260 82656 97276 82720
rect 97340 82656 97346 82720
rect 97030 82655 97346 82656
rect 4210 82176 4526 82177
rect 4210 82112 4216 82176
rect 4280 82112 4296 82176
rect 4360 82112 4376 82176
rect 4440 82112 4456 82176
rect 4520 82112 4526 82176
rect 4210 82111 4526 82112
rect 96370 82176 96686 82177
rect 96370 82112 96376 82176
rect 96440 82112 96456 82176
rect 96520 82112 96536 82176
rect 96600 82112 96616 82176
rect 96680 82112 96686 82176
rect 96370 82111 96686 82112
rect 8293 82106 8359 82109
rect 8293 82104 8402 82106
rect 8293 82048 8298 82104
rect 8354 82048 8402 82104
rect 8293 82043 8402 82048
rect 8342 81940 8402 82043
rect 97349 81970 97415 81973
rect 91908 81968 97415 81970
rect 91908 81912 97354 81968
rect 97410 81912 97415 81968
rect 91908 81910 97415 81912
rect 97349 81907 97415 81910
rect 841 81834 907 81837
rect 798 81832 907 81834
rect 798 81776 846 81832
rect 902 81776 907 81832
rect 798 81771 907 81776
rect 798 81728 858 81771
rect 0 81638 858 81728
rect 97533 81698 97599 81701
rect 98200 81698 99000 81728
rect 97533 81696 99000 81698
rect 97533 81640 97538 81696
rect 97594 81640 99000 81696
rect 97533 81638 99000 81640
rect 0 81608 800 81638
rect 97533 81635 97599 81638
rect 4870 81632 5186 81633
rect 4870 81568 4876 81632
rect 4940 81568 4956 81632
rect 5020 81568 5036 81632
rect 5100 81568 5116 81632
rect 5180 81568 5186 81632
rect 4870 81567 5186 81568
rect 97030 81632 97346 81633
rect 97030 81568 97036 81632
rect 97100 81568 97116 81632
rect 97180 81568 97196 81632
rect 97260 81568 97276 81632
rect 97340 81568 97346 81632
rect 98200 81608 99000 81638
rect 97030 81567 97346 81568
rect 8293 81290 8359 81293
rect 8293 81288 8402 81290
rect 8293 81232 8298 81288
rect 8354 81232 8402 81288
rect 8293 81227 8402 81232
rect 841 81154 907 81157
rect 798 81152 907 81154
rect 798 81096 846 81152
rect 902 81096 907 81152
rect 798 81091 907 81096
rect 798 81048 858 81091
rect 0 80958 858 81048
rect 4210 81088 4526 81089
rect 4210 81024 4216 81088
rect 4280 81024 4296 81088
rect 4360 81024 4376 81088
rect 4440 81024 4456 81088
rect 4520 81024 4526 81088
rect 4210 81023 4526 81024
rect 0 80928 800 80958
rect 8342 80852 8402 81227
rect 96370 81088 96686 81089
rect 96370 81024 96376 81088
rect 96440 81024 96456 81088
rect 96520 81024 96536 81088
rect 96600 81024 96616 81088
rect 96680 81024 96686 81088
rect 96370 81023 96686 81024
rect 97533 81018 97599 81021
rect 98200 81018 99000 81048
rect 97533 81016 99000 81018
rect 97533 80960 97538 81016
rect 97594 80960 99000 81016
rect 97533 80958 99000 80960
rect 97533 80955 97599 80958
rect 98200 80928 99000 80958
rect 97349 80882 97415 80885
rect 91908 80880 97415 80882
rect 91908 80824 97354 80880
rect 97410 80824 97415 80880
rect 91908 80822 97415 80824
rect 97349 80819 97415 80822
rect 4870 80544 5186 80545
rect 4870 80480 4876 80544
rect 4940 80480 4956 80544
rect 5020 80480 5036 80544
rect 5100 80480 5116 80544
rect 5180 80480 5186 80544
rect 4870 80479 5186 80480
rect 97030 80544 97346 80545
rect 97030 80480 97036 80544
rect 97100 80480 97116 80544
rect 97180 80480 97196 80544
rect 97260 80480 97276 80544
rect 97340 80480 97346 80544
rect 97030 80479 97346 80480
rect 4210 80000 4526 80001
rect 4210 79936 4216 80000
rect 4280 79936 4296 80000
rect 4360 79936 4376 80000
rect 4440 79936 4456 80000
rect 4520 79936 4526 80000
rect 4210 79935 4526 79936
rect 96370 80000 96686 80001
rect 96370 79936 96376 80000
rect 96440 79936 96456 80000
rect 96520 79936 96536 80000
rect 96600 79936 96616 80000
rect 96680 79936 96686 80000
rect 96370 79935 96686 79936
rect 8293 79930 8359 79933
rect 8293 79928 8402 79930
rect 8293 79872 8298 79928
rect 8354 79872 8402 79928
rect 8293 79867 8402 79872
rect 8342 79764 8402 79867
rect 97349 79794 97415 79797
rect 91908 79792 97415 79794
rect 91908 79736 97354 79792
rect 97410 79736 97415 79792
rect 91908 79734 97415 79736
rect 97349 79731 97415 79734
rect 0 79658 800 79688
rect 97533 79658 97599 79661
rect 98200 79658 99000 79688
rect 0 79568 858 79658
rect 97533 79656 99000 79658
rect 97533 79600 97538 79656
rect 97594 79600 99000 79656
rect 97533 79598 99000 79600
rect 97533 79595 97599 79598
rect 98200 79568 99000 79598
rect 798 79525 858 79568
rect 798 79520 907 79525
rect 798 79464 846 79520
rect 902 79464 907 79520
rect 798 79462 907 79464
rect 841 79459 907 79462
rect 4870 79456 5186 79457
rect 4870 79392 4876 79456
rect 4940 79392 4956 79456
rect 5020 79392 5036 79456
rect 5100 79392 5116 79456
rect 5180 79392 5186 79456
rect 4870 79391 5186 79392
rect 97030 79456 97346 79457
rect 97030 79392 97036 79456
rect 97100 79392 97116 79456
rect 97180 79392 97196 79456
rect 97260 79392 97276 79456
rect 97340 79392 97346 79456
rect 97030 79391 97346 79392
rect 841 79114 907 79117
rect 798 79112 907 79114
rect 798 79056 846 79112
rect 902 79056 907 79112
rect 798 79051 907 79056
rect 8293 79114 8359 79117
rect 8293 79112 8402 79114
rect 8293 79056 8298 79112
rect 8354 79056 8402 79112
rect 8293 79051 8402 79056
rect 798 79008 858 79051
rect 0 78918 858 79008
rect 0 78888 800 78918
rect 4210 78912 4526 78913
rect 4210 78848 4216 78912
rect 4280 78848 4296 78912
rect 4360 78848 4376 78912
rect 4440 78848 4456 78912
rect 4520 78848 4526 78912
rect 4210 78847 4526 78848
rect 8342 78676 8402 79051
rect 97441 78978 97507 78981
rect 98200 78978 99000 79008
rect 97441 78976 99000 78978
rect 97441 78920 97446 78976
rect 97502 78920 99000 78976
rect 97441 78918 99000 78920
rect 97441 78915 97507 78918
rect 96370 78912 96686 78913
rect 96370 78848 96376 78912
rect 96440 78848 96456 78912
rect 96520 78848 96536 78912
rect 96600 78848 96616 78912
rect 96680 78848 96686 78912
rect 98200 78888 99000 78918
rect 96370 78847 96686 78848
rect 97257 78706 97323 78709
rect 91908 78704 97323 78706
rect 91908 78648 97262 78704
rect 97318 78648 97323 78704
rect 91908 78646 97323 78648
rect 97257 78643 97323 78646
rect 4870 78368 5186 78369
rect 4870 78304 4876 78368
rect 4940 78304 4956 78368
rect 5020 78304 5036 78368
rect 5100 78304 5116 78368
rect 5180 78304 5186 78368
rect 4870 78303 5186 78304
rect 97030 78368 97346 78369
rect 97030 78304 97036 78368
rect 97100 78304 97116 78368
rect 97180 78304 97196 78368
rect 97260 78304 97276 78368
rect 97340 78304 97346 78368
rect 97030 78303 97346 78304
rect 8293 78026 8359 78029
rect 8293 78024 8402 78026
rect 8293 77968 8298 78024
rect 8354 77968 8402 78024
rect 8293 77963 8402 77968
rect 4210 77824 4526 77825
rect 4210 77760 4216 77824
rect 4280 77760 4296 77824
rect 4360 77760 4376 77824
rect 4440 77760 4456 77824
rect 4520 77760 4526 77824
rect 4210 77759 4526 77760
rect 841 77754 907 77757
rect 798 77752 907 77754
rect 798 77696 846 77752
rect 902 77696 907 77752
rect 798 77691 907 77696
rect 798 77648 858 77691
rect 0 77558 858 77648
rect 8342 77588 8402 77963
rect 96370 77824 96686 77825
rect 96370 77760 96376 77824
rect 96440 77760 96456 77824
rect 96520 77760 96536 77824
rect 96600 77760 96616 77824
rect 96680 77760 96686 77824
rect 96370 77759 96686 77760
rect 97349 77618 97415 77621
rect 91908 77616 97415 77618
rect 91908 77560 97354 77616
rect 97410 77560 97415 77616
rect 91908 77558 97415 77560
rect 0 77528 800 77558
rect 97349 77555 97415 77558
rect 97533 77618 97599 77621
rect 98200 77618 99000 77648
rect 97533 77616 99000 77618
rect 97533 77560 97538 77616
rect 97594 77560 99000 77616
rect 97533 77558 99000 77560
rect 97533 77555 97599 77558
rect 98200 77528 99000 77558
rect 4870 77280 5186 77281
rect 4870 77216 4876 77280
rect 4940 77216 4956 77280
rect 5020 77216 5036 77280
rect 5100 77216 5116 77280
rect 5180 77216 5186 77280
rect 4870 77215 5186 77216
rect 97030 77280 97346 77281
rect 97030 77216 97036 77280
rect 97100 77216 97116 77280
rect 97180 77216 97196 77280
rect 97260 77216 97276 77280
rect 97340 77216 97346 77280
rect 97030 77215 97346 77216
rect 4210 76736 4526 76737
rect 4210 76672 4216 76736
rect 4280 76672 4296 76736
rect 4360 76672 4376 76736
rect 4440 76672 4456 76736
rect 4520 76672 4526 76736
rect 4210 76671 4526 76672
rect 96370 76736 96686 76737
rect 96370 76672 96376 76736
rect 96440 76672 96456 76736
rect 96520 76672 96536 76736
rect 96600 76672 96616 76736
rect 96680 76672 96686 76736
rect 96370 76671 96686 76672
rect 8293 76666 8359 76669
rect 8293 76664 8402 76666
rect 8293 76608 8298 76664
rect 8354 76608 8402 76664
rect 8293 76603 8402 76608
rect 8342 76500 8402 76603
rect 97349 76530 97415 76533
rect 91908 76528 97415 76530
rect 91908 76472 97354 76528
rect 97410 76472 97415 76528
rect 91908 76470 97415 76472
rect 97349 76467 97415 76470
rect 841 76394 907 76397
rect 798 76392 907 76394
rect 798 76336 846 76392
rect 902 76336 907 76392
rect 798 76331 907 76336
rect 798 76288 858 76331
rect 0 76198 858 76288
rect 97533 76258 97599 76261
rect 98200 76258 99000 76288
rect 97533 76256 99000 76258
rect 97533 76200 97538 76256
rect 97594 76200 99000 76256
rect 97533 76198 99000 76200
rect 0 76168 800 76198
rect 97533 76195 97599 76198
rect 4870 76192 5186 76193
rect 4870 76128 4876 76192
rect 4940 76128 4956 76192
rect 5020 76128 5036 76192
rect 5100 76128 5116 76192
rect 5180 76128 5186 76192
rect 4870 76127 5186 76128
rect 97030 76192 97346 76193
rect 97030 76128 97036 76192
rect 97100 76128 97116 76192
rect 97180 76128 97196 76192
rect 97260 76128 97276 76192
rect 97340 76128 97346 76192
rect 98200 76168 99000 76198
rect 97030 76127 97346 76128
rect 841 75714 907 75717
rect 798 75712 907 75714
rect 798 75656 846 75712
rect 902 75656 907 75712
rect 798 75651 907 75656
rect 798 75608 858 75651
rect 0 75518 858 75608
rect 4210 75648 4526 75649
rect 4210 75584 4216 75648
rect 4280 75584 4296 75648
rect 4360 75584 4376 75648
rect 4440 75584 4456 75648
rect 4520 75584 4526 75648
rect 4210 75583 4526 75584
rect 96370 75648 96686 75649
rect 96370 75584 96376 75648
rect 96440 75584 96456 75648
rect 96520 75584 96536 75648
rect 96600 75584 96616 75648
rect 96680 75584 96686 75648
rect 96370 75583 96686 75584
rect 97533 75578 97599 75581
rect 98200 75578 99000 75608
rect 97533 75576 99000 75578
rect 97533 75520 97538 75576
rect 97594 75520 99000 75576
rect 97533 75518 99000 75520
rect 0 75488 800 75518
rect 97533 75515 97599 75518
rect 98200 75488 99000 75518
rect 1669 75442 1735 75445
rect 97349 75442 97415 75445
rect 1669 75440 8188 75442
rect 1669 75384 1674 75440
rect 1730 75384 8188 75440
rect 1669 75382 8188 75384
rect 91908 75440 97415 75442
rect 91908 75384 97354 75440
rect 97410 75384 97415 75440
rect 91908 75382 97415 75384
rect 1669 75379 1735 75382
rect 97349 75379 97415 75382
rect 4870 75104 5186 75105
rect 4870 75040 4876 75104
rect 4940 75040 4956 75104
rect 5020 75040 5036 75104
rect 5100 75040 5116 75104
rect 5180 75040 5186 75104
rect 4870 75039 5186 75040
rect 97030 75104 97346 75105
rect 97030 75040 97036 75104
rect 97100 75040 97116 75104
rect 97180 75040 97196 75104
rect 97260 75040 97276 75104
rect 97340 75040 97346 75104
rect 97030 75039 97346 75040
rect 4210 74560 4526 74561
rect 4210 74496 4216 74560
rect 4280 74496 4296 74560
rect 4360 74496 4376 74560
rect 4440 74496 4456 74560
rect 4520 74496 4526 74560
rect 4210 74495 4526 74496
rect 96370 74560 96686 74561
rect 96370 74496 96376 74560
rect 96440 74496 96456 74560
rect 96520 74496 96536 74560
rect 96600 74496 96616 74560
rect 96680 74496 96686 74560
rect 96370 74495 96686 74496
rect 8293 74490 8359 74493
rect 8293 74488 8402 74490
rect 8293 74432 8298 74488
rect 8354 74432 8402 74488
rect 8293 74427 8402 74432
rect 8342 74324 8402 74427
rect 97257 74354 97323 74357
rect 91908 74352 97323 74354
rect 91908 74296 97262 74352
rect 97318 74296 97323 74352
rect 91908 74294 97323 74296
rect 97257 74291 97323 74294
rect 0 74218 800 74248
rect 97441 74218 97507 74221
rect 98200 74218 99000 74248
rect 0 74128 858 74218
rect 97441 74216 99000 74218
rect 97441 74160 97446 74216
rect 97502 74160 99000 74216
rect 97441 74158 99000 74160
rect 97441 74155 97507 74158
rect 98200 74128 99000 74158
rect 798 74085 858 74128
rect 798 74080 907 74085
rect 798 74024 846 74080
rect 902 74024 907 74080
rect 798 74022 907 74024
rect 841 74019 907 74022
rect 4870 74016 5186 74017
rect 4870 73952 4876 74016
rect 4940 73952 4956 74016
rect 5020 73952 5036 74016
rect 5100 73952 5116 74016
rect 5180 73952 5186 74016
rect 4870 73951 5186 73952
rect 97030 74016 97346 74017
rect 97030 73952 97036 74016
rect 97100 73952 97116 74016
rect 97180 73952 97196 74016
rect 97260 73952 97276 74016
rect 97340 73952 97346 74016
rect 97030 73951 97346 73952
rect 841 73674 907 73677
rect 798 73672 907 73674
rect 798 73616 846 73672
rect 902 73616 907 73672
rect 798 73611 907 73616
rect 8293 73674 8359 73677
rect 8293 73672 8402 73674
rect 8293 73616 8298 73672
rect 8354 73616 8402 73672
rect 8293 73611 8402 73616
rect 798 73568 858 73611
rect 0 73478 858 73568
rect 0 73448 800 73478
rect 4210 73472 4526 73473
rect 4210 73408 4216 73472
rect 4280 73408 4296 73472
rect 4360 73408 4376 73472
rect 4440 73408 4456 73472
rect 4520 73408 4526 73472
rect 4210 73407 4526 73408
rect 8342 73236 8402 73611
rect 97533 73538 97599 73541
rect 98200 73538 99000 73568
rect 97533 73536 99000 73538
rect 97533 73480 97538 73536
rect 97594 73480 99000 73536
rect 97533 73478 99000 73480
rect 97533 73475 97599 73478
rect 96370 73472 96686 73473
rect 96370 73408 96376 73472
rect 96440 73408 96456 73472
rect 96520 73408 96536 73472
rect 96600 73408 96616 73472
rect 96680 73408 96686 73472
rect 98200 73448 99000 73478
rect 96370 73407 96686 73408
rect 97349 73266 97415 73269
rect 91908 73264 97415 73266
rect 91908 73208 97354 73264
rect 97410 73208 97415 73264
rect 91908 73206 97415 73208
rect 97349 73203 97415 73206
rect 4870 72928 5186 72929
rect 4870 72864 4876 72928
rect 4940 72864 4956 72928
rect 5020 72864 5036 72928
rect 5100 72864 5116 72928
rect 5180 72864 5186 72928
rect 4870 72863 5186 72864
rect 97030 72928 97346 72929
rect 97030 72864 97036 72928
rect 97100 72864 97116 72928
rect 97180 72864 97196 72928
rect 97260 72864 97276 72928
rect 97340 72864 97346 72928
rect 97030 72863 97346 72864
rect 8293 72586 8359 72589
rect 8293 72584 8402 72586
rect 8293 72528 8298 72584
rect 8354 72528 8402 72584
rect 8293 72523 8402 72528
rect 4210 72384 4526 72385
rect 4210 72320 4216 72384
rect 4280 72320 4296 72384
rect 4360 72320 4376 72384
rect 4440 72320 4456 72384
rect 4520 72320 4526 72384
rect 4210 72319 4526 72320
rect 841 72314 907 72317
rect 798 72312 907 72314
rect 798 72256 846 72312
rect 902 72256 907 72312
rect 798 72251 907 72256
rect 798 72208 858 72251
rect 0 72118 858 72208
rect 8342 72148 8402 72523
rect 96370 72384 96686 72385
rect 96370 72320 96376 72384
rect 96440 72320 96456 72384
rect 96520 72320 96536 72384
rect 96600 72320 96616 72384
rect 96680 72320 96686 72384
rect 96370 72319 96686 72320
rect 97257 72178 97323 72181
rect 91908 72176 97323 72178
rect 91908 72120 97262 72176
rect 97318 72120 97323 72176
rect 91908 72118 97323 72120
rect 0 72088 800 72118
rect 97257 72115 97323 72118
rect 97533 72178 97599 72181
rect 98200 72178 99000 72208
rect 97533 72176 99000 72178
rect 97533 72120 97538 72176
rect 97594 72120 99000 72176
rect 97533 72118 99000 72120
rect 97533 72115 97599 72118
rect 98200 72088 99000 72118
rect 4870 71840 5186 71841
rect 4870 71776 4876 71840
rect 4940 71776 4956 71840
rect 5020 71776 5036 71840
rect 5100 71776 5116 71840
rect 5180 71776 5186 71840
rect 4870 71775 5186 71776
rect 97030 71840 97346 71841
rect 97030 71776 97036 71840
rect 97100 71776 97116 71840
rect 97180 71776 97196 71840
rect 97260 71776 97276 71840
rect 97340 71776 97346 71840
rect 97030 71775 97346 71776
rect 4210 71296 4526 71297
rect 4210 71232 4216 71296
rect 4280 71232 4296 71296
rect 4360 71232 4376 71296
rect 4440 71232 4456 71296
rect 4520 71232 4526 71296
rect 4210 71231 4526 71232
rect 96370 71296 96686 71297
rect 96370 71232 96376 71296
rect 96440 71232 96456 71296
rect 96520 71232 96536 71296
rect 96600 71232 96616 71296
rect 96680 71232 96686 71296
rect 96370 71231 96686 71232
rect 8293 71226 8359 71229
rect 8293 71224 8402 71226
rect 8293 71168 8298 71224
rect 8354 71168 8402 71224
rect 8293 71163 8402 71168
rect 8342 71060 8402 71163
rect 97349 71090 97415 71093
rect 91908 71088 97415 71090
rect 91908 71032 97354 71088
rect 97410 71032 97415 71088
rect 91908 71030 97415 71032
rect 97349 71027 97415 71030
rect 841 70954 907 70957
rect 798 70952 907 70954
rect 798 70896 846 70952
rect 902 70896 907 70952
rect 798 70891 907 70896
rect 798 70848 858 70891
rect 0 70758 858 70848
rect 97533 70818 97599 70821
rect 98200 70818 99000 70848
rect 97533 70816 99000 70818
rect 97533 70760 97538 70816
rect 97594 70760 99000 70816
rect 97533 70758 99000 70760
rect 0 70728 800 70758
rect 97533 70755 97599 70758
rect 4870 70752 5186 70753
rect 4870 70688 4876 70752
rect 4940 70688 4956 70752
rect 5020 70688 5036 70752
rect 5100 70688 5116 70752
rect 5180 70688 5186 70752
rect 4870 70687 5186 70688
rect 97030 70752 97346 70753
rect 97030 70688 97036 70752
rect 97100 70688 97116 70752
rect 97180 70688 97196 70752
rect 97260 70688 97276 70752
rect 97340 70688 97346 70752
rect 98200 70728 99000 70758
rect 97030 70687 97346 70688
rect 4210 70208 4526 70209
rect 0 70138 800 70168
rect 4210 70144 4216 70208
rect 4280 70144 4296 70208
rect 4360 70144 4376 70208
rect 4440 70144 4456 70208
rect 4520 70144 4526 70208
rect 4210 70143 4526 70144
rect 96370 70208 96686 70209
rect 96370 70144 96376 70208
rect 96440 70144 96456 70208
rect 96520 70144 96536 70208
rect 96600 70144 96616 70208
rect 96680 70144 96686 70208
rect 96370 70143 96686 70144
rect 1301 70138 1367 70141
rect 0 70136 1367 70138
rect 0 70080 1306 70136
rect 1362 70080 1367 70136
rect 0 70078 1367 70080
rect 0 70048 800 70078
rect 1301 70075 1367 70078
rect 97441 70138 97507 70141
rect 98200 70138 99000 70168
rect 97441 70136 99000 70138
rect 97441 70080 97446 70136
rect 97502 70080 99000 70136
rect 97441 70078 99000 70080
rect 97441 70075 97507 70078
rect 98200 70048 99000 70078
rect 1577 70002 1643 70005
rect 97257 70002 97323 70005
rect 1577 70000 8188 70002
rect 1577 69944 1582 70000
rect 1638 69944 8188 70000
rect 1577 69942 8188 69944
rect 91908 70000 97323 70002
rect 91908 69944 97262 70000
rect 97318 69944 97323 70000
rect 91908 69942 97323 69944
rect 1577 69939 1643 69942
rect 97257 69939 97323 69942
rect 4870 69664 5186 69665
rect 4870 69600 4876 69664
rect 4940 69600 4956 69664
rect 5020 69600 5036 69664
rect 5100 69600 5116 69664
rect 5180 69600 5186 69664
rect 4870 69599 5186 69600
rect 97030 69664 97346 69665
rect 97030 69600 97036 69664
rect 97100 69600 97116 69664
rect 97180 69600 97196 69664
rect 97260 69600 97276 69664
rect 97340 69600 97346 69664
rect 97030 69599 97346 69600
rect 4210 69120 4526 69121
rect 4210 69056 4216 69120
rect 4280 69056 4296 69120
rect 4360 69056 4376 69120
rect 4440 69056 4456 69120
rect 4520 69056 4526 69120
rect 4210 69055 4526 69056
rect 96370 69120 96686 69121
rect 96370 69056 96376 69120
rect 96440 69056 96456 69120
rect 96520 69056 96536 69120
rect 96600 69056 96616 69120
rect 96680 69056 96686 69120
rect 96370 69055 96686 69056
rect 97257 68914 97323 68917
rect 91908 68912 97323 68914
rect 0 68778 800 68808
rect 1117 68778 1183 68781
rect 0 68776 1183 68778
rect 0 68720 1122 68776
rect 1178 68720 1183 68776
rect 0 68718 1183 68720
rect 0 68688 800 68718
rect 1117 68715 1183 68718
rect 8342 68645 8402 68884
rect 91908 68856 97262 68912
rect 97318 68856 97323 68912
rect 91908 68854 97323 68856
rect 97257 68851 97323 68854
rect 97441 68778 97507 68781
rect 98200 68778 99000 68808
rect 97441 68776 99000 68778
rect 97441 68720 97446 68776
rect 97502 68720 99000 68776
rect 97441 68718 99000 68720
rect 97441 68715 97507 68718
rect 98200 68688 99000 68718
rect 8293 68640 8402 68645
rect 8293 68584 8298 68640
rect 8354 68584 8402 68640
rect 8293 68582 8402 68584
rect 8293 68579 8359 68582
rect 4870 68576 5186 68577
rect 4870 68512 4876 68576
rect 4940 68512 4956 68576
rect 5020 68512 5036 68576
rect 5100 68512 5116 68576
rect 5180 68512 5186 68576
rect 4870 68511 5186 68512
rect 97030 68576 97346 68577
rect 97030 68512 97036 68576
rect 97100 68512 97116 68576
rect 97180 68512 97196 68576
rect 97260 68512 97276 68576
rect 97340 68512 97346 68576
rect 97030 68511 97346 68512
rect 0 68098 800 68128
rect 1301 68098 1367 68101
rect 0 68096 1367 68098
rect 0 68040 1306 68096
rect 1362 68040 1367 68096
rect 0 68038 1367 68040
rect 0 68008 800 68038
rect 1301 68035 1367 68038
rect 8293 68098 8359 68101
rect 97441 68098 97507 68101
rect 98200 68098 99000 68128
rect 8293 68096 8402 68098
rect 8293 68040 8298 68096
rect 8354 68040 8402 68096
rect 8293 68035 8402 68040
rect 97441 68096 99000 68098
rect 97441 68040 97446 68096
rect 97502 68040 99000 68096
rect 97441 68038 99000 68040
rect 97441 68035 97507 68038
rect 4210 68032 4526 68033
rect 4210 67968 4216 68032
rect 4280 67968 4296 68032
rect 4360 67968 4376 68032
rect 4440 67968 4456 68032
rect 4520 67968 4526 68032
rect 4210 67967 4526 67968
rect 8342 67796 8402 68035
rect 96370 68032 96686 68033
rect 96370 67968 96376 68032
rect 96440 67968 96456 68032
rect 96520 67968 96536 68032
rect 96600 67968 96616 68032
rect 96680 67968 96686 68032
rect 98200 68008 99000 68038
rect 96370 67967 96686 67968
rect 97257 67826 97323 67829
rect 91908 67824 97323 67826
rect 91908 67768 97262 67824
rect 97318 67768 97323 67824
rect 91908 67766 97323 67768
rect 97257 67763 97323 67766
rect 4870 67488 5186 67489
rect 4870 67424 4876 67488
rect 4940 67424 4956 67488
rect 5020 67424 5036 67488
rect 5100 67424 5116 67488
rect 5180 67424 5186 67488
rect 4870 67423 5186 67424
rect 97030 67488 97346 67489
rect 97030 67424 97036 67488
rect 97100 67424 97116 67488
rect 97180 67424 97196 67488
rect 97260 67424 97276 67488
rect 97340 67424 97346 67488
rect 97030 67423 97346 67424
rect 8293 67010 8359 67013
rect 8293 67008 8402 67010
rect 8293 66952 8298 67008
rect 8354 66952 8402 67008
rect 8293 66947 8402 66952
rect 4210 66944 4526 66945
rect 4210 66880 4216 66944
rect 4280 66880 4296 66944
rect 4360 66880 4376 66944
rect 4440 66880 4456 66944
rect 4520 66880 4526 66944
rect 4210 66879 4526 66880
rect 0 66738 800 66768
rect 1301 66738 1367 66741
rect 0 66736 1367 66738
rect 0 66680 1306 66736
rect 1362 66680 1367 66736
rect 8342 66708 8402 66947
rect 96370 66944 96686 66945
rect 96370 66880 96376 66944
rect 96440 66880 96456 66944
rect 96520 66880 96536 66944
rect 96600 66880 96616 66944
rect 96680 66880 96686 66944
rect 96370 66879 96686 66880
rect 97257 66738 97323 66741
rect 91908 66736 97323 66738
rect 0 66678 1367 66680
rect 91908 66680 97262 66736
rect 97318 66680 97323 66736
rect 91908 66678 97323 66680
rect 0 66648 800 66678
rect 1301 66675 1367 66678
rect 97257 66675 97323 66678
rect 97441 66738 97507 66741
rect 98200 66738 99000 66768
rect 97441 66736 99000 66738
rect 97441 66680 97446 66736
rect 97502 66680 99000 66736
rect 97441 66678 99000 66680
rect 97441 66675 97507 66678
rect 98200 66648 99000 66678
rect 4870 66400 5186 66401
rect 4870 66336 4876 66400
rect 4940 66336 4956 66400
rect 5020 66336 5036 66400
rect 5100 66336 5116 66400
rect 5180 66336 5186 66400
rect 4870 66335 5186 66336
rect 97030 66400 97346 66401
rect 97030 66336 97036 66400
rect 97100 66336 97116 66400
rect 97180 66336 97196 66400
rect 97260 66336 97276 66400
rect 97340 66336 97346 66400
rect 97030 66335 97346 66336
rect 4210 65856 4526 65857
rect 4210 65792 4216 65856
rect 4280 65792 4296 65856
rect 4360 65792 4376 65856
rect 4440 65792 4456 65856
rect 4520 65792 4526 65856
rect 4210 65791 4526 65792
rect 96370 65856 96686 65857
rect 96370 65792 96376 65856
rect 96440 65792 96456 65856
rect 96520 65792 96536 65856
rect 96600 65792 96616 65856
rect 96680 65792 96686 65856
rect 96370 65791 96686 65792
rect 8293 65786 8359 65789
rect 8293 65784 8402 65786
rect 8293 65728 8298 65784
rect 8354 65728 8402 65784
rect 8293 65723 8402 65728
rect 8342 65620 8402 65723
rect 97257 65650 97323 65653
rect 91908 65648 97323 65650
rect 91908 65592 97262 65648
rect 97318 65592 97323 65648
rect 91908 65590 97323 65592
rect 97257 65587 97323 65590
rect 0 65378 800 65408
rect 1117 65378 1183 65381
rect 0 65376 1183 65378
rect 0 65320 1122 65376
rect 1178 65320 1183 65376
rect 0 65318 1183 65320
rect 0 65288 800 65318
rect 1117 65315 1183 65318
rect 97441 65378 97507 65381
rect 98200 65378 99000 65408
rect 97441 65376 99000 65378
rect 97441 65320 97446 65376
rect 97502 65320 99000 65376
rect 97441 65318 99000 65320
rect 97441 65315 97507 65318
rect 4870 65312 5186 65313
rect 4870 65248 4876 65312
rect 4940 65248 4956 65312
rect 5020 65248 5036 65312
rect 5100 65248 5116 65312
rect 5180 65248 5186 65312
rect 4870 65247 5186 65248
rect 97030 65312 97346 65313
rect 97030 65248 97036 65312
rect 97100 65248 97116 65312
rect 97180 65248 97196 65312
rect 97260 65248 97276 65312
rect 97340 65248 97346 65312
rect 98200 65288 99000 65318
rect 97030 65247 97346 65248
rect 4210 64768 4526 64769
rect 0 64698 800 64728
rect 4210 64704 4216 64768
rect 4280 64704 4296 64768
rect 4360 64704 4376 64768
rect 4440 64704 4456 64768
rect 4520 64704 4526 64768
rect 4210 64703 4526 64704
rect 96370 64768 96686 64769
rect 96370 64704 96376 64768
rect 96440 64704 96456 64768
rect 96520 64704 96536 64768
rect 96600 64704 96616 64768
rect 96680 64704 96686 64768
rect 96370 64703 96686 64704
rect 1301 64698 1367 64701
rect 0 64696 1367 64698
rect 0 64640 1306 64696
rect 1362 64640 1367 64696
rect 0 64638 1367 64640
rect 0 64608 800 64638
rect 1301 64635 1367 64638
rect 97441 64698 97507 64701
rect 98200 64698 99000 64728
rect 97441 64696 99000 64698
rect 97441 64640 97446 64696
rect 97502 64640 99000 64696
rect 97441 64638 99000 64640
rect 97441 64635 97507 64638
rect 98200 64608 99000 64638
rect 1669 64562 1735 64565
rect 97257 64562 97323 64565
rect 1669 64560 8188 64562
rect 1669 64504 1674 64560
rect 1730 64504 8188 64560
rect 1669 64502 8188 64504
rect 91908 64560 97323 64562
rect 91908 64504 97262 64560
rect 97318 64504 97323 64560
rect 91908 64502 97323 64504
rect 1669 64499 1735 64502
rect 97257 64499 97323 64502
rect 4870 64224 5186 64225
rect 4870 64160 4876 64224
rect 4940 64160 4956 64224
rect 5020 64160 5036 64224
rect 5100 64160 5116 64224
rect 5180 64160 5186 64224
rect 4870 64159 5186 64160
rect 97030 64224 97346 64225
rect 97030 64160 97036 64224
rect 97100 64160 97116 64224
rect 97180 64160 97196 64224
rect 97260 64160 97276 64224
rect 97340 64160 97346 64224
rect 97030 64159 97346 64160
rect 4210 63680 4526 63681
rect 4210 63616 4216 63680
rect 4280 63616 4296 63680
rect 4360 63616 4376 63680
rect 4440 63616 4456 63680
rect 4520 63616 4526 63680
rect 4210 63615 4526 63616
rect 96370 63680 96686 63681
rect 96370 63616 96376 63680
rect 96440 63616 96456 63680
rect 96520 63616 96536 63680
rect 96600 63616 96616 63680
rect 96680 63616 96686 63680
rect 96370 63615 96686 63616
rect 97257 63474 97323 63477
rect 91908 63472 97323 63474
rect 0 63338 800 63368
rect 1117 63338 1183 63341
rect 0 63336 1183 63338
rect 0 63280 1122 63336
rect 1178 63280 1183 63336
rect 0 63278 1183 63280
rect 0 63248 800 63278
rect 1117 63275 1183 63278
rect 8342 63205 8402 63444
rect 91908 63416 97262 63472
rect 97318 63416 97323 63472
rect 91908 63414 97323 63416
rect 97257 63411 97323 63414
rect 97441 63338 97507 63341
rect 98200 63338 99000 63368
rect 97441 63336 99000 63338
rect 97441 63280 97446 63336
rect 97502 63280 99000 63336
rect 97441 63278 99000 63280
rect 97441 63275 97507 63278
rect 98200 63248 99000 63278
rect 8293 63200 8402 63205
rect 8293 63144 8298 63200
rect 8354 63144 8402 63200
rect 8293 63142 8402 63144
rect 8293 63139 8359 63142
rect 4870 63136 5186 63137
rect 4870 63072 4876 63136
rect 4940 63072 4956 63136
rect 5020 63072 5036 63136
rect 5100 63072 5116 63136
rect 5180 63072 5186 63136
rect 4870 63071 5186 63072
rect 97030 63136 97346 63137
rect 97030 63072 97036 63136
rect 97100 63072 97116 63136
rect 97180 63072 97196 63136
rect 97260 63072 97276 63136
rect 97340 63072 97346 63136
rect 97030 63071 97346 63072
rect 0 62658 800 62688
rect 1301 62658 1367 62661
rect 0 62656 1367 62658
rect 0 62600 1306 62656
rect 1362 62600 1367 62656
rect 0 62598 1367 62600
rect 0 62568 800 62598
rect 1301 62595 1367 62598
rect 8293 62658 8359 62661
rect 97441 62658 97507 62661
rect 98200 62658 99000 62688
rect 8293 62656 8402 62658
rect 8293 62600 8298 62656
rect 8354 62600 8402 62656
rect 8293 62595 8402 62600
rect 97441 62656 99000 62658
rect 97441 62600 97446 62656
rect 97502 62600 99000 62656
rect 97441 62598 99000 62600
rect 97441 62595 97507 62598
rect 4210 62592 4526 62593
rect 4210 62528 4216 62592
rect 4280 62528 4296 62592
rect 4360 62528 4376 62592
rect 4440 62528 4456 62592
rect 4520 62528 4526 62592
rect 4210 62527 4526 62528
rect 8342 62356 8402 62595
rect 96370 62592 96686 62593
rect 96370 62528 96376 62592
rect 96440 62528 96456 62592
rect 96520 62528 96536 62592
rect 96600 62528 96616 62592
rect 96680 62528 96686 62592
rect 98200 62568 99000 62598
rect 96370 62527 96686 62528
rect 97257 62386 97323 62389
rect 91908 62384 97323 62386
rect 91908 62328 97262 62384
rect 97318 62328 97323 62384
rect 91908 62326 97323 62328
rect 97257 62323 97323 62326
rect 4870 62048 5186 62049
rect 4870 61984 4876 62048
rect 4940 61984 4956 62048
rect 5020 61984 5036 62048
rect 5100 61984 5116 62048
rect 5180 61984 5186 62048
rect 4870 61983 5186 61984
rect 97030 62048 97346 62049
rect 97030 61984 97036 62048
rect 97100 61984 97116 62048
rect 97180 61984 97196 62048
rect 97260 61984 97276 62048
rect 97340 61984 97346 62048
rect 97030 61983 97346 61984
rect 8293 61570 8359 61573
rect 8293 61568 8402 61570
rect 8293 61512 8298 61568
rect 8354 61512 8402 61568
rect 8293 61507 8402 61512
rect 4210 61504 4526 61505
rect 4210 61440 4216 61504
rect 4280 61440 4296 61504
rect 4360 61440 4376 61504
rect 4440 61440 4456 61504
rect 4520 61440 4526 61504
rect 4210 61439 4526 61440
rect 0 61298 800 61328
rect 1301 61298 1367 61301
rect 0 61296 1367 61298
rect 0 61240 1306 61296
rect 1362 61240 1367 61296
rect 8342 61268 8402 61507
rect 96370 61504 96686 61505
rect 96370 61440 96376 61504
rect 96440 61440 96456 61504
rect 96520 61440 96536 61504
rect 96600 61440 96616 61504
rect 96680 61440 96686 61504
rect 96370 61439 96686 61440
rect 97257 61298 97323 61301
rect 91908 61296 97323 61298
rect 0 61238 1367 61240
rect 91908 61240 97262 61296
rect 97318 61240 97323 61296
rect 91908 61238 97323 61240
rect 0 61208 800 61238
rect 1301 61235 1367 61238
rect 97257 61235 97323 61238
rect 97441 61298 97507 61301
rect 98200 61298 99000 61328
rect 97441 61296 99000 61298
rect 97441 61240 97446 61296
rect 97502 61240 99000 61296
rect 97441 61238 99000 61240
rect 97441 61235 97507 61238
rect 98200 61208 99000 61238
rect 4870 60960 5186 60961
rect 4870 60896 4876 60960
rect 4940 60896 4956 60960
rect 5020 60896 5036 60960
rect 5100 60896 5116 60960
rect 5180 60896 5186 60960
rect 4870 60895 5186 60896
rect 97030 60960 97346 60961
rect 97030 60896 97036 60960
rect 97100 60896 97116 60960
rect 97180 60896 97196 60960
rect 97260 60896 97276 60960
rect 97340 60896 97346 60960
rect 97030 60895 97346 60896
rect 4210 60416 4526 60417
rect 4210 60352 4216 60416
rect 4280 60352 4296 60416
rect 4360 60352 4376 60416
rect 4440 60352 4456 60416
rect 4520 60352 4526 60416
rect 4210 60351 4526 60352
rect 96370 60416 96686 60417
rect 96370 60352 96376 60416
rect 96440 60352 96456 60416
rect 96520 60352 96536 60416
rect 96600 60352 96616 60416
rect 96680 60352 96686 60416
rect 96370 60351 96686 60352
rect 8293 60346 8359 60349
rect 8293 60344 8402 60346
rect 8293 60288 8298 60344
rect 8354 60288 8402 60344
rect 8293 60283 8402 60288
rect 8342 60180 8402 60283
rect 97257 60210 97323 60213
rect 91908 60208 97323 60210
rect 91908 60152 97262 60208
rect 97318 60152 97323 60208
rect 91908 60150 97323 60152
rect 97257 60147 97323 60150
rect 0 59938 800 59968
rect 1209 59938 1275 59941
rect 0 59936 1275 59938
rect 0 59880 1214 59936
rect 1270 59880 1275 59936
rect 0 59878 1275 59880
rect 0 59848 800 59878
rect 1209 59875 1275 59878
rect 97441 59938 97507 59941
rect 98200 59938 99000 59968
rect 97441 59936 99000 59938
rect 97441 59880 97446 59936
rect 97502 59880 99000 59936
rect 97441 59878 99000 59880
rect 97441 59875 97507 59878
rect 4870 59872 5186 59873
rect 4870 59808 4876 59872
rect 4940 59808 4956 59872
rect 5020 59808 5036 59872
rect 5100 59808 5116 59872
rect 5180 59808 5186 59872
rect 4870 59807 5186 59808
rect 97030 59872 97346 59873
rect 97030 59808 97036 59872
rect 97100 59808 97116 59872
rect 97180 59808 97196 59872
rect 97260 59808 97276 59872
rect 97340 59808 97346 59872
rect 98200 59848 99000 59878
rect 97030 59807 97346 59808
rect 4210 59328 4526 59329
rect 0 59258 800 59288
rect 4210 59264 4216 59328
rect 4280 59264 4296 59328
rect 4360 59264 4376 59328
rect 4440 59264 4456 59328
rect 4520 59264 4526 59328
rect 4210 59263 4526 59264
rect 96370 59328 96686 59329
rect 96370 59264 96376 59328
rect 96440 59264 96456 59328
rect 96520 59264 96536 59328
rect 96600 59264 96616 59328
rect 96680 59264 96686 59328
rect 96370 59263 96686 59264
rect 1209 59258 1275 59261
rect 0 59256 1275 59258
rect 0 59200 1214 59256
rect 1270 59200 1275 59256
rect 0 59198 1275 59200
rect 0 59168 800 59198
rect 1209 59195 1275 59198
rect 97441 59258 97507 59261
rect 98200 59258 99000 59288
rect 97441 59256 99000 59258
rect 97441 59200 97446 59256
rect 97502 59200 99000 59256
rect 97441 59198 99000 59200
rect 97441 59195 97507 59198
rect 98200 59168 99000 59198
rect 1577 59122 1643 59125
rect 97257 59122 97323 59125
rect 1577 59120 8188 59122
rect 1577 59064 1582 59120
rect 1638 59064 8188 59120
rect 1577 59062 8188 59064
rect 91908 59120 97323 59122
rect 91908 59064 97262 59120
rect 97318 59064 97323 59120
rect 91908 59062 97323 59064
rect 1577 59059 1643 59062
rect 97257 59059 97323 59062
rect 4870 58784 5186 58785
rect 4870 58720 4876 58784
rect 4940 58720 4956 58784
rect 5020 58720 5036 58784
rect 5100 58720 5116 58784
rect 5180 58720 5186 58784
rect 4870 58719 5186 58720
rect 97030 58784 97346 58785
rect 97030 58720 97036 58784
rect 97100 58720 97116 58784
rect 97180 58720 97196 58784
rect 97260 58720 97276 58784
rect 97340 58720 97346 58784
rect 97030 58719 97346 58720
rect 4210 58240 4526 58241
rect 4210 58176 4216 58240
rect 4280 58176 4296 58240
rect 4360 58176 4376 58240
rect 4440 58176 4456 58240
rect 4520 58176 4526 58240
rect 4210 58175 4526 58176
rect 96370 58240 96686 58241
rect 96370 58176 96376 58240
rect 96440 58176 96456 58240
rect 96520 58176 96536 58240
rect 96600 58176 96616 58240
rect 96680 58176 96686 58240
rect 96370 58175 96686 58176
rect 1577 58034 1643 58037
rect 97257 58034 97323 58037
rect 1577 58032 8188 58034
rect 1577 57976 1582 58032
rect 1638 57976 8188 58032
rect 1577 57974 8188 57976
rect 91908 58032 97323 58034
rect 91908 57976 97262 58032
rect 97318 57976 97323 58032
rect 91908 57974 97323 57976
rect 1577 57971 1643 57974
rect 97257 57971 97323 57974
rect 0 57898 800 57928
rect 1301 57898 1367 57901
rect 0 57896 1367 57898
rect 0 57840 1306 57896
rect 1362 57840 1367 57896
rect 0 57838 1367 57840
rect 0 57808 800 57838
rect 1301 57835 1367 57838
rect 97441 57898 97507 57901
rect 98200 57898 99000 57928
rect 97441 57896 99000 57898
rect 97441 57840 97446 57896
rect 97502 57840 99000 57896
rect 97441 57838 99000 57840
rect 97441 57835 97507 57838
rect 98200 57808 99000 57838
rect 4870 57696 5186 57697
rect 4870 57632 4876 57696
rect 4940 57632 4956 57696
rect 5020 57632 5036 57696
rect 5100 57632 5116 57696
rect 5180 57632 5186 57696
rect 4870 57631 5186 57632
rect 97030 57696 97346 57697
rect 97030 57632 97036 57696
rect 97100 57632 97116 57696
rect 97180 57632 97196 57696
rect 97260 57632 97276 57696
rect 97340 57632 97346 57696
rect 97030 57631 97346 57632
rect 0 57218 800 57248
rect 1301 57218 1367 57221
rect 0 57216 1367 57218
rect 0 57160 1306 57216
rect 1362 57160 1367 57216
rect 0 57158 1367 57160
rect 0 57128 800 57158
rect 1301 57155 1367 57158
rect 8293 57218 8359 57221
rect 97441 57218 97507 57221
rect 98200 57218 99000 57248
rect 8293 57216 8402 57218
rect 8293 57160 8298 57216
rect 8354 57160 8402 57216
rect 8293 57155 8402 57160
rect 97441 57216 99000 57218
rect 97441 57160 97446 57216
rect 97502 57160 99000 57216
rect 97441 57158 99000 57160
rect 97441 57155 97507 57158
rect 4210 57152 4526 57153
rect 4210 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4526 57152
rect 4210 57087 4526 57088
rect 8342 56916 8402 57155
rect 96370 57152 96686 57153
rect 96370 57088 96376 57152
rect 96440 57088 96456 57152
rect 96520 57088 96536 57152
rect 96600 57088 96616 57152
rect 96680 57088 96686 57152
rect 98200 57128 99000 57158
rect 96370 57087 96686 57088
rect 97257 56946 97323 56949
rect 91908 56944 97323 56946
rect 91908 56888 97262 56944
rect 97318 56888 97323 56944
rect 91908 56886 97323 56888
rect 97257 56883 97323 56886
rect 4870 56608 5186 56609
rect 4870 56544 4876 56608
rect 4940 56544 4956 56608
rect 5020 56544 5036 56608
rect 5100 56544 5116 56608
rect 5180 56544 5186 56608
rect 4870 56543 5186 56544
rect 97030 56608 97346 56609
rect 97030 56544 97036 56608
rect 97100 56544 97116 56608
rect 97180 56544 97196 56608
rect 97260 56544 97276 56608
rect 97340 56544 97346 56608
rect 97030 56543 97346 56544
rect 8293 56130 8359 56133
rect 8293 56128 8402 56130
rect 8293 56072 8298 56128
rect 8354 56072 8402 56128
rect 8293 56067 8402 56072
rect 4210 56064 4526 56065
rect 4210 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4526 56064
rect 4210 55999 4526 56000
rect 0 55858 800 55888
rect 1301 55858 1367 55861
rect 0 55856 1367 55858
rect 0 55800 1306 55856
rect 1362 55800 1367 55856
rect 8342 55828 8402 56067
rect 96370 56064 96686 56065
rect 96370 56000 96376 56064
rect 96440 56000 96456 56064
rect 96520 56000 96536 56064
rect 96600 56000 96616 56064
rect 96680 56000 96686 56064
rect 96370 55999 96686 56000
rect 97257 55858 97323 55861
rect 91908 55856 97323 55858
rect 0 55798 1367 55800
rect 91908 55800 97262 55856
rect 97318 55800 97323 55856
rect 91908 55798 97323 55800
rect 0 55768 800 55798
rect 1301 55795 1367 55798
rect 97257 55795 97323 55798
rect 97441 55858 97507 55861
rect 98200 55858 99000 55888
rect 97441 55856 99000 55858
rect 97441 55800 97446 55856
rect 97502 55800 99000 55856
rect 97441 55798 99000 55800
rect 97441 55795 97507 55798
rect 98200 55768 99000 55798
rect 4870 55520 5186 55521
rect 4870 55456 4876 55520
rect 4940 55456 4956 55520
rect 5020 55456 5036 55520
rect 5100 55456 5116 55520
rect 5180 55456 5186 55520
rect 4870 55455 5186 55456
rect 97030 55520 97346 55521
rect 97030 55456 97036 55520
rect 97100 55456 97116 55520
rect 97180 55456 97196 55520
rect 97260 55456 97276 55520
rect 97340 55456 97346 55520
rect 97030 55455 97346 55456
rect 4210 54976 4526 54977
rect 4210 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4526 54976
rect 4210 54911 4526 54912
rect 96370 54976 96686 54977
rect 96370 54912 96376 54976
rect 96440 54912 96456 54976
rect 96520 54912 96536 54976
rect 96600 54912 96616 54976
rect 96680 54912 96686 54976
rect 96370 54911 96686 54912
rect 8293 54906 8359 54909
rect 8293 54904 8402 54906
rect 8293 54848 8298 54904
rect 8354 54848 8402 54904
rect 8293 54843 8402 54848
rect 8342 54740 8402 54843
rect 97257 54770 97323 54773
rect 91908 54768 97323 54770
rect 91908 54712 97262 54768
rect 97318 54712 97323 54768
rect 91908 54710 97323 54712
rect 97257 54707 97323 54710
rect 0 54498 800 54528
rect 1301 54498 1367 54501
rect 0 54496 1367 54498
rect 0 54440 1306 54496
rect 1362 54440 1367 54496
rect 0 54438 1367 54440
rect 0 54408 800 54438
rect 1301 54435 1367 54438
rect 97441 54498 97507 54501
rect 98200 54498 99000 54528
rect 97441 54496 99000 54498
rect 97441 54440 97446 54496
rect 97502 54440 99000 54496
rect 97441 54438 99000 54440
rect 97441 54435 97507 54438
rect 4870 54432 5186 54433
rect 4870 54368 4876 54432
rect 4940 54368 4956 54432
rect 5020 54368 5036 54432
rect 5100 54368 5116 54432
rect 5180 54368 5186 54432
rect 4870 54367 5186 54368
rect 97030 54432 97346 54433
rect 97030 54368 97036 54432
rect 97100 54368 97116 54432
rect 97180 54368 97196 54432
rect 97260 54368 97276 54432
rect 97340 54368 97346 54432
rect 98200 54408 99000 54438
rect 97030 54367 97346 54368
rect 4210 53888 4526 53889
rect 0 53818 800 53848
rect 4210 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4526 53888
rect 4210 53823 4526 53824
rect 96370 53888 96686 53889
rect 96370 53824 96376 53888
rect 96440 53824 96456 53888
rect 96520 53824 96536 53888
rect 96600 53824 96616 53888
rect 96680 53824 96686 53888
rect 96370 53823 96686 53824
rect 1209 53818 1275 53821
rect 0 53816 1275 53818
rect 0 53760 1214 53816
rect 1270 53760 1275 53816
rect 0 53758 1275 53760
rect 0 53728 800 53758
rect 1209 53755 1275 53758
rect 97441 53818 97507 53821
rect 98200 53818 99000 53848
rect 97441 53816 99000 53818
rect 97441 53760 97446 53816
rect 97502 53760 99000 53816
rect 97441 53758 99000 53760
rect 97441 53755 97507 53758
rect 98200 53728 99000 53758
rect 1577 53682 1643 53685
rect 97257 53682 97323 53685
rect 1577 53680 8188 53682
rect 1577 53624 1582 53680
rect 1638 53624 8188 53680
rect 1577 53622 8188 53624
rect 91908 53680 97323 53682
rect 91908 53624 97262 53680
rect 97318 53624 97323 53680
rect 91908 53622 97323 53624
rect 1577 53619 1643 53622
rect 97257 53619 97323 53622
rect 4870 53344 5186 53345
rect 4870 53280 4876 53344
rect 4940 53280 4956 53344
rect 5020 53280 5036 53344
rect 5100 53280 5116 53344
rect 5180 53280 5186 53344
rect 4870 53279 5186 53280
rect 97030 53344 97346 53345
rect 97030 53280 97036 53344
rect 97100 53280 97116 53344
rect 97180 53280 97196 53344
rect 97260 53280 97276 53344
rect 97340 53280 97346 53344
rect 97030 53279 97346 53280
rect 4210 52800 4526 52801
rect 4210 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4526 52800
rect 4210 52735 4526 52736
rect 96370 52800 96686 52801
rect 96370 52736 96376 52800
rect 96440 52736 96456 52800
rect 96520 52736 96536 52800
rect 96600 52736 96616 52800
rect 96680 52736 96686 52800
rect 96370 52735 96686 52736
rect 4870 52256 5186 52257
rect 4870 52192 4876 52256
rect 4940 52192 4956 52256
rect 5020 52192 5036 52256
rect 5100 52192 5116 52256
rect 5180 52192 5186 52256
rect 4870 52191 5186 52192
rect 97030 52256 97346 52257
rect 97030 52192 97036 52256
rect 97100 52192 97116 52256
rect 97180 52192 97196 52256
rect 97260 52192 97276 52256
rect 97340 52192 97346 52256
rect 97030 52191 97346 52192
rect 4210 51712 4526 51713
rect 4210 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4526 51712
rect 4210 51647 4526 51648
rect 96370 51712 96686 51713
rect 96370 51648 96376 51712
rect 96440 51648 96456 51712
rect 96520 51648 96536 51712
rect 96600 51648 96616 51712
rect 96680 51648 96686 51712
rect 96370 51647 96686 51648
rect 4870 51168 5186 51169
rect 4870 51104 4876 51168
rect 4940 51104 4956 51168
rect 5020 51104 5036 51168
rect 5100 51104 5116 51168
rect 5180 51104 5186 51168
rect 4870 51103 5186 51104
rect 97030 51168 97346 51169
rect 97030 51104 97036 51168
rect 97100 51104 97116 51168
rect 97180 51104 97196 51168
rect 97260 51104 97276 51168
rect 97340 51104 97346 51168
rect 97030 51103 97346 51104
rect 4210 50624 4526 50625
rect 4210 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4526 50624
rect 4210 50559 4526 50560
rect 96370 50624 96686 50625
rect 96370 50560 96376 50624
rect 96440 50560 96456 50624
rect 96520 50560 96536 50624
rect 96600 50560 96616 50624
rect 96680 50560 96686 50624
rect 96370 50559 96686 50560
rect 4870 50080 5186 50081
rect 4870 50016 4876 50080
rect 4940 50016 4956 50080
rect 5020 50016 5036 50080
rect 5100 50016 5116 50080
rect 5180 50016 5186 50080
rect 4870 50015 5186 50016
rect 97030 50080 97346 50081
rect 97030 50016 97036 50080
rect 97100 50016 97116 50080
rect 97180 50016 97196 50080
rect 97260 50016 97276 50080
rect 97340 50016 97346 50080
rect 97030 50015 97346 50016
rect 4210 49536 4526 49537
rect 4210 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4526 49536
rect 4210 49471 4526 49472
rect 96370 49536 96686 49537
rect 96370 49472 96376 49536
rect 96440 49472 96456 49536
rect 96520 49472 96536 49536
rect 96600 49472 96616 49536
rect 96680 49472 96686 49536
rect 96370 49471 96686 49472
rect 4870 48992 5186 48993
rect 4870 48928 4876 48992
rect 4940 48928 4956 48992
rect 5020 48928 5036 48992
rect 5100 48928 5116 48992
rect 5180 48928 5186 48992
rect 4870 48927 5186 48928
rect 97030 48992 97346 48993
rect 97030 48928 97036 48992
rect 97100 48928 97116 48992
rect 97180 48928 97196 48992
rect 97260 48928 97276 48992
rect 97340 48928 97346 48992
rect 97030 48927 97346 48928
rect 4210 48448 4526 48449
rect 0 48378 800 48408
rect 4210 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4526 48448
rect 4210 48383 4526 48384
rect 96370 48448 96686 48449
rect 96370 48384 96376 48448
rect 96440 48384 96456 48448
rect 96520 48384 96536 48448
rect 96600 48384 96616 48448
rect 96680 48384 96686 48448
rect 96370 48383 96686 48384
rect 1209 48378 1275 48381
rect 0 48376 1275 48378
rect 0 48320 1214 48376
rect 1270 48320 1275 48376
rect 0 48318 1275 48320
rect 0 48288 800 48318
rect 1209 48315 1275 48318
rect 4870 47904 5186 47905
rect 4870 47840 4876 47904
rect 4940 47840 4956 47904
rect 5020 47840 5036 47904
rect 5100 47840 5116 47904
rect 5180 47840 5186 47904
rect 4870 47839 5186 47840
rect 97030 47904 97346 47905
rect 97030 47840 97036 47904
rect 97100 47840 97116 47904
rect 97180 47840 97196 47904
rect 97260 47840 97276 47904
rect 97340 47840 97346 47904
rect 97030 47839 97346 47840
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 96370 47360 96686 47361
rect 96370 47296 96376 47360
rect 96440 47296 96456 47360
rect 96520 47296 96536 47360
rect 96600 47296 96616 47360
rect 96680 47296 96686 47360
rect 96370 47295 96686 47296
rect 4870 46816 5186 46817
rect 4870 46752 4876 46816
rect 4940 46752 4956 46816
rect 5020 46752 5036 46816
rect 5100 46752 5116 46816
rect 5180 46752 5186 46816
rect 4870 46751 5186 46752
rect 97030 46816 97346 46817
rect 97030 46752 97036 46816
rect 97100 46752 97116 46816
rect 97180 46752 97196 46816
rect 97260 46752 97276 46816
rect 97340 46752 97346 46816
rect 97030 46751 97346 46752
rect 4210 46272 4526 46273
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 96370 46272 96686 46273
rect 96370 46208 96376 46272
rect 96440 46208 96456 46272
rect 96520 46208 96536 46272
rect 96600 46208 96616 46272
rect 96680 46208 96686 46272
rect 96370 46207 96686 46208
rect 841 45794 907 45797
rect 798 45792 907 45794
rect 798 45736 846 45792
rect 902 45736 907 45792
rect 798 45731 907 45736
rect 798 45688 858 45731
rect 0 45598 858 45688
rect 4870 45728 5186 45729
rect 4870 45664 4876 45728
rect 4940 45664 4956 45728
rect 5020 45664 5036 45728
rect 5100 45664 5116 45728
rect 5180 45664 5186 45728
rect 4870 45663 5186 45664
rect 97030 45728 97346 45729
rect 97030 45664 97036 45728
rect 97100 45664 97116 45728
rect 97180 45664 97196 45728
rect 97260 45664 97276 45728
rect 97340 45664 97346 45728
rect 97030 45663 97346 45664
rect 97533 45658 97599 45661
rect 98200 45658 99000 45688
rect 97533 45656 99000 45658
rect 97533 45600 97538 45656
rect 97594 45600 99000 45656
rect 97533 45598 99000 45600
rect 0 45568 800 45598
rect 97533 45595 97599 45598
rect 98200 45568 99000 45598
rect 1669 45386 1735 45389
rect 97441 45386 97507 45389
rect 1669 45384 8188 45386
rect 1669 45328 1674 45384
rect 1730 45328 8188 45384
rect 1669 45326 8188 45328
rect 91908 45384 97507 45386
rect 91908 45328 97446 45384
rect 97502 45328 97507 45384
rect 91908 45326 97507 45328
rect 1669 45323 1735 45326
rect 97441 45323 97507 45326
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 96370 45184 96686 45185
rect 96370 45120 96376 45184
rect 96440 45120 96456 45184
rect 96520 45120 96536 45184
rect 96600 45120 96616 45184
rect 96680 45120 96686 45184
rect 96370 45119 96686 45120
rect 4870 44640 5186 44641
rect 4870 44576 4876 44640
rect 4940 44576 4956 44640
rect 5020 44576 5036 44640
rect 5100 44576 5116 44640
rect 5180 44576 5186 44640
rect 4870 44575 5186 44576
rect 97030 44640 97346 44641
rect 97030 44576 97036 44640
rect 97100 44576 97116 44640
rect 97180 44576 97196 44640
rect 97260 44576 97276 44640
rect 97340 44576 97346 44640
rect 97030 44575 97346 44576
rect 841 44434 907 44437
rect 798 44432 907 44434
rect 798 44376 846 44432
rect 902 44376 907 44432
rect 798 44371 907 44376
rect 8293 44434 8359 44437
rect 8293 44432 8402 44434
rect 8293 44376 8298 44432
rect 8354 44376 8402 44432
rect 8293 44371 8402 44376
rect 798 44328 858 44371
rect 0 44238 858 44328
rect 8342 44268 8402 44371
rect 97349 44298 97415 44301
rect 91908 44296 97415 44298
rect 91908 44240 97354 44296
rect 97410 44240 97415 44296
rect 91908 44238 97415 44240
rect 0 44208 800 44238
rect 97349 44235 97415 44238
rect 97533 44298 97599 44301
rect 98200 44298 99000 44328
rect 97533 44296 99000 44298
rect 97533 44240 97538 44296
rect 97594 44240 99000 44296
rect 97533 44238 99000 44240
rect 97533 44235 97599 44238
rect 98200 44208 99000 44238
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 96370 44096 96686 44097
rect 96370 44032 96376 44096
rect 96440 44032 96456 44096
rect 96520 44032 96536 44096
rect 96600 44032 96616 44096
rect 96680 44032 96686 44096
rect 96370 44031 96686 44032
rect 4870 43552 5186 43553
rect 4870 43488 4876 43552
rect 4940 43488 4956 43552
rect 5020 43488 5036 43552
rect 5100 43488 5116 43552
rect 5180 43488 5186 43552
rect 4870 43487 5186 43488
rect 97030 43552 97346 43553
rect 97030 43488 97036 43552
rect 97100 43488 97116 43552
rect 97180 43488 97196 43552
rect 97260 43488 97276 43552
rect 97340 43488 97346 43552
rect 97030 43487 97346 43488
rect 8293 43346 8359 43349
rect 8293 43344 8402 43346
rect 8293 43288 8298 43344
rect 8354 43288 8402 43344
rect 8293 43283 8402 43288
rect 8342 43180 8402 43283
rect 97349 43210 97415 43213
rect 91908 43208 97415 43210
rect 91908 43152 97354 43208
rect 97410 43152 97415 43208
rect 91908 43150 97415 43152
rect 97349 43147 97415 43150
rect 841 43074 907 43077
rect 798 43072 907 43074
rect 798 43016 846 43072
rect 902 43016 907 43072
rect 798 43011 907 43016
rect 798 42968 858 43011
rect 0 42878 858 42968
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 96370 43008 96686 43009
rect 96370 42944 96376 43008
rect 96440 42944 96456 43008
rect 96520 42944 96536 43008
rect 96600 42944 96616 43008
rect 96680 42944 96686 43008
rect 96370 42943 96686 42944
rect 97533 42938 97599 42941
rect 98200 42938 99000 42968
rect 97533 42936 99000 42938
rect 97533 42880 97538 42936
rect 97594 42880 99000 42936
rect 97533 42878 99000 42880
rect 0 42848 800 42878
rect 97533 42875 97599 42878
rect 98200 42848 99000 42878
rect 8293 42666 8359 42669
rect 8293 42664 8402 42666
rect 8293 42608 8298 42664
rect 8354 42608 8402 42664
rect 8293 42603 8402 42608
rect 4870 42464 5186 42465
rect 4870 42400 4876 42464
rect 4940 42400 4956 42464
rect 5020 42400 5036 42464
rect 5100 42400 5116 42464
rect 5180 42400 5186 42464
rect 4870 42399 5186 42400
rect 841 42394 907 42397
rect 798 42392 907 42394
rect 798 42336 846 42392
rect 902 42336 907 42392
rect 798 42331 907 42336
rect 798 42288 858 42331
rect 0 42198 858 42288
rect 0 42168 800 42198
rect 8342 42092 8402 42603
rect 97030 42464 97346 42465
rect 97030 42400 97036 42464
rect 97100 42400 97116 42464
rect 97180 42400 97196 42464
rect 97260 42400 97276 42464
rect 97340 42400 97346 42464
rect 97030 42399 97346 42400
rect 97533 42258 97599 42261
rect 98200 42258 99000 42288
rect 97533 42256 99000 42258
rect 97533 42200 97538 42256
rect 97594 42200 99000 42256
rect 97533 42198 99000 42200
rect 97533 42195 97599 42198
rect 98200 42168 99000 42198
rect 97441 42122 97507 42125
rect 91908 42120 97507 42122
rect 91908 42064 97446 42120
rect 97502 42064 97507 42120
rect 91908 42062 97507 42064
rect 97441 42059 97507 42062
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 96370 41920 96686 41921
rect 96370 41856 96376 41920
rect 96440 41856 96456 41920
rect 96520 41856 96536 41920
rect 96600 41856 96616 41920
rect 96680 41856 96686 41920
rect 96370 41855 96686 41856
rect 4870 41376 5186 41377
rect 4870 41312 4876 41376
rect 4940 41312 4956 41376
rect 5020 41312 5036 41376
rect 5100 41312 5116 41376
rect 5180 41312 5186 41376
rect 4870 41311 5186 41312
rect 97030 41376 97346 41377
rect 97030 41312 97036 41376
rect 97100 41312 97116 41376
rect 97180 41312 97196 41376
rect 97260 41312 97276 41376
rect 97340 41312 97346 41376
rect 97030 41311 97346 41312
rect 8293 41170 8359 41173
rect 97349 41170 97415 41173
rect 8293 41168 8402 41170
rect 8293 41112 8298 41168
rect 8354 41112 8402 41168
rect 8293 41107 8402 41112
rect 841 41034 907 41037
rect 798 41032 907 41034
rect 798 40976 846 41032
rect 902 40976 907 41032
rect 8342 41004 8402 41107
rect 91878 41168 97415 41170
rect 91878 41112 97354 41168
rect 97410 41112 97415 41168
rect 91878 41110 97415 41112
rect 91878 41004 91938 41110
rect 97349 41107 97415 41110
rect 798 40971 907 40976
rect 798 40928 858 40971
rect 0 40838 858 40928
rect 97533 40898 97599 40901
rect 98200 40898 99000 40928
rect 97533 40896 99000 40898
rect 97533 40840 97538 40896
rect 97594 40840 99000 40896
rect 97533 40838 99000 40840
rect 0 40808 800 40838
rect 97533 40835 97599 40838
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 96370 40832 96686 40833
rect 96370 40768 96376 40832
rect 96440 40768 96456 40832
rect 96520 40768 96536 40832
rect 96600 40768 96616 40832
rect 96680 40768 96686 40832
rect 98200 40808 99000 40838
rect 96370 40767 96686 40768
rect 841 40354 907 40357
rect 798 40352 907 40354
rect 798 40296 846 40352
rect 902 40296 907 40352
rect 798 40291 907 40296
rect 798 40248 858 40291
rect 0 40158 858 40248
rect 4870 40288 5186 40289
rect 4870 40224 4876 40288
rect 4940 40224 4956 40288
rect 5020 40224 5036 40288
rect 5100 40224 5116 40288
rect 5180 40224 5186 40288
rect 4870 40223 5186 40224
rect 97030 40288 97346 40289
rect 97030 40224 97036 40288
rect 97100 40224 97116 40288
rect 97180 40224 97196 40288
rect 97260 40224 97276 40288
rect 97340 40224 97346 40288
rect 97030 40223 97346 40224
rect 97533 40218 97599 40221
rect 98200 40218 99000 40248
rect 97533 40216 99000 40218
rect 97533 40160 97538 40216
rect 97594 40160 99000 40216
rect 97533 40158 99000 40160
rect 0 40128 800 40158
rect 97533 40155 97599 40158
rect 98200 40128 99000 40158
rect 1669 39946 1735 39949
rect 97441 39946 97507 39949
rect 1669 39944 8188 39946
rect 1669 39888 1674 39944
rect 1730 39888 8188 39944
rect 1669 39886 8188 39888
rect 91908 39944 97507 39946
rect 91908 39888 97446 39944
rect 97502 39888 97507 39944
rect 91908 39886 97507 39888
rect 1669 39883 1735 39886
rect 97441 39883 97507 39886
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 96370 39744 96686 39745
rect 96370 39680 96376 39744
rect 96440 39680 96456 39744
rect 96520 39680 96536 39744
rect 96600 39680 96616 39744
rect 96680 39680 96686 39744
rect 96370 39679 96686 39680
rect 4870 39200 5186 39201
rect 4870 39136 4876 39200
rect 4940 39136 4956 39200
rect 5020 39136 5036 39200
rect 5100 39136 5116 39200
rect 5180 39136 5186 39200
rect 4870 39135 5186 39136
rect 97030 39200 97346 39201
rect 97030 39136 97036 39200
rect 97100 39136 97116 39200
rect 97180 39136 97196 39200
rect 97260 39136 97276 39200
rect 97340 39136 97346 39200
rect 97030 39135 97346 39136
rect 8293 38994 8359 38997
rect 97349 38994 97415 38997
rect 8293 38992 8402 38994
rect 8293 38936 8298 38992
rect 8354 38936 8402 38992
rect 8293 38931 8402 38936
rect 0 38858 800 38888
rect 0 38768 858 38858
rect 8342 38828 8402 38931
rect 91878 38992 97415 38994
rect 91878 38936 97354 38992
rect 97410 38936 97415 38992
rect 91878 38934 97415 38936
rect 91878 38828 91938 38934
rect 97349 38931 97415 38934
rect 97533 38858 97599 38861
rect 98200 38858 99000 38888
rect 97533 38856 99000 38858
rect 97533 38800 97538 38856
rect 97594 38800 99000 38856
rect 97533 38798 99000 38800
rect 97533 38795 97599 38798
rect 98200 38768 99000 38798
rect 798 38725 858 38768
rect 798 38720 907 38725
rect 798 38664 846 38720
rect 902 38664 907 38720
rect 798 38662 907 38664
rect 841 38659 907 38662
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 96370 38656 96686 38657
rect 96370 38592 96376 38656
rect 96440 38592 96456 38656
rect 96520 38592 96536 38656
rect 96600 38592 96616 38656
rect 96680 38592 96686 38656
rect 96370 38591 96686 38592
rect 4870 38112 5186 38113
rect 4870 38048 4876 38112
rect 4940 38048 4956 38112
rect 5020 38048 5036 38112
rect 5100 38048 5116 38112
rect 5180 38048 5186 38112
rect 4870 38047 5186 38048
rect 97030 38112 97346 38113
rect 97030 38048 97036 38112
rect 97100 38048 97116 38112
rect 97180 38048 97196 38112
rect 97260 38048 97276 38112
rect 97340 38048 97346 38112
rect 97030 38047 97346 38048
rect 8293 37906 8359 37909
rect 97349 37906 97415 37909
rect 8293 37904 8402 37906
rect 8293 37848 8298 37904
rect 8354 37848 8402 37904
rect 8293 37843 8402 37848
rect 8342 37740 8402 37843
rect 91878 37904 97415 37906
rect 91878 37848 97354 37904
rect 97410 37848 97415 37904
rect 91878 37846 97415 37848
rect 91878 37740 91938 37846
rect 97349 37843 97415 37846
rect 841 37634 907 37637
rect 798 37632 907 37634
rect 798 37576 846 37632
rect 902 37576 907 37632
rect 798 37571 907 37576
rect 798 37528 858 37571
rect 0 37438 858 37528
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 96370 37568 96686 37569
rect 96370 37504 96376 37568
rect 96440 37504 96456 37568
rect 96520 37504 96536 37568
rect 96600 37504 96616 37568
rect 96680 37504 96686 37568
rect 96370 37503 96686 37504
rect 97533 37498 97599 37501
rect 98200 37498 99000 37528
rect 97533 37496 99000 37498
rect 97533 37440 97538 37496
rect 97594 37440 99000 37496
rect 97533 37438 99000 37440
rect 0 37408 800 37438
rect 97533 37435 97599 37438
rect 98200 37408 99000 37438
rect 8293 37226 8359 37229
rect 8293 37224 8402 37226
rect 8293 37168 8298 37224
rect 8354 37168 8402 37224
rect 8293 37163 8402 37168
rect 4870 37024 5186 37025
rect 4870 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5186 37024
rect 4870 36959 5186 36960
rect 841 36954 907 36957
rect 798 36952 907 36954
rect 798 36896 846 36952
rect 902 36896 907 36952
rect 798 36891 907 36896
rect 798 36848 858 36891
rect 0 36758 858 36848
rect 0 36728 800 36758
rect 8342 36652 8402 37163
rect 97030 37024 97346 37025
rect 97030 36960 97036 37024
rect 97100 36960 97116 37024
rect 97180 36960 97196 37024
rect 97260 36960 97276 37024
rect 97340 36960 97346 37024
rect 97030 36959 97346 36960
rect 96613 36818 96679 36821
rect 91878 36816 96679 36818
rect 91878 36760 96618 36816
rect 96674 36760 96679 36816
rect 91878 36758 96679 36760
rect 91878 36652 91938 36758
rect 96613 36755 96679 36758
rect 97441 36818 97507 36821
rect 98200 36818 99000 36848
rect 97441 36816 99000 36818
rect 97441 36760 97446 36816
rect 97502 36760 99000 36816
rect 97441 36758 99000 36760
rect 97441 36755 97507 36758
rect 98200 36728 99000 36758
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 96370 36480 96686 36481
rect 96370 36416 96376 36480
rect 96440 36416 96456 36480
rect 96520 36416 96536 36480
rect 96600 36416 96616 36480
rect 96680 36416 96686 36480
rect 96370 36415 96686 36416
rect 4870 35936 5186 35937
rect 4870 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5186 35936
rect 4870 35871 5186 35872
rect 97030 35936 97346 35937
rect 97030 35872 97036 35936
rect 97100 35872 97116 35936
rect 97180 35872 97196 35936
rect 97260 35872 97276 35936
rect 97340 35872 97346 35936
rect 97030 35871 97346 35872
rect 8293 35730 8359 35733
rect 97349 35730 97415 35733
rect 8293 35728 8402 35730
rect 8293 35672 8298 35728
rect 8354 35672 8402 35728
rect 8293 35667 8402 35672
rect 841 35594 907 35597
rect 798 35592 907 35594
rect 798 35536 846 35592
rect 902 35536 907 35592
rect 8342 35564 8402 35667
rect 91878 35728 97415 35730
rect 91878 35672 97354 35728
rect 97410 35672 97415 35728
rect 91878 35670 97415 35672
rect 91878 35564 91938 35670
rect 97349 35667 97415 35670
rect 798 35531 907 35536
rect 798 35488 858 35531
rect 0 35398 858 35488
rect 97533 35458 97599 35461
rect 98200 35458 99000 35488
rect 97533 35456 99000 35458
rect 97533 35400 97538 35456
rect 97594 35400 99000 35456
rect 97533 35398 99000 35400
rect 0 35368 800 35398
rect 97533 35395 97599 35398
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 96370 35392 96686 35393
rect 96370 35328 96376 35392
rect 96440 35328 96456 35392
rect 96520 35328 96536 35392
rect 96600 35328 96616 35392
rect 96680 35328 96686 35392
rect 98200 35368 99000 35398
rect 96370 35327 96686 35328
rect 841 34914 907 34917
rect 798 34912 907 34914
rect 798 34856 846 34912
rect 902 34856 907 34912
rect 798 34851 907 34856
rect 798 34808 858 34851
rect 0 34718 858 34808
rect 4870 34848 5186 34849
rect 4870 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5186 34848
rect 4870 34783 5186 34784
rect 97030 34848 97346 34849
rect 97030 34784 97036 34848
rect 97100 34784 97116 34848
rect 97180 34784 97196 34848
rect 97260 34784 97276 34848
rect 97340 34784 97346 34848
rect 97030 34783 97346 34784
rect 97533 34778 97599 34781
rect 98200 34778 99000 34808
rect 97533 34776 99000 34778
rect 97533 34720 97538 34776
rect 97594 34720 99000 34776
rect 97533 34718 99000 34720
rect 0 34688 800 34718
rect 97533 34715 97599 34718
rect 98200 34688 99000 34718
rect 1669 34506 1735 34509
rect 97441 34506 97507 34509
rect 1669 34504 8188 34506
rect 1669 34448 1674 34504
rect 1730 34448 8188 34504
rect 1669 34446 8188 34448
rect 91908 34504 97507 34506
rect 91908 34448 97446 34504
rect 97502 34448 97507 34504
rect 91908 34446 97507 34448
rect 1669 34443 1735 34446
rect 97441 34443 97507 34446
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 96370 34304 96686 34305
rect 96370 34240 96376 34304
rect 96440 34240 96456 34304
rect 96520 34240 96536 34304
rect 96600 34240 96616 34304
rect 96680 34240 96686 34304
rect 96370 34239 96686 34240
rect 4870 33760 5186 33761
rect 4870 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5186 33760
rect 4870 33695 5186 33696
rect 97030 33760 97346 33761
rect 97030 33696 97036 33760
rect 97100 33696 97116 33760
rect 97180 33696 97196 33760
rect 97260 33696 97276 33760
rect 97340 33696 97346 33760
rect 97030 33695 97346 33696
rect 8293 33554 8359 33557
rect 97349 33554 97415 33557
rect 8293 33552 8402 33554
rect 8293 33496 8298 33552
rect 8354 33496 8402 33552
rect 8293 33491 8402 33496
rect 0 33418 800 33448
rect 0 33328 858 33418
rect 8342 33388 8402 33491
rect 91878 33552 97415 33554
rect 91878 33496 97354 33552
rect 97410 33496 97415 33552
rect 91878 33494 97415 33496
rect 91878 33388 91938 33494
rect 97349 33491 97415 33494
rect 97533 33418 97599 33421
rect 98200 33418 99000 33448
rect 97533 33416 99000 33418
rect 97533 33360 97538 33416
rect 97594 33360 99000 33416
rect 97533 33358 99000 33360
rect 97533 33355 97599 33358
rect 98200 33328 99000 33358
rect 798 33285 858 33328
rect 798 33280 907 33285
rect 798 33224 846 33280
rect 902 33224 907 33280
rect 798 33222 907 33224
rect 841 33219 907 33222
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 96370 33216 96686 33217
rect 96370 33152 96376 33216
rect 96440 33152 96456 33216
rect 96520 33152 96536 33216
rect 96600 33152 96616 33216
rect 96680 33152 96686 33216
rect 96370 33151 96686 33152
rect 4870 32672 5186 32673
rect 4870 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5186 32672
rect 4870 32607 5186 32608
rect 97030 32672 97346 32673
rect 97030 32608 97036 32672
rect 97100 32608 97116 32672
rect 97180 32608 97196 32672
rect 97260 32608 97276 32672
rect 97340 32608 97346 32672
rect 97030 32607 97346 32608
rect 8293 32466 8359 32469
rect 97257 32466 97323 32469
rect 8293 32464 8402 32466
rect 8293 32408 8298 32464
rect 8354 32408 8402 32464
rect 8293 32403 8402 32408
rect 8342 32300 8402 32403
rect 91878 32464 97323 32466
rect 91878 32408 97262 32464
rect 97318 32408 97323 32464
rect 91878 32406 97323 32408
rect 91878 32300 91938 32406
rect 97257 32403 97323 32406
rect 841 32194 907 32197
rect 798 32192 907 32194
rect 798 32136 846 32192
rect 902 32136 907 32192
rect 798 32131 907 32136
rect 798 32088 858 32131
rect 0 31998 858 32088
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 96370 32128 96686 32129
rect 96370 32064 96376 32128
rect 96440 32064 96456 32128
rect 96520 32064 96536 32128
rect 96600 32064 96616 32128
rect 96680 32064 96686 32128
rect 96370 32063 96686 32064
rect 97441 32058 97507 32061
rect 98200 32058 99000 32088
rect 97441 32056 99000 32058
rect 97441 32000 97446 32056
rect 97502 32000 99000 32056
rect 97441 31998 99000 32000
rect 0 31968 800 31998
rect 97441 31995 97507 31998
rect 98200 31968 99000 31998
rect 4870 31584 5186 31585
rect 4870 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5186 31584
rect 4870 31519 5186 31520
rect 97030 31584 97346 31585
rect 97030 31520 97036 31584
rect 97100 31520 97116 31584
rect 97180 31520 97196 31584
rect 97260 31520 97276 31584
rect 97340 31520 97346 31584
rect 97030 31519 97346 31520
rect 841 31514 907 31517
rect 798 31512 907 31514
rect 798 31456 846 31512
rect 902 31456 907 31512
rect 798 31451 907 31456
rect 798 31408 858 31451
rect 0 31318 858 31408
rect 96613 31378 96679 31381
rect 91878 31376 96679 31378
rect 91878 31320 96618 31376
rect 96674 31320 96679 31376
rect 91878 31318 96679 31320
rect 0 31288 800 31318
rect 1669 31242 1735 31245
rect 1669 31240 8188 31242
rect 1669 31184 1674 31240
rect 1730 31184 8188 31240
rect 91878 31212 91938 31318
rect 96613 31315 96679 31318
rect 97533 31378 97599 31381
rect 98200 31378 99000 31408
rect 97533 31376 99000 31378
rect 97533 31320 97538 31376
rect 97594 31320 99000 31376
rect 97533 31318 99000 31320
rect 97533 31315 97599 31318
rect 98200 31288 99000 31318
rect 1669 31182 8188 31184
rect 1669 31179 1735 31182
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 96370 31040 96686 31041
rect 96370 30976 96376 31040
rect 96440 30976 96456 31040
rect 96520 30976 96536 31040
rect 96600 30976 96616 31040
rect 96680 30976 96686 31040
rect 96370 30975 96686 30976
rect 4870 30496 5186 30497
rect 4870 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5186 30496
rect 4870 30431 5186 30432
rect 97030 30496 97346 30497
rect 97030 30432 97036 30496
rect 97100 30432 97116 30496
rect 97180 30432 97196 30496
rect 97260 30432 97276 30496
rect 97340 30432 97346 30496
rect 97030 30431 97346 30432
rect 8293 30290 8359 30293
rect 97257 30290 97323 30293
rect 8293 30288 8402 30290
rect 8293 30232 8298 30288
rect 8354 30232 8402 30288
rect 8293 30227 8402 30232
rect 841 30154 907 30157
rect 798 30152 907 30154
rect 798 30096 846 30152
rect 902 30096 907 30152
rect 8342 30124 8402 30227
rect 91878 30288 97323 30290
rect 91878 30232 97262 30288
rect 97318 30232 97323 30288
rect 91878 30230 97323 30232
rect 91878 30124 91938 30230
rect 97257 30227 97323 30230
rect 798 30091 907 30096
rect 798 30048 858 30091
rect 0 29958 858 30048
rect 97533 30018 97599 30021
rect 98200 30018 99000 30048
rect 97533 30016 99000 30018
rect 97533 29960 97538 30016
rect 97594 29960 99000 30016
rect 97533 29958 99000 29960
rect 0 29928 800 29958
rect 97533 29955 97599 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 96370 29952 96686 29953
rect 96370 29888 96376 29952
rect 96440 29888 96456 29952
rect 96520 29888 96536 29952
rect 96600 29888 96616 29952
rect 96680 29888 96686 29952
rect 98200 29928 99000 29958
rect 96370 29887 96686 29888
rect 8293 29610 8359 29613
rect 8293 29608 8402 29610
rect 8293 29552 8298 29608
rect 8354 29552 8402 29608
rect 8293 29547 8402 29552
rect 841 29474 907 29477
rect 798 29472 907 29474
rect 798 29416 846 29472
rect 902 29416 907 29472
rect 798 29411 907 29416
rect 798 29368 858 29411
rect 0 29278 858 29368
rect 4870 29408 5186 29409
rect 4870 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5186 29408
rect 4870 29343 5186 29344
rect 0 29248 800 29278
rect 8342 29036 8402 29547
rect 97030 29408 97346 29409
rect 97030 29344 97036 29408
rect 97100 29344 97116 29408
rect 97180 29344 97196 29408
rect 97260 29344 97276 29408
rect 97340 29344 97346 29408
rect 97030 29343 97346 29344
rect 97533 29338 97599 29341
rect 98200 29338 99000 29368
rect 97533 29336 99000 29338
rect 97533 29280 97538 29336
rect 97594 29280 99000 29336
rect 97533 29278 99000 29280
rect 97533 29275 97599 29278
rect 98200 29248 99000 29278
rect 97441 29202 97507 29205
rect 91878 29200 97507 29202
rect 91878 29144 97446 29200
rect 97502 29144 97507 29200
rect 91878 29142 97507 29144
rect 91878 29036 91938 29142
rect 97441 29139 97507 29142
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 96370 28864 96686 28865
rect 96370 28800 96376 28864
rect 96440 28800 96456 28864
rect 96520 28800 96536 28864
rect 96600 28800 96616 28864
rect 96680 28800 96686 28864
rect 96370 28799 96686 28800
rect 4870 28320 5186 28321
rect 4870 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5186 28320
rect 4870 28255 5186 28256
rect 97030 28320 97346 28321
rect 97030 28256 97036 28320
rect 97100 28256 97116 28320
rect 97180 28256 97196 28320
rect 97260 28256 97276 28320
rect 97340 28256 97346 28320
rect 97030 28255 97346 28256
rect 8293 28114 8359 28117
rect 97257 28114 97323 28117
rect 8293 28112 8402 28114
rect 8293 28056 8298 28112
rect 8354 28056 8402 28112
rect 8293 28051 8402 28056
rect 0 27978 800 28008
rect 1301 27978 1367 27981
rect 0 27976 1367 27978
rect 0 27920 1306 27976
rect 1362 27920 1367 27976
rect 8342 27948 8402 28051
rect 91878 28112 97323 28114
rect 91878 28056 97262 28112
rect 97318 28056 97323 28112
rect 91878 28054 97323 28056
rect 91878 27948 91938 28054
rect 97257 28051 97323 28054
rect 97441 27978 97507 27981
rect 98200 27978 99000 28008
rect 97441 27976 99000 27978
rect 0 27918 1367 27920
rect 0 27888 800 27918
rect 1301 27915 1367 27918
rect 97441 27920 97446 27976
rect 97502 27920 99000 27976
rect 97441 27918 99000 27920
rect 97441 27915 97507 27918
rect 98200 27888 99000 27918
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 96370 27776 96686 27777
rect 96370 27712 96376 27776
rect 96440 27712 96456 27776
rect 96520 27712 96536 27776
rect 96600 27712 96616 27776
rect 96680 27712 96686 27776
rect 96370 27711 96686 27712
rect 4870 27232 5186 27233
rect 4870 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5186 27232
rect 4870 27167 5186 27168
rect 97030 27232 97346 27233
rect 97030 27168 97036 27232
rect 97100 27168 97116 27232
rect 97180 27168 97196 27232
rect 97260 27168 97276 27232
rect 97340 27168 97346 27232
rect 97030 27167 97346 27168
rect 8293 27026 8359 27029
rect 97257 27026 97323 27029
rect 8293 27024 8402 27026
rect 8293 26968 8298 27024
rect 8354 26968 8402 27024
rect 8293 26963 8402 26968
rect 8342 26860 8402 26963
rect 91878 27024 97323 27026
rect 91878 26968 97262 27024
rect 97318 26968 97323 27024
rect 91878 26966 97323 26968
rect 91878 26860 91938 26966
rect 97257 26963 97323 26966
rect 4210 26688 4526 26689
rect 0 26618 800 26648
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 96370 26688 96686 26689
rect 96370 26624 96376 26688
rect 96440 26624 96456 26688
rect 96520 26624 96536 26688
rect 96600 26624 96616 26688
rect 96680 26624 96686 26688
rect 96370 26623 96686 26624
rect 1301 26618 1367 26621
rect 0 26616 1367 26618
rect 0 26560 1306 26616
rect 1362 26560 1367 26616
rect 0 26558 1367 26560
rect 0 26528 800 26558
rect 1301 26555 1367 26558
rect 97441 26618 97507 26621
rect 98200 26618 99000 26648
rect 97441 26616 99000 26618
rect 97441 26560 97446 26616
rect 97502 26560 99000 26616
rect 97441 26558 99000 26560
rect 97441 26555 97507 26558
rect 98200 26528 99000 26558
rect 4870 26144 5186 26145
rect 4870 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5186 26144
rect 4870 26079 5186 26080
rect 97030 26144 97346 26145
rect 97030 26080 97036 26144
rect 97100 26080 97116 26144
rect 97180 26080 97196 26144
rect 97260 26080 97276 26144
rect 97340 26080 97346 26144
rect 97030 26079 97346 26080
rect 0 25938 800 25968
rect 1301 25938 1367 25941
rect 96889 25938 96955 25941
rect 0 25936 1367 25938
rect 0 25880 1306 25936
rect 1362 25880 1367 25936
rect 0 25878 1367 25880
rect 0 25848 800 25878
rect 1301 25875 1367 25878
rect 91878 25936 96955 25938
rect 91878 25880 96894 25936
rect 96950 25880 96955 25936
rect 91878 25878 96955 25880
rect 1669 25802 1735 25805
rect 1669 25800 8188 25802
rect 1669 25744 1674 25800
rect 1730 25744 8188 25800
rect 91878 25772 91938 25878
rect 96889 25875 96955 25878
rect 97441 25938 97507 25941
rect 98200 25938 99000 25968
rect 97441 25936 99000 25938
rect 97441 25880 97446 25936
rect 97502 25880 99000 25936
rect 97441 25878 99000 25880
rect 97441 25875 97507 25878
rect 98200 25848 99000 25878
rect 1669 25742 8188 25744
rect 1669 25739 1735 25742
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 96370 25600 96686 25601
rect 96370 25536 96376 25600
rect 96440 25536 96456 25600
rect 96520 25536 96536 25600
rect 96600 25536 96616 25600
rect 96680 25536 96686 25600
rect 96370 25535 96686 25536
rect 4870 25056 5186 25057
rect 4870 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5186 25056
rect 4870 24991 5186 24992
rect 97030 25056 97346 25057
rect 97030 24992 97036 25056
rect 97100 24992 97116 25056
rect 97180 24992 97196 25056
rect 97260 24992 97276 25056
rect 97340 24992 97346 25056
rect 97030 24991 97346 24992
rect 8293 24850 8359 24853
rect 97257 24850 97323 24853
rect 8293 24848 8402 24850
rect 8293 24792 8298 24848
rect 8354 24792 8402 24848
rect 8293 24787 8402 24792
rect 8342 24684 8402 24787
rect 91878 24848 97323 24850
rect 91878 24792 97262 24848
rect 97318 24792 97323 24848
rect 91878 24790 97323 24792
rect 91878 24684 91938 24790
rect 97257 24787 97323 24790
rect 0 24578 800 24608
rect 1301 24578 1367 24581
rect 0 24576 1367 24578
rect 0 24520 1306 24576
rect 1362 24520 1367 24576
rect 0 24518 1367 24520
rect 0 24488 800 24518
rect 1301 24515 1367 24518
rect 97441 24578 97507 24581
rect 98200 24578 99000 24608
rect 97441 24576 99000 24578
rect 97441 24520 97446 24576
rect 97502 24520 99000 24576
rect 97441 24518 99000 24520
rect 97441 24515 97507 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 96370 24512 96686 24513
rect 96370 24448 96376 24512
rect 96440 24448 96456 24512
rect 96520 24448 96536 24512
rect 96600 24448 96616 24512
rect 96680 24448 96686 24512
rect 98200 24488 99000 24518
rect 96370 24447 96686 24448
rect 8293 24034 8359 24037
rect 8293 24032 8402 24034
rect 8293 23976 8298 24032
rect 8354 23976 8402 24032
rect 8293 23971 8402 23976
rect 4870 23968 5186 23969
rect 0 23898 800 23928
rect 4870 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5186 23968
rect 4870 23903 5186 23904
rect 1301 23898 1367 23901
rect 0 23896 1367 23898
rect 0 23840 1306 23896
rect 1362 23840 1367 23896
rect 0 23838 1367 23840
rect 0 23808 800 23838
rect 1301 23835 1367 23838
rect 8342 23596 8402 23971
rect 97030 23968 97346 23969
rect 97030 23904 97036 23968
rect 97100 23904 97116 23968
rect 97180 23904 97196 23968
rect 97260 23904 97276 23968
rect 97340 23904 97346 23968
rect 97030 23903 97346 23904
rect 97441 23898 97507 23901
rect 98200 23898 99000 23928
rect 97441 23896 99000 23898
rect 97441 23840 97446 23896
rect 97502 23840 99000 23896
rect 97441 23838 99000 23840
rect 97441 23835 97507 23838
rect 98200 23808 99000 23838
rect 96613 23762 96679 23765
rect 91878 23760 96679 23762
rect 91878 23704 96618 23760
rect 96674 23704 96679 23760
rect 91878 23702 96679 23704
rect 91878 23596 91938 23702
rect 96613 23699 96679 23702
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 96370 23424 96686 23425
rect 96370 23360 96376 23424
rect 96440 23360 96456 23424
rect 96520 23360 96536 23424
rect 96600 23360 96616 23424
rect 96680 23360 96686 23424
rect 96370 23359 96686 23360
rect 4870 22880 5186 22881
rect 4870 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5186 22880
rect 4870 22815 5186 22816
rect 97030 22880 97346 22881
rect 97030 22816 97036 22880
rect 97100 22816 97116 22880
rect 97180 22816 97196 22880
rect 97260 22816 97276 22880
rect 97340 22816 97346 22880
rect 97030 22815 97346 22816
rect 8293 22674 8359 22677
rect 97257 22674 97323 22677
rect 8293 22672 8402 22674
rect 8293 22616 8298 22672
rect 8354 22616 8402 22672
rect 8293 22611 8402 22616
rect 0 22538 800 22568
rect 1117 22538 1183 22541
rect 0 22536 1183 22538
rect 0 22480 1122 22536
rect 1178 22480 1183 22536
rect 8342 22508 8402 22611
rect 91878 22672 97323 22674
rect 91878 22616 97262 22672
rect 97318 22616 97323 22672
rect 91878 22614 97323 22616
rect 91878 22508 91938 22614
rect 97257 22611 97323 22614
rect 97441 22538 97507 22541
rect 98200 22538 99000 22568
rect 97441 22536 99000 22538
rect 0 22478 1183 22480
rect 0 22448 800 22478
rect 1117 22475 1183 22478
rect 97441 22480 97446 22536
rect 97502 22480 99000 22536
rect 97441 22478 99000 22480
rect 97441 22475 97507 22478
rect 98200 22448 99000 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 96370 22336 96686 22337
rect 96370 22272 96376 22336
rect 96440 22272 96456 22336
rect 96520 22272 96536 22336
rect 96600 22272 96616 22336
rect 96680 22272 96686 22336
rect 96370 22271 96686 22272
rect 4870 21792 5186 21793
rect 4870 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5186 21792
rect 4870 21727 5186 21728
rect 97030 21792 97346 21793
rect 97030 21728 97036 21792
rect 97100 21728 97116 21792
rect 97180 21728 97196 21792
rect 97260 21728 97276 21792
rect 97340 21728 97346 21792
rect 97030 21727 97346 21728
rect 8293 21586 8359 21589
rect 97257 21586 97323 21589
rect 8293 21584 8402 21586
rect 8293 21528 8298 21584
rect 8354 21528 8402 21584
rect 8293 21523 8402 21528
rect 8342 21420 8402 21523
rect 91878 21584 97323 21586
rect 91878 21528 97262 21584
rect 97318 21528 97323 21584
rect 91878 21526 97323 21528
rect 91878 21420 91938 21526
rect 97257 21523 97323 21526
rect 4210 21248 4526 21249
rect 0 21178 800 21208
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 96370 21248 96686 21249
rect 96370 21184 96376 21248
rect 96440 21184 96456 21248
rect 96520 21184 96536 21248
rect 96600 21184 96616 21248
rect 96680 21184 96686 21248
rect 96370 21183 96686 21184
rect 1301 21178 1367 21181
rect 0 21176 1367 21178
rect 0 21120 1306 21176
rect 1362 21120 1367 21176
rect 0 21118 1367 21120
rect 0 21088 800 21118
rect 1301 21115 1367 21118
rect 97441 21178 97507 21181
rect 98200 21178 99000 21208
rect 97441 21176 99000 21178
rect 97441 21120 97446 21176
rect 97502 21120 99000 21176
rect 97441 21118 99000 21120
rect 97441 21115 97507 21118
rect 98200 21088 99000 21118
rect 4870 20704 5186 20705
rect 4870 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5186 20704
rect 4870 20639 5186 20640
rect 97030 20704 97346 20705
rect 97030 20640 97036 20704
rect 97100 20640 97116 20704
rect 97180 20640 97196 20704
rect 97260 20640 97276 20704
rect 97340 20640 97346 20704
rect 97030 20639 97346 20640
rect 0 20498 800 20528
rect 1301 20498 1367 20501
rect 96613 20498 96679 20501
rect 0 20496 1367 20498
rect 0 20440 1306 20496
rect 1362 20440 1367 20496
rect 0 20438 1367 20440
rect 0 20408 800 20438
rect 1301 20435 1367 20438
rect 91878 20496 96679 20498
rect 91878 20440 96618 20496
rect 96674 20440 96679 20496
rect 91878 20438 96679 20440
rect 1853 20362 1919 20365
rect 1853 20360 8188 20362
rect 1853 20304 1858 20360
rect 1914 20304 8188 20360
rect 91878 20332 91938 20438
rect 96613 20435 96679 20438
rect 97441 20498 97507 20501
rect 98200 20498 99000 20528
rect 97441 20496 99000 20498
rect 97441 20440 97446 20496
rect 97502 20440 99000 20496
rect 97441 20438 99000 20440
rect 97441 20435 97507 20438
rect 98200 20408 99000 20438
rect 1853 20302 8188 20304
rect 1853 20299 1919 20302
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 96370 20160 96686 20161
rect 96370 20096 96376 20160
rect 96440 20096 96456 20160
rect 96520 20096 96536 20160
rect 96600 20096 96616 20160
rect 96680 20096 96686 20160
rect 96370 20095 96686 20096
rect 4870 19616 5186 19617
rect 4870 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5186 19616
rect 4870 19551 5186 19552
rect 97030 19616 97346 19617
rect 97030 19552 97036 19616
rect 97100 19552 97116 19616
rect 97180 19552 97196 19616
rect 97260 19552 97276 19616
rect 97340 19552 97346 19616
rect 97030 19551 97346 19552
rect 97257 19274 97323 19277
rect 91908 19272 97323 19274
rect 0 19138 800 19168
rect 1485 19138 1551 19141
rect 0 19136 1551 19138
rect 0 19080 1490 19136
rect 1546 19080 1551 19136
rect 0 19078 1551 19080
rect 0 19048 800 19078
rect 1485 19075 1551 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 8342 19005 8402 19244
rect 91908 19216 97262 19272
rect 97318 19216 97323 19272
rect 91908 19214 97323 19216
rect 97257 19211 97323 19214
rect 97441 19138 97507 19141
rect 98200 19138 99000 19168
rect 97441 19136 99000 19138
rect 97441 19080 97446 19136
rect 97502 19080 99000 19136
rect 97441 19078 99000 19080
rect 97441 19075 97507 19078
rect 96370 19072 96686 19073
rect 96370 19008 96376 19072
rect 96440 19008 96456 19072
rect 96520 19008 96536 19072
rect 96600 19008 96616 19072
rect 96680 19008 96686 19072
rect 98200 19048 99000 19078
rect 96370 19007 96686 19008
rect 8293 19000 8402 19005
rect 8293 18944 8298 19000
rect 8354 18944 8402 19000
rect 8293 18942 8402 18944
rect 8293 18939 8359 18942
rect 8293 18594 8359 18597
rect 8293 18592 8402 18594
rect 8293 18536 8298 18592
rect 8354 18536 8402 18592
rect 8293 18531 8402 18536
rect 4870 18528 5186 18529
rect 0 18458 800 18488
rect 4870 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5186 18528
rect 4870 18463 5186 18464
rect 1301 18458 1367 18461
rect 0 18456 1367 18458
rect 0 18400 1306 18456
rect 1362 18400 1367 18456
rect 0 18398 1367 18400
rect 0 18368 800 18398
rect 1301 18395 1367 18398
rect 8342 18156 8402 18531
rect 97030 18528 97346 18529
rect 97030 18464 97036 18528
rect 97100 18464 97116 18528
rect 97180 18464 97196 18528
rect 97260 18464 97276 18528
rect 97340 18464 97346 18528
rect 97030 18463 97346 18464
rect 97441 18458 97507 18461
rect 98200 18458 99000 18488
rect 97441 18456 99000 18458
rect 97441 18400 97446 18456
rect 97502 18400 99000 18456
rect 97441 18398 99000 18400
rect 97441 18395 97507 18398
rect 98200 18368 99000 18398
rect 96613 18322 96679 18325
rect 91878 18320 96679 18322
rect 91878 18264 96618 18320
rect 96674 18264 96679 18320
rect 91878 18262 96679 18264
rect 91878 18156 91938 18262
rect 96613 18259 96679 18262
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 96370 17984 96686 17985
rect 96370 17920 96376 17984
rect 96440 17920 96456 17984
rect 96520 17920 96536 17984
rect 96600 17920 96616 17984
rect 96680 17920 96686 17984
rect 96370 17919 96686 17920
rect 4870 17440 5186 17441
rect 4870 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5186 17440
rect 4870 17375 5186 17376
rect 97030 17440 97346 17441
rect 97030 17376 97036 17440
rect 97100 17376 97116 17440
rect 97180 17376 97196 17440
rect 97260 17376 97276 17440
rect 97340 17376 97346 17440
rect 97030 17375 97346 17376
rect 8293 17234 8359 17237
rect 97257 17234 97323 17237
rect 8293 17232 8402 17234
rect 8293 17176 8298 17232
rect 8354 17176 8402 17232
rect 8293 17171 8402 17176
rect 0 17098 800 17128
rect 1117 17098 1183 17101
rect 0 17096 1183 17098
rect 0 17040 1122 17096
rect 1178 17040 1183 17096
rect 8342 17068 8402 17171
rect 91878 17232 97323 17234
rect 91878 17176 97262 17232
rect 97318 17176 97323 17232
rect 91878 17174 97323 17176
rect 91878 17068 91938 17174
rect 97257 17171 97323 17174
rect 97441 17098 97507 17101
rect 98200 17098 99000 17128
rect 97441 17096 99000 17098
rect 0 17038 1183 17040
rect 0 17008 800 17038
rect 1117 17035 1183 17038
rect 97441 17040 97446 17096
rect 97502 17040 99000 17096
rect 97441 17038 99000 17040
rect 97441 17035 97507 17038
rect 98200 17008 99000 17038
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 96370 16896 96686 16897
rect 96370 16832 96376 16896
rect 96440 16832 96456 16896
rect 96520 16832 96536 16896
rect 96600 16832 96616 16896
rect 96680 16832 96686 16896
rect 96370 16831 96686 16832
rect 4870 16352 5186 16353
rect 4870 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5186 16352
rect 4870 16287 5186 16288
rect 97030 16352 97346 16353
rect 97030 16288 97036 16352
rect 97100 16288 97116 16352
rect 97180 16288 97196 16352
rect 97260 16288 97276 16352
rect 97340 16288 97346 16352
rect 97030 16287 97346 16288
rect 8293 16146 8359 16149
rect 97257 16146 97323 16149
rect 8293 16144 8402 16146
rect 8293 16088 8298 16144
rect 8354 16088 8402 16144
rect 8293 16083 8402 16088
rect 8342 15980 8402 16083
rect 91878 16144 97323 16146
rect 91878 16088 97262 16144
rect 97318 16088 97323 16144
rect 91878 16086 97323 16088
rect 91878 15980 91938 16086
rect 97257 16083 97323 16086
rect 4210 15808 4526 15809
rect 0 15738 800 15768
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 96370 15808 96686 15809
rect 96370 15744 96376 15808
rect 96440 15744 96456 15808
rect 96520 15744 96536 15808
rect 96600 15744 96616 15808
rect 96680 15744 96686 15808
rect 96370 15743 96686 15744
rect 1209 15738 1275 15741
rect 0 15736 1275 15738
rect 0 15680 1214 15736
rect 1270 15680 1275 15736
rect 0 15678 1275 15680
rect 0 15648 800 15678
rect 1209 15675 1275 15678
rect 97441 15738 97507 15741
rect 98200 15738 99000 15768
rect 97441 15736 99000 15738
rect 97441 15680 97446 15736
rect 97502 15680 99000 15736
rect 97441 15678 99000 15680
rect 97441 15675 97507 15678
rect 98200 15648 99000 15678
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 97030 15264 97346 15265
rect 97030 15200 97036 15264
rect 97100 15200 97116 15264
rect 97180 15200 97196 15264
rect 97260 15200 97276 15264
rect 97340 15200 97346 15264
rect 97030 15199 97346 15200
rect 0 15058 800 15088
rect 1301 15058 1367 15061
rect 96613 15058 96679 15061
rect 0 15056 1367 15058
rect 0 15000 1306 15056
rect 1362 15000 1367 15056
rect 0 14998 1367 15000
rect 0 14968 800 14998
rect 1301 14995 1367 14998
rect 91878 15056 96679 15058
rect 91878 15000 96618 15056
rect 96674 15000 96679 15056
rect 91878 14998 96679 15000
rect 1853 14922 1919 14925
rect 1853 14920 8188 14922
rect 1853 14864 1858 14920
rect 1914 14864 8188 14920
rect 91878 14892 91938 14998
rect 96613 14995 96679 14998
rect 97441 15058 97507 15061
rect 98200 15058 99000 15088
rect 97441 15056 99000 15058
rect 97441 15000 97446 15056
rect 97502 15000 99000 15056
rect 97441 14998 99000 15000
rect 97441 14995 97507 14998
rect 98200 14968 99000 14998
rect 1853 14862 8188 14864
rect 1853 14859 1919 14862
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 96370 14720 96686 14721
rect 96370 14656 96376 14720
rect 96440 14656 96456 14720
rect 96520 14656 96536 14720
rect 96600 14656 96616 14720
rect 96680 14656 96686 14720
rect 96370 14655 96686 14656
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 97030 14176 97346 14177
rect 97030 14112 97036 14176
rect 97100 14112 97116 14176
rect 97180 14112 97196 14176
rect 97260 14112 97276 14176
rect 97340 14112 97346 14176
rect 97030 14111 97346 14112
rect 8293 13970 8359 13973
rect 97257 13970 97323 13973
rect 8293 13968 8402 13970
rect 8293 13912 8298 13968
rect 8354 13912 8402 13968
rect 8293 13907 8402 13912
rect 8342 13804 8402 13907
rect 91878 13968 97323 13970
rect 91878 13912 97262 13968
rect 97318 13912 97323 13968
rect 91878 13910 97323 13912
rect 91878 13804 91938 13910
rect 97257 13907 97323 13910
rect 0 13698 800 13728
rect 1301 13698 1367 13701
rect 0 13696 1367 13698
rect 0 13640 1306 13696
rect 1362 13640 1367 13696
rect 0 13638 1367 13640
rect 0 13608 800 13638
rect 1301 13635 1367 13638
rect 97441 13698 97507 13701
rect 98200 13698 99000 13728
rect 97441 13696 99000 13698
rect 97441 13640 97446 13696
rect 97502 13640 99000 13696
rect 97441 13638 99000 13640
rect 97441 13635 97507 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 96370 13632 96686 13633
rect 96370 13568 96376 13632
rect 96440 13568 96456 13632
rect 96520 13568 96536 13632
rect 96600 13568 96616 13632
rect 96680 13568 96686 13632
rect 98200 13608 99000 13638
rect 96370 13567 96686 13568
rect 8293 13290 8359 13293
rect 8293 13288 8402 13290
rect 8293 13232 8298 13288
rect 8354 13232 8402 13288
rect 8293 13227 8402 13232
rect 4870 13088 5186 13089
rect 0 13018 800 13048
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 1301 13018 1367 13021
rect 0 13016 1367 13018
rect 0 12960 1306 13016
rect 1362 12960 1367 13016
rect 0 12958 1367 12960
rect 0 12928 800 12958
rect 1301 12955 1367 12958
rect 8342 12716 8402 13227
rect 97030 13088 97346 13089
rect 97030 13024 97036 13088
rect 97100 13024 97116 13088
rect 97180 13024 97196 13088
rect 97260 13024 97276 13088
rect 97340 13024 97346 13088
rect 97030 13023 97346 13024
rect 97441 13018 97507 13021
rect 98200 13018 99000 13048
rect 97441 13016 99000 13018
rect 97441 12960 97446 13016
rect 97502 12960 99000 13016
rect 97441 12958 99000 12960
rect 97441 12955 97507 12958
rect 98200 12928 99000 12958
rect 96613 12882 96679 12885
rect 91878 12880 96679 12882
rect 91878 12824 96618 12880
rect 96674 12824 96679 12880
rect 91878 12822 96679 12824
rect 91878 12716 91938 12822
rect 96613 12819 96679 12822
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 96370 12544 96686 12545
rect 96370 12480 96376 12544
rect 96440 12480 96456 12544
rect 96520 12480 96536 12544
rect 96600 12480 96616 12544
rect 96680 12480 96686 12544
rect 96370 12479 96686 12480
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 97030 12000 97346 12001
rect 97030 11936 97036 12000
rect 97100 11936 97116 12000
rect 97180 11936 97196 12000
rect 97260 11936 97276 12000
rect 97340 11936 97346 12000
rect 97030 11935 97346 11936
rect 8293 11794 8359 11797
rect 97257 11794 97323 11797
rect 8293 11792 8402 11794
rect 8293 11736 8298 11792
rect 8354 11736 8402 11792
rect 8293 11731 8402 11736
rect 0 11658 800 11688
rect 1117 11658 1183 11661
rect 0 11656 1183 11658
rect 0 11600 1122 11656
rect 1178 11600 1183 11656
rect 8342 11628 8402 11731
rect 91878 11792 97323 11794
rect 91878 11736 97262 11792
rect 97318 11736 97323 11792
rect 91878 11734 97323 11736
rect 91878 11628 91938 11734
rect 97257 11731 97323 11734
rect 97441 11658 97507 11661
rect 98200 11658 99000 11688
rect 97441 11656 99000 11658
rect 0 11598 1183 11600
rect 0 11568 800 11598
rect 1117 11595 1183 11598
rect 97441 11600 97446 11656
rect 97502 11600 99000 11656
rect 97441 11598 99000 11600
rect 97441 11595 97507 11598
rect 98200 11568 99000 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 96370 11456 96686 11457
rect 96370 11392 96376 11456
rect 96440 11392 96456 11456
rect 96520 11392 96536 11456
rect 96600 11392 96616 11456
rect 96680 11392 96686 11456
rect 96370 11391 96686 11392
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 4870 10847 5186 10848
rect 97030 10912 97346 10913
rect 97030 10848 97036 10912
rect 97100 10848 97116 10912
rect 97180 10848 97196 10912
rect 97260 10848 97276 10912
rect 97340 10848 97346 10912
rect 97030 10847 97346 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 96370 10368 96686 10369
rect 96370 10304 96376 10368
rect 96440 10304 96456 10368
rect 96520 10304 96536 10368
rect 96600 10304 96616 10368
rect 96680 10304 96686 10368
rect 96370 10303 96686 10304
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 97030 9824 97346 9825
rect 97030 9760 97036 9824
rect 97100 9760 97116 9824
rect 97180 9760 97196 9824
rect 97260 9760 97276 9824
rect 97340 9760 97346 9824
rect 97030 9759 97346 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 96370 9280 96686 9281
rect 96370 9216 96376 9280
rect 96440 9216 96456 9280
rect 96520 9216 96536 9280
rect 96600 9216 96616 9280
rect 96680 9216 96686 9280
rect 96370 9215 96686 9216
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 97030 8736 97346 8737
rect 97030 8672 97036 8736
rect 97100 8672 97116 8736
rect 97180 8672 97196 8736
rect 97260 8672 97276 8736
rect 97340 8672 97346 8736
rect 97030 8671 97346 8672
rect 50843 8668 50909 8669
rect 50838 8666 50844 8668
rect 50756 8606 50844 8666
rect 50838 8604 50844 8606
rect 50908 8604 50914 8668
rect 50843 8603 50909 8604
rect 97533 8258 97599 8261
rect 98200 8258 99000 8288
rect 97533 8256 99000 8258
rect 97533 8200 97538 8256
rect 97594 8200 99000 8256
rect 97533 8198 99000 8200
rect 97533 8195 97599 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 96370 8192 96686 8193
rect 96370 8128 96376 8192
rect 96440 8128 96456 8192
rect 96520 8128 96536 8192
rect 96600 8128 96616 8192
rect 96680 8128 96686 8192
rect 98200 8168 99000 8198
rect 96370 8127 96686 8128
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 97030 7648 97346 7649
rect 97030 7584 97036 7648
rect 97100 7584 97116 7648
rect 97180 7584 97196 7648
rect 97260 7584 97276 7648
rect 97340 7584 97346 7648
rect 97030 7583 97346 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 96370 7104 96686 7105
rect 96370 7040 96376 7104
rect 96440 7040 96456 7104
rect 96520 7040 96536 7104
rect 96600 7040 96616 7104
rect 96680 7040 96686 7104
rect 96370 7039 96686 7040
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 97030 6560 97346 6561
rect 97030 6496 97036 6560
rect 97100 6496 97116 6560
rect 97180 6496 97196 6560
rect 97260 6496 97276 6560
rect 97340 6496 97346 6560
rect 97030 6495 97346 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 65650 6016 65966 6017
rect 65650 5952 65656 6016
rect 65720 5952 65736 6016
rect 65800 5952 65816 6016
rect 65880 5952 65896 6016
rect 65960 5952 65966 6016
rect 65650 5951 65966 5952
rect 96370 6016 96686 6017
rect 96370 5952 96376 6016
rect 96440 5952 96456 6016
rect 96520 5952 96536 6016
rect 96600 5952 96616 6016
rect 96680 5952 96686 6016
rect 96370 5951 96686 5952
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 4870 5407 5186 5408
rect 35590 5472 35906 5473
rect 35590 5408 35596 5472
rect 35660 5408 35676 5472
rect 35740 5408 35756 5472
rect 35820 5408 35836 5472
rect 35900 5408 35906 5472
rect 35590 5407 35906 5408
rect 66310 5472 66626 5473
rect 66310 5408 66316 5472
rect 66380 5408 66396 5472
rect 66460 5408 66476 5472
rect 66540 5408 66556 5472
rect 66620 5408 66626 5472
rect 66310 5407 66626 5408
rect 97030 5472 97346 5473
rect 97030 5408 97036 5472
rect 97100 5408 97116 5472
rect 97180 5408 97196 5472
rect 97260 5408 97276 5472
rect 97340 5408 97346 5472
rect 97030 5407 97346 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 65650 4928 65966 4929
rect 65650 4864 65656 4928
rect 65720 4864 65736 4928
rect 65800 4864 65816 4928
rect 65880 4864 65896 4928
rect 65960 4864 65966 4928
rect 65650 4863 65966 4864
rect 96370 4928 96686 4929
rect 96370 4864 96376 4928
rect 96440 4864 96456 4928
rect 96520 4864 96536 4928
rect 96600 4864 96616 4928
rect 96680 4864 96686 4928
rect 96370 4863 96686 4864
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 35590 4384 35906 4385
rect 35590 4320 35596 4384
rect 35660 4320 35676 4384
rect 35740 4320 35756 4384
rect 35820 4320 35836 4384
rect 35900 4320 35906 4384
rect 35590 4319 35906 4320
rect 66310 4384 66626 4385
rect 66310 4320 66316 4384
rect 66380 4320 66396 4384
rect 66460 4320 66476 4384
rect 66540 4320 66556 4384
rect 66620 4320 66626 4384
rect 66310 4319 66626 4320
rect 97030 4384 97346 4385
rect 97030 4320 97036 4384
rect 97100 4320 97116 4384
rect 97180 4320 97196 4384
rect 97260 4320 97276 4384
rect 97340 4320 97346 4384
rect 97030 4319 97346 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 65650 3840 65966 3841
rect 65650 3776 65656 3840
rect 65720 3776 65736 3840
rect 65800 3776 65816 3840
rect 65880 3776 65896 3840
rect 65960 3776 65966 3840
rect 65650 3775 65966 3776
rect 96370 3840 96686 3841
rect 96370 3776 96376 3840
rect 96440 3776 96456 3840
rect 96520 3776 96536 3840
rect 96600 3776 96616 3840
rect 96680 3776 96686 3840
rect 96370 3775 96686 3776
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 35590 3296 35906 3297
rect 35590 3232 35596 3296
rect 35660 3232 35676 3296
rect 35740 3232 35756 3296
rect 35820 3232 35836 3296
rect 35900 3232 35906 3296
rect 35590 3231 35906 3232
rect 66310 3296 66626 3297
rect 66310 3232 66316 3296
rect 66380 3232 66396 3296
rect 66460 3232 66476 3296
rect 66540 3232 66556 3296
rect 66620 3232 66626 3296
rect 66310 3231 66626 3232
rect 97030 3296 97346 3297
rect 97030 3232 97036 3296
rect 97100 3232 97116 3296
rect 97180 3232 97196 3296
rect 97260 3232 97276 3296
rect 97340 3232 97346 3296
rect 97030 3231 97346 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 65650 2752 65966 2753
rect 65650 2688 65656 2752
rect 65720 2688 65736 2752
rect 65800 2688 65816 2752
rect 65880 2688 65896 2752
rect 65960 2688 65966 2752
rect 65650 2687 65966 2688
rect 96370 2752 96686 2753
rect 96370 2688 96376 2752
rect 96440 2688 96456 2752
rect 96520 2688 96536 2752
rect 96600 2688 96616 2752
rect 96680 2688 96686 2752
rect 96370 2687 96686 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
rect 35590 2208 35906 2209
rect 35590 2144 35596 2208
rect 35660 2144 35676 2208
rect 35740 2144 35756 2208
rect 35820 2144 35836 2208
rect 35900 2144 35906 2208
rect 35590 2143 35906 2144
rect 66310 2208 66626 2209
rect 66310 2144 66316 2208
rect 66380 2144 66396 2208
rect 66460 2144 66476 2208
rect 66540 2144 66556 2208
rect 66620 2144 66626 2208
rect 66310 2143 66626 2144
rect 97030 2208 97346 2209
rect 97030 2144 97036 2208
rect 97100 2144 97116 2208
rect 97180 2144 97196 2208
rect 97260 2144 97276 2208
rect 97340 2144 97346 2208
rect 97030 2143 97346 2144
<< via3 >>
rect 4876 95772 4940 95776
rect 4876 95716 4880 95772
rect 4880 95716 4936 95772
rect 4936 95716 4940 95772
rect 4876 95712 4940 95716
rect 4956 95772 5020 95776
rect 4956 95716 4960 95772
rect 4960 95716 5016 95772
rect 5016 95716 5020 95772
rect 4956 95712 5020 95716
rect 5036 95772 5100 95776
rect 5036 95716 5040 95772
rect 5040 95716 5096 95772
rect 5096 95716 5100 95772
rect 5036 95712 5100 95716
rect 5116 95772 5180 95776
rect 5116 95716 5120 95772
rect 5120 95716 5176 95772
rect 5176 95716 5180 95772
rect 5116 95712 5180 95716
rect 35596 95772 35660 95776
rect 35596 95716 35600 95772
rect 35600 95716 35656 95772
rect 35656 95716 35660 95772
rect 35596 95712 35660 95716
rect 35676 95772 35740 95776
rect 35676 95716 35680 95772
rect 35680 95716 35736 95772
rect 35736 95716 35740 95772
rect 35676 95712 35740 95716
rect 35756 95772 35820 95776
rect 35756 95716 35760 95772
rect 35760 95716 35816 95772
rect 35816 95716 35820 95772
rect 35756 95712 35820 95716
rect 35836 95772 35900 95776
rect 35836 95716 35840 95772
rect 35840 95716 35896 95772
rect 35896 95716 35900 95772
rect 35836 95712 35900 95716
rect 66316 95772 66380 95776
rect 66316 95716 66320 95772
rect 66320 95716 66376 95772
rect 66376 95716 66380 95772
rect 66316 95712 66380 95716
rect 66396 95772 66460 95776
rect 66396 95716 66400 95772
rect 66400 95716 66456 95772
rect 66456 95716 66460 95772
rect 66396 95712 66460 95716
rect 66476 95772 66540 95776
rect 66476 95716 66480 95772
rect 66480 95716 66536 95772
rect 66536 95716 66540 95772
rect 66476 95712 66540 95716
rect 66556 95772 66620 95776
rect 66556 95716 66560 95772
rect 66560 95716 66616 95772
rect 66616 95716 66620 95772
rect 66556 95712 66620 95716
rect 97036 95772 97100 95776
rect 97036 95716 97040 95772
rect 97040 95716 97096 95772
rect 97096 95716 97100 95772
rect 97036 95712 97100 95716
rect 97116 95772 97180 95776
rect 97116 95716 97120 95772
rect 97120 95716 97176 95772
rect 97176 95716 97180 95772
rect 97116 95712 97180 95716
rect 97196 95772 97260 95776
rect 97196 95716 97200 95772
rect 97200 95716 97256 95772
rect 97256 95716 97260 95772
rect 97196 95712 97260 95716
rect 97276 95772 97340 95776
rect 97276 95716 97280 95772
rect 97280 95716 97336 95772
rect 97336 95716 97340 95772
rect 97276 95712 97340 95716
rect 4216 95228 4280 95232
rect 4216 95172 4220 95228
rect 4220 95172 4276 95228
rect 4276 95172 4280 95228
rect 4216 95168 4280 95172
rect 4296 95228 4360 95232
rect 4296 95172 4300 95228
rect 4300 95172 4356 95228
rect 4356 95172 4360 95228
rect 4296 95168 4360 95172
rect 4376 95228 4440 95232
rect 4376 95172 4380 95228
rect 4380 95172 4436 95228
rect 4436 95172 4440 95228
rect 4376 95168 4440 95172
rect 4456 95228 4520 95232
rect 4456 95172 4460 95228
rect 4460 95172 4516 95228
rect 4516 95172 4520 95228
rect 4456 95168 4520 95172
rect 34936 95228 35000 95232
rect 34936 95172 34940 95228
rect 34940 95172 34996 95228
rect 34996 95172 35000 95228
rect 34936 95168 35000 95172
rect 35016 95228 35080 95232
rect 35016 95172 35020 95228
rect 35020 95172 35076 95228
rect 35076 95172 35080 95228
rect 35016 95168 35080 95172
rect 35096 95228 35160 95232
rect 35096 95172 35100 95228
rect 35100 95172 35156 95228
rect 35156 95172 35160 95228
rect 35096 95168 35160 95172
rect 35176 95228 35240 95232
rect 35176 95172 35180 95228
rect 35180 95172 35236 95228
rect 35236 95172 35240 95228
rect 35176 95168 35240 95172
rect 65656 95228 65720 95232
rect 65656 95172 65660 95228
rect 65660 95172 65716 95228
rect 65716 95172 65720 95228
rect 65656 95168 65720 95172
rect 65736 95228 65800 95232
rect 65736 95172 65740 95228
rect 65740 95172 65796 95228
rect 65796 95172 65800 95228
rect 65736 95168 65800 95172
rect 65816 95228 65880 95232
rect 65816 95172 65820 95228
rect 65820 95172 65876 95228
rect 65876 95172 65880 95228
rect 65816 95168 65880 95172
rect 65896 95228 65960 95232
rect 65896 95172 65900 95228
rect 65900 95172 65956 95228
rect 65956 95172 65960 95228
rect 65896 95168 65960 95172
rect 96376 95228 96440 95232
rect 96376 95172 96380 95228
rect 96380 95172 96436 95228
rect 96436 95172 96440 95228
rect 96376 95168 96440 95172
rect 96456 95228 96520 95232
rect 96456 95172 96460 95228
rect 96460 95172 96516 95228
rect 96516 95172 96520 95228
rect 96456 95168 96520 95172
rect 96536 95228 96600 95232
rect 96536 95172 96540 95228
rect 96540 95172 96596 95228
rect 96596 95172 96600 95228
rect 96536 95168 96600 95172
rect 96616 95228 96680 95232
rect 96616 95172 96620 95228
rect 96620 95172 96676 95228
rect 96676 95172 96680 95228
rect 96616 95168 96680 95172
rect 4876 94684 4940 94688
rect 4876 94628 4880 94684
rect 4880 94628 4936 94684
rect 4936 94628 4940 94684
rect 4876 94624 4940 94628
rect 4956 94684 5020 94688
rect 4956 94628 4960 94684
rect 4960 94628 5016 94684
rect 5016 94628 5020 94684
rect 4956 94624 5020 94628
rect 5036 94684 5100 94688
rect 5036 94628 5040 94684
rect 5040 94628 5096 94684
rect 5096 94628 5100 94684
rect 5036 94624 5100 94628
rect 5116 94684 5180 94688
rect 5116 94628 5120 94684
rect 5120 94628 5176 94684
rect 5176 94628 5180 94684
rect 5116 94624 5180 94628
rect 35596 94684 35660 94688
rect 35596 94628 35600 94684
rect 35600 94628 35656 94684
rect 35656 94628 35660 94684
rect 35596 94624 35660 94628
rect 35676 94684 35740 94688
rect 35676 94628 35680 94684
rect 35680 94628 35736 94684
rect 35736 94628 35740 94684
rect 35676 94624 35740 94628
rect 35756 94684 35820 94688
rect 35756 94628 35760 94684
rect 35760 94628 35816 94684
rect 35816 94628 35820 94684
rect 35756 94624 35820 94628
rect 35836 94684 35900 94688
rect 35836 94628 35840 94684
rect 35840 94628 35896 94684
rect 35896 94628 35900 94684
rect 35836 94624 35900 94628
rect 66316 94684 66380 94688
rect 66316 94628 66320 94684
rect 66320 94628 66376 94684
rect 66376 94628 66380 94684
rect 66316 94624 66380 94628
rect 66396 94684 66460 94688
rect 66396 94628 66400 94684
rect 66400 94628 66456 94684
rect 66456 94628 66460 94684
rect 66396 94624 66460 94628
rect 66476 94684 66540 94688
rect 66476 94628 66480 94684
rect 66480 94628 66536 94684
rect 66536 94628 66540 94684
rect 66476 94624 66540 94628
rect 66556 94684 66620 94688
rect 66556 94628 66560 94684
rect 66560 94628 66616 94684
rect 66616 94628 66620 94684
rect 66556 94624 66620 94628
rect 97036 94684 97100 94688
rect 97036 94628 97040 94684
rect 97040 94628 97096 94684
rect 97096 94628 97100 94684
rect 97036 94624 97100 94628
rect 97116 94684 97180 94688
rect 97116 94628 97120 94684
rect 97120 94628 97176 94684
rect 97176 94628 97180 94684
rect 97116 94624 97180 94628
rect 97196 94684 97260 94688
rect 97196 94628 97200 94684
rect 97200 94628 97256 94684
rect 97256 94628 97260 94684
rect 97196 94624 97260 94628
rect 97276 94684 97340 94688
rect 97276 94628 97280 94684
rect 97280 94628 97336 94684
rect 97336 94628 97340 94684
rect 97276 94624 97340 94628
rect 4216 94140 4280 94144
rect 4216 94084 4220 94140
rect 4220 94084 4276 94140
rect 4276 94084 4280 94140
rect 4216 94080 4280 94084
rect 4296 94140 4360 94144
rect 4296 94084 4300 94140
rect 4300 94084 4356 94140
rect 4356 94084 4360 94140
rect 4296 94080 4360 94084
rect 4376 94140 4440 94144
rect 4376 94084 4380 94140
rect 4380 94084 4436 94140
rect 4436 94084 4440 94140
rect 4376 94080 4440 94084
rect 4456 94140 4520 94144
rect 4456 94084 4460 94140
rect 4460 94084 4516 94140
rect 4516 94084 4520 94140
rect 4456 94080 4520 94084
rect 34936 94140 35000 94144
rect 34936 94084 34940 94140
rect 34940 94084 34996 94140
rect 34996 94084 35000 94140
rect 34936 94080 35000 94084
rect 35016 94140 35080 94144
rect 35016 94084 35020 94140
rect 35020 94084 35076 94140
rect 35076 94084 35080 94140
rect 35016 94080 35080 94084
rect 35096 94140 35160 94144
rect 35096 94084 35100 94140
rect 35100 94084 35156 94140
rect 35156 94084 35160 94140
rect 35096 94080 35160 94084
rect 35176 94140 35240 94144
rect 35176 94084 35180 94140
rect 35180 94084 35236 94140
rect 35236 94084 35240 94140
rect 35176 94080 35240 94084
rect 65656 94140 65720 94144
rect 65656 94084 65660 94140
rect 65660 94084 65716 94140
rect 65716 94084 65720 94140
rect 65656 94080 65720 94084
rect 65736 94140 65800 94144
rect 65736 94084 65740 94140
rect 65740 94084 65796 94140
rect 65796 94084 65800 94140
rect 65736 94080 65800 94084
rect 65816 94140 65880 94144
rect 65816 94084 65820 94140
rect 65820 94084 65876 94140
rect 65876 94084 65880 94140
rect 65816 94080 65880 94084
rect 65896 94140 65960 94144
rect 65896 94084 65900 94140
rect 65900 94084 65956 94140
rect 65956 94084 65960 94140
rect 65896 94080 65960 94084
rect 96376 94140 96440 94144
rect 96376 94084 96380 94140
rect 96380 94084 96436 94140
rect 96436 94084 96440 94140
rect 96376 94080 96440 94084
rect 96456 94140 96520 94144
rect 96456 94084 96460 94140
rect 96460 94084 96516 94140
rect 96516 94084 96520 94140
rect 96456 94080 96520 94084
rect 96536 94140 96600 94144
rect 96536 94084 96540 94140
rect 96540 94084 96596 94140
rect 96596 94084 96600 94140
rect 96536 94080 96600 94084
rect 96616 94140 96680 94144
rect 96616 94084 96620 94140
rect 96620 94084 96676 94140
rect 96676 94084 96680 94140
rect 96616 94080 96680 94084
rect 4876 93596 4940 93600
rect 4876 93540 4880 93596
rect 4880 93540 4936 93596
rect 4936 93540 4940 93596
rect 4876 93536 4940 93540
rect 4956 93596 5020 93600
rect 4956 93540 4960 93596
rect 4960 93540 5016 93596
rect 5016 93540 5020 93596
rect 4956 93536 5020 93540
rect 5036 93596 5100 93600
rect 5036 93540 5040 93596
rect 5040 93540 5096 93596
rect 5096 93540 5100 93596
rect 5036 93536 5100 93540
rect 5116 93596 5180 93600
rect 5116 93540 5120 93596
rect 5120 93540 5176 93596
rect 5176 93540 5180 93596
rect 5116 93536 5180 93540
rect 35596 93596 35660 93600
rect 35596 93540 35600 93596
rect 35600 93540 35656 93596
rect 35656 93540 35660 93596
rect 35596 93536 35660 93540
rect 35676 93596 35740 93600
rect 35676 93540 35680 93596
rect 35680 93540 35736 93596
rect 35736 93540 35740 93596
rect 35676 93536 35740 93540
rect 35756 93596 35820 93600
rect 35756 93540 35760 93596
rect 35760 93540 35816 93596
rect 35816 93540 35820 93596
rect 35756 93536 35820 93540
rect 35836 93596 35900 93600
rect 35836 93540 35840 93596
rect 35840 93540 35896 93596
rect 35896 93540 35900 93596
rect 35836 93536 35900 93540
rect 66316 93596 66380 93600
rect 66316 93540 66320 93596
rect 66320 93540 66376 93596
rect 66376 93540 66380 93596
rect 66316 93536 66380 93540
rect 66396 93596 66460 93600
rect 66396 93540 66400 93596
rect 66400 93540 66456 93596
rect 66456 93540 66460 93596
rect 66396 93536 66460 93540
rect 66476 93596 66540 93600
rect 66476 93540 66480 93596
rect 66480 93540 66536 93596
rect 66536 93540 66540 93596
rect 66476 93536 66540 93540
rect 66556 93596 66620 93600
rect 66556 93540 66560 93596
rect 66560 93540 66616 93596
rect 66616 93540 66620 93596
rect 66556 93536 66620 93540
rect 97036 93596 97100 93600
rect 97036 93540 97040 93596
rect 97040 93540 97096 93596
rect 97096 93540 97100 93596
rect 97036 93536 97100 93540
rect 97116 93596 97180 93600
rect 97116 93540 97120 93596
rect 97120 93540 97176 93596
rect 97176 93540 97180 93596
rect 97116 93536 97180 93540
rect 97196 93596 97260 93600
rect 97196 93540 97200 93596
rect 97200 93540 97256 93596
rect 97256 93540 97260 93596
rect 97196 93536 97260 93540
rect 97276 93596 97340 93600
rect 97276 93540 97280 93596
rect 97280 93540 97336 93596
rect 97336 93540 97340 93596
rect 97276 93536 97340 93540
rect 4216 93052 4280 93056
rect 4216 92996 4220 93052
rect 4220 92996 4276 93052
rect 4276 92996 4280 93052
rect 4216 92992 4280 92996
rect 4296 93052 4360 93056
rect 4296 92996 4300 93052
rect 4300 92996 4356 93052
rect 4356 92996 4360 93052
rect 4296 92992 4360 92996
rect 4376 93052 4440 93056
rect 4376 92996 4380 93052
rect 4380 92996 4436 93052
rect 4436 92996 4440 93052
rect 4376 92992 4440 92996
rect 4456 93052 4520 93056
rect 4456 92996 4460 93052
rect 4460 92996 4516 93052
rect 4516 92996 4520 93052
rect 4456 92992 4520 92996
rect 34936 93052 35000 93056
rect 34936 92996 34940 93052
rect 34940 92996 34996 93052
rect 34996 92996 35000 93052
rect 34936 92992 35000 92996
rect 35016 93052 35080 93056
rect 35016 92996 35020 93052
rect 35020 92996 35076 93052
rect 35076 92996 35080 93052
rect 35016 92992 35080 92996
rect 35096 93052 35160 93056
rect 35096 92996 35100 93052
rect 35100 92996 35156 93052
rect 35156 92996 35160 93052
rect 35096 92992 35160 92996
rect 35176 93052 35240 93056
rect 35176 92996 35180 93052
rect 35180 92996 35236 93052
rect 35236 92996 35240 93052
rect 35176 92992 35240 92996
rect 65656 93052 65720 93056
rect 65656 92996 65660 93052
rect 65660 92996 65716 93052
rect 65716 92996 65720 93052
rect 65656 92992 65720 92996
rect 65736 93052 65800 93056
rect 65736 92996 65740 93052
rect 65740 92996 65796 93052
rect 65796 92996 65800 93052
rect 65736 92992 65800 92996
rect 65816 93052 65880 93056
rect 65816 92996 65820 93052
rect 65820 92996 65876 93052
rect 65876 92996 65880 93052
rect 65816 92992 65880 92996
rect 65896 93052 65960 93056
rect 65896 92996 65900 93052
rect 65900 92996 65956 93052
rect 65956 92996 65960 93052
rect 65896 92992 65960 92996
rect 96376 93052 96440 93056
rect 96376 92996 96380 93052
rect 96380 92996 96436 93052
rect 96436 92996 96440 93052
rect 96376 92992 96440 92996
rect 96456 93052 96520 93056
rect 96456 92996 96460 93052
rect 96460 92996 96516 93052
rect 96516 92996 96520 93052
rect 96456 92992 96520 92996
rect 96536 93052 96600 93056
rect 96536 92996 96540 93052
rect 96540 92996 96596 93052
rect 96596 92996 96600 93052
rect 96536 92992 96600 92996
rect 96616 93052 96680 93056
rect 96616 92996 96620 93052
rect 96620 92996 96676 93052
rect 96676 92996 96680 93052
rect 96616 92992 96680 92996
rect 4876 92508 4940 92512
rect 4876 92452 4880 92508
rect 4880 92452 4936 92508
rect 4936 92452 4940 92508
rect 4876 92448 4940 92452
rect 4956 92508 5020 92512
rect 4956 92452 4960 92508
rect 4960 92452 5016 92508
rect 5016 92452 5020 92508
rect 4956 92448 5020 92452
rect 5036 92508 5100 92512
rect 5036 92452 5040 92508
rect 5040 92452 5096 92508
rect 5096 92452 5100 92508
rect 5036 92448 5100 92452
rect 5116 92508 5180 92512
rect 5116 92452 5120 92508
rect 5120 92452 5176 92508
rect 5176 92452 5180 92508
rect 5116 92448 5180 92452
rect 97036 92508 97100 92512
rect 97036 92452 97040 92508
rect 97040 92452 97096 92508
rect 97096 92452 97100 92508
rect 97036 92448 97100 92452
rect 97116 92508 97180 92512
rect 97116 92452 97120 92508
rect 97120 92452 97176 92508
rect 97176 92452 97180 92508
rect 97116 92448 97180 92452
rect 97196 92508 97260 92512
rect 97196 92452 97200 92508
rect 97200 92452 97256 92508
rect 97256 92452 97260 92508
rect 97196 92448 97260 92452
rect 97276 92508 97340 92512
rect 97276 92452 97280 92508
rect 97280 92452 97336 92508
rect 97336 92452 97340 92508
rect 97276 92448 97340 92452
rect 4216 91964 4280 91968
rect 4216 91908 4220 91964
rect 4220 91908 4276 91964
rect 4276 91908 4280 91964
rect 4216 91904 4280 91908
rect 4296 91964 4360 91968
rect 4296 91908 4300 91964
rect 4300 91908 4356 91964
rect 4356 91908 4360 91964
rect 4296 91904 4360 91908
rect 4376 91964 4440 91968
rect 4376 91908 4380 91964
rect 4380 91908 4436 91964
rect 4436 91908 4440 91964
rect 4376 91904 4440 91908
rect 4456 91964 4520 91968
rect 4456 91908 4460 91964
rect 4460 91908 4516 91964
rect 4516 91908 4520 91964
rect 4456 91904 4520 91908
rect 96376 91964 96440 91968
rect 96376 91908 96380 91964
rect 96380 91908 96436 91964
rect 96436 91908 96440 91964
rect 96376 91904 96440 91908
rect 96456 91964 96520 91968
rect 96456 91908 96460 91964
rect 96460 91908 96516 91964
rect 96516 91908 96520 91964
rect 96456 91904 96520 91908
rect 96536 91964 96600 91968
rect 96536 91908 96540 91964
rect 96540 91908 96596 91964
rect 96596 91908 96600 91964
rect 96536 91904 96600 91908
rect 96616 91964 96680 91968
rect 96616 91908 96620 91964
rect 96620 91908 96676 91964
rect 96676 91908 96680 91964
rect 96616 91904 96680 91908
rect 4876 91420 4940 91424
rect 4876 91364 4880 91420
rect 4880 91364 4936 91420
rect 4936 91364 4940 91420
rect 4876 91360 4940 91364
rect 4956 91420 5020 91424
rect 4956 91364 4960 91420
rect 4960 91364 5016 91420
rect 5016 91364 5020 91420
rect 4956 91360 5020 91364
rect 5036 91420 5100 91424
rect 5036 91364 5040 91420
rect 5040 91364 5096 91420
rect 5096 91364 5100 91420
rect 5036 91360 5100 91364
rect 5116 91420 5180 91424
rect 5116 91364 5120 91420
rect 5120 91364 5176 91420
rect 5176 91364 5180 91420
rect 5116 91360 5180 91364
rect 97036 91420 97100 91424
rect 97036 91364 97040 91420
rect 97040 91364 97096 91420
rect 97096 91364 97100 91420
rect 97036 91360 97100 91364
rect 97116 91420 97180 91424
rect 97116 91364 97120 91420
rect 97120 91364 97176 91420
rect 97176 91364 97180 91420
rect 97116 91360 97180 91364
rect 97196 91420 97260 91424
rect 97196 91364 97200 91420
rect 97200 91364 97256 91420
rect 97256 91364 97260 91420
rect 97196 91360 97260 91364
rect 97276 91420 97340 91424
rect 97276 91364 97280 91420
rect 97280 91364 97336 91420
rect 97336 91364 97340 91420
rect 97276 91360 97340 91364
rect 4216 90876 4280 90880
rect 4216 90820 4220 90876
rect 4220 90820 4276 90876
rect 4276 90820 4280 90876
rect 4216 90816 4280 90820
rect 4296 90876 4360 90880
rect 4296 90820 4300 90876
rect 4300 90820 4356 90876
rect 4356 90820 4360 90876
rect 4296 90816 4360 90820
rect 4376 90876 4440 90880
rect 4376 90820 4380 90876
rect 4380 90820 4436 90876
rect 4436 90820 4440 90876
rect 4376 90816 4440 90820
rect 4456 90876 4520 90880
rect 4456 90820 4460 90876
rect 4460 90820 4516 90876
rect 4516 90820 4520 90876
rect 4456 90816 4520 90820
rect 96376 90876 96440 90880
rect 96376 90820 96380 90876
rect 96380 90820 96436 90876
rect 96436 90820 96440 90876
rect 96376 90816 96440 90820
rect 96456 90876 96520 90880
rect 96456 90820 96460 90876
rect 96460 90820 96516 90876
rect 96516 90820 96520 90876
rect 96456 90816 96520 90820
rect 96536 90876 96600 90880
rect 96536 90820 96540 90876
rect 96540 90820 96596 90876
rect 96596 90820 96600 90876
rect 96536 90816 96600 90820
rect 96616 90876 96680 90880
rect 96616 90820 96620 90876
rect 96620 90820 96676 90876
rect 96676 90820 96680 90876
rect 96616 90816 96680 90820
rect 50844 90476 50908 90540
rect 4876 90332 4940 90336
rect 4876 90276 4880 90332
rect 4880 90276 4936 90332
rect 4936 90276 4940 90332
rect 4876 90272 4940 90276
rect 4956 90332 5020 90336
rect 4956 90276 4960 90332
rect 4960 90276 5016 90332
rect 5016 90276 5020 90332
rect 4956 90272 5020 90276
rect 5036 90332 5100 90336
rect 5036 90276 5040 90332
rect 5040 90276 5096 90332
rect 5096 90276 5100 90332
rect 5036 90272 5100 90276
rect 5116 90332 5180 90336
rect 5116 90276 5120 90332
rect 5120 90276 5176 90332
rect 5176 90276 5180 90332
rect 5116 90272 5180 90276
rect 97036 90332 97100 90336
rect 97036 90276 97040 90332
rect 97040 90276 97096 90332
rect 97096 90276 97100 90332
rect 97036 90272 97100 90276
rect 97116 90332 97180 90336
rect 97116 90276 97120 90332
rect 97120 90276 97176 90332
rect 97176 90276 97180 90332
rect 97116 90272 97180 90276
rect 97196 90332 97260 90336
rect 97196 90276 97200 90332
rect 97200 90276 97256 90332
rect 97256 90276 97260 90332
rect 97196 90272 97260 90276
rect 97276 90332 97340 90336
rect 97276 90276 97280 90332
rect 97280 90276 97336 90332
rect 97336 90276 97340 90332
rect 97276 90272 97340 90276
rect 4216 89788 4280 89792
rect 4216 89732 4220 89788
rect 4220 89732 4276 89788
rect 4276 89732 4280 89788
rect 4216 89728 4280 89732
rect 4296 89788 4360 89792
rect 4296 89732 4300 89788
rect 4300 89732 4356 89788
rect 4356 89732 4360 89788
rect 4296 89728 4360 89732
rect 4376 89788 4440 89792
rect 4376 89732 4380 89788
rect 4380 89732 4436 89788
rect 4436 89732 4440 89788
rect 4376 89728 4440 89732
rect 4456 89788 4520 89792
rect 4456 89732 4460 89788
rect 4460 89732 4516 89788
rect 4516 89732 4520 89788
rect 4456 89728 4520 89732
rect 96376 89788 96440 89792
rect 96376 89732 96380 89788
rect 96380 89732 96436 89788
rect 96436 89732 96440 89788
rect 96376 89728 96440 89732
rect 96456 89788 96520 89792
rect 96456 89732 96460 89788
rect 96460 89732 96516 89788
rect 96516 89732 96520 89788
rect 96456 89728 96520 89732
rect 96536 89788 96600 89792
rect 96536 89732 96540 89788
rect 96540 89732 96596 89788
rect 96596 89732 96600 89788
rect 96536 89728 96600 89732
rect 96616 89788 96680 89792
rect 96616 89732 96620 89788
rect 96620 89732 96676 89788
rect 96676 89732 96680 89788
rect 96616 89728 96680 89732
rect 4876 89244 4940 89248
rect 4876 89188 4880 89244
rect 4880 89188 4936 89244
rect 4936 89188 4940 89244
rect 4876 89184 4940 89188
rect 4956 89244 5020 89248
rect 4956 89188 4960 89244
rect 4960 89188 5016 89244
rect 5016 89188 5020 89244
rect 4956 89184 5020 89188
rect 5036 89244 5100 89248
rect 5036 89188 5040 89244
rect 5040 89188 5096 89244
rect 5096 89188 5100 89244
rect 5036 89184 5100 89188
rect 5116 89244 5180 89248
rect 5116 89188 5120 89244
rect 5120 89188 5176 89244
rect 5176 89188 5180 89244
rect 5116 89184 5180 89188
rect 97036 89244 97100 89248
rect 97036 89188 97040 89244
rect 97040 89188 97096 89244
rect 97096 89188 97100 89244
rect 97036 89184 97100 89188
rect 97116 89244 97180 89248
rect 97116 89188 97120 89244
rect 97120 89188 97176 89244
rect 97176 89188 97180 89244
rect 97116 89184 97180 89188
rect 97196 89244 97260 89248
rect 97196 89188 97200 89244
rect 97200 89188 97256 89244
rect 97256 89188 97260 89244
rect 97196 89184 97260 89188
rect 97276 89244 97340 89248
rect 97276 89188 97280 89244
rect 97280 89188 97336 89244
rect 97336 89188 97340 89244
rect 97276 89184 97340 89188
rect 4216 88700 4280 88704
rect 4216 88644 4220 88700
rect 4220 88644 4276 88700
rect 4276 88644 4280 88700
rect 4216 88640 4280 88644
rect 4296 88700 4360 88704
rect 4296 88644 4300 88700
rect 4300 88644 4356 88700
rect 4356 88644 4360 88700
rect 4296 88640 4360 88644
rect 4376 88700 4440 88704
rect 4376 88644 4380 88700
rect 4380 88644 4436 88700
rect 4436 88644 4440 88700
rect 4376 88640 4440 88644
rect 4456 88700 4520 88704
rect 4456 88644 4460 88700
rect 4460 88644 4516 88700
rect 4516 88644 4520 88700
rect 4456 88640 4520 88644
rect 96376 88700 96440 88704
rect 96376 88644 96380 88700
rect 96380 88644 96436 88700
rect 96436 88644 96440 88700
rect 96376 88640 96440 88644
rect 96456 88700 96520 88704
rect 96456 88644 96460 88700
rect 96460 88644 96516 88700
rect 96516 88644 96520 88700
rect 96456 88640 96520 88644
rect 96536 88700 96600 88704
rect 96536 88644 96540 88700
rect 96540 88644 96596 88700
rect 96596 88644 96600 88700
rect 96536 88640 96600 88644
rect 96616 88700 96680 88704
rect 96616 88644 96620 88700
rect 96620 88644 96676 88700
rect 96676 88644 96680 88700
rect 96616 88640 96680 88644
rect 4876 88156 4940 88160
rect 4876 88100 4880 88156
rect 4880 88100 4936 88156
rect 4936 88100 4940 88156
rect 4876 88096 4940 88100
rect 4956 88156 5020 88160
rect 4956 88100 4960 88156
rect 4960 88100 5016 88156
rect 5016 88100 5020 88156
rect 4956 88096 5020 88100
rect 5036 88156 5100 88160
rect 5036 88100 5040 88156
rect 5040 88100 5096 88156
rect 5096 88100 5100 88156
rect 5036 88096 5100 88100
rect 5116 88156 5180 88160
rect 5116 88100 5120 88156
rect 5120 88100 5176 88156
rect 5176 88100 5180 88156
rect 5116 88096 5180 88100
rect 97036 88156 97100 88160
rect 97036 88100 97040 88156
rect 97040 88100 97096 88156
rect 97096 88100 97100 88156
rect 97036 88096 97100 88100
rect 97116 88156 97180 88160
rect 97116 88100 97120 88156
rect 97120 88100 97176 88156
rect 97176 88100 97180 88156
rect 97116 88096 97180 88100
rect 97196 88156 97260 88160
rect 97196 88100 97200 88156
rect 97200 88100 97256 88156
rect 97256 88100 97260 88156
rect 97196 88096 97260 88100
rect 97276 88156 97340 88160
rect 97276 88100 97280 88156
rect 97280 88100 97336 88156
rect 97336 88100 97340 88156
rect 97276 88096 97340 88100
rect 4216 87612 4280 87616
rect 4216 87556 4220 87612
rect 4220 87556 4276 87612
rect 4276 87556 4280 87612
rect 4216 87552 4280 87556
rect 4296 87612 4360 87616
rect 4296 87556 4300 87612
rect 4300 87556 4356 87612
rect 4356 87556 4360 87612
rect 4296 87552 4360 87556
rect 4376 87612 4440 87616
rect 4376 87556 4380 87612
rect 4380 87556 4436 87612
rect 4436 87556 4440 87612
rect 4376 87552 4440 87556
rect 4456 87612 4520 87616
rect 4456 87556 4460 87612
rect 4460 87556 4516 87612
rect 4516 87556 4520 87612
rect 4456 87552 4520 87556
rect 96376 87612 96440 87616
rect 96376 87556 96380 87612
rect 96380 87556 96436 87612
rect 96436 87556 96440 87612
rect 96376 87552 96440 87556
rect 96456 87612 96520 87616
rect 96456 87556 96460 87612
rect 96460 87556 96516 87612
rect 96516 87556 96520 87612
rect 96456 87552 96520 87556
rect 96536 87612 96600 87616
rect 96536 87556 96540 87612
rect 96540 87556 96596 87612
rect 96596 87556 96600 87612
rect 96536 87552 96600 87556
rect 96616 87612 96680 87616
rect 96616 87556 96620 87612
rect 96620 87556 96676 87612
rect 96676 87556 96680 87612
rect 96616 87552 96680 87556
rect 4876 87068 4940 87072
rect 4876 87012 4880 87068
rect 4880 87012 4936 87068
rect 4936 87012 4940 87068
rect 4876 87008 4940 87012
rect 4956 87068 5020 87072
rect 4956 87012 4960 87068
rect 4960 87012 5016 87068
rect 5016 87012 5020 87068
rect 4956 87008 5020 87012
rect 5036 87068 5100 87072
rect 5036 87012 5040 87068
rect 5040 87012 5096 87068
rect 5096 87012 5100 87068
rect 5036 87008 5100 87012
rect 5116 87068 5180 87072
rect 5116 87012 5120 87068
rect 5120 87012 5176 87068
rect 5176 87012 5180 87068
rect 5116 87008 5180 87012
rect 97036 87068 97100 87072
rect 97036 87012 97040 87068
rect 97040 87012 97096 87068
rect 97096 87012 97100 87068
rect 97036 87008 97100 87012
rect 97116 87068 97180 87072
rect 97116 87012 97120 87068
rect 97120 87012 97176 87068
rect 97176 87012 97180 87068
rect 97116 87008 97180 87012
rect 97196 87068 97260 87072
rect 97196 87012 97200 87068
rect 97200 87012 97256 87068
rect 97256 87012 97260 87068
rect 97196 87008 97260 87012
rect 97276 87068 97340 87072
rect 97276 87012 97280 87068
rect 97280 87012 97336 87068
rect 97336 87012 97340 87068
rect 97276 87008 97340 87012
rect 4216 86524 4280 86528
rect 4216 86468 4220 86524
rect 4220 86468 4276 86524
rect 4276 86468 4280 86524
rect 4216 86464 4280 86468
rect 4296 86524 4360 86528
rect 4296 86468 4300 86524
rect 4300 86468 4356 86524
rect 4356 86468 4360 86524
rect 4296 86464 4360 86468
rect 4376 86524 4440 86528
rect 4376 86468 4380 86524
rect 4380 86468 4436 86524
rect 4436 86468 4440 86524
rect 4376 86464 4440 86468
rect 4456 86524 4520 86528
rect 4456 86468 4460 86524
rect 4460 86468 4516 86524
rect 4516 86468 4520 86524
rect 4456 86464 4520 86468
rect 96376 86524 96440 86528
rect 96376 86468 96380 86524
rect 96380 86468 96436 86524
rect 96436 86468 96440 86524
rect 96376 86464 96440 86468
rect 96456 86524 96520 86528
rect 96456 86468 96460 86524
rect 96460 86468 96516 86524
rect 96516 86468 96520 86524
rect 96456 86464 96520 86468
rect 96536 86524 96600 86528
rect 96536 86468 96540 86524
rect 96540 86468 96596 86524
rect 96596 86468 96600 86524
rect 96536 86464 96600 86468
rect 96616 86524 96680 86528
rect 96616 86468 96620 86524
rect 96620 86468 96676 86524
rect 96676 86468 96680 86524
rect 96616 86464 96680 86468
rect 4876 85980 4940 85984
rect 4876 85924 4880 85980
rect 4880 85924 4936 85980
rect 4936 85924 4940 85980
rect 4876 85920 4940 85924
rect 4956 85980 5020 85984
rect 4956 85924 4960 85980
rect 4960 85924 5016 85980
rect 5016 85924 5020 85980
rect 4956 85920 5020 85924
rect 5036 85980 5100 85984
rect 5036 85924 5040 85980
rect 5040 85924 5096 85980
rect 5096 85924 5100 85980
rect 5036 85920 5100 85924
rect 5116 85980 5180 85984
rect 5116 85924 5120 85980
rect 5120 85924 5176 85980
rect 5176 85924 5180 85980
rect 5116 85920 5180 85924
rect 97036 85980 97100 85984
rect 97036 85924 97040 85980
rect 97040 85924 97096 85980
rect 97096 85924 97100 85980
rect 97036 85920 97100 85924
rect 97116 85980 97180 85984
rect 97116 85924 97120 85980
rect 97120 85924 97176 85980
rect 97176 85924 97180 85980
rect 97116 85920 97180 85924
rect 97196 85980 97260 85984
rect 97196 85924 97200 85980
rect 97200 85924 97256 85980
rect 97256 85924 97260 85980
rect 97196 85920 97260 85924
rect 97276 85980 97340 85984
rect 97276 85924 97280 85980
rect 97280 85924 97336 85980
rect 97336 85924 97340 85980
rect 97276 85920 97340 85924
rect 4216 85436 4280 85440
rect 4216 85380 4220 85436
rect 4220 85380 4276 85436
rect 4276 85380 4280 85436
rect 4216 85376 4280 85380
rect 4296 85436 4360 85440
rect 4296 85380 4300 85436
rect 4300 85380 4356 85436
rect 4356 85380 4360 85436
rect 4296 85376 4360 85380
rect 4376 85436 4440 85440
rect 4376 85380 4380 85436
rect 4380 85380 4436 85436
rect 4436 85380 4440 85436
rect 4376 85376 4440 85380
rect 4456 85436 4520 85440
rect 4456 85380 4460 85436
rect 4460 85380 4516 85436
rect 4516 85380 4520 85436
rect 4456 85376 4520 85380
rect 96376 85436 96440 85440
rect 96376 85380 96380 85436
rect 96380 85380 96436 85436
rect 96436 85380 96440 85436
rect 96376 85376 96440 85380
rect 96456 85436 96520 85440
rect 96456 85380 96460 85436
rect 96460 85380 96516 85436
rect 96516 85380 96520 85436
rect 96456 85376 96520 85380
rect 96536 85436 96600 85440
rect 96536 85380 96540 85436
rect 96540 85380 96596 85436
rect 96596 85380 96600 85436
rect 96536 85376 96600 85380
rect 96616 85436 96680 85440
rect 96616 85380 96620 85436
rect 96620 85380 96676 85436
rect 96676 85380 96680 85436
rect 96616 85376 96680 85380
rect 4876 84892 4940 84896
rect 4876 84836 4880 84892
rect 4880 84836 4936 84892
rect 4936 84836 4940 84892
rect 4876 84832 4940 84836
rect 4956 84892 5020 84896
rect 4956 84836 4960 84892
rect 4960 84836 5016 84892
rect 5016 84836 5020 84892
rect 4956 84832 5020 84836
rect 5036 84892 5100 84896
rect 5036 84836 5040 84892
rect 5040 84836 5096 84892
rect 5096 84836 5100 84892
rect 5036 84832 5100 84836
rect 5116 84892 5180 84896
rect 5116 84836 5120 84892
rect 5120 84836 5176 84892
rect 5176 84836 5180 84892
rect 5116 84832 5180 84836
rect 97036 84892 97100 84896
rect 97036 84836 97040 84892
rect 97040 84836 97096 84892
rect 97096 84836 97100 84892
rect 97036 84832 97100 84836
rect 97116 84892 97180 84896
rect 97116 84836 97120 84892
rect 97120 84836 97176 84892
rect 97176 84836 97180 84892
rect 97116 84832 97180 84836
rect 97196 84892 97260 84896
rect 97196 84836 97200 84892
rect 97200 84836 97256 84892
rect 97256 84836 97260 84892
rect 97196 84832 97260 84836
rect 97276 84892 97340 84896
rect 97276 84836 97280 84892
rect 97280 84836 97336 84892
rect 97336 84836 97340 84892
rect 97276 84832 97340 84836
rect 4216 84348 4280 84352
rect 4216 84292 4220 84348
rect 4220 84292 4276 84348
rect 4276 84292 4280 84348
rect 4216 84288 4280 84292
rect 4296 84348 4360 84352
rect 4296 84292 4300 84348
rect 4300 84292 4356 84348
rect 4356 84292 4360 84348
rect 4296 84288 4360 84292
rect 4376 84348 4440 84352
rect 4376 84292 4380 84348
rect 4380 84292 4436 84348
rect 4436 84292 4440 84348
rect 4376 84288 4440 84292
rect 4456 84348 4520 84352
rect 4456 84292 4460 84348
rect 4460 84292 4516 84348
rect 4516 84292 4520 84348
rect 4456 84288 4520 84292
rect 96376 84348 96440 84352
rect 96376 84292 96380 84348
rect 96380 84292 96436 84348
rect 96436 84292 96440 84348
rect 96376 84288 96440 84292
rect 96456 84348 96520 84352
rect 96456 84292 96460 84348
rect 96460 84292 96516 84348
rect 96516 84292 96520 84348
rect 96456 84288 96520 84292
rect 96536 84348 96600 84352
rect 96536 84292 96540 84348
rect 96540 84292 96596 84348
rect 96596 84292 96600 84348
rect 96536 84288 96600 84292
rect 96616 84348 96680 84352
rect 96616 84292 96620 84348
rect 96620 84292 96676 84348
rect 96676 84292 96680 84348
rect 96616 84288 96680 84292
rect 4876 83804 4940 83808
rect 4876 83748 4880 83804
rect 4880 83748 4936 83804
rect 4936 83748 4940 83804
rect 4876 83744 4940 83748
rect 4956 83804 5020 83808
rect 4956 83748 4960 83804
rect 4960 83748 5016 83804
rect 5016 83748 5020 83804
rect 4956 83744 5020 83748
rect 5036 83804 5100 83808
rect 5036 83748 5040 83804
rect 5040 83748 5096 83804
rect 5096 83748 5100 83804
rect 5036 83744 5100 83748
rect 5116 83804 5180 83808
rect 5116 83748 5120 83804
rect 5120 83748 5176 83804
rect 5176 83748 5180 83804
rect 5116 83744 5180 83748
rect 97036 83804 97100 83808
rect 97036 83748 97040 83804
rect 97040 83748 97096 83804
rect 97096 83748 97100 83804
rect 97036 83744 97100 83748
rect 97116 83804 97180 83808
rect 97116 83748 97120 83804
rect 97120 83748 97176 83804
rect 97176 83748 97180 83804
rect 97116 83744 97180 83748
rect 97196 83804 97260 83808
rect 97196 83748 97200 83804
rect 97200 83748 97256 83804
rect 97256 83748 97260 83804
rect 97196 83744 97260 83748
rect 97276 83804 97340 83808
rect 97276 83748 97280 83804
rect 97280 83748 97336 83804
rect 97336 83748 97340 83804
rect 97276 83744 97340 83748
rect 4216 83260 4280 83264
rect 4216 83204 4220 83260
rect 4220 83204 4276 83260
rect 4276 83204 4280 83260
rect 4216 83200 4280 83204
rect 4296 83260 4360 83264
rect 4296 83204 4300 83260
rect 4300 83204 4356 83260
rect 4356 83204 4360 83260
rect 4296 83200 4360 83204
rect 4376 83260 4440 83264
rect 4376 83204 4380 83260
rect 4380 83204 4436 83260
rect 4436 83204 4440 83260
rect 4376 83200 4440 83204
rect 4456 83260 4520 83264
rect 4456 83204 4460 83260
rect 4460 83204 4516 83260
rect 4516 83204 4520 83260
rect 4456 83200 4520 83204
rect 96376 83260 96440 83264
rect 96376 83204 96380 83260
rect 96380 83204 96436 83260
rect 96436 83204 96440 83260
rect 96376 83200 96440 83204
rect 96456 83260 96520 83264
rect 96456 83204 96460 83260
rect 96460 83204 96516 83260
rect 96516 83204 96520 83260
rect 96456 83200 96520 83204
rect 96536 83260 96600 83264
rect 96536 83204 96540 83260
rect 96540 83204 96596 83260
rect 96596 83204 96600 83260
rect 96536 83200 96600 83204
rect 96616 83260 96680 83264
rect 96616 83204 96620 83260
rect 96620 83204 96676 83260
rect 96676 83204 96680 83260
rect 96616 83200 96680 83204
rect 4876 82716 4940 82720
rect 4876 82660 4880 82716
rect 4880 82660 4936 82716
rect 4936 82660 4940 82716
rect 4876 82656 4940 82660
rect 4956 82716 5020 82720
rect 4956 82660 4960 82716
rect 4960 82660 5016 82716
rect 5016 82660 5020 82716
rect 4956 82656 5020 82660
rect 5036 82716 5100 82720
rect 5036 82660 5040 82716
rect 5040 82660 5096 82716
rect 5096 82660 5100 82716
rect 5036 82656 5100 82660
rect 5116 82716 5180 82720
rect 5116 82660 5120 82716
rect 5120 82660 5176 82716
rect 5176 82660 5180 82716
rect 5116 82656 5180 82660
rect 97036 82716 97100 82720
rect 97036 82660 97040 82716
rect 97040 82660 97096 82716
rect 97096 82660 97100 82716
rect 97036 82656 97100 82660
rect 97116 82716 97180 82720
rect 97116 82660 97120 82716
rect 97120 82660 97176 82716
rect 97176 82660 97180 82716
rect 97116 82656 97180 82660
rect 97196 82716 97260 82720
rect 97196 82660 97200 82716
rect 97200 82660 97256 82716
rect 97256 82660 97260 82716
rect 97196 82656 97260 82660
rect 97276 82716 97340 82720
rect 97276 82660 97280 82716
rect 97280 82660 97336 82716
rect 97336 82660 97340 82716
rect 97276 82656 97340 82660
rect 4216 82172 4280 82176
rect 4216 82116 4220 82172
rect 4220 82116 4276 82172
rect 4276 82116 4280 82172
rect 4216 82112 4280 82116
rect 4296 82172 4360 82176
rect 4296 82116 4300 82172
rect 4300 82116 4356 82172
rect 4356 82116 4360 82172
rect 4296 82112 4360 82116
rect 4376 82172 4440 82176
rect 4376 82116 4380 82172
rect 4380 82116 4436 82172
rect 4436 82116 4440 82172
rect 4376 82112 4440 82116
rect 4456 82172 4520 82176
rect 4456 82116 4460 82172
rect 4460 82116 4516 82172
rect 4516 82116 4520 82172
rect 4456 82112 4520 82116
rect 96376 82172 96440 82176
rect 96376 82116 96380 82172
rect 96380 82116 96436 82172
rect 96436 82116 96440 82172
rect 96376 82112 96440 82116
rect 96456 82172 96520 82176
rect 96456 82116 96460 82172
rect 96460 82116 96516 82172
rect 96516 82116 96520 82172
rect 96456 82112 96520 82116
rect 96536 82172 96600 82176
rect 96536 82116 96540 82172
rect 96540 82116 96596 82172
rect 96596 82116 96600 82172
rect 96536 82112 96600 82116
rect 96616 82172 96680 82176
rect 96616 82116 96620 82172
rect 96620 82116 96676 82172
rect 96676 82116 96680 82172
rect 96616 82112 96680 82116
rect 4876 81628 4940 81632
rect 4876 81572 4880 81628
rect 4880 81572 4936 81628
rect 4936 81572 4940 81628
rect 4876 81568 4940 81572
rect 4956 81628 5020 81632
rect 4956 81572 4960 81628
rect 4960 81572 5016 81628
rect 5016 81572 5020 81628
rect 4956 81568 5020 81572
rect 5036 81628 5100 81632
rect 5036 81572 5040 81628
rect 5040 81572 5096 81628
rect 5096 81572 5100 81628
rect 5036 81568 5100 81572
rect 5116 81628 5180 81632
rect 5116 81572 5120 81628
rect 5120 81572 5176 81628
rect 5176 81572 5180 81628
rect 5116 81568 5180 81572
rect 97036 81628 97100 81632
rect 97036 81572 97040 81628
rect 97040 81572 97096 81628
rect 97096 81572 97100 81628
rect 97036 81568 97100 81572
rect 97116 81628 97180 81632
rect 97116 81572 97120 81628
rect 97120 81572 97176 81628
rect 97176 81572 97180 81628
rect 97116 81568 97180 81572
rect 97196 81628 97260 81632
rect 97196 81572 97200 81628
rect 97200 81572 97256 81628
rect 97256 81572 97260 81628
rect 97196 81568 97260 81572
rect 97276 81628 97340 81632
rect 97276 81572 97280 81628
rect 97280 81572 97336 81628
rect 97336 81572 97340 81628
rect 97276 81568 97340 81572
rect 4216 81084 4280 81088
rect 4216 81028 4220 81084
rect 4220 81028 4276 81084
rect 4276 81028 4280 81084
rect 4216 81024 4280 81028
rect 4296 81084 4360 81088
rect 4296 81028 4300 81084
rect 4300 81028 4356 81084
rect 4356 81028 4360 81084
rect 4296 81024 4360 81028
rect 4376 81084 4440 81088
rect 4376 81028 4380 81084
rect 4380 81028 4436 81084
rect 4436 81028 4440 81084
rect 4376 81024 4440 81028
rect 4456 81084 4520 81088
rect 4456 81028 4460 81084
rect 4460 81028 4516 81084
rect 4516 81028 4520 81084
rect 4456 81024 4520 81028
rect 96376 81084 96440 81088
rect 96376 81028 96380 81084
rect 96380 81028 96436 81084
rect 96436 81028 96440 81084
rect 96376 81024 96440 81028
rect 96456 81084 96520 81088
rect 96456 81028 96460 81084
rect 96460 81028 96516 81084
rect 96516 81028 96520 81084
rect 96456 81024 96520 81028
rect 96536 81084 96600 81088
rect 96536 81028 96540 81084
rect 96540 81028 96596 81084
rect 96596 81028 96600 81084
rect 96536 81024 96600 81028
rect 96616 81084 96680 81088
rect 96616 81028 96620 81084
rect 96620 81028 96676 81084
rect 96676 81028 96680 81084
rect 96616 81024 96680 81028
rect 4876 80540 4940 80544
rect 4876 80484 4880 80540
rect 4880 80484 4936 80540
rect 4936 80484 4940 80540
rect 4876 80480 4940 80484
rect 4956 80540 5020 80544
rect 4956 80484 4960 80540
rect 4960 80484 5016 80540
rect 5016 80484 5020 80540
rect 4956 80480 5020 80484
rect 5036 80540 5100 80544
rect 5036 80484 5040 80540
rect 5040 80484 5096 80540
rect 5096 80484 5100 80540
rect 5036 80480 5100 80484
rect 5116 80540 5180 80544
rect 5116 80484 5120 80540
rect 5120 80484 5176 80540
rect 5176 80484 5180 80540
rect 5116 80480 5180 80484
rect 97036 80540 97100 80544
rect 97036 80484 97040 80540
rect 97040 80484 97096 80540
rect 97096 80484 97100 80540
rect 97036 80480 97100 80484
rect 97116 80540 97180 80544
rect 97116 80484 97120 80540
rect 97120 80484 97176 80540
rect 97176 80484 97180 80540
rect 97116 80480 97180 80484
rect 97196 80540 97260 80544
rect 97196 80484 97200 80540
rect 97200 80484 97256 80540
rect 97256 80484 97260 80540
rect 97196 80480 97260 80484
rect 97276 80540 97340 80544
rect 97276 80484 97280 80540
rect 97280 80484 97336 80540
rect 97336 80484 97340 80540
rect 97276 80480 97340 80484
rect 4216 79996 4280 80000
rect 4216 79940 4220 79996
rect 4220 79940 4276 79996
rect 4276 79940 4280 79996
rect 4216 79936 4280 79940
rect 4296 79996 4360 80000
rect 4296 79940 4300 79996
rect 4300 79940 4356 79996
rect 4356 79940 4360 79996
rect 4296 79936 4360 79940
rect 4376 79996 4440 80000
rect 4376 79940 4380 79996
rect 4380 79940 4436 79996
rect 4436 79940 4440 79996
rect 4376 79936 4440 79940
rect 4456 79996 4520 80000
rect 4456 79940 4460 79996
rect 4460 79940 4516 79996
rect 4516 79940 4520 79996
rect 4456 79936 4520 79940
rect 96376 79996 96440 80000
rect 96376 79940 96380 79996
rect 96380 79940 96436 79996
rect 96436 79940 96440 79996
rect 96376 79936 96440 79940
rect 96456 79996 96520 80000
rect 96456 79940 96460 79996
rect 96460 79940 96516 79996
rect 96516 79940 96520 79996
rect 96456 79936 96520 79940
rect 96536 79996 96600 80000
rect 96536 79940 96540 79996
rect 96540 79940 96596 79996
rect 96596 79940 96600 79996
rect 96536 79936 96600 79940
rect 96616 79996 96680 80000
rect 96616 79940 96620 79996
rect 96620 79940 96676 79996
rect 96676 79940 96680 79996
rect 96616 79936 96680 79940
rect 4876 79452 4940 79456
rect 4876 79396 4880 79452
rect 4880 79396 4936 79452
rect 4936 79396 4940 79452
rect 4876 79392 4940 79396
rect 4956 79452 5020 79456
rect 4956 79396 4960 79452
rect 4960 79396 5016 79452
rect 5016 79396 5020 79452
rect 4956 79392 5020 79396
rect 5036 79452 5100 79456
rect 5036 79396 5040 79452
rect 5040 79396 5096 79452
rect 5096 79396 5100 79452
rect 5036 79392 5100 79396
rect 5116 79452 5180 79456
rect 5116 79396 5120 79452
rect 5120 79396 5176 79452
rect 5176 79396 5180 79452
rect 5116 79392 5180 79396
rect 97036 79452 97100 79456
rect 97036 79396 97040 79452
rect 97040 79396 97096 79452
rect 97096 79396 97100 79452
rect 97036 79392 97100 79396
rect 97116 79452 97180 79456
rect 97116 79396 97120 79452
rect 97120 79396 97176 79452
rect 97176 79396 97180 79452
rect 97116 79392 97180 79396
rect 97196 79452 97260 79456
rect 97196 79396 97200 79452
rect 97200 79396 97256 79452
rect 97256 79396 97260 79452
rect 97196 79392 97260 79396
rect 97276 79452 97340 79456
rect 97276 79396 97280 79452
rect 97280 79396 97336 79452
rect 97336 79396 97340 79452
rect 97276 79392 97340 79396
rect 4216 78908 4280 78912
rect 4216 78852 4220 78908
rect 4220 78852 4276 78908
rect 4276 78852 4280 78908
rect 4216 78848 4280 78852
rect 4296 78908 4360 78912
rect 4296 78852 4300 78908
rect 4300 78852 4356 78908
rect 4356 78852 4360 78908
rect 4296 78848 4360 78852
rect 4376 78908 4440 78912
rect 4376 78852 4380 78908
rect 4380 78852 4436 78908
rect 4436 78852 4440 78908
rect 4376 78848 4440 78852
rect 4456 78908 4520 78912
rect 4456 78852 4460 78908
rect 4460 78852 4516 78908
rect 4516 78852 4520 78908
rect 4456 78848 4520 78852
rect 96376 78908 96440 78912
rect 96376 78852 96380 78908
rect 96380 78852 96436 78908
rect 96436 78852 96440 78908
rect 96376 78848 96440 78852
rect 96456 78908 96520 78912
rect 96456 78852 96460 78908
rect 96460 78852 96516 78908
rect 96516 78852 96520 78908
rect 96456 78848 96520 78852
rect 96536 78908 96600 78912
rect 96536 78852 96540 78908
rect 96540 78852 96596 78908
rect 96596 78852 96600 78908
rect 96536 78848 96600 78852
rect 96616 78908 96680 78912
rect 96616 78852 96620 78908
rect 96620 78852 96676 78908
rect 96676 78852 96680 78908
rect 96616 78848 96680 78852
rect 4876 78364 4940 78368
rect 4876 78308 4880 78364
rect 4880 78308 4936 78364
rect 4936 78308 4940 78364
rect 4876 78304 4940 78308
rect 4956 78364 5020 78368
rect 4956 78308 4960 78364
rect 4960 78308 5016 78364
rect 5016 78308 5020 78364
rect 4956 78304 5020 78308
rect 5036 78364 5100 78368
rect 5036 78308 5040 78364
rect 5040 78308 5096 78364
rect 5096 78308 5100 78364
rect 5036 78304 5100 78308
rect 5116 78364 5180 78368
rect 5116 78308 5120 78364
rect 5120 78308 5176 78364
rect 5176 78308 5180 78364
rect 5116 78304 5180 78308
rect 97036 78364 97100 78368
rect 97036 78308 97040 78364
rect 97040 78308 97096 78364
rect 97096 78308 97100 78364
rect 97036 78304 97100 78308
rect 97116 78364 97180 78368
rect 97116 78308 97120 78364
rect 97120 78308 97176 78364
rect 97176 78308 97180 78364
rect 97116 78304 97180 78308
rect 97196 78364 97260 78368
rect 97196 78308 97200 78364
rect 97200 78308 97256 78364
rect 97256 78308 97260 78364
rect 97196 78304 97260 78308
rect 97276 78364 97340 78368
rect 97276 78308 97280 78364
rect 97280 78308 97336 78364
rect 97336 78308 97340 78364
rect 97276 78304 97340 78308
rect 4216 77820 4280 77824
rect 4216 77764 4220 77820
rect 4220 77764 4276 77820
rect 4276 77764 4280 77820
rect 4216 77760 4280 77764
rect 4296 77820 4360 77824
rect 4296 77764 4300 77820
rect 4300 77764 4356 77820
rect 4356 77764 4360 77820
rect 4296 77760 4360 77764
rect 4376 77820 4440 77824
rect 4376 77764 4380 77820
rect 4380 77764 4436 77820
rect 4436 77764 4440 77820
rect 4376 77760 4440 77764
rect 4456 77820 4520 77824
rect 4456 77764 4460 77820
rect 4460 77764 4516 77820
rect 4516 77764 4520 77820
rect 4456 77760 4520 77764
rect 96376 77820 96440 77824
rect 96376 77764 96380 77820
rect 96380 77764 96436 77820
rect 96436 77764 96440 77820
rect 96376 77760 96440 77764
rect 96456 77820 96520 77824
rect 96456 77764 96460 77820
rect 96460 77764 96516 77820
rect 96516 77764 96520 77820
rect 96456 77760 96520 77764
rect 96536 77820 96600 77824
rect 96536 77764 96540 77820
rect 96540 77764 96596 77820
rect 96596 77764 96600 77820
rect 96536 77760 96600 77764
rect 96616 77820 96680 77824
rect 96616 77764 96620 77820
rect 96620 77764 96676 77820
rect 96676 77764 96680 77820
rect 96616 77760 96680 77764
rect 4876 77276 4940 77280
rect 4876 77220 4880 77276
rect 4880 77220 4936 77276
rect 4936 77220 4940 77276
rect 4876 77216 4940 77220
rect 4956 77276 5020 77280
rect 4956 77220 4960 77276
rect 4960 77220 5016 77276
rect 5016 77220 5020 77276
rect 4956 77216 5020 77220
rect 5036 77276 5100 77280
rect 5036 77220 5040 77276
rect 5040 77220 5096 77276
rect 5096 77220 5100 77276
rect 5036 77216 5100 77220
rect 5116 77276 5180 77280
rect 5116 77220 5120 77276
rect 5120 77220 5176 77276
rect 5176 77220 5180 77276
rect 5116 77216 5180 77220
rect 97036 77276 97100 77280
rect 97036 77220 97040 77276
rect 97040 77220 97096 77276
rect 97096 77220 97100 77276
rect 97036 77216 97100 77220
rect 97116 77276 97180 77280
rect 97116 77220 97120 77276
rect 97120 77220 97176 77276
rect 97176 77220 97180 77276
rect 97116 77216 97180 77220
rect 97196 77276 97260 77280
rect 97196 77220 97200 77276
rect 97200 77220 97256 77276
rect 97256 77220 97260 77276
rect 97196 77216 97260 77220
rect 97276 77276 97340 77280
rect 97276 77220 97280 77276
rect 97280 77220 97336 77276
rect 97336 77220 97340 77276
rect 97276 77216 97340 77220
rect 4216 76732 4280 76736
rect 4216 76676 4220 76732
rect 4220 76676 4276 76732
rect 4276 76676 4280 76732
rect 4216 76672 4280 76676
rect 4296 76732 4360 76736
rect 4296 76676 4300 76732
rect 4300 76676 4356 76732
rect 4356 76676 4360 76732
rect 4296 76672 4360 76676
rect 4376 76732 4440 76736
rect 4376 76676 4380 76732
rect 4380 76676 4436 76732
rect 4436 76676 4440 76732
rect 4376 76672 4440 76676
rect 4456 76732 4520 76736
rect 4456 76676 4460 76732
rect 4460 76676 4516 76732
rect 4516 76676 4520 76732
rect 4456 76672 4520 76676
rect 96376 76732 96440 76736
rect 96376 76676 96380 76732
rect 96380 76676 96436 76732
rect 96436 76676 96440 76732
rect 96376 76672 96440 76676
rect 96456 76732 96520 76736
rect 96456 76676 96460 76732
rect 96460 76676 96516 76732
rect 96516 76676 96520 76732
rect 96456 76672 96520 76676
rect 96536 76732 96600 76736
rect 96536 76676 96540 76732
rect 96540 76676 96596 76732
rect 96596 76676 96600 76732
rect 96536 76672 96600 76676
rect 96616 76732 96680 76736
rect 96616 76676 96620 76732
rect 96620 76676 96676 76732
rect 96676 76676 96680 76732
rect 96616 76672 96680 76676
rect 4876 76188 4940 76192
rect 4876 76132 4880 76188
rect 4880 76132 4936 76188
rect 4936 76132 4940 76188
rect 4876 76128 4940 76132
rect 4956 76188 5020 76192
rect 4956 76132 4960 76188
rect 4960 76132 5016 76188
rect 5016 76132 5020 76188
rect 4956 76128 5020 76132
rect 5036 76188 5100 76192
rect 5036 76132 5040 76188
rect 5040 76132 5096 76188
rect 5096 76132 5100 76188
rect 5036 76128 5100 76132
rect 5116 76188 5180 76192
rect 5116 76132 5120 76188
rect 5120 76132 5176 76188
rect 5176 76132 5180 76188
rect 5116 76128 5180 76132
rect 97036 76188 97100 76192
rect 97036 76132 97040 76188
rect 97040 76132 97096 76188
rect 97096 76132 97100 76188
rect 97036 76128 97100 76132
rect 97116 76188 97180 76192
rect 97116 76132 97120 76188
rect 97120 76132 97176 76188
rect 97176 76132 97180 76188
rect 97116 76128 97180 76132
rect 97196 76188 97260 76192
rect 97196 76132 97200 76188
rect 97200 76132 97256 76188
rect 97256 76132 97260 76188
rect 97196 76128 97260 76132
rect 97276 76188 97340 76192
rect 97276 76132 97280 76188
rect 97280 76132 97336 76188
rect 97336 76132 97340 76188
rect 97276 76128 97340 76132
rect 4216 75644 4280 75648
rect 4216 75588 4220 75644
rect 4220 75588 4276 75644
rect 4276 75588 4280 75644
rect 4216 75584 4280 75588
rect 4296 75644 4360 75648
rect 4296 75588 4300 75644
rect 4300 75588 4356 75644
rect 4356 75588 4360 75644
rect 4296 75584 4360 75588
rect 4376 75644 4440 75648
rect 4376 75588 4380 75644
rect 4380 75588 4436 75644
rect 4436 75588 4440 75644
rect 4376 75584 4440 75588
rect 4456 75644 4520 75648
rect 4456 75588 4460 75644
rect 4460 75588 4516 75644
rect 4516 75588 4520 75644
rect 4456 75584 4520 75588
rect 96376 75644 96440 75648
rect 96376 75588 96380 75644
rect 96380 75588 96436 75644
rect 96436 75588 96440 75644
rect 96376 75584 96440 75588
rect 96456 75644 96520 75648
rect 96456 75588 96460 75644
rect 96460 75588 96516 75644
rect 96516 75588 96520 75644
rect 96456 75584 96520 75588
rect 96536 75644 96600 75648
rect 96536 75588 96540 75644
rect 96540 75588 96596 75644
rect 96596 75588 96600 75644
rect 96536 75584 96600 75588
rect 96616 75644 96680 75648
rect 96616 75588 96620 75644
rect 96620 75588 96676 75644
rect 96676 75588 96680 75644
rect 96616 75584 96680 75588
rect 4876 75100 4940 75104
rect 4876 75044 4880 75100
rect 4880 75044 4936 75100
rect 4936 75044 4940 75100
rect 4876 75040 4940 75044
rect 4956 75100 5020 75104
rect 4956 75044 4960 75100
rect 4960 75044 5016 75100
rect 5016 75044 5020 75100
rect 4956 75040 5020 75044
rect 5036 75100 5100 75104
rect 5036 75044 5040 75100
rect 5040 75044 5096 75100
rect 5096 75044 5100 75100
rect 5036 75040 5100 75044
rect 5116 75100 5180 75104
rect 5116 75044 5120 75100
rect 5120 75044 5176 75100
rect 5176 75044 5180 75100
rect 5116 75040 5180 75044
rect 97036 75100 97100 75104
rect 97036 75044 97040 75100
rect 97040 75044 97096 75100
rect 97096 75044 97100 75100
rect 97036 75040 97100 75044
rect 97116 75100 97180 75104
rect 97116 75044 97120 75100
rect 97120 75044 97176 75100
rect 97176 75044 97180 75100
rect 97116 75040 97180 75044
rect 97196 75100 97260 75104
rect 97196 75044 97200 75100
rect 97200 75044 97256 75100
rect 97256 75044 97260 75100
rect 97196 75040 97260 75044
rect 97276 75100 97340 75104
rect 97276 75044 97280 75100
rect 97280 75044 97336 75100
rect 97336 75044 97340 75100
rect 97276 75040 97340 75044
rect 4216 74556 4280 74560
rect 4216 74500 4220 74556
rect 4220 74500 4276 74556
rect 4276 74500 4280 74556
rect 4216 74496 4280 74500
rect 4296 74556 4360 74560
rect 4296 74500 4300 74556
rect 4300 74500 4356 74556
rect 4356 74500 4360 74556
rect 4296 74496 4360 74500
rect 4376 74556 4440 74560
rect 4376 74500 4380 74556
rect 4380 74500 4436 74556
rect 4436 74500 4440 74556
rect 4376 74496 4440 74500
rect 4456 74556 4520 74560
rect 4456 74500 4460 74556
rect 4460 74500 4516 74556
rect 4516 74500 4520 74556
rect 4456 74496 4520 74500
rect 96376 74556 96440 74560
rect 96376 74500 96380 74556
rect 96380 74500 96436 74556
rect 96436 74500 96440 74556
rect 96376 74496 96440 74500
rect 96456 74556 96520 74560
rect 96456 74500 96460 74556
rect 96460 74500 96516 74556
rect 96516 74500 96520 74556
rect 96456 74496 96520 74500
rect 96536 74556 96600 74560
rect 96536 74500 96540 74556
rect 96540 74500 96596 74556
rect 96596 74500 96600 74556
rect 96536 74496 96600 74500
rect 96616 74556 96680 74560
rect 96616 74500 96620 74556
rect 96620 74500 96676 74556
rect 96676 74500 96680 74556
rect 96616 74496 96680 74500
rect 4876 74012 4940 74016
rect 4876 73956 4880 74012
rect 4880 73956 4936 74012
rect 4936 73956 4940 74012
rect 4876 73952 4940 73956
rect 4956 74012 5020 74016
rect 4956 73956 4960 74012
rect 4960 73956 5016 74012
rect 5016 73956 5020 74012
rect 4956 73952 5020 73956
rect 5036 74012 5100 74016
rect 5036 73956 5040 74012
rect 5040 73956 5096 74012
rect 5096 73956 5100 74012
rect 5036 73952 5100 73956
rect 5116 74012 5180 74016
rect 5116 73956 5120 74012
rect 5120 73956 5176 74012
rect 5176 73956 5180 74012
rect 5116 73952 5180 73956
rect 97036 74012 97100 74016
rect 97036 73956 97040 74012
rect 97040 73956 97096 74012
rect 97096 73956 97100 74012
rect 97036 73952 97100 73956
rect 97116 74012 97180 74016
rect 97116 73956 97120 74012
rect 97120 73956 97176 74012
rect 97176 73956 97180 74012
rect 97116 73952 97180 73956
rect 97196 74012 97260 74016
rect 97196 73956 97200 74012
rect 97200 73956 97256 74012
rect 97256 73956 97260 74012
rect 97196 73952 97260 73956
rect 97276 74012 97340 74016
rect 97276 73956 97280 74012
rect 97280 73956 97336 74012
rect 97336 73956 97340 74012
rect 97276 73952 97340 73956
rect 4216 73468 4280 73472
rect 4216 73412 4220 73468
rect 4220 73412 4276 73468
rect 4276 73412 4280 73468
rect 4216 73408 4280 73412
rect 4296 73468 4360 73472
rect 4296 73412 4300 73468
rect 4300 73412 4356 73468
rect 4356 73412 4360 73468
rect 4296 73408 4360 73412
rect 4376 73468 4440 73472
rect 4376 73412 4380 73468
rect 4380 73412 4436 73468
rect 4436 73412 4440 73468
rect 4376 73408 4440 73412
rect 4456 73468 4520 73472
rect 4456 73412 4460 73468
rect 4460 73412 4516 73468
rect 4516 73412 4520 73468
rect 4456 73408 4520 73412
rect 96376 73468 96440 73472
rect 96376 73412 96380 73468
rect 96380 73412 96436 73468
rect 96436 73412 96440 73468
rect 96376 73408 96440 73412
rect 96456 73468 96520 73472
rect 96456 73412 96460 73468
rect 96460 73412 96516 73468
rect 96516 73412 96520 73468
rect 96456 73408 96520 73412
rect 96536 73468 96600 73472
rect 96536 73412 96540 73468
rect 96540 73412 96596 73468
rect 96596 73412 96600 73468
rect 96536 73408 96600 73412
rect 96616 73468 96680 73472
rect 96616 73412 96620 73468
rect 96620 73412 96676 73468
rect 96676 73412 96680 73468
rect 96616 73408 96680 73412
rect 4876 72924 4940 72928
rect 4876 72868 4880 72924
rect 4880 72868 4936 72924
rect 4936 72868 4940 72924
rect 4876 72864 4940 72868
rect 4956 72924 5020 72928
rect 4956 72868 4960 72924
rect 4960 72868 5016 72924
rect 5016 72868 5020 72924
rect 4956 72864 5020 72868
rect 5036 72924 5100 72928
rect 5036 72868 5040 72924
rect 5040 72868 5096 72924
rect 5096 72868 5100 72924
rect 5036 72864 5100 72868
rect 5116 72924 5180 72928
rect 5116 72868 5120 72924
rect 5120 72868 5176 72924
rect 5176 72868 5180 72924
rect 5116 72864 5180 72868
rect 97036 72924 97100 72928
rect 97036 72868 97040 72924
rect 97040 72868 97096 72924
rect 97096 72868 97100 72924
rect 97036 72864 97100 72868
rect 97116 72924 97180 72928
rect 97116 72868 97120 72924
rect 97120 72868 97176 72924
rect 97176 72868 97180 72924
rect 97116 72864 97180 72868
rect 97196 72924 97260 72928
rect 97196 72868 97200 72924
rect 97200 72868 97256 72924
rect 97256 72868 97260 72924
rect 97196 72864 97260 72868
rect 97276 72924 97340 72928
rect 97276 72868 97280 72924
rect 97280 72868 97336 72924
rect 97336 72868 97340 72924
rect 97276 72864 97340 72868
rect 4216 72380 4280 72384
rect 4216 72324 4220 72380
rect 4220 72324 4276 72380
rect 4276 72324 4280 72380
rect 4216 72320 4280 72324
rect 4296 72380 4360 72384
rect 4296 72324 4300 72380
rect 4300 72324 4356 72380
rect 4356 72324 4360 72380
rect 4296 72320 4360 72324
rect 4376 72380 4440 72384
rect 4376 72324 4380 72380
rect 4380 72324 4436 72380
rect 4436 72324 4440 72380
rect 4376 72320 4440 72324
rect 4456 72380 4520 72384
rect 4456 72324 4460 72380
rect 4460 72324 4516 72380
rect 4516 72324 4520 72380
rect 4456 72320 4520 72324
rect 96376 72380 96440 72384
rect 96376 72324 96380 72380
rect 96380 72324 96436 72380
rect 96436 72324 96440 72380
rect 96376 72320 96440 72324
rect 96456 72380 96520 72384
rect 96456 72324 96460 72380
rect 96460 72324 96516 72380
rect 96516 72324 96520 72380
rect 96456 72320 96520 72324
rect 96536 72380 96600 72384
rect 96536 72324 96540 72380
rect 96540 72324 96596 72380
rect 96596 72324 96600 72380
rect 96536 72320 96600 72324
rect 96616 72380 96680 72384
rect 96616 72324 96620 72380
rect 96620 72324 96676 72380
rect 96676 72324 96680 72380
rect 96616 72320 96680 72324
rect 4876 71836 4940 71840
rect 4876 71780 4880 71836
rect 4880 71780 4936 71836
rect 4936 71780 4940 71836
rect 4876 71776 4940 71780
rect 4956 71836 5020 71840
rect 4956 71780 4960 71836
rect 4960 71780 5016 71836
rect 5016 71780 5020 71836
rect 4956 71776 5020 71780
rect 5036 71836 5100 71840
rect 5036 71780 5040 71836
rect 5040 71780 5096 71836
rect 5096 71780 5100 71836
rect 5036 71776 5100 71780
rect 5116 71836 5180 71840
rect 5116 71780 5120 71836
rect 5120 71780 5176 71836
rect 5176 71780 5180 71836
rect 5116 71776 5180 71780
rect 97036 71836 97100 71840
rect 97036 71780 97040 71836
rect 97040 71780 97096 71836
rect 97096 71780 97100 71836
rect 97036 71776 97100 71780
rect 97116 71836 97180 71840
rect 97116 71780 97120 71836
rect 97120 71780 97176 71836
rect 97176 71780 97180 71836
rect 97116 71776 97180 71780
rect 97196 71836 97260 71840
rect 97196 71780 97200 71836
rect 97200 71780 97256 71836
rect 97256 71780 97260 71836
rect 97196 71776 97260 71780
rect 97276 71836 97340 71840
rect 97276 71780 97280 71836
rect 97280 71780 97336 71836
rect 97336 71780 97340 71836
rect 97276 71776 97340 71780
rect 4216 71292 4280 71296
rect 4216 71236 4220 71292
rect 4220 71236 4276 71292
rect 4276 71236 4280 71292
rect 4216 71232 4280 71236
rect 4296 71292 4360 71296
rect 4296 71236 4300 71292
rect 4300 71236 4356 71292
rect 4356 71236 4360 71292
rect 4296 71232 4360 71236
rect 4376 71292 4440 71296
rect 4376 71236 4380 71292
rect 4380 71236 4436 71292
rect 4436 71236 4440 71292
rect 4376 71232 4440 71236
rect 4456 71292 4520 71296
rect 4456 71236 4460 71292
rect 4460 71236 4516 71292
rect 4516 71236 4520 71292
rect 4456 71232 4520 71236
rect 96376 71292 96440 71296
rect 96376 71236 96380 71292
rect 96380 71236 96436 71292
rect 96436 71236 96440 71292
rect 96376 71232 96440 71236
rect 96456 71292 96520 71296
rect 96456 71236 96460 71292
rect 96460 71236 96516 71292
rect 96516 71236 96520 71292
rect 96456 71232 96520 71236
rect 96536 71292 96600 71296
rect 96536 71236 96540 71292
rect 96540 71236 96596 71292
rect 96596 71236 96600 71292
rect 96536 71232 96600 71236
rect 96616 71292 96680 71296
rect 96616 71236 96620 71292
rect 96620 71236 96676 71292
rect 96676 71236 96680 71292
rect 96616 71232 96680 71236
rect 4876 70748 4940 70752
rect 4876 70692 4880 70748
rect 4880 70692 4936 70748
rect 4936 70692 4940 70748
rect 4876 70688 4940 70692
rect 4956 70748 5020 70752
rect 4956 70692 4960 70748
rect 4960 70692 5016 70748
rect 5016 70692 5020 70748
rect 4956 70688 5020 70692
rect 5036 70748 5100 70752
rect 5036 70692 5040 70748
rect 5040 70692 5096 70748
rect 5096 70692 5100 70748
rect 5036 70688 5100 70692
rect 5116 70748 5180 70752
rect 5116 70692 5120 70748
rect 5120 70692 5176 70748
rect 5176 70692 5180 70748
rect 5116 70688 5180 70692
rect 97036 70748 97100 70752
rect 97036 70692 97040 70748
rect 97040 70692 97096 70748
rect 97096 70692 97100 70748
rect 97036 70688 97100 70692
rect 97116 70748 97180 70752
rect 97116 70692 97120 70748
rect 97120 70692 97176 70748
rect 97176 70692 97180 70748
rect 97116 70688 97180 70692
rect 97196 70748 97260 70752
rect 97196 70692 97200 70748
rect 97200 70692 97256 70748
rect 97256 70692 97260 70748
rect 97196 70688 97260 70692
rect 97276 70748 97340 70752
rect 97276 70692 97280 70748
rect 97280 70692 97336 70748
rect 97336 70692 97340 70748
rect 97276 70688 97340 70692
rect 4216 70204 4280 70208
rect 4216 70148 4220 70204
rect 4220 70148 4276 70204
rect 4276 70148 4280 70204
rect 4216 70144 4280 70148
rect 4296 70204 4360 70208
rect 4296 70148 4300 70204
rect 4300 70148 4356 70204
rect 4356 70148 4360 70204
rect 4296 70144 4360 70148
rect 4376 70204 4440 70208
rect 4376 70148 4380 70204
rect 4380 70148 4436 70204
rect 4436 70148 4440 70204
rect 4376 70144 4440 70148
rect 4456 70204 4520 70208
rect 4456 70148 4460 70204
rect 4460 70148 4516 70204
rect 4516 70148 4520 70204
rect 4456 70144 4520 70148
rect 96376 70204 96440 70208
rect 96376 70148 96380 70204
rect 96380 70148 96436 70204
rect 96436 70148 96440 70204
rect 96376 70144 96440 70148
rect 96456 70204 96520 70208
rect 96456 70148 96460 70204
rect 96460 70148 96516 70204
rect 96516 70148 96520 70204
rect 96456 70144 96520 70148
rect 96536 70204 96600 70208
rect 96536 70148 96540 70204
rect 96540 70148 96596 70204
rect 96596 70148 96600 70204
rect 96536 70144 96600 70148
rect 96616 70204 96680 70208
rect 96616 70148 96620 70204
rect 96620 70148 96676 70204
rect 96676 70148 96680 70204
rect 96616 70144 96680 70148
rect 4876 69660 4940 69664
rect 4876 69604 4880 69660
rect 4880 69604 4936 69660
rect 4936 69604 4940 69660
rect 4876 69600 4940 69604
rect 4956 69660 5020 69664
rect 4956 69604 4960 69660
rect 4960 69604 5016 69660
rect 5016 69604 5020 69660
rect 4956 69600 5020 69604
rect 5036 69660 5100 69664
rect 5036 69604 5040 69660
rect 5040 69604 5096 69660
rect 5096 69604 5100 69660
rect 5036 69600 5100 69604
rect 5116 69660 5180 69664
rect 5116 69604 5120 69660
rect 5120 69604 5176 69660
rect 5176 69604 5180 69660
rect 5116 69600 5180 69604
rect 97036 69660 97100 69664
rect 97036 69604 97040 69660
rect 97040 69604 97096 69660
rect 97096 69604 97100 69660
rect 97036 69600 97100 69604
rect 97116 69660 97180 69664
rect 97116 69604 97120 69660
rect 97120 69604 97176 69660
rect 97176 69604 97180 69660
rect 97116 69600 97180 69604
rect 97196 69660 97260 69664
rect 97196 69604 97200 69660
rect 97200 69604 97256 69660
rect 97256 69604 97260 69660
rect 97196 69600 97260 69604
rect 97276 69660 97340 69664
rect 97276 69604 97280 69660
rect 97280 69604 97336 69660
rect 97336 69604 97340 69660
rect 97276 69600 97340 69604
rect 4216 69116 4280 69120
rect 4216 69060 4220 69116
rect 4220 69060 4276 69116
rect 4276 69060 4280 69116
rect 4216 69056 4280 69060
rect 4296 69116 4360 69120
rect 4296 69060 4300 69116
rect 4300 69060 4356 69116
rect 4356 69060 4360 69116
rect 4296 69056 4360 69060
rect 4376 69116 4440 69120
rect 4376 69060 4380 69116
rect 4380 69060 4436 69116
rect 4436 69060 4440 69116
rect 4376 69056 4440 69060
rect 4456 69116 4520 69120
rect 4456 69060 4460 69116
rect 4460 69060 4516 69116
rect 4516 69060 4520 69116
rect 4456 69056 4520 69060
rect 96376 69116 96440 69120
rect 96376 69060 96380 69116
rect 96380 69060 96436 69116
rect 96436 69060 96440 69116
rect 96376 69056 96440 69060
rect 96456 69116 96520 69120
rect 96456 69060 96460 69116
rect 96460 69060 96516 69116
rect 96516 69060 96520 69116
rect 96456 69056 96520 69060
rect 96536 69116 96600 69120
rect 96536 69060 96540 69116
rect 96540 69060 96596 69116
rect 96596 69060 96600 69116
rect 96536 69056 96600 69060
rect 96616 69116 96680 69120
rect 96616 69060 96620 69116
rect 96620 69060 96676 69116
rect 96676 69060 96680 69116
rect 96616 69056 96680 69060
rect 4876 68572 4940 68576
rect 4876 68516 4880 68572
rect 4880 68516 4936 68572
rect 4936 68516 4940 68572
rect 4876 68512 4940 68516
rect 4956 68572 5020 68576
rect 4956 68516 4960 68572
rect 4960 68516 5016 68572
rect 5016 68516 5020 68572
rect 4956 68512 5020 68516
rect 5036 68572 5100 68576
rect 5036 68516 5040 68572
rect 5040 68516 5096 68572
rect 5096 68516 5100 68572
rect 5036 68512 5100 68516
rect 5116 68572 5180 68576
rect 5116 68516 5120 68572
rect 5120 68516 5176 68572
rect 5176 68516 5180 68572
rect 5116 68512 5180 68516
rect 97036 68572 97100 68576
rect 97036 68516 97040 68572
rect 97040 68516 97096 68572
rect 97096 68516 97100 68572
rect 97036 68512 97100 68516
rect 97116 68572 97180 68576
rect 97116 68516 97120 68572
rect 97120 68516 97176 68572
rect 97176 68516 97180 68572
rect 97116 68512 97180 68516
rect 97196 68572 97260 68576
rect 97196 68516 97200 68572
rect 97200 68516 97256 68572
rect 97256 68516 97260 68572
rect 97196 68512 97260 68516
rect 97276 68572 97340 68576
rect 97276 68516 97280 68572
rect 97280 68516 97336 68572
rect 97336 68516 97340 68572
rect 97276 68512 97340 68516
rect 4216 68028 4280 68032
rect 4216 67972 4220 68028
rect 4220 67972 4276 68028
rect 4276 67972 4280 68028
rect 4216 67968 4280 67972
rect 4296 68028 4360 68032
rect 4296 67972 4300 68028
rect 4300 67972 4356 68028
rect 4356 67972 4360 68028
rect 4296 67968 4360 67972
rect 4376 68028 4440 68032
rect 4376 67972 4380 68028
rect 4380 67972 4436 68028
rect 4436 67972 4440 68028
rect 4376 67968 4440 67972
rect 4456 68028 4520 68032
rect 4456 67972 4460 68028
rect 4460 67972 4516 68028
rect 4516 67972 4520 68028
rect 4456 67968 4520 67972
rect 96376 68028 96440 68032
rect 96376 67972 96380 68028
rect 96380 67972 96436 68028
rect 96436 67972 96440 68028
rect 96376 67968 96440 67972
rect 96456 68028 96520 68032
rect 96456 67972 96460 68028
rect 96460 67972 96516 68028
rect 96516 67972 96520 68028
rect 96456 67968 96520 67972
rect 96536 68028 96600 68032
rect 96536 67972 96540 68028
rect 96540 67972 96596 68028
rect 96596 67972 96600 68028
rect 96536 67968 96600 67972
rect 96616 68028 96680 68032
rect 96616 67972 96620 68028
rect 96620 67972 96676 68028
rect 96676 67972 96680 68028
rect 96616 67968 96680 67972
rect 4876 67484 4940 67488
rect 4876 67428 4880 67484
rect 4880 67428 4936 67484
rect 4936 67428 4940 67484
rect 4876 67424 4940 67428
rect 4956 67484 5020 67488
rect 4956 67428 4960 67484
rect 4960 67428 5016 67484
rect 5016 67428 5020 67484
rect 4956 67424 5020 67428
rect 5036 67484 5100 67488
rect 5036 67428 5040 67484
rect 5040 67428 5096 67484
rect 5096 67428 5100 67484
rect 5036 67424 5100 67428
rect 5116 67484 5180 67488
rect 5116 67428 5120 67484
rect 5120 67428 5176 67484
rect 5176 67428 5180 67484
rect 5116 67424 5180 67428
rect 97036 67484 97100 67488
rect 97036 67428 97040 67484
rect 97040 67428 97096 67484
rect 97096 67428 97100 67484
rect 97036 67424 97100 67428
rect 97116 67484 97180 67488
rect 97116 67428 97120 67484
rect 97120 67428 97176 67484
rect 97176 67428 97180 67484
rect 97116 67424 97180 67428
rect 97196 67484 97260 67488
rect 97196 67428 97200 67484
rect 97200 67428 97256 67484
rect 97256 67428 97260 67484
rect 97196 67424 97260 67428
rect 97276 67484 97340 67488
rect 97276 67428 97280 67484
rect 97280 67428 97336 67484
rect 97336 67428 97340 67484
rect 97276 67424 97340 67428
rect 4216 66940 4280 66944
rect 4216 66884 4220 66940
rect 4220 66884 4276 66940
rect 4276 66884 4280 66940
rect 4216 66880 4280 66884
rect 4296 66940 4360 66944
rect 4296 66884 4300 66940
rect 4300 66884 4356 66940
rect 4356 66884 4360 66940
rect 4296 66880 4360 66884
rect 4376 66940 4440 66944
rect 4376 66884 4380 66940
rect 4380 66884 4436 66940
rect 4436 66884 4440 66940
rect 4376 66880 4440 66884
rect 4456 66940 4520 66944
rect 4456 66884 4460 66940
rect 4460 66884 4516 66940
rect 4516 66884 4520 66940
rect 4456 66880 4520 66884
rect 96376 66940 96440 66944
rect 96376 66884 96380 66940
rect 96380 66884 96436 66940
rect 96436 66884 96440 66940
rect 96376 66880 96440 66884
rect 96456 66940 96520 66944
rect 96456 66884 96460 66940
rect 96460 66884 96516 66940
rect 96516 66884 96520 66940
rect 96456 66880 96520 66884
rect 96536 66940 96600 66944
rect 96536 66884 96540 66940
rect 96540 66884 96596 66940
rect 96596 66884 96600 66940
rect 96536 66880 96600 66884
rect 96616 66940 96680 66944
rect 96616 66884 96620 66940
rect 96620 66884 96676 66940
rect 96676 66884 96680 66940
rect 96616 66880 96680 66884
rect 4876 66396 4940 66400
rect 4876 66340 4880 66396
rect 4880 66340 4936 66396
rect 4936 66340 4940 66396
rect 4876 66336 4940 66340
rect 4956 66396 5020 66400
rect 4956 66340 4960 66396
rect 4960 66340 5016 66396
rect 5016 66340 5020 66396
rect 4956 66336 5020 66340
rect 5036 66396 5100 66400
rect 5036 66340 5040 66396
rect 5040 66340 5096 66396
rect 5096 66340 5100 66396
rect 5036 66336 5100 66340
rect 5116 66396 5180 66400
rect 5116 66340 5120 66396
rect 5120 66340 5176 66396
rect 5176 66340 5180 66396
rect 5116 66336 5180 66340
rect 97036 66396 97100 66400
rect 97036 66340 97040 66396
rect 97040 66340 97096 66396
rect 97096 66340 97100 66396
rect 97036 66336 97100 66340
rect 97116 66396 97180 66400
rect 97116 66340 97120 66396
rect 97120 66340 97176 66396
rect 97176 66340 97180 66396
rect 97116 66336 97180 66340
rect 97196 66396 97260 66400
rect 97196 66340 97200 66396
rect 97200 66340 97256 66396
rect 97256 66340 97260 66396
rect 97196 66336 97260 66340
rect 97276 66396 97340 66400
rect 97276 66340 97280 66396
rect 97280 66340 97336 66396
rect 97336 66340 97340 66396
rect 97276 66336 97340 66340
rect 4216 65852 4280 65856
rect 4216 65796 4220 65852
rect 4220 65796 4276 65852
rect 4276 65796 4280 65852
rect 4216 65792 4280 65796
rect 4296 65852 4360 65856
rect 4296 65796 4300 65852
rect 4300 65796 4356 65852
rect 4356 65796 4360 65852
rect 4296 65792 4360 65796
rect 4376 65852 4440 65856
rect 4376 65796 4380 65852
rect 4380 65796 4436 65852
rect 4436 65796 4440 65852
rect 4376 65792 4440 65796
rect 4456 65852 4520 65856
rect 4456 65796 4460 65852
rect 4460 65796 4516 65852
rect 4516 65796 4520 65852
rect 4456 65792 4520 65796
rect 96376 65852 96440 65856
rect 96376 65796 96380 65852
rect 96380 65796 96436 65852
rect 96436 65796 96440 65852
rect 96376 65792 96440 65796
rect 96456 65852 96520 65856
rect 96456 65796 96460 65852
rect 96460 65796 96516 65852
rect 96516 65796 96520 65852
rect 96456 65792 96520 65796
rect 96536 65852 96600 65856
rect 96536 65796 96540 65852
rect 96540 65796 96596 65852
rect 96596 65796 96600 65852
rect 96536 65792 96600 65796
rect 96616 65852 96680 65856
rect 96616 65796 96620 65852
rect 96620 65796 96676 65852
rect 96676 65796 96680 65852
rect 96616 65792 96680 65796
rect 4876 65308 4940 65312
rect 4876 65252 4880 65308
rect 4880 65252 4936 65308
rect 4936 65252 4940 65308
rect 4876 65248 4940 65252
rect 4956 65308 5020 65312
rect 4956 65252 4960 65308
rect 4960 65252 5016 65308
rect 5016 65252 5020 65308
rect 4956 65248 5020 65252
rect 5036 65308 5100 65312
rect 5036 65252 5040 65308
rect 5040 65252 5096 65308
rect 5096 65252 5100 65308
rect 5036 65248 5100 65252
rect 5116 65308 5180 65312
rect 5116 65252 5120 65308
rect 5120 65252 5176 65308
rect 5176 65252 5180 65308
rect 5116 65248 5180 65252
rect 97036 65308 97100 65312
rect 97036 65252 97040 65308
rect 97040 65252 97096 65308
rect 97096 65252 97100 65308
rect 97036 65248 97100 65252
rect 97116 65308 97180 65312
rect 97116 65252 97120 65308
rect 97120 65252 97176 65308
rect 97176 65252 97180 65308
rect 97116 65248 97180 65252
rect 97196 65308 97260 65312
rect 97196 65252 97200 65308
rect 97200 65252 97256 65308
rect 97256 65252 97260 65308
rect 97196 65248 97260 65252
rect 97276 65308 97340 65312
rect 97276 65252 97280 65308
rect 97280 65252 97336 65308
rect 97336 65252 97340 65308
rect 97276 65248 97340 65252
rect 4216 64764 4280 64768
rect 4216 64708 4220 64764
rect 4220 64708 4276 64764
rect 4276 64708 4280 64764
rect 4216 64704 4280 64708
rect 4296 64764 4360 64768
rect 4296 64708 4300 64764
rect 4300 64708 4356 64764
rect 4356 64708 4360 64764
rect 4296 64704 4360 64708
rect 4376 64764 4440 64768
rect 4376 64708 4380 64764
rect 4380 64708 4436 64764
rect 4436 64708 4440 64764
rect 4376 64704 4440 64708
rect 4456 64764 4520 64768
rect 4456 64708 4460 64764
rect 4460 64708 4516 64764
rect 4516 64708 4520 64764
rect 4456 64704 4520 64708
rect 96376 64764 96440 64768
rect 96376 64708 96380 64764
rect 96380 64708 96436 64764
rect 96436 64708 96440 64764
rect 96376 64704 96440 64708
rect 96456 64764 96520 64768
rect 96456 64708 96460 64764
rect 96460 64708 96516 64764
rect 96516 64708 96520 64764
rect 96456 64704 96520 64708
rect 96536 64764 96600 64768
rect 96536 64708 96540 64764
rect 96540 64708 96596 64764
rect 96596 64708 96600 64764
rect 96536 64704 96600 64708
rect 96616 64764 96680 64768
rect 96616 64708 96620 64764
rect 96620 64708 96676 64764
rect 96676 64708 96680 64764
rect 96616 64704 96680 64708
rect 4876 64220 4940 64224
rect 4876 64164 4880 64220
rect 4880 64164 4936 64220
rect 4936 64164 4940 64220
rect 4876 64160 4940 64164
rect 4956 64220 5020 64224
rect 4956 64164 4960 64220
rect 4960 64164 5016 64220
rect 5016 64164 5020 64220
rect 4956 64160 5020 64164
rect 5036 64220 5100 64224
rect 5036 64164 5040 64220
rect 5040 64164 5096 64220
rect 5096 64164 5100 64220
rect 5036 64160 5100 64164
rect 5116 64220 5180 64224
rect 5116 64164 5120 64220
rect 5120 64164 5176 64220
rect 5176 64164 5180 64220
rect 5116 64160 5180 64164
rect 97036 64220 97100 64224
rect 97036 64164 97040 64220
rect 97040 64164 97096 64220
rect 97096 64164 97100 64220
rect 97036 64160 97100 64164
rect 97116 64220 97180 64224
rect 97116 64164 97120 64220
rect 97120 64164 97176 64220
rect 97176 64164 97180 64220
rect 97116 64160 97180 64164
rect 97196 64220 97260 64224
rect 97196 64164 97200 64220
rect 97200 64164 97256 64220
rect 97256 64164 97260 64220
rect 97196 64160 97260 64164
rect 97276 64220 97340 64224
rect 97276 64164 97280 64220
rect 97280 64164 97336 64220
rect 97336 64164 97340 64220
rect 97276 64160 97340 64164
rect 4216 63676 4280 63680
rect 4216 63620 4220 63676
rect 4220 63620 4276 63676
rect 4276 63620 4280 63676
rect 4216 63616 4280 63620
rect 4296 63676 4360 63680
rect 4296 63620 4300 63676
rect 4300 63620 4356 63676
rect 4356 63620 4360 63676
rect 4296 63616 4360 63620
rect 4376 63676 4440 63680
rect 4376 63620 4380 63676
rect 4380 63620 4436 63676
rect 4436 63620 4440 63676
rect 4376 63616 4440 63620
rect 4456 63676 4520 63680
rect 4456 63620 4460 63676
rect 4460 63620 4516 63676
rect 4516 63620 4520 63676
rect 4456 63616 4520 63620
rect 96376 63676 96440 63680
rect 96376 63620 96380 63676
rect 96380 63620 96436 63676
rect 96436 63620 96440 63676
rect 96376 63616 96440 63620
rect 96456 63676 96520 63680
rect 96456 63620 96460 63676
rect 96460 63620 96516 63676
rect 96516 63620 96520 63676
rect 96456 63616 96520 63620
rect 96536 63676 96600 63680
rect 96536 63620 96540 63676
rect 96540 63620 96596 63676
rect 96596 63620 96600 63676
rect 96536 63616 96600 63620
rect 96616 63676 96680 63680
rect 96616 63620 96620 63676
rect 96620 63620 96676 63676
rect 96676 63620 96680 63676
rect 96616 63616 96680 63620
rect 4876 63132 4940 63136
rect 4876 63076 4880 63132
rect 4880 63076 4936 63132
rect 4936 63076 4940 63132
rect 4876 63072 4940 63076
rect 4956 63132 5020 63136
rect 4956 63076 4960 63132
rect 4960 63076 5016 63132
rect 5016 63076 5020 63132
rect 4956 63072 5020 63076
rect 5036 63132 5100 63136
rect 5036 63076 5040 63132
rect 5040 63076 5096 63132
rect 5096 63076 5100 63132
rect 5036 63072 5100 63076
rect 5116 63132 5180 63136
rect 5116 63076 5120 63132
rect 5120 63076 5176 63132
rect 5176 63076 5180 63132
rect 5116 63072 5180 63076
rect 97036 63132 97100 63136
rect 97036 63076 97040 63132
rect 97040 63076 97096 63132
rect 97096 63076 97100 63132
rect 97036 63072 97100 63076
rect 97116 63132 97180 63136
rect 97116 63076 97120 63132
rect 97120 63076 97176 63132
rect 97176 63076 97180 63132
rect 97116 63072 97180 63076
rect 97196 63132 97260 63136
rect 97196 63076 97200 63132
rect 97200 63076 97256 63132
rect 97256 63076 97260 63132
rect 97196 63072 97260 63076
rect 97276 63132 97340 63136
rect 97276 63076 97280 63132
rect 97280 63076 97336 63132
rect 97336 63076 97340 63132
rect 97276 63072 97340 63076
rect 4216 62588 4280 62592
rect 4216 62532 4220 62588
rect 4220 62532 4276 62588
rect 4276 62532 4280 62588
rect 4216 62528 4280 62532
rect 4296 62588 4360 62592
rect 4296 62532 4300 62588
rect 4300 62532 4356 62588
rect 4356 62532 4360 62588
rect 4296 62528 4360 62532
rect 4376 62588 4440 62592
rect 4376 62532 4380 62588
rect 4380 62532 4436 62588
rect 4436 62532 4440 62588
rect 4376 62528 4440 62532
rect 4456 62588 4520 62592
rect 4456 62532 4460 62588
rect 4460 62532 4516 62588
rect 4516 62532 4520 62588
rect 4456 62528 4520 62532
rect 96376 62588 96440 62592
rect 96376 62532 96380 62588
rect 96380 62532 96436 62588
rect 96436 62532 96440 62588
rect 96376 62528 96440 62532
rect 96456 62588 96520 62592
rect 96456 62532 96460 62588
rect 96460 62532 96516 62588
rect 96516 62532 96520 62588
rect 96456 62528 96520 62532
rect 96536 62588 96600 62592
rect 96536 62532 96540 62588
rect 96540 62532 96596 62588
rect 96596 62532 96600 62588
rect 96536 62528 96600 62532
rect 96616 62588 96680 62592
rect 96616 62532 96620 62588
rect 96620 62532 96676 62588
rect 96676 62532 96680 62588
rect 96616 62528 96680 62532
rect 4876 62044 4940 62048
rect 4876 61988 4880 62044
rect 4880 61988 4936 62044
rect 4936 61988 4940 62044
rect 4876 61984 4940 61988
rect 4956 62044 5020 62048
rect 4956 61988 4960 62044
rect 4960 61988 5016 62044
rect 5016 61988 5020 62044
rect 4956 61984 5020 61988
rect 5036 62044 5100 62048
rect 5036 61988 5040 62044
rect 5040 61988 5096 62044
rect 5096 61988 5100 62044
rect 5036 61984 5100 61988
rect 5116 62044 5180 62048
rect 5116 61988 5120 62044
rect 5120 61988 5176 62044
rect 5176 61988 5180 62044
rect 5116 61984 5180 61988
rect 97036 62044 97100 62048
rect 97036 61988 97040 62044
rect 97040 61988 97096 62044
rect 97096 61988 97100 62044
rect 97036 61984 97100 61988
rect 97116 62044 97180 62048
rect 97116 61988 97120 62044
rect 97120 61988 97176 62044
rect 97176 61988 97180 62044
rect 97116 61984 97180 61988
rect 97196 62044 97260 62048
rect 97196 61988 97200 62044
rect 97200 61988 97256 62044
rect 97256 61988 97260 62044
rect 97196 61984 97260 61988
rect 97276 62044 97340 62048
rect 97276 61988 97280 62044
rect 97280 61988 97336 62044
rect 97336 61988 97340 62044
rect 97276 61984 97340 61988
rect 4216 61500 4280 61504
rect 4216 61444 4220 61500
rect 4220 61444 4276 61500
rect 4276 61444 4280 61500
rect 4216 61440 4280 61444
rect 4296 61500 4360 61504
rect 4296 61444 4300 61500
rect 4300 61444 4356 61500
rect 4356 61444 4360 61500
rect 4296 61440 4360 61444
rect 4376 61500 4440 61504
rect 4376 61444 4380 61500
rect 4380 61444 4436 61500
rect 4436 61444 4440 61500
rect 4376 61440 4440 61444
rect 4456 61500 4520 61504
rect 4456 61444 4460 61500
rect 4460 61444 4516 61500
rect 4516 61444 4520 61500
rect 4456 61440 4520 61444
rect 96376 61500 96440 61504
rect 96376 61444 96380 61500
rect 96380 61444 96436 61500
rect 96436 61444 96440 61500
rect 96376 61440 96440 61444
rect 96456 61500 96520 61504
rect 96456 61444 96460 61500
rect 96460 61444 96516 61500
rect 96516 61444 96520 61500
rect 96456 61440 96520 61444
rect 96536 61500 96600 61504
rect 96536 61444 96540 61500
rect 96540 61444 96596 61500
rect 96596 61444 96600 61500
rect 96536 61440 96600 61444
rect 96616 61500 96680 61504
rect 96616 61444 96620 61500
rect 96620 61444 96676 61500
rect 96676 61444 96680 61500
rect 96616 61440 96680 61444
rect 4876 60956 4940 60960
rect 4876 60900 4880 60956
rect 4880 60900 4936 60956
rect 4936 60900 4940 60956
rect 4876 60896 4940 60900
rect 4956 60956 5020 60960
rect 4956 60900 4960 60956
rect 4960 60900 5016 60956
rect 5016 60900 5020 60956
rect 4956 60896 5020 60900
rect 5036 60956 5100 60960
rect 5036 60900 5040 60956
rect 5040 60900 5096 60956
rect 5096 60900 5100 60956
rect 5036 60896 5100 60900
rect 5116 60956 5180 60960
rect 5116 60900 5120 60956
rect 5120 60900 5176 60956
rect 5176 60900 5180 60956
rect 5116 60896 5180 60900
rect 97036 60956 97100 60960
rect 97036 60900 97040 60956
rect 97040 60900 97096 60956
rect 97096 60900 97100 60956
rect 97036 60896 97100 60900
rect 97116 60956 97180 60960
rect 97116 60900 97120 60956
rect 97120 60900 97176 60956
rect 97176 60900 97180 60956
rect 97116 60896 97180 60900
rect 97196 60956 97260 60960
rect 97196 60900 97200 60956
rect 97200 60900 97256 60956
rect 97256 60900 97260 60956
rect 97196 60896 97260 60900
rect 97276 60956 97340 60960
rect 97276 60900 97280 60956
rect 97280 60900 97336 60956
rect 97336 60900 97340 60956
rect 97276 60896 97340 60900
rect 4216 60412 4280 60416
rect 4216 60356 4220 60412
rect 4220 60356 4276 60412
rect 4276 60356 4280 60412
rect 4216 60352 4280 60356
rect 4296 60412 4360 60416
rect 4296 60356 4300 60412
rect 4300 60356 4356 60412
rect 4356 60356 4360 60412
rect 4296 60352 4360 60356
rect 4376 60412 4440 60416
rect 4376 60356 4380 60412
rect 4380 60356 4436 60412
rect 4436 60356 4440 60412
rect 4376 60352 4440 60356
rect 4456 60412 4520 60416
rect 4456 60356 4460 60412
rect 4460 60356 4516 60412
rect 4516 60356 4520 60412
rect 4456 60352 4520 60356
rect 96376 60412 96440 60416
rect 96376 60356 96380 60412
rect 96380 60356 96436 60412
rect 96436 60356 96440 60412
rect 96376 60352 96440 60356
rect 96456 60412 96520 60416
rect 96456 60356 96460 60412
rect 96460 60356 96516 60412
rect 96516 60356 96520 60412
rect 96456 60352 96520 60356
rect 96536 60412 96600 60416
rect 96536 60356 96540 60412
rect 96540 60356 96596 60412
rect 96596 60356 96600 60412
rect 96536 60352 96600 60356
rect 96616 60412 96680 60416
rect 96616 60356 96620 60412
rect 96620 60356 96676 60412
rect 96676 60356 96680 60412
rect 96616 60352 96680 60356
rect 4876 59868 4940 59872
rect 4876 59812 4880 59868
rect 4880 59812 4936 59868
rect 4936 59812 4940 59868
rect 4876 59808 4940 59812
rect 4956 59868 5020 59872
rect 4956 59812 4960 59868
rect 4960 59812 5016 59868
rect 5016 59812 5020 59868
rect 4956 59808 5020 59812
rect 5036 59868 5100 59872
rect 5036 59812 5040 59868
rect 5040 59812 5096 59868
rect 5096 59812 5100 59868
rect 5036 59808 5100 59812
rect 5116 59868 5180 59872
rect 5116 59812 5120 59868
rect 5120 59812 5176 59868
rect 5176 59812 5180 59868
rect 5116 59808 5180 59812
rect 97036 59868 97100 59872
rect 97036 59812 97040 59868
rect 97040 59812 97096 59868
rect 97096 59812 97100 59868
rect 97036 59808 97100 59812
rect 97116 59868 97180 59872
rect 97116 59812 97120 59868
rect 97120 59812 97176 59868
rect 97176 59812 97180 59868
rect 97116 59808 97180 59812
rect 97196 59868 97260 59872
rect 97196 59812 97200 59868
rect 97200 59812 97256 59868
rect 97256 59812 97260 59868
rect 97196 59808 97260 59812
rect 97276 59868 97340 59872
rect 97276 59812 97280 59868
rect 97280 59812 97336 59868
rect 97336 59812 97340 59868
rect 97276 59808 97340 59812
rect 4216 59324 4280 59328
rect 4216 59268 4220 59324
rect 4220 59268 4276 59324
rect 4276 59268 4280 59324
rect 4216 59264 4280 59268
rect 4296 59324 4360 59328
rect 4296 59268 4300 59324
rect 4300 59268 4356 59324
rect 4356 59268 4360 59324
rect 4296 59264 4360 59268
rect 4376 59324 4440 59328
rect 4376 59268 4380 59324
rect 4380 59268 4436 59324
rect 4436 59268 4440 59324
rect 4376 59264 4440 59268
rect 4456 59324 4520 59328
rect 4456 59268 4460 59324
rect 4460 59268 4516 59324
rect 4516 59268 4520 59324
rect 4456 59264 4520 59268
rect 96376 59324 96440 59328
rect 96376 59268 96380 59324
rect 96380 59268 96436 59324
rect 96436 59268 96440 59324
rect 96376 59264 96440 59268
rect 96456 59324 96520 59328
rect 96456 59268 96460 59324
rect 96460 59268 96516 59324
rect 96516 59268 96520 59324
rect 96456 59264 96520 59268
rect 96536 59324 96600 59328
rect 96536 59268 96540 59324
rect 96540 59268 96596 59324
rect 96596 59268 96600 59324
rect 96536 59264 96600 59268
rect 96616 59324 96680 59328
rect 96616 59268 96620 59324
rect 96620 59268 96676 59324
rect 96676 59268 96680 59324
rect 96616 59264 96680 59268
rect 4876 58780 4940 58784
rect 4876 58724 4880 58780
rect 4880 58724 4936 58780
rect 4936 58724 4940 58780
rect 4876 58720 4940 58724
rect 4956 58780 5020 58784
rect 4956 58724 4960 58780
rect 4960 58724 5016 58780
rect 5016 58724 5020 58780
rect 4956 58720 5020 58724
rect 5036 58780 5100 58784
rect 5036 58724 5040 58780
rect 5040 58724 5096 58780
rect 5096 58724 5100 58780
rect 5036 58720 5100 58724
rect 5116 58780 5180 58784
rect 5116 58724 5120 58780
rect 5120 58724 5176 58780
rect 5176 58724 5180 58780
rect 5116 58720 5180 58724
rect 97036 58780 97100 58784
rect 97036 58724 97040 58780
rect 97040 58724 97096 58780
rect 97096 58724 97100 58780
rect 97036 58720 97100 58724
rect 97116 58780 97180 58784
rect 97116 58724 97120 58780
rect 97120 58724 97176 58780
rect 97176 58724 97180 58780
rect 97116 58720 97180 58724
rect 97196 58780 97260 58784
rect 97196 58724 97200 58780
rect 97200 58724 97256 58780
rect 97256 58724 97260 58780
rect 97196 58720 97260 58724
rect 97276 58780 97340 58784
rect 97276 58724 97280 58780
rect 97280 58724 97336 58780
rect 97336 58724 97340 58780
rect 97276 58720 97340 58724
rect 4216 58236 4280 58240
rect 4216 58180 4220 58236
rect 4220 58180 4276 58236
rect 4276 58180 4280 58236
rect 4216 58176 4280 58180
rect 4296 58236 4360 58240
rect 4296 58180 4300 58236
rect 4300 58180 4356 58236
rect 4356 58180 4360 58236
rect 4296 58176 4360 58180
rect 4376 58236 4440 58240
rect 4376 58180 4380 58236
rect 4380 58180 4436 58236
rect 4436 58180 4440 58236
rect 4376 58176 4440 58180
rect 4456 58236 4520 58240
rect 4456 58180 4460 58236
rect 4460 58180 4516 58236
rect 4516 58180 4520 58236
rect 4456 58176 4520 58180
rect 96376 58236 96440 58240
rect 96376 58180 96380 58236
rect 96380 58180 96436 58236
rect 96436 58180 96440 58236
rect 96376 58176 96440 58180
rect 96456 58236 96520 58240
rect 96456 58180 96460 58236
rect 96460 58180 96516 58236
rect 96516 58180 96520 58236
rect 96456 58176 96520 58180
rect 96536 58236 96600 58240
rect 96536 58180 96540 58236
rect 96540 58180 96596 58236
rect 96596 58180 96600 58236
rect 96536 58176 96600 58180
rect 96616 58236 96680 58240
rect 96616 58180 96620 58236
rect 96620 58180 96676 58236
rect 96676 58180 96680 58236
rect 96616 58176 96680 58180
rect 4876 57692 4940 57696
rect 4876 57636 4880 57692
rect 4880 57636 4936 57692
rect 4936 57636 4940 57692
rect 4876 57632 4940 57636
rect 4956 57692 5020 57696
rect 4956 57636 4960 57692
rect 4960 57636 5016 57692
rect 5016 57636 5020 57692
rect 4956 57632 5020 57636
rect 5036 57692 5100 57696
rect 5036 57636 5040 57692
rect 5040 57636 5096 57692
rect 5096 57636 5100 57692
rect 5036 57632 5100 57636
rect 5116 57692 5180 57696
rect 5116 57636 5120 57692
rect 5120 57636 5176 57692
rect 5176 57636 5180 57692
rect 5116 57632 5180 57636
rect 97036 57692 97100 57696
rect 97036 57636 97040 57692
rect 97040 57636 97096 57692
rect 97096 57636 97100 57692
rect 97036 57632 97100 57636
rect 97116 57692 97180 57696
rect 97116 57636 97120 57692
rect 97120 57636 97176 57692
rect 97176 57636 97180 57692
rect 97116 57632 97180 57636
rect 97196 57692 97260 57696
rect 97196 57636 97200 57692
rect 97200 57636 97256 57692
rect 97256 57636 97260 57692
rect 97196 57632 97260 57636
rect 97276 57692 97340 57696
rect 97276 57636 97280 57692
rect 97280 57636 97336 57692
rect 97336 57636 97340 57692
rect 97276 57632 97340 57636
rect 4216 57148 4280 57152
rect 4216 57092 4220 57148
rect 4220 57092 4276 57148
rect 4276 57092 4280 57148
rect 4216 57088 4280 57092
rect 4296 57148 4360 57152
rect 4296 57092 4300 57148
rect 4300 57092 4356 57148
rect 4356 57092 4360 57148
rect 4296 57088 4360 57092
rect 4376 57148 4440 57152
rect 4376 57092 4380 57148
rect 4380 57092 4436 57148
rect 4436 57092 4440 57148
rect 4376 57088 4440 57092
rect 4456 57148 4520 57152
rect 4456 57092 4460 57148
rect 4460 57092 4516 57148
rect 4516 57092 4520 57148
rect 4456 57088 4520 57092
rect 96376 57148 96440 57152
rect 96376 57092 96380 57148
rect 96380 57092 96436 57148
rect 96436 57092 96440 57148
rect 96376 57088 96440 57092
rect 96456 57148 96520 57152
rect 96456 57092 96460 57148
rect 96460 57092 96516 57148
rect 96516 57092 96520 57148
rect 96456 57088 96520 57092
rect 96536 57148 96600 57152
rect 96536 57092 96540 57148
rect 96540 57092 96596 57148
rect 96596 57092 96600 57148
rect 96536 57088 96600 57092
rect 96616 57148 96680 57152
rect 96616 57092 96620 57148
rect 96620 57092 96676 57148
rect 96676 57092 96680 57148
rect 96616 57088 96680 57092
rect 4876 56604 4940 56608
rect 4876 56548 4880 56604
rect 4880 56548 4936 56604
rect 4936 56548 4940 56604
rect 4876 56544 4940 56548
rect 4956 56604 5020 56608
rect 4956 56548 4960 56604
rect 4960 56548 5016 56604
rect 5016 56548 5020 56604
rect 4956 56544 5020 56548
rect 5036 56604 5100 56608
rect 5036 56548 5040 56604
rect 5040 56548 5096 56604
rect 5096 56548 5100 56604
rect 5036 56544 5100 56548
rect 5116 56604 5180 56608
rect 5116 56548 5120 56604
rect 5120 56548 5176 56604
rect 5176 56548 5180 56604
rect 5116 56544 5180 56548
rect 97036 56604 97100 56608
rect 97036 56548 97040 56604
rect 97040 56548 97096 56604
rect 97096 56548 97100 56604
rect 97036 56544 97100 56548
rect 97116 56604 97180 56608
rect 97116 56548 97120 56604
rect 97120 56548 97176 56604
rect 97176 56548 97180 56604
rect 97116 56544 97180 56548
rect 97196 56604 97260 56608
rect 97196 56548 97200 56604
rect 97200 56548 97256 56604
rect 97256 56548 97260 56604
rect 97196 56544 97260 56548
rect 97276 56604 97340 56608
rect 97276 56548 97280 56604
rect 97280 56548 97336 56604
rect 97336 56548 97340 56604
rect 97276 56544 97340 56548
rect 4216 56060 4280 56064
rect 4216 56004 4220 56060
rect 4220 56004 4276 56060
rect 4276 56004 4280 56060
rect 4216 56000 4280 56004
rect 4296 56060 4360 56064
rect 4296 56004 4300 56060
rect 4300 56004 4356 56060
rect 4356 56004 4360 56060
rect 4296 56000 4360 56004
rect 4376 56060 4440 56064
rect 4376 56004 4380 56060
rect 4380 56004 4436 56060
rect 4436 56004 4440 56060
rect 4376 56000 4440 56004
rect 4456 56060 4520 56064
rect 4456 56004 4460 56060
rect 4460 56004 4516 56060
rect 4516 56004 4520 56060
rect 4456 56000 4520 56004
rect 96376 56060 96440 56064
rect 96376 56004 96380 56060
rect 96380 56004 96436 56060
rect 96436 56004 96440 56060
rect 96376 56000 96440 56004
rect 96456 56060 96520 56064
rect 96456 56004 96460 56060
rect 96460 56004 96516 56060
rect 96516 56004 96520 56060
rect 96456 56000 96520 56004
rect 96536 56060 96600 56064
rect 96536 56004 96540 56060
rect 96540 56004 96596 56060
rect 96596 56004 96600 56060
rect 96536 56000 96600 56004
rect 96616 56060 96680 56064
rect 96616 56004 96620 56060
rect 96620 56004 96676 56060
rect 96676 56004 96680 56060
rect 96616 56000 96680 56004
rect 4876 55516 4940 55520
rect 4876 55460 4880 55516
rect 4880 55460 4936 55516
rect 4936 55460 4940 55516
rect 4876 55456 4940 55460
rect 4956 55516 5020 55520
rect 4956 55460 4960 55516
rect 4960 55460 5016 55516
rect 5016 55460 5020 55516
rect 4956 55456 5020 55460
rect 5036 55516 5100 55520
rect 5036 55460 5040 55516
rect 5040 55460 5096 55516
rect 5096 55460 5100 55516
rect 5036 55456 5100 55460
rect 5116 55516 5180 55520
rect 5116 55460 5120 55516
rect 5120 55460 5176 55516
rect 5176 55460 5180 55516
rect 5116 55456 5180 55460
rect 97036 55516 97100 55520
rect 97036 55460 97040 55516
rect 97040 55460 97096 55516
rect 97096 55460 97100 55516
rect 97036 55456 97100 55460
rect 97116 55516 97180 55520
rect 97116 55460 97120 55516
rect 97120 55460 97176 55516
rect 97176 55460 97180 55516
rect 97116 55456 97180 55460
rect 97196 55516 97260 55520
rect 97196 55460 97200 55516
rect 97200 55460 97256 55516
rect 97256 55460 97260 55516
rect 97196 55456 97260 55460
rect 97276 55516 97340 55520
rect 97276 55460 97280 55516
rect 97280 55460 97336 55516
rect 97336 55460 97340 55516
rect 97276 55456 97340 55460
rect 4216 54972 4280 54976
rect 4216 54916 4220 54972
rect 4220 54916 4276 54972
rect 4276 54916 4280 54972
rect 4216 54912 4280 54916
rect 4296 54972 4360 54976
rect 4296 54916 4300 54972
rect 4300 54916 4356 54972
rect 4356 54916 4360 54972
rect 4296 54912 4360 54916
rect 4376 54972 4440 54976
rect 4376 54916 4380 54972
rect 4380 54916 4436 54972
rect 4436 54916 4440 54972
rect 4376 54912 4440 54916
rect 4456 54972 4520 54976
rect 4456 54916 4460 54972
rect 4460 54916 4516 54972
rect 4516 54916 4520 54972
rect 4456 54912 4520 54916
rect 96376 54972 96440 54976
rect 96376 54916 96380 54972
rect 96380 54916 96436 54972
rect 96436 54916 96440 54972
rect 96376 54912 96440 54916
rect 96456 54972 96520 54976
rect 96456 54916 96460 54972
rect 96460 54916 96516 54972
rect 96516 54916 96520 54972
rect 96456 54912 96520 54916
rect 96536 54972 96600 54976
rect 96536 54916 96540 54972
rect 96540 54916 96596 54972
rect 96596 54916 96600 54972
rect 96536 54912 96600 54916
rect 96616 54972 96680 54976
rect 96616 54916 96620 54972
rect 96620 54916 96676 54972
rect 96676 54916 96680 54972
rect 96616 54912 96680 54916
rect 4876 54428 4940 54432
rect 4876 54372 4880 54428
rect 4880 54372 4936 54428
rect 4936 54372 4940 54428
rect 4876 54368 4940 54372
rect 4956 54428 5020 54432
rect 4956 54372 4960 54428
rect 4960 54372 5016 54428
rect 5016 54372 5020 54428
rect 4956 54368 5020 54372
rect 5036 54428 5100 54432
rect 5036 54372 5040 54428
rect 5040 54372 5096 54428
rect 5096 54372 5100 54428
rect 5036 54368 5100 54372
rect 5116 54428 5180 54432
rect 5116 54372 5120 54428
rect 5120 54372 5176 54428
rect 5176 54372 5180 54428
rect 5116 54368 5180 54372
rect 97036 54428 97100 54432
rect 97036 54372 97040 54428
rect 97040 54372 97096 54428
rect 97096 54372 97100 54428
rect 97036 54368 97100 54372
rect 97116 54428 97180 54432
rect 97116 54372 97120 54428
rect 97120 54372 97176 54428
rect 97176 54372 97180 54428
rect 97116 54368 97180 54372
rect 97196 54428 97260 54432
rect 97196 54372 97200 54428
rect 97200 54372 97256 54428
rect 97256 54372 97260 54428
rect 97196 54368 97260 54372
rect 97276 54428 97340 54432
rect 97276 54372 97280 54428
rect 97280 54372 97336 54428
rect 97336 54372 97340 54428
rect 97276 54368 97340 54372
rect 4216 53884 4280 53888
rect 4216 53828 4220 53884
rect 4220 53828 4276 53884
rect 4276 53828 4280 53884
rect 4216 53824 4280 53828
rect 4296 53884 4360 53888
rect 4296 53828 4300 53884
rect 4300 53828 4356 53884
rect 4356 53828 4360 53884
rect 4296 53824 4360 53828
rect 4376 53884 4440 53888
rect 4376 53828 4380 53884
rect 4380 53828 4436 53884
rect 4436 53828 4440 53884
rect 4376 53824 4440 53828
rect 4456 53884 4520 53888
rect 4456 53828 4460 53884
rect 4460 53828 4516 53884
rect 4516 53828 4520 53884
rect 4456 53824 4520 53828
rect 96376 53884 96440 53888
rect 96376 53828 96380 53884
rect 96380 53828 96436 53884
rect 96436 53828 96440 53884
rect 96376 53824 96440 53828
rect 96456 53884 96520 53888
rect 96456 53828 96460 53884
rect 96460 53828 96516 53884
rect 96516 53828 96520 53884
rect 96456 53824 96520 53828
rect 96536 53884 96600 53888
rect 96536 53828 96540 53884
rect 96540 53828 96596 53884
rect 96596 53828 96600 53884
rect 96536 53824 96600 53828
rect 96616 53884 96680 53888
rect 96616 53828 96620 53884
rect 96620 53828 96676 53884
rect 96676 53828 96680 53884
rect 96616 53824 96680 53828
rect 4876 53340 4940 53344
rect 4876 53284 4880 53340
rect 4880 53284 4936 53340
rect 4936 53284 4940 53340
rect 4876 53280 4940 53284
rect 4956 53340 5020 53344
rect 4956 53284 4960 53340
rect 4960 53284 5016 53340
rect 5016 53284 5020 53340
rect 4956 53280 5020 53284
rect 5036 53340 5100 53344
rect 5036 53284 5040 53340
rect 5040 53284 5096 53340
rect 5096 53284 5100 53340
rect 5036 53280 5100 53284
rect 5116 53340 5180 53344
rect 5116 53284 5120 53340
rect 5120 53284 5176 53340
rect 5176 53284 5180 53340
rect 5116 53280 5180 53284
rect 97036 53340 97100 53344
rect 97036 53284 97040 53340
rect 97040 53284 97096 53340
rect 97096 53284 97100 53340
rect 97036 53280 97100 53284
rect 97116 53340 97180 53344
rect 97116 53284 97120 53340
rect 97120 53284 97176 53340
rect 97176 53284 97180 53340
rect 97116 53280 97180 53284
rect 97196 53340 97260 53344
rect 97196 53284 97200 53340
rect 97200 53284 97256 53340
rect 97256 53284 97260 53340
rect 97196 53280 97260 53284
rect 97276 53340 97340 53344
rect 97276 53284 97280 53340
rect 97280 53284 97336 53340
rect 97336 53284 97340 53340
rect 97276 53280 97340 53284
rect 4216 52796 4280 52800
rect 4216 52740 4220 52796
rect 4220 52740 4276 52796
rect 4276 52740 4280 52796
rect 4216 52736 4280 52740
rect 4296 52796 4360 52800
rect 4296 52740 4300 52796
rect 4300 52740 4356 52796
rect 4356 52740 4360 52796
rect 4296 52736 4360 52740
rect 4376 52796 4440 52800
rect 4376 52740 4380 52796
rect 4380 52740 4436 52796
rect 4436 52740 4440 52796
rect 4376 52736 4440 52740
rect 4456 52796 4520 52800
rect 4456 52740 4460 52796
rect 4460 52740 4516 52796
rect 4516 52740 4520 52796
rect 4456 52736 4520 52740
rect 96376 52796 96440 52800
rect 96376 52740 96380 52796
rect 96380 52740 96436 52796
rect 96436 52740 96440 52796
rect 96376 52736 96440 52740
rect 96456 52796 96520 52800
rect 96456 52740 96460 52796
rect 96460 52740 96516 52796
rect 96516 52740 96520 52796
rect 96456 52736 96520 52740
rect 96536 52796 96600 52800
rect 96536 52740 96540 52796
rect 96540 52740 96596 52796
rect 96596 52740 96600 52796
rect 96536 52736 96600 52740
rect 96616 52796 96680 52800
rect 96616 52740 96620 52796
rect 96620 52740 96676 52796
rect 96676 52740 96680 52796
rect 96616 52736 96680 52740
rect 4876 52252 4940 52256
rect 4876 52196 4880 52252
rect 4880 52196 4936 52252
rect 4936 52196 4940 52252
rect 4876 52192 4940 52196
rect 4956 52252 5020 52256
rect 4956 52196 4960 52252
rect 4960 52196 5016 52252
rect 5016 52196 5020 52252
rect 4956 52192 5020 52196
rect 5036 52252 5100 52256
rect 5036 52196 5040 52252
rect 5040 52196 5096 52252
rect 5096 52196 5100 52252
rect 5036 52192 5100 52196
rect 5116 52252 5180 52256
rect 5116 52196 5120 52252
rect 5120 52196 5176 52252
rect 5176 52196 5180 52252
rect 5116 52192 5180 52196
rect 97036 52252 97100 52256
rect 97036 52196 97040 52252
rect 97040 52196 97096 52252
rect 97096 52196 97100 52252
rect 97036 52192 97100 52196
rect 97116 52252 97180 52256
rect 97116 52196 97120 52252
rect 97120 52196 97176 52252
rect 97176 52196 97180 52252
rect 97116 52192 97180 52196
rect 97196 52252 97260 52256
rect 97196 52196 97200 52252
rect 97200 52196 97256 52252
rect 97256 52196 97260 52252
rect 97196 52192 97260 52196
rect 97276 52252 97340 52256
rect 97276 52196 97280 52252
rect 97280 52196 97336 52252
rect 97336 52196 97340 52252
rect 97276 52192 97340 52196
rect 4216 51708 4280 51712
rect 4216 51652 4220 51708
rect 4220 51652 4276 51708
rect 4276 51652 4280 51708
rect 4216 51648 4280 51652
rect 4296 51708 4360 51712
rect 4296 51652 4300 51708
rect 4300 51652 4356 51708
rect 4356 51652 4360 51708
rect 4296 51648 4360 51652
rect 4376 51708 4440 51712
rect 4376 51652 4380 51708
rect 4380 51652 4436 51708
rect 4436 51652 4440 51708
rect 4376 51648 4440 51652
rect 4456 51708 4520 51712
rect 4456 51652 4460 51708
rect 4460 51652 4516 51708
rect 4516 51652 4520 51708
rect 4456 51648 4520 51652
rect 96376 51708 96440 51712
rect 96376 51652 96380 51708
rect 96380 51652 96436 51708
rect 96436 51652 96440 51708
rect 96376 51648 96440 51652
rect 96456 51708 96520 51712
rect 96456 51652 96460 51708
rect 96460 51652 96516 51708
rect 96516 51652 96520 51708
rect 96456 51648 96520 51652
rect 96536 51708 96600 51712
rect 96536 51652 96540 51708
rect 96540 51652 96596 51708
rect 96596 51652 96600 51708
rect 96536 51648 96600 51652
rect 96616 51708 96680 51712
rect 96616 51652 96620 51708
rect 96620 51652 96676 51708
rect 96676 51652 96680 51708
rect 96616 51648 96680 51652
rect 4876 51164 4940 51168
rect 4876 51108 4880 51164
rect 4880 51108 4936 51164
rect 4936 51108 4940 51164
rect 4876 51104 4940 51108
rect 4956 51164 5020 51168
rect 4956 51108 4960 51164
rect 4960 51108 5016 51164
rect 5016 51108 5020 51164
rect 4956 51104 5020 51108
rect 5036 51164 5100 51168
rect 5036 51108 5040 51164
rect 5040 51108 5096 51164
rect 5096 51108 5100 51164
rect 5036 51104 5100 51108
rect 5116 51164 5180 51168
rect 5116 51108 5120 51164
rect 5120 51108 5176 51164
rect 5176 51108 5180 51164
rect 5116 51104 5180 51108
rect 97036 51164 97100 51168
rect 97036 51108 97040 51164
rect 97040 51108 97096 51164
rect 97096 51108 97100 51164
rect 97036 51104 97100 51108
rect 97116 51164 97180 51168
rect 97116 51108 97120 51164
rect 97120 51108 97176 51164
rect 97176 51108 97180 51164
rect 97116 51104 97180 51108
rect 97196 51164 97260 51168
rect 97196 51108 97200 51164
rect 97200 51108 97256 51164
rect 97256 51108 97260 51164
rect 97196 51104 97260 51108
rect 97276 51164 97340 51168
rect 97276 51108 97280 51164
rect 97280 51108 97336 51164
rect 97336 51108 97340 51164
rect 97276 51104 97340 51108
rect 4216 50620 4280 50624
rect 4216 50564 4220 50620
rect 4220 50564 4276 50620
rect 4276 50564 4280 50620
rect 4216 50560 4280 50564
rect 4296 50620 4360 50624
rect 4296 50564 4300 50620
rect 4300 50564 4356 50620
rect 4356 50564 4360 50620
rect 4296 50560 4360 50564
rect 4376 50620 4440 50624
rect 4376 50564 4380 50620
rect 4380 50564 4436 50620
rect 4436 50564 4440 50620
rect 4376 50560 4440 50564
rect 4456 50620 4520 50624
rect 4456 50564 4460 50620
rect 4460 50564 4516 50620
rect 4516 50564 4520 50620
rect 4456 50560 4520 50564
rect 96376 50620 96440 50624
rect 96376 50564 96380 50620
rect 96380 50564 96436 50620
rect 96436 50564 96440 50620
rect 96376 50560 96440 50564
rect 96456 50620 96520 50624
rect 96456 50564 96460 50620
rect 96460 50564 96516 50620
rect 96516 50564 96520 50620
rect 96456 50560 96520 50564
rect 96536 50620 96600 50624
rect 96536 50564 96540 50620
rect 96540 50564 96596 50620
rect 96596 50564 96600 50620
rect 96536 50560 96600 50564
rect 96616 50620 96680 50624
rect 96616 50564 96620 50620
rect 96620 50564 96676 50620
rect 96676 50564 96680 50620
rect 96616 50560 96680 50564
rect 4876 50076 4940 50080
rect 4876 50020 4880 50076
rect 4880 50020 4936 50076
rect 4936 50020 4940 50076
rect 4876 50016 4940 50020
rect 4956 50076 5020 50080
rect 4956 50020 4960 50076
rect 4960 50020 5016 50076
rect 5016 50020 5020 50076
rect 4956 50016 5020 50020
rect 5036 50076 5100 50080
rect 5036 50020 5040 50076
rect 5040 50020 5096 50076
rect 5096 50020 5100 50076
rect 5036 50016 5100 50020
rect 5116 50076 5180 50080
rect 5116 50020 5120 50076
rect 5120 50020 5176 50076
rect 5176 50020 5180 50076
rect 5116 50016 5180 50020
rect 97036 50076 97100 50080
rect 97036 50020 97040 50076
rect 97040 50020 97096 50076
rect 97096 50020 97100 50076
rect 97036 50016 97100 50020
rect 97116 50076 97180 50080
rect 97116 50020 97120 50076
rect 97120 50020 97176 50076
rect 97176 50020 97180 50076
rect 97116 50016 97180 50020
rect 97196 50076 97260 50080
rect 97196 50020 97200 50076
rect 97200 50020 97256 50076
rect 97256 50020 97260 50076
rect 97196 50016 97260 50020
rect 97276 50076 97340 50080
rect 97276 50020 97280 50076
rect 97280 50020 97336 50076
rect 97336 50020 97340 50076
rect 97276 50016 97340 50020
rect 4216 49532 4280 49536
rect 4216 49476 4220 49532
rect 4220 49476 4276 49532
rect 4276 49476 4280 49532
rect 4216 49472 4280 49476
rect 4296 49532 4360 49536
rect 4296 49476 4300 49532
rect 4300 49476 4356 49532
rect 4356 49476 4360 49532
rect 4296 49472 4360 49476
rect 4376 49532 4440 49536
rect 4376 49476 4380 49532
rect 4380 49476 4436 49532
rect 4436 49476 4440 49532
rect 4376 49472 4440 49476
rect 4456 49532 4520 49536
rect 4456 49476 4460 49532
rect 4460 49476 4516 49532
rect 4516 49476 4520 49532
rect 4456 49472 4520 49476
rect 96376 49532 96440 49536
rect 96376 49476 96380 49532
rect 96380 49476 96436 49532
rect 96436 49476 96440 49532
rect 96376 49472 96440 49476
rect 96456 49532 96520 49536
rect 96456 49476 96460 49532
rect 96460 49476 96516 49532
rect 96516 49476 96520 49532
rect 96456 49472 96520 49476
rect 96536 49532 96600 49536
rect 96536 49476 96540 49532
rect 96540 49476 96596 49532
rect 96596 49476 96600 49532
rect 96536 49472 96600 49476
rect 96616 49532 96680 49536
rect 96616 49476 96620 49532
rect 96620 49476 96676 49532
rect 96676 49476 96680 49532
rect 96616 49472 96680 49476
rect 4876 48988 4940 48992
rect 4876 48932 4880 48988
rect 4880 48932 4936 48988
rect 4936 48932 4940 48988
rect 4876 48928 4940 48932
rect 4956 48988 5020 48992
rect 4956 48932 4960 48988
rect 4960 48932 5016 48988
rect 5016 48932 5020 48988
rect 4956 48928 5020 48932
rect 5036 48988 5100 48992
rect 5036 48932 5040 48988
rect 5040 48932 5096 48988
rect 5096 48932 5100 48988
rect 5036 48928 5100 48932
rect 5116 48988 5180 48992
rect 5116 48932 5120 48988
rect 5120 48932 5176 48988
rect 5176 48932 5180 48988
rect 5116 48928 5180 48932
rect 97036 48988 97100 48992
rect 97036 48932 97040 48988
rect 97040 48932 97096 48988
rect 97096 48932 97100 48988
rect 97036 48928 97100 48932
rect 97116 48988 97180 48992
rect 97116 48932 97120 48988
rect 97120 48932 97176 48988
rect 97176 48932 97180 48988
rect 97116 48928 97180 48932
rect 97196 48988 97260 48992
rect 97196 48932 97200 48988
rect 97200 48932 97256 48988
rect 97256 48932 97260 48988
rect 97196 48928 97260 48932
rect 97276 48988 97340 48992
rect 97276 48932 97280 48988
rect 97280 48932 97336 48988
rect 97336 48932 97340 48988
rect 97276 48928 97340 48932
rect 4216 48444 4280 48448
rect 4216 48388 4220 48444
rect 4220 48388 4276 48444
rect 4276 48388 4280 48444
rect 4216 48384 4280 48388
rect 4296 48444 4360 48448
rect 4296 48388 4300 48444
rect 4300 48388 4356 48444
rect 4356 48388 4360 48444
rect 4296 48384 4360 48388
rect 4376 48444 4440 48448
rect 4376 48388 4380 48444
rect 4380 48388 4436 48444
rect 4436 48388 4440 48444
rect 4376 48384 4440 48388
rect 4456 48444 4520 48448
rect 4456 48388 4460 48444
rect 4460 48388 4516 48444
rect 4516 48388 4520 48444
rect 4456 48384 4520 48388
rect 96376 48444 96440 48448
rect 96376 48388 96380 48444
rect 96380 48388 96436 48444
rect 96436 48388 96440 48444
rect 96376 48384 96440 48388
rect 96456 48444 96520 48448
rect 96456 48388 96460 48444
rect 96460 48388 96516 48444
rect 96516 48388 96520 48444
rect 96456 48384 96520 48388
rect 96536 48444 96600 48448
rect 96536 48388 96540 48444
rect 96540 48388 96596 48444
rect 96596 48388 96600 48444
rect 96536 48384 96600 48388
rect 96616 48444 96680 48448
rect 96616 48388 96620 48444
rect 96620 48388 96676 48444
rect 96676 48388 96680 48444
rect 96616 48384 96680 48388
rect 4876 47900 4940 47904
rect 4876 47844 4880 47900
rect 4880 47844 4936 47900
rect 4936 47844 4940 47900
rect 4876 47840 4940 47844
rect 4956 47900 5020 47904
rect 4956 47844 4960 47900
rect 4960 47844 5016 47900
rect 5016 47844 5020 47900
rect 4956 47840 5020 47844
rect 5036 47900 5100 47904
rect 5036 47844 5040 47900
rect 5040 47844 5096 47900
rect 5096 47844 5100 47900
rect 5036 47840 5100 47844
rect 5116 47900 5180 47904
rect 5116 47844 5120 47900
rect 5120 47844 5176 47900
rect 5176 47844 5180 47900
rect 5116 47840 5180 47844
rect 97036 47900 97100 47904
rect 97036 47844 97040 47900
rect 97040 47844 97096 47900
rect 97096 47844 97100 47900
rect 97036 47840 97100 47844
rect 97116 47900 97180 47904
rect 97116 47844 97120 47900
rect 97120 47844 97176 47900
rect 97176 47844 97180 47900
rect 97116 47840 97180 47844
rect 97196 47900 97260 47904
rect 97196 47844 97200 47900
rect 97200 47844 97256 47900
rect 97256 47844 97260 47900
rect 97196 47840 97260 47844
rect 97276 47900 97340 47904
rect 97276 47844 97280 47900
rect 97280 47844 97336 47900
rect 97336 47844 97340 47900
rect 97276 47840 97340 47844
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 96376 47356 96440 47360
rect 96376 47300 96380 47356
rect 96380 47300 96436 47356
rect 96436 47300 96440 47356
rect 96376 47296 96440 47300
rect 96456 47356 96520 47360
rect 96456 47300 96460 47356
rect 96460 47300 96516 47356
rect 96516 47300 96520 47356
rect 96456 47296 96520 47300
rect 96536 47356 96600 47360
rect 96536 47300 96540 47356
rect 96540 47300 96596 47356
rect 96596 47300 96600 47356
rect 96536 47296 96600 47300
rect 96616 47356 96680 47360
rect 96616 47300 96620 47356
rect 96620 47300 96676 47356
rect 96676 47300 96680 47356
rect 96616 47296 96680 47300
rect 4876 46812 4940 46816
rect 4876 46756 4880 46812
rect 4880 46756 4936 46812
rect 4936 46756 4940 46812
rect 4876 46752 4940 46756
rect 4956 46812 5020 46816
rect 4956 46756 4960 46812
rect 4960 46756 5016 46812
rect 5016 46756 5020 46812
rect 4956 46752 5020 46756
rect 5036 46812 5100 46816
rect 5036 46756 5040 46812
rect 5040 46756 5096 46812
rect 5096 46756 5100 46812
rect 5036 46752 5100 46756
rect 5116 46812 5180 46816
rect 5116 46756 5120 46812
rect 5120 46756 5176 46812
rect 5176 46756 5180 46812
rect 5116 46752 5180 46756
rect 97036 46812 97100 46816
rect 97036 46756 97040 46812
rect 97040 46756 97096 46812
rect 97096 46756 97100 46812
rect 97036 46752 97100 46756
rect 97116 46812 97180 46816
rect 97116 46756 97120 46812
rect 97120 46756 97176 46812
rect 97176 46756 97180 46812
rect 97116 46752 97180 46756
rect 97196 46812 97260 46816
rect 97196 46756 97200 46812
rect 97200 46756 97256 46812
rect 97256 46756 97260 46812
rect 97196 46752 97260 46756
rect 97276 46812 97340 46816
rect 97276 46756 97280 46812
rect 97280 46756 97336 46812
rect 97336 46756 97340 46812
rect 97276 46752 97340 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 96376 46268 96440 46272
rect 96376 46212 96380 46268
rect 96380 46212 96436 46268
rect 96436 46212 96440 46268
rect 96376 46208 96440 46212
rect 96456 46268 96520 46272
rect 96456 46212 96460 46268
rect 96460 46212 96516 46268
rect 96516 46212 96520 46268
rect 96456 46208 96520 46212
rect 96536 46268 96600 46272
rect 96536 46212 96540 46268
rect 96540 46212 96596 46268
rect 96596 46212 96600 46268
rect 96536 46208 96600 46212
rect 96616 46268 96680 46272
rect 96616 46212 96620 46268
rect 96620 46212 96676 46268
rect 96676 46212 96680 46268
rect 96616 46208 96680 46212
rect 4876 45724 4940 45728
rect 4876 45668 4880 45724
rect 4880 45668 4936 45724
rect 4936 45668 4940 45724
rect 4876 45664 4940 45668
rect 4956 45724 5020 45728
rect 4956 45668 4960 45724
rect 4960 45668 5016 45724
rect 5016 45668 5020 45724
rect 4956 45664 5020 45668
rect 5036 45724 5100 45728
rect 5036 45668 5040 45724
rect 5040 45668 5096 45724
rect 5096 45668 5100 45724
rect 5036 45664 5100 45668
rect 5116 45724 5180 45728
rect 5116 45668 5120 45724
rect 5120 45668 5176 45724
rect 5176 45668 5180 45724
rect 5116 45664 5180 45668
rect 97036 45724 97100 45728
rect 97036 45668 97040 45724
rect 97040 45668 97096 45724
rect 97096 45668 97100 45724
rect 97036 45664 97100 45668
rect 97116 45724 97180 45728
rect 97116 45668 97120 45724
rect 97120 45668 97176 45724
rect 97176 45668 97180 45724
rect 97116 45664 97180 45668
rect 97196 45724 97260 45728
rect 97196 45668 97200 45724
rect 97200 45668 97256 45724
rect 97256 45668 97260 45724
rect 97196 45664 97260 45668
rect 97276 45724 97340 45728
rect 97276 45668 97280 45724
rect 97280 45668 97336 45724
rect 97336 45668 97340 45724
rect 97276 45664 97340 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 96376 45180 96440 45184
rect 96376 45124 96380 45180
rect 96380 45124 96436 45180
rect 96436 45124 96440 45180
rect 96376 45120 96440 45124
rect 96456 45180 96520 45184
rect 96456 45124 96460 45180
rect 96460 45124 96516 45180
rect 96516 45124 96520 45180
rect 96456 45120 96520 45124
rect 96536 45180 96600 45184
rect 96536 45124 96540 45180
rect 96540 45124 96596 45180
rect 96596 45124 96600 45180
rect 96536 45120 96600 45124
rect 96616 45180 96680 45184
rect 96616 45124 96620 45180
rect 96620 45124 96676 45180
rect 96676 45124 96680 45180
rect 96616 45120 96680 45124
rect 4876 44636 4940 44640
rect 4876 44580 4880 44636
rect 4880 44580 4936 44636
rect 4936 44580 4940 44636
rect 4876 44576 4940 44580
rect 4956 44636 5020 44640
rect 4956 44580 4960 44636
rect 4960 44580 5016 44636
rect 5016 44580 5020 44636
rect 4956 44576 5020 44580
rect 5036 44636 5100 44640
rect 5036 44580 5040 44636
rect 5040 44580 5096 44636
rect 5096 44580 5100 44636
rect 5036 44576 5100 44580
rect 5116 44636 5180 44640
rect 5116 44580 5120 44636
rect 5120 44580 5176 44636
rect 5176 44580 5180 44636
rect 5116 44576 5180 44580
rect 97036 44636 97100 44640
rect 97036 44580 97040 44636
rect 97040 44580 97096 44636
rect 97096 44580 97100 44636
rect 97036 44576 97100 44580
rect 97116 44636 97180 44640
rect 97116 44580 97120 44636
rect 97120 44580 97176 44636
rect 97176 44580 97180 44636
rect 97116 44576 97180 44580
rect 97196 44636 97260 44640
rect 97196 44580 97200 44636
rect 97200 44580 97256 44636
rect 97256 44580 97260 44636
rect 97196 44576 97260 44580
rect 97276 44636 97340 44640
rect 97276 44580 97280 44636
rect 97280 44580 97336 44636
rect 97336 44580 97340 44636
rect 97276 44576 97340 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 96376 44092 96440 44096
rect 96376 44036 96380 44092
rect 96380 44036 96436 44092
rect 96436 44036 96440 44092
rect 96376 44032 96440 44036
rect 96456 44092 96520 44096
rect 96456 44036 96460 44092
rect 96460 44036 96516 44092
rect 96516 44036 96520 44092
rect 96456 44032 96520 44036
rect 96536 44092 96600 44096
rect 96536 44036 96540 44092
rect 96540 44036 96596 44092
rect 96596 44036 96600 44092
rect 96536 44032 96600 44036
rect 96616 44092 96680 44096
rect 96616 44036 96620 44092
rect 96620 44036 96676 44092
rect 96676 44036 96680 44092
rect 96616 44032 96680 44036
rect 4876 43548 4940 43552
rect 4876 43492 4880 43548
rect 4880 43492 4936 43548
rect 4936 43492 4940 43548
rect 4876 43488 4940 43492
rect 4956 43548 5020 43552
rect 4956 43492 4960 43548
rect 4960 43492 5016 43548
rect 5016 43492 5020 43548
rect 4956 43488 5020 43492
rect 5036 43548 5100 43552
rect 5036 43492 5040 43548
rect 5040 43492 5096 43548
rect 5096 43492 5100 43548
rect 5036 43488 5100 43492
rect 5116 43548 5180 43552
rect 5116 43492 5120 43548
rect 5120 43492 5176 43548
rect 5176 43492 5180 43548
rect 5116 43488 5180 43492
rect 97036 43548 97100 43552
rect 97036 43492 97040 43548
rect 97040 43492 97096 43548
rect 97096 43492 97100 43548
rect 97036 43488 97100 43492
rect 97116 43548 97180 43552
rect 97116 43492 97120 43548
rect 97120 43492 97176 43548
rect 97176 43492 97180 43548
rect 97116 43488 97180 43492
rect 97196 43548 97260 43552
rect 97196 43492 97200 43548
rect 97200 43492 97256 43548
rect 97256 43492 97260 43548
rect 97196 43488 97260 43492
rect 97276 43548 97340 43552
rect 97276 43492 97280 43548
rect 97280 43492 97336 43548
rect 97336 43492 97340 43548
rect 97276 43488 97340 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 96376 43004 96440 43008
rect 96376 42948 96380 43004
rect 96380 42948 96436 43004
rect 96436 42948 96440 43004
rect 96376 42944 96440 42948
rect 96456 43004 96520 43008
rect 96456 42948 96460 43004
rect 96460 42948 96516 43004
rect 96516 42948 96520 43004
rect 96456 42944 96520 42948
rect 96536 43004 96600 43008
rect 96536 42948 96540 43004
rect 96540 42948 96596 43004
rect 96596 42948 96600 43004
rect 96536 42944 96600 42948
rect 96616 43004 96680 43008
rect 96616 42948 96620 43004
rect 96620 42948 96676 43004
rect 96676 42948 96680 43004
rect 96616 42944 96680 42948
rect 4876 42460 4940 42464
rect 4876 42404 4880 42460
rect 4880 42404 4936 42460
rect 4936 42404 4940 42460
rect 4876 42400 4940 42404
rect 4956 42460 5020 42464
rect 4956 42404 4960 42460
rect 4960 42404 5016 42460
rect 5016 42404 5020 42460
rect 4956 42400 5020 42404
rect 5036 42460 5100 42464
rect 5036 42404 5040 42460
rect 5040 42404 5096 42460
rect 5096 42404 5100 42460
rect 5036 42400 5100 42404
rect 5116 42460 5180 42464
rect 5116 42404 5120 42460
rect 5120 42404 5176 42460
rect 5176 42404 5180 42460
rect 5116 42400 5180 42404
rect 97036 42460 97100 42464
rect 97036 42404 97040 42460
rect 97040 42404 97096 42460
rect 97096 42404 97100 42460
rect 97036 42400 97100 42404
rect 97116 42460 97180 42464
rect 97116 42404 97120 42460
rect 97120 42404 97176 42460
rect 97176 42404 97180 42460
rect 97116 42400 97180 42404
rect 97196 42460 97260 42464
rect 97196 42404 97200 42460
rect 97200 42404 97256 42460
rect 97256 42404 97260 42460
rect 97196 42400 97260 42404
rect 97276 42460 97340 42464
rect 97276 42404 97280 42460
rect 97280 42404 97336 42460
rect 97336 42404 97340 42460
rect 97276 42400 97340 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 96376 41916 96440 41920
rect 96376 41860 96380 41916
rect 96380 41860 96436 41916
rect 96436 41860 96440 41916
rect 96376 41856 96440 41860
rect 96456 41916 96520 41920
rect 96456 41860 96460 41916
rect 96460 41860 96516 41916
rect 96516 41860 96520 41916
rect 96456 41856 96520 41860
rect 96536 41916 96600 41920
rect 96536 41860 96540 41916
rect 96540 41860 96596 41916
rect 96596 41860 96600 41916
rect 96536 41856 96600 41860
rect 96616 41916 96680 41920
rect 96616 41860 96620 41916
rect 96620 41860 96676 41916
rect 96676 41860 96680 41916
rect 96616 41856 96680 41860
rect 4876 41372 4940 41376
rect 4876 41316 4880 41372
rect 4880 41316 4936 41372
rect 4936 41316 4940 41372
rect 4876 41312 4940 41316
rect 4956 41372 5020 41376
rect 4956 41316 4960 41372
rect 4960 41316 5016 41372
rect 5016 41316 5020 41372
rect 4956 41312 5020 41316
rect 5036 41372 5100 41376
rect 5036 41316 5040 41372
rect 5040 41316 5096 41372
rect 5096 41316 5100 41372
rect 5036 41312 5100 41316
rect 5116 41372 5180 41376
rect 5116 41316 5120 41372
rect 5120 41316 5176 41372
rect 5176 41316 5180 41372
rect 5116 41312 5180 41316
rect 97036 41372 97100 41376
rect 97036 41316 97040 41372
rect 97040 41316 97096 41372
rect 97096 41316 97100 41372
rect 97036 41312 97100 41316
rect 97116 41372 97180 41376
rect 97116 41316 97120 41372
rect 97120 41316 97176 41372
rect 97176 41316 97180 41372
rect 97116 41312 97180 41316
rect 97196 41372 97260 41376
rect 97196 41316 97200 41372
rect 97200 41316 97256 41372
rect 97256 41316 97260 41372
rect 97196 41312 97260 41316
rect 97276 41372 97340 41376
rect 97276 41316 97280 41372
rect 97280 41316 97336 41372
rect 97336 41316 97340 41372
rect 97276 41312 97340 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 96376 40828 96440 40832
rect 96376 40772 96380 40828
rect 96380 40772 96436 40828
rect 96436 40772 96440 40828
rect 96376 40768 96440 40772
rect 96456 40828 96520 40832
rect 96456 40772 96460 40828
rect 96460 40772 96516 40828
rect 96516 40772 96520 40828
rect 96456 40768 96520 40772
rect 96536 40828 96600 40832
rect 96536 40772 96540 40828
rect 96540 40772 96596 40828
rect 96596 40772 96600 40828
rect 96536 40768 96600 40772
rect 96616 40828 96680 40832
rect 96616 40772 96620 40828
rect 96620 40772 96676 40828
rect 96676 40772 96680 40828
rect 96616 40768 96680 40772
rect 4876 40284 4940 40288
rect 4876 40228 4880 40284
rect 4880 40228 4936 40284
rect 4936 40228 4940 40284
rect 4876 40224 4940 40228
rect 4956 40284 5020 40288
rect 4956 40228 4960 40284
rect 4960 40228 5016 40284
rect 5016 40228 5020 40284
rect 4956 40224 5020 40228
rect 5036 40284 5100 40288
rect 5036 40228 5040 40284
rect 5040 40228 5096 40284
rect 5096 40228 5100 40284
rect 5036 40224 5100 40228
rect 5116 40284 5180 40288
rect 5116 40228 5120 40284
rect 5120 40228 5176 40284
rect 5176 40228 5180 40284
rect 5116 40224 5180 40228
rect 97036 40284 97100 40288
rect 97036 40228 97040 40284
rect 97040 40228 97096 40284
rect 97096 40228 97100 40284
rect 97036 40224 97100 40228
rect 97116 40284 97180 40288
rect 97116 40228 97120 40284
rect 97120 40228 97176 40284
rect 97176 40228 97180 40284
rect 97116 40224 97180 40228
rect 97196 40284 97260 40288
rect 97196 40228 97200 40284
rect 97200 40228 97256 40284
rect 97256 40228 97260 40284
rect 97196 40224 97260 40228
rect 97276 40284 97340 40288
rect 97276 40228 97280 40284
rect 97280 40228 97336 40284
rect 97336 40228 97340 40284
rect 97276 40224 97340 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 96376 39740 96440 39744
rect 96376 39684 96380 39740
rect 96380 39684 96436 39740
rect 96436 39684 96440 39740
rect 96376 39680 96440 39684
rect 96456 39740 96520 39744
rect 96456 39684 96460 39740
rect 96460 39684 96516 39740
rect 96516 39684 96520 39740
rect 96456 39680 96520 39684
rect 96536 39740 96600 39744
rect 96536 39684 96540 39740
rect 96540 39684 96596 39740
rect 96596 39684 96600 39740
rect 96536 39680 96600 39684
rect 96616 39740 96680 39744
rect 96616 39684 96620 39740
rect 96620 39684 96676 39740
rect 96676 39684 96680 39740
rect 96616 39680 96680 39684
rect 4876 39196 4940 39200
rect 4876 39140 4880 39196
rect 4880 39140 4936 39196
rect 4936 39140 4940 39196
rect 4876 39136 4940 39140
rect 4956 39196 5020 39200
rect 4956 39140 4960 39196
rect 4960 39140 5016 39196
rect 5016 39140 5020 39196
rect 4956 39136 5020 39140
rect 5036 39196 5100 39200
rect 5036 39140 5040 39196
rect 5040 39140 5096 39196
rect 5096 39140 5100 39196
rect 5036 39136 5100 39140
rect 5116 39196 5180 39200
rect 5116 39140 5120 39196
rect 5120 39140 5176 39196
rect 5176 39140 5180 39196
rect 5116 39136 5180 39140
rect 97036 39196 97100 39200
rect 97036 39140 97040 39196
rect 97040 39140 97096 39196
rect 97096 39140 97100 39196
rect 97036 39136 97100 39140
rect 97116 39196 97180 39200
rect 97116 39140 97120 39196
rect 97120 39140 97176 39196
rect 97176 39140 97180 39196
rect 97116 39136 97180 39140
rect 97196 39196 97260 39200
rect 97196 39140 97200 39196
rect 97200 39140 97256 39196
rect 97256 39140 97260 39196
rect 97196 39136 97260 39140
rect 97276 39196 97340 39200
rect 97276 39140 97280 39196
rect 97280 39140 97336 39196
rect 97336 39140 97340 39196
rect 97276 39136 97340 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 96376 38652 96440 38656
rect 96376 38596 96380 38652
rect 96380 38596 96436 38652
rect 96436 38596 96440 38652
rect 96376 38592 96440 38596
rect 96456 38652 96520 38656
rect 96456 38596 96460 38652
rect 96460 38596 96516 38652
rect 96516 38596 96520 38652
rect 96456 38592 96520 38596
rect 96536 38652 96600 38656
rect 96536 38596 96540 38652
rect 96540 38596 96596 38652
rect 96596 38596 96600 38652
rect 96536 38592 96600 38596
rect 96616 38652 96680 38656
rect 96616 38596 96620 38652
rect 96620 38596 96676 38652
rect 96676 38596 96680 38652
rect 96616 38592 96680 38596
rect 4876 38108 4940 38112
rect 4876 38052 4880 38108
rect 4880 38052 4936 38108
rect 4936 38052 4940 38108
rect 4876 38048 4940 38052
rect 4956 38108 5020 38112
rect 4956 38052 4960 38108
rect 4960 38052 5016 38108
rect 5016 38052 5020 38108
rect 4956 38048 5020 38052
rect 5036 38108 5100 38112
rect 5036 38052 5040 38108
rect 5040 38052 5096 38108
rect 5096 38052 5100 38108
rect 5036 38048 5100 38052
rect 5116 38108 5180 38112
rect 5116 38052 5120 38108
rect 5120 38052 5176 38108
rect 5176 38052 5180 38108
rect 5116 38048 5180 38052
rect 97036 38108 97100 38112
rect 97036 38052 97040 38108
rect 97040 38052 97096 38108
rect 97096 38052 97100 38108
rect 97036 38048 97100 38052
rect 97116 38108 97180 38112
rect 97116 38052 97120 38108
rect 97120 38052 97176 38108
rect 97176 38052 97180 38108
rect 97116 38048 97180 38052
rect 97196 38108 97260 38112
rect 97196 38052 97200 38108
rect 97200 38052 97256 38108
rect 97256 38052 97260 38108
rect 97196 38048 97260 38052
rect 97276 38108 97340 38112
rect 97276 38052 97280 38108
rect 97280 38052 97336 38108
rect 97336 38052 97340 38108
rect 97276 38048 97340 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 96376 37564 96440 37568
rect 96376 37508 96380 37564
rect 96380 37508 96436 37564
rect 96436 37508 96440 37564
rect 96376 37504 96440 37508
rect 96456 37564 96520 37568
rect 96456 37508 96460 37564
rect 96460 37508 96516 37564
rect 96516 37508 96520 37564
rect 96456 37504 96520 37508
rect 96536 37564 96600 37568
rect 96536 37508 96540 37564
rect 96540 37508 96596 37564
rect 96596 37508 96600 37564
rect 96536 37504 96600 37508
rect 96616 37564 96680 37568
rect 96616 37508 96620 37564
rect 96620 37508 96676 37564
rect 96676 37508 96680 37564
rect 96616 37504 96680 37508
rect 4876 37020 4940 37024
rect 4876 36964 4880 37020
rect 4880 36964 4936 37020
rect 4936 36964 4940 37020
rect 4876 36960 4940 36964
rect 4956 37020 5020 37024
rect 4956 36964 4960 37020
rect 4960 36964 5016 37020
rect 5016 36964 5020 37020
rect 4956 36960 5020 36964
rect 5036 37020 5100 37024
rect 5036 36964 5040 37020
rect 5040 36964 5096 37020
rect 5096 36964 5100 37020
rect 5036 36960 5100 36964
rect 5116 37020 5180 37024
rect 5116 36964 5120 37020
rect 5120 36964 5176 37020
rect 5176 36964 5180 37020
rect 5116 36960 5180 36964
rect 97036 37020 97100 37024
rect 97036 36964 97040 37020
rect 97040 36964 97096 37020
rect 97096 36964 97100 37020
rect 97036 36960 97100 36964
rect 97116 37020 97180 37024
rect 97116 36964 97120 37020
rect 97120 36964 97176 37020
rect 97176 36964 97180 37020
rect 97116 36960 97180 36964
rect 97196 37020 97260 37024
rect 97196 36964 97200 37020
rect 97200 36964 97256 37020
rect 97256 36964 97260 37020
rect 97196 36960 97260 36964
rect 97276 37020 97340 37024
rect 97276 36964 97280 37020
rect 97280 36964 97336 37020
rect 97336 36964 97340 37020
rect 97276 36960 97340 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 96376 36476 96440 36480
rect 96376 36420 96380 36476
rect 96380 36420 96436 36476
rect 96436 36420 96440 36476
rect 96376 36416 96440 36420
rect 96456 36476 96520 36480
rect 96456 36420 96460 36476
rect 96460 36420 96516 36476
rect 96516 36420 96520 36476
rect 96456 36416 96520 36420
rect 96536 36476 96600 36480
rect 96536 36420 96540 36476
rect 96540 36420 96596 36476
rect 96596 36420 96600 36476
rect 96536 36416 96600 36420
rect 96616 36476 96680 36480
rect 96616 36420 96620 36476
rect 96620 36420 96676 36476
rect 96676 36420 96680 36476
rect 96616 36416 96680 36420
rect 4876 35932 4940 35936
rect 4876 35876 4880 35932
rect 4880 35876 4936 35932
rect 4936 35876 4940 35932
rect 4876 35872 4940 35876
rect 4956 35932 5020 35936
rect 4956 35876 4960 35932
rect 4960 35876 5016 35932
rect 5016 35876 5020 35932
rect 4956 35872 5020 35876
rect 5036 35932 5100 35936
rect 5036 35876 5040 35932
rect 5040 35876 5096 35932
rect 5096 35876 5100 35932
rect 5036 35872 5100 35876
rect 5116 35932 5180 35936
rect 5116 35876 5120 35932
rect 5120 35876 5176 35932
rect 5176 35876 5180 35932
rect 5116 35872 5180 35876
rect 97036 35932 97100 35936
rect 97036 35876 97040 35932
rect 97040 35876 97096 35932
rect 97096 35876 97100 35932
rect 97036 35872 97100 35876
rect 97116 35932 97180 35936
rect 97116 35876 97120 35932
rect 97120 35876 97176 35932
rect 97176 35876 97180 35932
rect 97116 35872 97180 35876
rect 97196 35932 97260 35936
rect 97196 35876 97200 35932
rect 97200 35876 97256 35932
rect 97256 35876 97260 35932
rect 97196 35872 97260 35876
rect 97276 35932 97340 35936
rect 97276 35876 97280 35932
rect 97280 35876 97336 35932
rect 97336 35876 97340 35932
rect 97276 35872 97340 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 96376 35388 96440 35392
rect 96376 35332 96380 35388
rect 96380 35332 96436 35388
rect 96436 35332 96440 35388
rect 96376 35328 96440 35332
rect 96456 35388 96520 35392
rect 96456 35332 96460 35388
rect 96460 35332 96516 35388
rect 96516 35332 96520 35388
rect 96456 35328 96520 35332
rect 96536 35388 96600 35392
rect 96536 35332 96540 35388
rect 96540 35332 96596 35388
rect 96596 35332 96600 35388
rect 96536 35328 96600 35332
rect 96616 35388 96680 35392
rect 96616 35332 96620 35388
rect 96620 35332 96676 35388
rect 96676 35332 96680 35388
rect 96616 35328 96680 35332
rect 4876 34844 4940 34848
rect 4876 34788 4880 34844
rect 4880 34788 4936 34844
rect 4936 34788 4940 34844
rect 4876 34784 4940 34788
rect 4956 34844 5020 34848
rect 4956 34788 4960 34844
rect 4960 34788 5016 34844
rect 5016 34788 5020 34844
rect 4956 34784 5020 34788
rect 5036 34844 5100 34848
rect 5036 34788 5040 34844
rect 5040 34788 5096 34844
rect 5096 34788 5100 34844
rect 5036 34784 5100 34788
rect 5116 34844 5180 34848
rect 5116 34788 5120 34844
rect 5120 34788 5176 34844
rect 5176 34788 5180 34844
rect 5116 34784 5180 34788
rect 97036 34844 97100 34848
rect 97036 34788 97040 34844
rect 97040 34788 97096 34844
rect 97096 34788 97100 34844
rect 97036 34784 97100 34788
rect 97116 34844 97180 34848
rect 97116 34788 97120 34844
rect 97120 34788 97176 34844
rect 97176 34788 97180 34844
rect 97116 34784 97180 34788
rect 97196 34844 97260 34848
rect 97196 34788 97200 34844
rect 97200 34788 97256 34844
rect 97256 34788 97260 34844
rect 97196 34784 97260 34788
rect 97276 34844 97340 34848
rect 97276 34788 97280 34844
rect 97280 34788 97336 34844
rect 97336 34788 97340 34844
rect 97276 34784 97340 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 96376 34300 96440 34304
rect 96376 34244 96380 34300
rect 96380 34244 96436 34300
rect 96436 34244 96440 34300
rect 96376 34240 96440 34244
rect 96456 34300 96520 34304
rect 96456 34244 96460 34300
rect 96460 34244 96516 34300
rect 96516 34244 96520 34300
rect 96456 34240 96520 34244
rect 96536 34300 96600 34304
rect 96536 34244 96540 34300
rect 96540 34244 96596 34300
rect 96596 34244 96600 34300
rect 96536 34240 96600 34244
rect 96616 34300 96680 34304
rect 96616 34244 96620 34300
rect 96620 34244 96676 34300
rect 96676 34244 96680 34300
rect 96616 34240 96680 34244
rect 4876 33756 4940 33760
rect 4876 33700 4880 33756
rect 4880 33700 4936 33756
rect 4936 33700 4940 33756
rect 4876 33696 4940 33700
rect 4956 33756 5020 33760
rect 4956 33700 4960 33756
rect 4960 33700 5016 33756
rect 5016 33700 5020 33756
rect 4956 33696 5020 33700
rect 5036 33756 5100 33760
rect 5036 33700 5040 33756
rect 5040 33700 5096 33756
rect 5096 33700 5100 33756
rect 5036 33696 5100 33700
rect 5116 33756 5180 33760
rect 5116 33700 5120 33756
rect 5120 33700 5176 33756
rect 5176 33700 5180 33756
rect 5116 33696 5180 33700
rect 97036 33756 97100 33760
rect 97036 33700 97040 33756
rect 97040 33700 97096 33756
rect 97096 33700 97100 33756
rect 97036 33696 97100 33700
rect 97116 33756 97180 33760
rect 97116 33700 97120 33756
rect 97120 33700 97176 33756
rect 97176 33700 97180 33756
rect 97116 33696 97180 33700
rect 97196 33756 97260 33760
rect 97196 33700 97200 33756
rect 97200 33700 97256 33756
rect 97256 33700 97260 33756
rect 97196 33696 97260 33700
rect 97276 33756 97340 33760
rect 97276 33700 97280 33756
rect 97280 33700 97336 33756
rect 97336 33700 97340 33756
rect 97276 33696 97340 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 96376 33212 96440 33216
rect 96376 33156 96380 33212
rect 96380 33156 96436 33212
rect 96436 33156 96440 33212
rect 96376 33152 96440 33156
rect 96456 33212 96520 33216
rect 96456 33156 96460 33212
rect 96460 33156 96516 33212
rect 96516 33156 96520 33212
rect 96456 33152 96520 33156
rect 96536 33212 96600 33216
rect 96536 33156 96540 33212
rect 96540 33156 96596 33212
rect 96596 33156 96600 33212
rect 96536 33152 96600 33156
rect 96616 33212 96680 33216
rect 96616 33156 96620 33212
rect 96620 33156 96676 33212
rect 96676 33156 96680 33212
rect 96616 33152 96680 33156
rect 4876 32668 4940 32672
rect 4876 32612 4880 32668
rect 4880 32612 4936 32668
rect 4936 32612 4940 32668
rect 4876 32608 4940 32612
rect 4956 32668 5020 32672
rect 4956 32612 4960 32668
rect 4960 32612 5016 32668
rect 5016 32612 5020 32668
rect 4956 32608 5020 32612
rect 5036 32668 5100 32672
rect 5036 32612 5040 32668
rect 5040 32612 5096 32668
rect 5096 32612 5100 32668
rect 5036 32608 5100 32612
rect 5116 32668 5180 32672
rect 5116 32612 5120 32668
rect 5120 32612 5176 32668
rect 5176 32612 5180 32668
rect 5116 32608 5180 32612
rect 97036 32668 97100 32672
rect 97036 32612 97040 32668
rect 97040 32612 97096 32668
rect 97096 32612 97100 32668
rect 97036 32608 97100 32612
rect 97116 32668 97180 32672
rect 97116 32612 97120 32668
rect 97120 32612 97176 32668
rect 97176 32612 97180 32668
rect 97116 32608 97180 32612
rect 97196 32668 97260 32672
rect 97196 32612 97200 32668
rect 97200 32612 97256 32668
rect 97256 32612 97260 32668
rect 97196 32608 97260 32612
rect 97276 32668 97340 32672
rect 97276 32612 97280 32668
rect 97280 32612 97336 32668
rect 97336 32612 97340 32668
rect 97276 32608 97340 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 96376 32124 96440 32128
rect 96376 32068 96380 32124
rect 96380 32068 96436 32124
rect 96436 32068 96440 32124
rect 96376 32064 96440 32068
rect 96456 32124 96520 32128
rect 96456 32068 96460 32124
rect 96460 32068 96516 32124
rect 96516 32068 96520 32124
rect 96456 32064 96520 32068
rect 96536 32124 96600 32128
rect 96536 32068 96540 32124
rect 96540 32068 96596 32124
rect 96596 32068 96600 32124
rect 96536 32064 96600 32068
rect 96616 32124 96680 32128
rect 96616 32068 96620 32124
rect 96620 32068 96676 32124
rect 96676 32068 96680 32124
rect 96616 32064 96680 32068
rect 4876 31580 4940 31584
rect 4876 31524 4880 31580
rect 4880 31524 4936 31580
rect 4936 31524 4940 31580
rect 4876 31520 4940 31524
rect 4956 31580 5020 31584
rect 4956 31524 4960 31580
rect 4960 31524 5016 31580
rect 5016 31524 5020 31580
rect 4956 31520 5020 31524
rect 5036 31580 5100 31584
rect 5036 31524 5040 31580
rect 5040 31524 5096 31580
rect 5096 31524 5100 31580
rect 5036 31520 5100 31524
rect 5116 31580 5180 31584
rect 5116 31524 5120 31580
rect 5120 31524 5176 31580
rect 5176 31524 5180 31580
rect 5116 31520 5180 31524
rect 97036 31580 97100 31584
rect 97036 31524 97040 31580
rect 97040 31524 97096 31580
rect 97096 31524 97100 31580
rect 97036 31520 97100 31524
rect 97116 31580 97180 31584
rect 97116 31524 97120 31580
rect 97120 31524 97176 31580
rect 97176 31524 97180 31580
rect 97116 31520 97180 31524
rect 97196 31580 97260 31584
rect 97196 31524 97200 31580
rect 97200 31524 97256 31580
rect 97256 31524 97260 31580
rect 97196 31520 97260 31524
rect 97276 31580 97340 31584
rect 97276 31524 97280 31580
rect 97280 31524 97336 31580
rect 97336 31524 97340 31580
rect 97276 31520 97340 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 96376 31036 96440 31040
rect 96376 30980 96380 31036
rect 96380 30980 96436 31036
rect 96436 30980 96440 31036
rect 96376 30976 96440 30980
rect 96456 31036 96520 31040
rect 96456 30980 96460 31036
rect 96460 30980 96516 31036
rect 96516 30980 96520 31036
rect 96456 30976 96520 30980
rect 96536 31036 96600 31040
rect 96536 30980 96540 31036
rect 96540 30980 96596 31036
rect 96596 30980 96600 31036
rect 96536 30976 96600 30980
rect 96616 31036 96680 31040
rect 96616 30980 96620 31036
rect 96620 30980 96676 31036
rect 96676 30980 96680 31036
rect 96616 30976 96680 30980
rect 4876 30492 4940 30496
rect 4876 30436 4880 30492
rect 4880 30436 4936 30492
rect 4936 30436 4940 30492
rect 4876 30432 4940 30436
rect 4956 30492 5020 30496
rect 4956 30436 4960 30492
rect 4960 30436 5016 30492
rect 5016 30436 5020 30492
rect 4956 30432 5020 30436
rect 5036 30492 5100 30496
rect 5036 30436 5040 30492
rect 5040 30436 5096 30492
rect 5096 30436 5100 30492
rect 5036 30432 5100 30436
rect 5116 30492 5180 30496
rect 5116 30436 5120 30492
rect 5120 30436 5176 30492
rect 5176 30436 5180 30492
rect 5116 30432 5180 30436
rect 97036 30492 97100 30496
rect 97036 30436 97040 30492
rect 97040 30436 97096 30492
rect 97096 30436 97100 30492
rect 97036 30432 97100 30436
rect 97116 30492 97180 30496
rect 97116 30436 97120 30492
rect 97120 30436 97176 30492
rect 97176 30436 97180 30492
rect 97116 30432 97180 30436
rect 97196 30492 97260 30496
rect 97196 30436 97200 30492
rect 97200 30436 97256 30492
rect 97256 30436 97260 30492
rect 97196 30432 97260 30436
rect 97276 30492 97340 30496
rect 97276 30436 97280 30492
rect 97280 30436 97336 30492
rect 97336 30436 97340 30492
rect 97276 30432 97340 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 96376 29948 96440 29952
rect 96376 29892 96380 29948
rect 96380 29892 96436 29948
rect 96436 29892 96440 29948
rect 96376 29888 96440 29892
rect 96456 29948 96520 29952
rect 96456 29892 96460 29948
rect 96460 29892 96516 29948
rect 96516 29892 96520 29948
rect 96456 29888 96520 29892
rect 96536 29948 96600 29952
rect 96536 29892 96540 29948
rect 96540 29892 96596 29948
rect 96596 29892 96600 29948
rect 96536 29888 96600 29892
rect 96616 29948 96680 29952
rect 96616 29892 96620 29948
rect 96620 29892 96676 29948
rect 96676 29892 96680 29948
rect 96616 29888 96680 29892
rect 4876 29404 4940 29408
rect 4876 29348 4880 29404
rect 4880 29348 4936 29404
rect 4936 29348 4940 29404
rect 4876 29344 4940 29348
rect 4956 29404 5020 29408
rect 4956 29348 4960 29404
rect 4960 29348 5016 29404
rect 5016 29348 5020 29404
rect 4956 29344 5020 29348
rect 5036 29404 5100 29408
rect 5036 29348 5040 29404
rect 5040 29348 5096 29404
rect 5096 29348 5100 29404
rect 5036 29344 5100 29348
rect 5116 29404 5180 29408
rect 5116 29348 5120 29404
rect 5120 29348 5176 29404
rect 5176 29348 5180 29404
rect 5116 29344 5180 29348
rect 97036 29404 97100 29408
rect 97036 29348 97040 29404
rect 97040 29348 97096 29404
rect 97096 29348 97100 29404
rect 97036 29344 97100 29348
rect 97116 29404 97180 29408
rect 97116 29348 97120 29404
rect 97120 29348 97176 29404
rect 97176 29348 97180 29404
rect 97116 29344 97180 29348
rect 97196 29404 97260 29408
rect 97196 29348 97200 29404
rect 97200 29348 97256 29404
rect 97256 29348 97260 29404
rect 97196 29344 97260 29348
rect 97276 29404 97340 29408
rect 97276 29348 97280 29404
rect 97280 29348 97336 29404
rect 97336 29348 97340 29404
rect 97276 29344 97340 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 96376 28860 96440 28864
rect 96376 28804 96380 28860
rect 96380 28804 96436 28860
rect 96436 28804 96440 28860
rect 96376 28800 96440 28804
rect 96456 28860 96520 28864
rect 96456 28804 96460 28860
rect 96460 28804 96516 28860
rect 96516 28804 96520 28860
rect 96456 28800 96520 28804
rect 96536 28860 96600 28864
rect 96536 28804 96540 28860
rect 96540 28804 96596 28860
rect 96596 28804 96600 28860
rect 96536 28800 96600 28804
rect 96616 28860 96680 28864
rect 96616 28804 96620 28860
rect 96620 28804 96676 28860
rect 96676 28804 96680 28860
rect 96616 28800 96680 28804
rect 4876 28316 4940 28320
rect 4876 28260 4880 28316
rect 4880 28260 4936 28316
rect 4936 28260 4940 28316
rect 4876 28256 4940 28260
rect 4956 28316 5020 28320
rect 4956 28260 4960 28316
rect 4960 28260 5016 28316
rect 5016 28260 5020 28316
rect 4956 28256 5020 28260
rect 5036 28316 5100 28320
rect 5036 28260 5040 28316
rect 5040 28260 5096 28316
rect 5096 28260 5100 28316
rect 5036 28256 5100 28260
rect 5116 28316 5180 28320
rect 5116 28260 5120 28316
rect 5120 28260 5176 28316
rect 5176 28260 5180 28316
rect 5116 28256 5180 28260
rect 97036 28316 97100 28320
rect 97036 28260 97040 28316
rect 97040 28260 97096 28316
rect 97096 28260 97100 28316
rect 97036 28256 97100 28260
rect 97116 28316 97180 28320
rect 97116 28260 97120 28316
rect 97120 28260 97176 28316
rect 97176 28260 97180 28316
rect 97116 28256 97180 28260
rect 97196 28316 97260 28320
rect 97196 28260 97200 28316
rect 97200 28260 97256 28316
rect 97256 28260 97260 28316
rect 97196 28256 97260 28260
rect 97276 28316 97340 28320
rect 97276 28260 97280 28316
rect 97280 28260 97336 28316
rect 97336 28260 97340 28316
rect 97276 28256 97340 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 96376 27772 96440 27776
rect 96376 27716 96380 27772
rect 96380 27716 96436 27772
rect 96436 27716 96440 27772
rect 96376 27712 96440 27716
rect 96456 27772 96520 27776
rect 96456 27716 96460 27772
rect 96460 27716 96516 27772
rect 96516 27716 96520 27772
rect 96456 27712 96520 27716
rect 96536 27772 96600 27776
rect 96536 27716 96540 27772
rect 96540 27716 96596 27772
rect 96596 27716 96600 27772
rect 96536 27712 96600 27716
rect 96616 27772 96680 27776
rect 96616 27716 96620 27772
rect 96620 27716 96676 27772
rect 96676 27716 96680 27772
rect 96616 27712 96680 27716
rect 4876 27228 4940 27232
rect 4876 27172 4880 27228
rect 4880 27172 4936 27228
rect 4936 27172 4940 27228
rect 4876 27168 4940 27172
rect 4956 27228 5020 27232
rect 4956 27172 4960 27228
rect 4960 27172 5016 27228
rect 5016 27172 5020 27228
rect 4956 27168 5020 27172
rect 5036 27228 5100 27232
rect 5036 27172 5040 27228
rect 5040 27172 5096 27228
rect 5096 27172 5100 27228
rect 5036 27168 5100 27172
rect 5116 27228 5180 27232
rect 5116 27172 5120 27228
rect 5120 27172 5176 27228
rect 5176 27172 5180 27228
rect 5116 27168 5180 27172
rect 97036 27228 97100 27232
rect 97036 27172 97040 27228
rect 97040 27172 97096 27228
rect 97096 27172 97100 27228
rect 97036 27168 97100 27172
rect 97116 27228 97180 27232
rect 97116 27172 97120 27228
rect 97120 27172 97176 27228
rect 97176 27172 97180 27228
rect 97116 27168 97180 27172
rect 97196 27228 97260 27232
rect 97196 27172 97200 27228
rect 97200 27172 97256 27228
rect 97256 27172 97260 27228
rect 97196 27168 97260 27172
rect 97276 27228 97340 27232
rect 97276 27172 97280 27228
rect 97280 27172 97336 27228
rect 97336 27172 97340 27228
rect 97276 27168 97340 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 96376 26684 96440 26688
rect 96376 26628 96380 26684
rect 96380 26628 96436 26684
rect 96436 26628 96440 26684
rect 96376 26624 96440 26628
rect 96456 26684 96520 26688
rect 96456 26628 96460 26684
rect 96460 26628 96516 26684
rect 96516 26628 96520 26684
rect 96456 26624 96520 26628
rect 96536 26684 96600 26688
rect 96536 26628 96540 26684
rect 96540 26628 96596 26684
rect 96596 26628 96600 26684
rect 96536 26624 96600 26628
rect 96616 26684 96680 26688
rect 96616 26628 96620 26684
rect 96620 26628 96676 26684
rect 96676 26628 96680 26684
rect 96616 26624 96680 26628
rect 4876 26140 4940 26144
rect 4876 26084 4880 26140
rect 4880 26084 4936 26140
rect 4936 26084 4940 26140
rect 4876 26080 4940 26084
rect 4956 26140 5020 26144
rect 4956 26084 4960 26140
rect 4960 26084 5016 26140
rect 5016 26084 5020 26140
rect 4956 26080 5020 26084
rect 5036 26140 5100 26144
rect 5036 26084 5040 26140
rect 5040 26084 5096 26140
rect 5096 26084 5100 26140
rect 5036 26080 5100 26084
rect 5116 26140 5180 26144
rect 5116 26084 5120 26140
rect 5120 26084 5176 26140
rect 5176 26084 5180 26140
rect 5116 26080 5180 26084
rect 97036 26140 97100 26144
rect 97036 26084 97040 26140
rect 97040 26084 97096 26140
rect 97096 26084 97100 26140
rect 97036 26080 97100 26084
rect 97116 26140 97180 26144
rect 97116 26084 97120 26140
rect 97120 26084 97176 26140
rect 97176 26084 97180 26140
rect 97116 26080 97180 26084
rect 97196 26140 97260 26144
rect 97196 26084 97200 26140
rect 97200 26084 97256 26140
rect 97256 26084 97260 26140
rect 97196 26080 97260 26084
rect 97276 26140 97340 26144
rect 97276 26084 97280 26140
rect 97280 26084 97336 26140
rect 97336 26084 97340 26140
rect 97276 26080 97340 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 96376 25596 96440 25600
rect 96376 25540 96380 25596
rect 96380 25540 96436 25596
rect 96436 25540 96440 25596
rect 96376 25536 96440 25540
rect 96456 25596 96520 25600
rect 96456 25540 96460 25596
rect 96460 25540 96516 25596
rect 96516 25540 96520 25596
rect 96456 25536 96520 25540
rect 96536 25596 96600 25600
rect 96536 25540 96540 25596
rect 96540 25540 96596 25596
rect 96596 25540 96600 25596
rect 96536 25536 96600 25540
rect 96616 25596 96680 25600
rect 96616 25540 96620 25596
rect 96620 25540 96676 25596
rect 96676 25540 96680 25596
rect 96616 25536 96680 25540
rect 4876 25052 4940 25056
rect 4876 24996 4880 25052
rect 4880 24996 4936 25052
rect 4936 24996 4940 25052
rect 4876 24992 4940 24996
rect 4956 25052 5020 25056
rect 4956 24996 4960 25052
rect 4960 24996 5016 25052
rect 5016 24996 5020 25052
rect 4956 24992 5020 24996
rect 5036 25052 5100 25056
rect 5036 24996 5040 25052
rect 5040 24996 5096 25052
rect 5096 24996 5100 25052
rect 5036 24992 5100 24996
rect 5116 25052 5180 25056
rect 5116 24996 5120 25052
rect 5120 24996 5176 25052
rect 5176 24996 5180 25052
rect 5116 24992 5180 24996
rect 97036 25052 97100 25056
rect 97036 24996 97040 25052
rect 97040 24996 97096 25052
rect 97096 24996 97100 25052
rect 97036 24992 97100 24996
rect 97116 25052 97180 25056
rect 97116 24996 97120 25052
rect 97120 24996 97176 25052
rect 97176 24996 97180 25052
rect 97116 24992 97180 24996
rect 97196 25052 97260 25056
rect 97196 24996 97200 25052
rect 97200 24996 97256 25052
rect 97256 24996 97260 25052
rect 97196 24992 97260 24996
rect 97276 25052 97340 25056
rect 97276 24996 97280 25052
rect 97280 24996 97336 25052
rect 97336 24996 97340 25052
rect 97276 24992 97340 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 96376 24508 96440 24512
rect 96376 24452 96380 24508
rect 96380 24452 96436 24508
rect 96436 24452 96440 24508
rect 96376 24448 96440 24452
rect 96456 24508 96520 24512
rect 96456 24452 96460 24508
rect 96460 24452 96516 24508
rect 96516 24452 96520 24508
rect 96456 24448 96520 24452
rect 96536 24508 96600 24512
rect 96536 24452 96540 24508
rect 96540 24452 96596 24508
rect 96596 24452 96600 24508
rect 96536 24448 96600 24452
rect 96616 24508 96680 24512
rect 96616 24452 96620 24508
rect 96620 24452 96676 24508
rect 96676 24452 96680 24508
rect 96616 24448 96680 24452
rect 4876 23964 4940 23968
rect 4876 23908 4880 23964
rect 4880 23908 4936 23964
rect 4936 23908 4940 23964
rect 4876 23904 4940 23908
rect 4956 23964 5020 23968
rect 4956 23908 4960 23964
rect 4960 23908 5016 23964
rect 5016 23908 5020 23964
rect 4956 23904 5020 23908
rect 5036 23964 5100 23968
rect 5036 23908 5040 23964
rect 5040 23908 5096 23964
rect 5096 23908 5100 23964
rect 5036 23904 5100 23908
rect 5116 23964 5180 23968
rect 5116 23908 5120 23964
rect 5120 23908 5176 23964
rect 5176 23908 5180 23964
rect 5116 23904 5180 23908
rect 97036 23964 97100 23968
rect 97036 23908 97040 23964
rect 97040 23908 97096 23964
rect 97096 23908 97100 23964
rect 97036 23904 97100 23908
rect 97116 23964 97180 23968
rect 97116 23908 97120 23964
rect 97120 23908 97176 23964
rect 97176 23908 97180 23964
rect 97116 23904 97180 23908
rect 97196 23964 97260 23968
rect 97196 23908 97200 23964
rect 97200 23908 97256 23964
rect 97256 23908 97260 23964
rect 97196 23904 97260 23908
rect 97276 23964 97340 23968
rect 97276 23908 97280 23964
rect 97280 23908 97336 23964
rect 97336 23908 97340 23964
rect 97276 23904 97340 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 96376 23420 96440 23424
rect 96376 23364 96380 23420
rect 96380 23364 96436 23420
rect 96436 23364 96440 23420
rect 96376 23360 96440 23364
rect 96456 23420 96520 23424
rect 96456 23364 96460 23420
rect 96460 23364 96516 23420
rect 96516 23364 96520 23420
rect 96456 23360 96520 23364
rect 96536 23420 96600 23424
rect 96536 23364 96540 23420
rect 96540 23364 96596 23420
rect 96596 23364 96600 23420
rect 96536 23360 96600 23364
rect 96616 23420 96680 23424
rect 96616 23364 96620 23420
rect 96620 23364 96676 23420
rect 96676 23364 96680 23420
rect 96616 23360 96680 23364
rect 4876 22876 4940 22880
rect 4876 22820 4880 22876
rect 4880 22820 4936 22876
rect 4936 22820 4940 22876
rect 4876 22816 4940 22820
rect 4956 22876 5020 22880
rect 4956 22820 4960 22876
rect 4960 22820 5016 22876
rect 5016 22820 5020 22876
rect 4956 22816 5020 22820
rect 5036 22876 5100 22880
rect 5036 22820 5040 22876
rect 5040 22820 5096 22876
rect 5096 22820 5100 22876
rect 5036 22816 5100 22820
rect 5116 22876 5180 22880
rect 5116 22820 5120 22876
rect 5120 22820 5176 22876
rect 5176 22820 5180 22876
rect 5116 22816 5180 22820
rect 97036 22876 97100 22880
rect 97036 22820 97040 22876
rect 97040 22820 97096 22876
rect 97096 22820 97100 22876
rect 97036 22816 97100 22820
rect 97116 22876 97180 22880
rect 97116 22820 97120 22876
rect 97120 22820 97176 22876
rect 97176 22820 97180 22876
rect 97116 22816 97180 22820
rect 97196 22876 97260 22880
rect 97196 22820 97200 22876
rect 97200 22820 97256 22876
rect 97256 22820 97260 22876
rect 97196 22816 97260 22820
rect 97276 22876 97340 22880
rect 97276 22820 97280 22876
rect 97280 22820 97336 22876
rect 97336 22820 97340 22876
rect 97276 22816 97340 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 96376 22332 96440 22336
rect 96376 22276 96380 22332
rect 96380 22276 96436 22332
rect 96436 22276 96440 22332
rect 96376 22272 96440 22276
rect 96456 22332 96520 22336
rect 96456 22276 96460 22332
rect 96460 22276 96516 22332
rect 96516 22276 96520 22332
rect 96456 22272 96520 22276
rect 96536 22332 96600 22336
rect 96536 22276 96540 22332
rect 96540 22276 96596 22332
rect 96596 22276 96600 22332
rect 96536 22272 96600 22276
rect 96616 22332 96680 22336
rect 96616 22276 96620 22332
rect 96620 22276 96676 22332
rect 96676 22276 96680 22332
rect 96616 22272 96680 22276
rect 4876 21788 4940 21792
rect 4876 21732 4880 21788
rect 4880 21732 4936 21788
rect 4936 21732 4940 21788
rect 4876 21728 4940 21732
rect 4956 21788 5020 21792
rect 4956 21732 4960 21788
rect 4960 21732 5016 21788
rect 5016 21732 5020 21788
rect 4956 21728 5020 21732
rect 5036 21788 5100 21792
rect 5036 21732 5040 21788
rect 5040 21732 5096 21788
rect 5096 21732 5100 21788
rect 5036 21728 5100 21732
rect 5116 21788 5180 21792
rect 5116 21732 5120 21788
rect 5120 21732 5176 21788
rect 5176 21732 5180 21788
rect 5116 21728 5180 21732
rect 97036 21788 97100 21792
rect 97036 21732 97040 21788
rect 97040 21732 97096 21788
rect 97096 21732 97100 21788
rect 97036 21728 97100 21732
rect 97116 21788 97180 21792
rect 97116 21732 97120 21788
rect 97120 21732 97176 21788
rect 97176 21732 97180 21788
rect 97116 21728 97180 21732
rect 97196 21788 97260 21792
rect 97196 21732 97200 21788
rect 97200 21732 97256 21788
rect 97256 21732 97260 21788
rect 97196 21728 97260 21732
rect 97276 21788 97340 21792
rect 97276 21732 97280 21788
rect 97280 21732 97336 21788
rect 97336 21732 97340 21788
rect 97276 21728 97340 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 96376 21244 96440 21248
rect 96376 21188 96380 21244
rect 96380 21188 96436 21244
rect 96436 21188 96440 21244
rect 96376 21184 96440 21188
rect 96456 21244 96520 21248
rect 96456 21188 96460 21244
rect 96460 21188 96516 21244
rect 96516 21188 96520 21244
rect 96456 21184 96520 21188
rect 96536 21244 96600 21248
rect 96536 21188 96540 21244
rect 96540 21188 96596 21244
rect 96596 21188 96600 21244
rect 96536 21184 96600 21188
rect 96616 21244 96680 21248
rect 96616 21188 96620 21244
rect 96620 21188 96676 21244
rect 96676 21188 96680 21244
rect 96616 21184 96680 21188
rect 4876 20700 4940 20704
rect 4876 20644 4880 20700
rect 4880 20644 4936 20700
rect 4936 20644 4940 20700
rect 4876 20640 4940 20644
rect 4956 20700 5020 20704
rect 4956 20644 4960 20700
rect 4960 20644 5016 20700
rect 5016 20644 5020 20700
rect 4956 20640 5020 20644
rect 5036 20700 5100 20704
rect 5036 20644 5040 20700
rect 5040 20644 5096 20700
rect 5096 20644 5100 20700
rect 5036 20640 5100 20644
rect 5116 20700 5180 20704
rect 5116 20644 5120 20700
rect 5120 20644 5176 20700
rect 5176 20644 5180 20700
rect 5116 20640 5180 20644
rect 97036 20700 97100 20704
rect 97036 20644 97040 20700
rect 97040 20644 97096 20700
rect 97096 20644 97100 20700
rect 97036 20640 97100 20644
rect 97116 20700 97180 20704
rect 97116 20644 97120 20700
rect 97120 20644 97176 20700
rect 97176 20644 97180 20700
rect 97116 20640 97180 20644
rect 97196 20700 97260 20704
rect 97196 20644 97200 20700
rect 97200 20644 97256 20700
rect 97256 20644 97260 20700
rect 97196 20640 97260 20644
rect 97276 20700 97340 20704
rect 97276 20644 97280 20700
rect 97280 20644 97336 20700
rect 97336 20644 97340 20700
rect 97276 20640 97340 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 96376 20156 96440 20160
rect 96376 20100 96380 20156
rect 96380 20100 96436 20156
rect 96436 20100 96440 20156
rect 96376 20096 96440 20100
rect 96456 20156 96520 20160
rect 96456 20100 96460 20156
rect 96460 20100 96516 20156
rect 96516 20100 96520 20156
rect 96456 20096 96520 20100
rect 96536 20156 96600 20160
rect 96536 20100 96540 20156
rect 96540 20100 96596 20156
rect 96596 20100 96600 20156
rect 96536 20096 96600 20100
rect 96616 20156 96680 20160
rect 96616 20100 96620 20156
rect 96620 20100 96676 20156
rect 96676 20100 96680 20156
rect 96616 20096 96680 20100
rect 4876 19612 4940 19616
rect 4876 19556 4880 19612
rect 4880 19556 4936 19612
rect 4936 19556 4940 19612
rect 4876 19552 4940 19556
rect 4956 19612 5020 19616
rect 4956 19556 4960 19612
rect 4960 19556 5016 19612
rect 5016 19556 5020 19612
rect 4956 19552 5020 19556
rect 5036 19612 5100 19616
rect 5036 19556 5040 19612
rect 5040 19556 5096 19612
rect 5096 19556 5100 19612
rect 5036 19552 5100 19556
rect 5116 19612 5180 19616
rect 5116 19556 5120 19612
rect 5120 19556 5176 19612
rect 5176 19556 5180 19612
rect 5116 19552 5180 19556
rect 97036 19612 97100 19616
rect 97036 19556 97040 19612
rect 97040 19556 97096 19612
rect 97096 19556 97100 19612
rect 97036 19552 97100 19556
rect 97116 19612 97180 19616
rect 97116 19556 97120 19612
rect 97120 19556 97176 19612
rect 97176 19556 97180 19612
rect 97116 19552 97180 19556
rect 97196 19612 97260 19616
rect 97196 19556 97200 19612
rect 97200 19556 97256 19612
rect 97256 19556 97260 19612
rect 97196 19552 97260 19556
rect 97276 19612 97340 19616
rect 97276 19556 97280 19612
rect 97280 19556 97336 19612
rect 97336 19556 97340 19612
rect 97276 19552 97340 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 96376 19068 96440 19072
rect 96376 19012 96380 19068
rect 96380 19012 96436 19068
rect 96436 19012 96440 19068
rect 96376 19008 96440 19012
rect 96456 19068 96520 19072
rect 96456 19012 96460 19068
rect 96460 19012 96516 19068
rect 96516 19012 96520 19068
rect 96456 19008 96520 19012
rect 96536 19068 96600 19072
rect 96536 19012 96540 19068
rect 96540 19012 96596 19068
rect 96596 19012 96600 19068
rect 96536 19008 96600 19012
rect 96616 19068 96680 19072
rect 96616 19012 96620 19068
rect 96620 19012 96676 19068
rect 96676 19012 96680 19068
rect 96616 19008 96680 19012
rect 4876 18524 4940 18528
rect 4876 18468 4880 18524
rect 4880 18468 4936 18524
rect 4936 18468 4940 18524
rect 4876 18464 4940 18468
rect 4956 18524 5020 18528
rect 4956 18468 4960 18524
rect 4960 18468 5016 18524
rect 5016 18468 5020 18524
rect 4956 18464 5020 18468
rect 5036 18524 5100 18528
rect 5036 18468 5040 18524
rect 5040 18468 5096 18524
rect 5096 18468 5100 18524
rect 5036 18464 5100 18468
rect 5116 18524 5180 18528
rect 5116 18468 5120 18524
rect 5120 18468 5176 18524
rect 5176 18468 5180 18524
rect 5116 18464 5180 18468
rect 97036 18524 97100 18528
rect 97036 18468 97040 18524
rect 97040 18468 97096 18524
rect 97096 18468 97100 18524
rect 97036 18464 97100 18468
rect 97116 18524 97180 18528
rect 97116 18468 97120 18524
rect 97120 18468 97176 18524
rect 97176 18468 97180 18524
rect 97116 18464 97180 18468
rect 97196 18524 97260 18528
rect 97196 18468 97200 18524
rect 97200 18468 97256 18524
rect 97256 18468 97260 18524
rect 97196 18464 97260 18468
rect 97276 18524 97340 18528
rect 97276 18468 97280 18524
rect 97280 18468 97336 18524
rect 97336 18468 97340 18524
rect 97276 18464 97340 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 96376 17980 96440 17984
rect 96376 17924 96380 17980
rect 96380 17924 96436 17980
rect 96436 17924 96440 17980
rect 96376 17920 96440 17924
rect 96456 17980 96520 17984
rect 96456 17924 96460 17980
rect 96460 17924 96516 17980
rect 96516 17924 96520 17980
rect 96456 17920 96520 17924
rect 96536 17980 96600 17984
rect 96536 17924 96540 17980
rect 96540 17924 96596 17980
rect 96596 17924 96600 17980
rect 96536 17920 96600 17924
rect 96616 17980 96680 17984
rect 96616 17924 96620 17980
rect 96620 17924 96676 17980
rect 96676 17924 96680 17980
rect 96616 17920 96680 17924
rect 4876 17436 4940 17440
rect 4876 17380 4880 17436
rect 4880 17380 4936 17436
rect 4936 17380 4940 17436
rect 4876 17376 4940 17380
rect 4956 17436 5020 17440
rect 4956 17380 4960 17436
rect 4960 17380 5016 17436
rect 5016 17380 5020 17436
rect 4956 17376 5020 17380
rect 5036 17436 5100 17440
rect 5036 17380 5040 17436
rect 5040 17380 5096 17436
rect 5096 17380 5100 17436
rect 5036 17376 5100 17380
rect 5116 17436 5180 17440
rect 5116 17380 5120 17436
rect 5120 17380 5176 17436
rect 5176 17380 5180 17436
rect 5116 17376 5180 17380
rect 97036 17436 97100 17440
rect 97036 17380 97040 17436
rect 97040 17380 97096 17436
rect 97096 17380 97100 17436
rect 97036 17376 97100 17380
rect 97116 17436 97180 17440
rect 97116 17380 97120 17436
rect 97120 17380 97176 17436
rect 97176 17380 97180 17436
rect 97116 17376 97180 17380
rect 97196 17436 97260 17440
rect 97196 17380 97200 17436
rect 97200 17380 97256 17436
rect 97256 17380 97260 17436
rect 97196 17376 97260 17380
rect 97276 17436 97340 17440
rect 97276 17380 97280 17436
rect 97280 17380 97336 17436
rect 97336 17380 97340 17436
rect 97276 17376 97340 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 96376 16892 96440 16896
rect 96376 16836 96380 16892
rect 96380 16836 96436 16892
rect 96436 16836 96440 16892
rect 96376 16832 96440 16836
rect 96456 16892 96520 16896
rect 96456 16836 96460 16892
rect 96460 16836 96516 16892
rect 96516 16836 96520 16892
rect 96456 16832 96520 16836
rect 96536 16892 96600 16896
rect 96536 16836 96540 16892
rect 96540 16836 96596 16892
rect 96596 16836 96600 16892
rect 96536 16832 96600 16836
rect 96616 16892 96680 16896
rect 96616 16836 96620 16892
rect 96620 16836 96676 16892
rect 96676 16836 96680 16892
rect 96616 16832 96680 16836
rect 4876 16348 4940 16352
rect 4876 16292 4880 16348
rect 4880 16292 4936 16348
rect 4936 16292 4940 16348
rect 4876 16288 4940 16292
rect 4956 16348 5020 16352
rect 4956 16292 4960 16348
rect 4960 16292 5016 16348
rect 5016 16292 5020 16348
rect 4956 16288 5020 16292
rect 5036 16348 5100 16352
rect 5036 16292 5040 16348
rect 5040 16292 5096 16348
rect 5096 16292 5100 16348
rect 5036 16288 5100 16292
rect 5116 16348 5180 16352
rect 5116 16292 5120 16348
rect 5120 16292 5176 16348
rect 5176 16292 5180 16348
rect 5116 16288 5180 16292
rect 97036 16348 97100 16352
rect 97036 16292 97040 16348
rect 97040 16292 97096 16348
rect 97096 16292 97100 16348
rect 97036 16288 97100 16292
rect 97116 16348 97180 16352
rect 97116 16292 97120 16348
rect 97120 16292 97176 16348
rect 97176 16292 97180 16348
rect 97116 16288 97180 16292
rect 97196 16348 97260 16352
rect 97196 16292 97200 16348
rect 97200 16292 97256 16348
rect 97256 16292 97260 16348
rect 97196 16288 97260 16292
rect 97276 16348 97340 16352
rect 97276 16292 97280 16348
rect 97280 16292 97336 16348
rect 97336 16292 97340 16348
rect 97276 16288 97340 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 96376 15804 96440 15808
rect 96376 15748 96380 15804
rect 96380 15748 96436 15804
rect 96436 15748 96440 15804
rect 96376 15744 96440 15748
rect 96456 15804 96520 15808
rect 96456 15748 96460 15804
rect 96460 15748 96516 15804
rect 96516 15748 96520 15804
rect 96456 15744 96520 15748
rect 96536 15804 96600 15808
rect 96536 15748 96540 15804
rect 96540 15748 96596 15804
rect 96596 15748 96600 15804
rect 96536 15744 96600 15748
rect 96616 15804 96680 15808
rect 96616 15748 96620 15804
rect 96620 15748 96676 15804
rect 96676 15748 96680 15804
rect 96616 15744 96680 15748
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 97036 15260 97100 15264
rect 97036 15204 97040 15260
rect 97040 15204 97096 15260
rect 97096 15204 97100 15260
rect 97036 15200 97100 15204
rect 97116 15260 97180 15264
rect 97116 15204 97120 15260
rect 97120 15204 97176 15260
rect 97176 15204 97180 15260
rect 97116 15200 97180 15204
rect 97196 15260 97260 15264
rect 97196 15204 97200 15260
rect 97200 15204 97256 15260
rect 97256 15204 97260 15260
rect 97196 15200 97260 15204
rect 97276 15260 97340 15264
rect 97276 15204 97280 15260
rect 97280 15204 97336 15260
rect 97336 15204 97340 15260
rect 97276 15200 97340 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 96376 14716 96440 14720
rect 96376 14660 96380 14716
rect 96380 14660 96436 14716
rect 96436 14660 96440 14716
rect 96376 14656 96440 14660
rect 96456 14716 96520 14720
rect 96456 14660 96460 14716
rect 96460 14660 96516 14716
rect 96516 14660 96520 14716
rect 96456 14656 96520 14660
rect 96536 14716 96600 14720
rect 96536 14660 96540 14716
rect 96540 14660 96596 14716
rect 96596 14660 96600 14716
rect 96536 14656 96600 14660
rect 96616 14716 96680 14720
rect 96616 14660 96620 14716
rect 96620 14660 96676 14716
rect 96676 14660 96680 14716
rect 96616 14656 96680 14660
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 97036 14172 97100 14176
rect 97036 14116 97040 14172
rect 97040 14116 97096 14172
rect 97096 14116 97100 14172
rect 97036 14112 97100 14116
rect 97116 14172 97180 14176
rect 97116 14116 97120 14172
rect 97120 14116 97176 14172
rect 97176 14116 97180 14172
rect 97116 14112 97180 14116
rect 97196 14172 97260 14176
rect 97196 14116 97200 14172
rect 97200 14116 97256 14172
rect 97256 14116 97260 14172
rect 97196 14112 97260 14116
rect 97276 14172 97340 14176
rect 97276 14116 97280 14172
rect 97280 14116 97336 14172
rect 97336 14116 97340 14172
rect 97276 14112 97340 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 96376 13628 96440 13632
rect 96376 13572 96380 13628
rect 96380 13572 96436 13628
rect 96436 13572 96440 13628
rect 96376 13568 96440 13572
rect 96456 13628 96520 13632
rect 96456 13572 96460 13628
rect 96460 13572 96516 13628
rect 96516 13572 96520 13628
rect 96456 13568 96520 13572
rect 96536 13628 96600 13632
rect 96536 13572 96540 13628
rect 96540 13572 96596 13628
rect 96596 13572 96600 13628
rect 96536 13568 96600 13572
rect 96616 13628 96680 13632
rect 96616 13572 96620 13628
rect 96620 13572 96676 13628
rect 96676 13572 96680 13628
rect 96616 13568 96680 13572
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 97036 13084 97100 13088
rect 97036 13028 97040 13084
rect 97040 13028 97096 13084
rect 97096 13028 97100 13084
rect 97036 13024 97100 13028
rect 97116 13084 97180 13088
rect 97116 13028 97120 13084
rect 97120 13028 97176 13084
rect 97176 13028 97180 13084
rect 97116 13024 97180 13028
rect 97196 13084 97260 13088
rect 97196 13028 97200 13084
rect 97200 13028 97256 13084
rect 97256 13028 97260 13084
rect 97196 13024 97260 13028
rect 97276 13084 97340 13088
rect 97276 13028 97280 13084
rect 97280 13028 97336 13084
rect 97336 13028 97340 13084
rect 97276 13024 97340 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 96376 12540 96440 12544
rect 96376 12484 96380 12540
rect 96380 12484 96436 12540
rect 96436 12484 96440 12540
rect 96376 12480 96440 12484
rect 96456 12540 96520 12544
rect 96456 12484 96460 12540
rect 96460 12484 96516 12540
rect 96516 12484 96520 12540
rect 96456 12480 96520 12484
rect 96536 12540 96600 12544
rect 96536 12484 96540 12540
rect 96540 12484 96596 12540
rect 96596 12484 96600 12540
rect 96536 12480 96600 12484
rect 96616 12540 96680 12544
rect 96616 12484 96620 12540
rect 96620 12484 96676 12540
rect 96676 12484 96680 12540
rect 96616 12480 96680 12484
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 97036 11996 97100 12000
rect 97036 11940 97040 11996
rect 97040 11940 97096 11996
rect 97096 11940 97100 11996
rect 97036 11936 97100 11940
rect 97116 11996 97180 12000
rect 97116 11940 97120 11996
rect 97120 11940 97176 11996
rect 97176 11940 97180 11996
rect 97116 11936 97180 11940
rect 97196 11996 97260 12000
rect 97196 11940 97200 11996
rect 97200 11940 97256 11996
rect 97256 11940 97260 11996
rect 97196 11936 97260 11940
rect 97276 11996 97340 12000
rect 97276 11940 97280 11996
rect 97280 11940 97336 11996
rect 97336 11940 97340 11996
rect 97276 11936 97340 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 96376 11452 96440 11456
rect 96376 11396 96380 11452
rect 96380 11396 96436 11452
rect 96436 11396 96440 11452
rect 96376 11392 96440 11396
rect 96456 11452 96520 11456
rect 96456 11396 96460 11452
rect 96460 11396 96516 11452
rect 96516 11396 96520 11452
rect 96456 11392 96520 11396
rect 96536 11452 96600 11456
rect 96536 11396 96540 11452
rect 96540 11396 96596 11452
rect 96596 11396 96600 11452
rect 96536 11392 96600 11396
rect 96616 11452 96680 11456
rect 96616 11396 96620 11452
rect 96620 11396 96676 11452
rect 96676 11396 96680 11452
rect 96616 11392 96680 11396
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 97036 10908 97100 10912
rect 97036 10852 97040 10908
rect 97040 10852 97096 10908
rect 97096 10852 97100 10908
rect 97036 10848 97100 10852
rect 97116 10908 97180 10912
rect 97116 10852 97120 10908
rect 97120 10852 97176 10908
rect 97176 10852 97180 10908
rect 97116 10848 97180 10852
rect 97196 10908 97260 10912
rect 97196 10852 97200 10908
rect 97200 10852 97256 10908
rect 97256 10852 97260 10908
rect 97196 10848 97260 10852
rect 97276 10908 97340 10912
rect 97276 10852 97280 10908
rect 97280 10852 97336 10908
rect 97336 10852 97340 10908
rect 97276 10848 97340 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 96376 10364 96440 10368
rect 96376 10308 96380 10364
rect 96380 10308 96436 10364
rect 96436 10308 96440 10364
rect 96376 10304 96440 10308
rect 96456 10364 96520 10368
rect 96456 10308 96460 10364
rect 96460 10308 96516 10364
rect 96516 10308 96520 10364
rect 96456 10304 96520 10308
rect 96536 10364 96600 10368
rect 96536 10308 96540 10364
rect 96540 10308 96596 10364
rect 96596 10308 96600 10364
rect 96536 10304 96600 10308
rect 96616 10364 96680 10368
rect 96616 10308 96620 10364
rect 96620 10308 96676 10364
rect 96676 10308 96680 10364
rect 96616 10304 96680 10308
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 97036 9820 97100 9824
rect 97036 9764 97040 9820
rect 97040 9764 97096 9820
rect 97096 9764 97100 9820
rect 97036 9760 97100 9764
rect 97116 9820 97180 9824
rect 97116 9764 97120 9820
rect 97120 9764 97176 9820
rect 97176 9764 97180 9820
rect 97116 9760 97180 9764
rect 97196 9820 97260 9824
rect 97196 9764 97200 9820
rect 97200 9764 97256 9820
rect 97256 9764 97260 9820
rect 97196 9760 97260 9764
rect 97276 9820 97340 9824
rect 97276 9764 97280 9820
rect 97280 9764 97336 9820
rect 97336 9764 97340 9820
rect 97276 9760 97340 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 96376 9276 96440 9280
rect 96376 9220 96380 9276
rect 96380 9220 96436 9276
rect 96436 9220 96440 9276
rect 96376 9216 96440 9220
rect 96456 9276 96520 9280
rect 96456 9220 96460 9276
rect 96460 9220 96516 9276
rect 96516 9220 96520 9276
rect 96456 9216 96520 9220
rect 96536 9276 96600 9280
rect 96536 9220 96540 9276
rect 96540 9220 96596 9276
rect 96596 9220 96600 9276
rect 96536 9216 96600 9220
rect 96616 9276 96680 9280
rect 96616 9220 96620 9276
rect 96620 9220 96676 9276
rect 96676 9220 96680 9276
rect 96616 9216 96680 9220
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 97036 8732 97100 8736
rect 97036 8676 97040 8732
rect 97040 8676 97096 8732
rect 97096 8676 97100 8732
rect 97036 8672 97100 8676
rect 97116 8732 97180 8736
rect 97116 8676 97120 8732
rect 97120 8676 97176 8732
rect 97176 8676 97180 8732
rect 97116 8672 97180 8676
rect 97196 8732 97260 8736
rect 97196 8676 97200 8732
rect 97200 8676 97256 8732
rect 97256 8676 97260 8732
rect 97196 8672 97260 8676
rect 97276 8732 97340 8736
rect 97276 8676 97280 8732
rect 97280 8676 97336 8732
rect 97336 8676 97340 8732
rect 97276 8672 97340 8676
rect 50844 8664 50908 8668
rect 50844 8608 50848 8664
rect 50848 8608 50904 8664
rect 50904 8608 50908 8664
rect 50844 8604 50908 8608
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 96376 8188 96440 8192
rect 96376 8132 96380 8188
rect 96380 8132 96436 8188
rect 96436 8132 96440 8188
rect 96376 8128 96440 8132
rect 96456 8188 96520 8192
rect 96456 8132 96460 8188
rect 96460 8132 96516 8188
rect 96516 8132 96520 8188
rect 96456 8128 96520 8132
rect 96536 8188 96600 8192
rect 96536 8132 96540 8188
rect 96540 8132 96596 8188
rect 96596 8132 96600 8188
rect 96536 8128 96600 8132
rect 96616 8188 96680 8192
rect 96616 8132 96620 8188
rect 96620 8132 96676 8188
rect 96676 8132 96680 8188
rect 96616 8128 96680 8132
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 97036 7644 97100 7648
rect 97036 7588 97040 7644
rect 97040 7588 97096 7644
rect 97096 7588 97100 7644
rect 97036 7584 97100 7588
rect 97116 7644 97180 7648
rect 97116 7588 97120 7644
rect 97120 7588 97176 7644
rect 97176 7588 97180 7644
rect 97116 7584 97180 7588
rect 97196 7644 97260 7648
rect 97196 7588 97200 7644
rect 97200 7588 97256 7644
rect 97256 7588 97260 7644
rect 97196 7584 97260 7588
rect 97276 7644 97340 7648
rect 97276 7588 97280 7644
rect 97280 7588 97336 7644
rect 97336 7588 97340 7644
rect 97276 7584 97340 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 96376 7100 96440 7104
rect 96376 7044 96380 7100
rect 96380 7044 96436 7100
rect 96436 7044 96440 7100
rect 96376 7040 96440 7044
rect 96456 7100 96520 7104
rect 96456 7044 96460 7100
rect 96460 7044 96516 7100
rect 96516 7044 96520 7100
rect 96456 7040 96520 7044
rect 96536 7100 96600 7104
rect 96536 7044 96540 7100
rect 96540 7044 96596 7100
rect 96596 7044 96600 7100
rect 96536 7040 96600 7044
rect 96616 7100 96680 7104
rect 96616 7044 96620 7100
rect 96620 7044 96676 7100
rect 96676 7044 96680 7100
rect 96616 7040 96680 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 97036 6556 97100 6560
rect 97036 6500 97040 6556
rect 97040 6500 97096 6556
rect 97096 6500 97100 6556
rect 97036 6496 97100 6500
rect 97116 6556 97180 6560
rect 97116 6500 97120 6556
rect 97120 6500 97176 6556
rect 97176 6500 97180 6556
rect 97116 6496 97180 6500
rect 97196 6556 97260 6560
rect 97196 6500 97200 6556
rect 97200 6500 97256 6556
rect 97256 6500 97260 6556
rect 97196 6496 97260 6500
rect 97276 6556 97340 6560
rect 97276 6500 97280 6556
rect 97280 6500 97336 6556
rect 97336 6500 97340 6556
rect 97276 6496 97340 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 65656 6012 65720 6016
rect 65656 5956 65660 6012
rect 65660 5956 65716 6012
rect 65716 5956 65720 6012
rect 65656 5952 65720 5956
rect 65736 6012 65800 6016
rect 65736 5956 65740 6012
rect 65740 5956 65796 6012
rect 65796 5956 65800 6012
rect 65736 5952 65800 5956
rect 65816 6012 65880 6016
rect 65816 5956 65820 6012
rect 65820 5956 65876 6012
rect 65876 5956 65880 6012
rect 65816 5952 65880 5956
rect 65896 6012 65960 6016
rect 65896 5956 65900 6012
rect 65900 5956 65956 6012
rect 65956 5956 65960 6012
rect 65896 5952 65960 5956
rect 96376 6012 96440 6016
rect 96376 5956 96380 6012
rect 96380 5956 96436 6012
rect 96436 5956 96440 6012
rect 96376 5952 96440 5956
rect 96456 6012 96520 6016
rect 96456 5956 96460 6012
rect 96460 5956 96516 6012
rect 96516 5956 96520 6012
rect 96456 5952 96520 5956
rect 96536 6012 96600 6016
rect 96536 5956 96540 6012
rect 96540 5956 96596 6012
rect 96596 5956 96600 6012
rect 96536 5952 96600 5956
rect 96616 6012 96680 6016
rect 96616 5956 96620 6012
rect 96620 5956 96676 6012
rect 96676 5956 96680 6012
rect 96616 5952 96680 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 35596 5468 35660 5472
rect 35596 5412 35600 5468
rect 35600 5412 35656 5468
rect 35656 5412 35660 5468
rect 35596 5408 35660 5412
rect 35676 5468 35740 5472
rect 35676 5412 35680 5468
rect 35680 5412 35736 5468
rect 35736 5412 35740 5468
rect 35676 5408 35740 5412
rect 35756 5468 35820 5472
rect 35756 5412 35760 5468
rect 35760 5412 35816 5468
rect 35816 5412 35820 5468
rect 35756 5408 35820 5412
rect 35836 5468 35900 5472
rect 35836 5412 35840 5468
rect 35840 5412 35896 5468
rect 35896 5412 35900 5468
rect 35836 5408 35900 5412
rect 66316 5468 66380 5472
rect 66316 5412 66320 5468
rect 66320 5412 66376 5468
rect 66376 5412 66380 5468
rect 66316 5408 66380 5412
rect 66396 5468 66460 5472
rect 66396 5412 66400 5468
rect 66400 5412 66456 5468
rect 66456 5412 66460 5468
rect 66396 5408 66460 5412
rect 66476 5468 66540 5472
rect 66476 5412 66480 5468
rect 66480 5412 66536 5468
rect 66536 5412 66540 5468
rect 66476 5408 66540 5412
rect 66556 5468 66620 5472
rect 66556 5412 66560 5468
rect 66560 5412 66616 5468
rect 66616 5412 66620 5468
rect 66556 5408 66620 5412
rect 97036 5468 97100 5472
rect 97036 5412 97040 5468
rect 97040 5412 97096 5468
rect 97096 5412 97100 5468
rect 97036 5408 97100 5412
rect 97116 5468 97180 5472
rect 97116 5412 97120 5468
rect 97120 5412 97176 5468
rect 97176 5412 97180 5468
rect 97116 5408 97180 5412
rect 97196 5468 97260 5472
rect 97196 5412 97200 5468
rect 97200 5412 97256 5468
rect 97256 5412 97260 5468
rect 97196 5408 97260 5412
rect 97276 5468 97340 5472
rect 97276 5412 97280 5468
rect 97280 5412 97336 5468
rect 97336 5412 97340 5468
rect 97276 5408 97340 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 65656 4924 65720 4928
rect 65656 4868 65660 4924
rect 65660 4868 65716 4924
rect 65716 4868 65720 4924
rect 65656 4864 65720 4868
rect 65736 4924 65800 4928
rect 65736 4868 65740 4924
rect 65740 4868 65796 4924
rect 65796 4868 65800 4924
rect 65736 4864 65800 4868
rect 65816 4924 65880 4928
rect 65816 4868 65820 4924
rect 65820 4868 65876 4924
rect 65876 4868 65880 4924
rect 65816 4864 65880 4868
rect 65896 4924 65960 4928
rect 65896 4868 65900 4924
rect 65900 4868 65956 4924
rect 65956 4868 65960 4924
rect 65896 4864 65960 4868
rect 96376 4924 96440 4928
rect 96376 4868 96380 4924
rect 96380 4868 96436 4924
rect 96436 4868 96440 4924
rect 96376 4864 96440 4868
rect 96456 4924 96520 4928
rect 96456 4868 96460 4924
rect 96460 4868 96516 4924
rect 96516 4868 96520 4924
rect 96456 4864 96520 4868
rect 96536 4924 96600 4928
rect 96536 4868 96540 4924
rect 96540 4868 96596 4924
rect 96596 4868 96600 4924
rect 96536 4864 96600 4868
rect 96616 4924 96680 4928
rect 96616 4868 96620 4924
rect 96620 4868 96676 4924
rect 96676 4868 96680 4924
rect 96616 4864 96680 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 35596 4380 35660 4384
rect 35596 4324 35600 4380
rect 35600 4324 35656 4380
rect 35656 4324 35660 4380
rect 35596 4320 35660 4324
rect 35676 4380 35740 4384
rect 35676 4324 35680 4380
rect 35680 4324 35736 4380
rect 35736 4324 35740 4380
rect 35676 4320 35740 4324
rect 35756 4380 35820 4384
rect 35756 4324 35760 4380
rect 35760 4324 35816 4380
rect 35816 4324 35820 4380
rect 35756 4320 35820 4324
rect 35836 4380 35900 4384
rect 35836 4324 35840 4380
rect 35840 4324 35896 4380
rect 35896 4324 35900 4380
rect 35836 4320 35900 4324
rect 66316 4380 66380 4384
rect 66316 4324 66320 4380
rect 66320 4324 66376 4380
rect 66376 4324 66380 4380
rect 66316 4320 66380 4324
rect 66396 4380 66460 4384
rect 66396 4324 66400 4380
rect 66400 4324 66456 4380
rect 66456 4324 66460 4380
rect 66396 4320 66460 4324
rect 66476 4380 66540 4384
rect 66476 4324 66480 4380
rect 66480 4324 66536 4380
rect 66536 4324 66540 4380
rect 66476 4320 66540 4324
rect 66556 4380 66620 4384
rect 66556 4324 66560 4380
rect 66560 4324 66616 4380
rect 66616 4324 66620 4380
rect 66556 4320 66620 4324
rect 97036 4380 97100 4384
rect 97036 4324 97040 4380
rect 97040 4324 97096 4380
rect 97096 4324 97100 4380
rect 97036 4320 97100 4324
rect 97116 4380 97180 4384
rect 97116 4324 97120 4380
rect 97120 4324 97176 4380
rect 97176 4324 97180 4380
rect 97116 4320 97180 4324
rect 97196 4380 97260 4384
rect 97196 4324 97200 4380
rect 97200 4324 97256 4380
rect 97256 4324 97260 4380
rect 97196 4320 97260 4324
rect 97276 4380 97340 4384
rect 97276 4324 97280 4380
rect 97280 4324 97336 4380
rect 97336 4324 97340 4380
rect 97276 4320 97340 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 65656 3836 65720 3840
rect 65656 3780 65660 3836
rect 65660 3780 65716 3836
rect 65716 3780 65720 3836
rect 65656 3776 65720 3780
rect 65736 3836 65800 3840
rect 65736 3780 65740 3836
rect 65740 3780 65796 3836
rect 65796 3780 65800 3836
rect 65736 3776 65800 3780
rect 65816 3836 65880 3840
rect 65816 3780 65820 3836
rect 65820 3780 65876 3836
rect 65876 3780 65880 3836
rect 65816 3776 65880 3780
rect 65896 3836 65960 3840
rect 65896 3780 65900 3836
rect 65900 3780 65956 3836
rect 65956 3780 65960 3836
rect 65896 3776 65960 3780
rect 96376 3836 96440 3840
rect 96376 3780 96380 3836
rect 96380 3780 96436 3836
rect 96436 3780 96440 3836
rect 96376 3776 96440 3780
rect 96456 3836 96520 3840
rect 96456 3780 96460 3836
rect 96460 3780 96516 3836
rect 96516 3780 96520 3836
rect 96456 3776 96520 3780
rect 96536 3836 96600 3840
rect 96536 3780 96540 3836
rect 96540 3780 96596 3836
rect 96596 3780 96600 3836
rect 96536 3776 96600 3780
rect 96616 3836 96680 3840
rect 96616 3780 96620 3836
rect 96620 3780 96676 3836
rect 96676 3780 96680 3836
rect 96616 3776 96680 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 35596 3292 35660 3296
rect 35596 3236 35600 3292
rect 35600 3236 35656 3292
rect 35656 3236 35660 3292
rect 35596 3232 35660 3236
rect 35676 3292 35740 3296
rect 35676 3236 35680 3292
rect 35680 3236 35736 3292
rect 35736 3236 35740 3292
rect 35676 3232 35740 3236
rect 35756 3292 35820 3296
rect 35756 3236 35760 3292
rect 35760 3236 35816 3292
rect 35816 3236 35820 3292
rect 35756 3232 35820 3236
rect 35836 3292 35900 3296
rect 35836 3236 35840 3292
rect 35840 3236 35896 3292
rect 35896 3236 35900 3292
rect 35836 3232 35900 3236
rect 66316 3292 66380 3296
rect 66316 3236 66320 3292
rect 66320 3236 66376 3292
rect 66376 3236 66380 3292
rect 66316 3232 66380 3236
rect 66396 3292 66460 3296
rect 66396 3236 66400 3292
rect 66400 3236 66456 3292
rect 66456 3236 66460 3292
rect 66396 3232 66460 3236
rect 66476 3292 66540 3296
rect 66476 3236 66480 3292
rect 66480 3236 66536 3292
rect 66536 3236 66540 3292
rect 66476 3232 66540 3236
rect 66556 3292 66620 3296
rect 66556 3236 66560 3292
rect 66560 3236 66616 3292
rect 66616 3236 66620 3292
rect 66556 3232 66620 3236
rect 97036 3292 97100 3296
rect 97036 3236 97040 3292
rect 97040 3236 97096 3292
rect 97096 3236 97100 3292
rect 97036 3232 97100 3236
rect 97116 3292 97180 3296
rect 97116 3236 97120 3292
rect 97120 3236 97176 3292
rect 97176 3236 97180 3292
rect 97116 3232 97180 3236
rect 97196 3292 97260 3296
rect 97196 3236 97200 3292
rect 97200 3236 97256 3292
rect 97256 3236 97260 3292
rect 97196 3232 97260 3236
rect 97276 3292 97340 3296
rect 97276 3236 97280 3292
rect 97280 3236 97336 3292
rect 97336 3236 97340 3292
rect 97276 3232 97340 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 65656 2748 65720 2752
rect 65656 2692 65660 2748
rect 65660 2692 65716 2748
rect 65716 2692 65720 2748
rect 65656 2688 65720 2692
rect 65736 2748 65800 2752
rect 65736 2692 65740 2748
rect 65740 2692 65796 2748
rect 65796 2692 65800 2748
rect 65736 2688 65800 2692
rect 65816 2748 65880 2752
rect 65816 2692 65820 2748
rect 65820 2692 65876 2748
rect 65876 2692 65880 2748
rect 65816 2688 65880 2692
rect 65896 2748 65960 2752
rect 65896 2692 65900 2748
rect 65900 2692 65956 2748
rect 65956 2692 65960 2748
rect 65896 2688 65960 2692
rect 96376 2748 96440 2752
rect 96376 2692 96380 2748
rect 96380 2692 96436 2748
rect 96436 2692 96440 2748
rect 96376 2688 96440 2692
rect 96456 2748 96520 2752
rect 96456 2692 96460 2748
rect 96460 2692 96516 2748
rect 96516 2692 96520 2748
rect 96456 2688 96520 2692
rect 96536 2748 96600 2752
rect 96536 2692 96540 2748
rect 96540 2692 96596 2748
rect 96596 2692 96600 2748
rect 96536 2688 96600 2692
rect 96616 2748 96680 2752
rect 96616 2692 96620 2748
rect 96620 2692 96676 2748
rect 96676 2692 96680 2748
rect 96616 2688 96680 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
rect 35596 2204 35660 2208
rect 35596 2148 35600 2204
rect 35600 2148 35656 2204
rect 35656 2148 35660 2204
rect 35596 2144 35660 2148
rect 35676 2204 35740 2208
rect 35676 2148 35680 2204
rect 35680 2148 35736 2204
rect 35736 2148 35740 2204
rect 35676 2144 35740 2148
rect 35756 2204 35820 2208
rect 35756 2148 35760 2204
rect 35760 2148 35816 2204
rect 35816 2148 35820 2204
rect 35756 2144 35820 2148
rect 35836 2204 35900 2208
rect 35836 2148 35840 2204
rect 35840 2148 35896 2204
rect 35896 2148 35900 2204
rect 35836 2144 35900 2148
rect 66316 2204 66380 2208
rect 66316 2148 66320 2204
rect 66320 2148 66376 2204
rect 66376 2148 66380 2204
rect 66316 2144 66380 2148
rect 66396 2204 66460 2208
rect 66396 2148 66400 2204
rect 66400 2148 66456 2204
rect 66456 2148 66460 2204
rect 66396 2144 66460 2148
rect 66476 2204 66540 2208
rect 66476 2148 66480 2204
rect 66480 2148 66536 2204
rect 66536 2148 66540 2204
rect 66476 2144 66540 2148
rect 66556 2204 66620 2208
rect 66556 2148 66560 2204
rect 66560 2148 66616 2204
rect 66616 2148 66620 2204
rect 66556 2144 66620 2148
rect 97036 2204 97100 2208
rect 97036 2148 97040 2204
rect 97040 2148 97096 2204
rect 97096 2148 97100 2204
rect 97036 2144 97100 2148
rect 97116 2204 97180 2208
rect 97116 2148 97120 2204
rect 97120 2148 97176 2204
rect 97176 2148 97180 2204
rect 97116 2144 97180 2148
rect 97196 2204 97260 2208
rect 97196 2148 97200 2204
rect 97200 2148 97256 2204
rect 97256 2148 97260 2204
rect 97196 2144 97260 2148
rect 97276 2204 97340 2208
rect 97276 2148 97280 2204
rect 97280 2148 97336 2204
rect 97336 2148 97340 2204
rect 97276 2144 97340 2148
<< metal4 >>
rect -1076 97882 -756 97924
rect -1076 97646 -1034 97882
rect -798 97646 -756 97882
rect -1076 67556 -756 97646
rect -1076 67320 -1034 67556
rect -798 67320 -756 67556
rect -1076 36920 -756 67320
rect -1076 36684 -1034 36920
rect -798 36684 -756 36920
rect -1076 6284 -756 36684
rect -1076 6048 -1034 6284
rect -798 6048 -756 6284
rect -1076 274 -756 6048
rect -416 97222 -96 97264
rect -416 96986 -374 97222
rect -138 96986 -96 97222
rect -416 66896 -96 96986
rect -416 66660 -374 66896
rect -138 66660 -96 66896
rect -416 36260 -96 66660
rect -416 36024 -374 36260
rect -138 36024 -96 36260
rect -416 5624 -96 36024
rect -416 5388 -374 5624
rect -138 5388 -96 5624
rect -416 934 -96 5388
rect -416 698 -374 934
rect -138 698 -96 934
rect -416 656 -96 698
rect 4208 97222 4528 97924
rect 4208 96986 4250 97222
rect 4486 96986 4528 97222
rect 4208 95232 4528 96986
rect 4208 95168 4216 95232
rect 4280 95168 4296 95232
rect 4360 95168 4376 95232
rect 4440 95168 4456 95232
rect 4520 95168 4528 95232
rect 4208 94144 4528 95168
rect 4208 94080 4216 94144
rect 4280 94080 4296 94144
rect 4360 94080 4376 94144
rect 4440 94080 4456 94144
rect 4520 94080 4528 94144
rect 4208 93056 4528 94080
rect 4208 92992 4216 93056
rect 4280 92992 4296 93056
rect 4360 92992 4376 93056
rect 4440 92992 4456 93056
rect 4520 92992 4528 93056
rect 4208 91968 4528 92992
rect 4208 91904 4216 91968
rect 4280 91904 4296 91968
rect 4360 91904 4376 91968
rect 4440 91904 4456 91968
rect 4520 91904 4528 91968
rect 4208 90880 4528 91904
rect 4208 90816 4216 90880
rect 4280 90816 4296 90880
rect 4360 90816 4376 90880
rect 4440 90816 4456 90880
rect 4520 90816 4528 90880
rect 4208 89792 4528 90816
rect 4208 89728 4216 89792
rect 4280 89728 4296 89792
rect 4360 89728 4376 89792
rect 4440 89728 4456 89792
rect 4520 89728 4528 89792
rect 4208 88704 4528 89728
rect 4208 88640 4216 88704
rect 4280 88640 4296 88704
rect 4360 88640 4376 88704
rect 4440 88640 4456 88704
rect 4520 88640 4528 88704
rect 4208 87616 4528 88640
rect 4208 87552 4216 87616
rect 4280 87552 4296 87616
rect 4360 87552 4376 87616
rect 4440 87552 4456 87616
rect 4520 87552 4528 87616
rect 4208 86528 4528 87552
rect 4208 86464 4216 86528
rect 4280 86464 4296 86528
rect 4360 86464 4376 86528
rect 4440 86464 4456 86528
rect 4520 86464 4528 86528
rect 4208 85440 4528 86464
rect 4208 85376 4216 85440
rect 4280 85376 4296 85440
rect 4360 85376 4376 85440
rect 4440 85376 4456 85440
rect 4520 85376 4528 85440
rect 4208 84352 4528 85376
rect 4208 84288 4216 84352
rect 4280 84288 4296 84352
rect 4360 84288 4376 84352
rect 4440 84288 4456 84352
rect 4520 84288 4528 84352
rect 4208 83264 4528 84288
rect 4208 83200 4216 83264
rect 4280 83200 4296 83264
rect 4360 83200 4376 83264
rect 4440 83200 4456 83264
rect 4520 83200 4528 83264
rect 4208 82176 4528 83200
rect 4208 82112 4216 82176
rect 4280 82112 4296 82176
rect 4360 82112 4376 82176
rect 4440 82112 4456 82176
rect 4520 82112 4528 82176
rect 4208 81088 4528 82112
rect 4208 81024 4216 81088
rect 4280 81024 4296 81088
rect 4360 81024 4376 81088
rect 4440 81024 4456 81088
rect 4520 81024 4528 81088
rect 4208 80000 4528 81024
rect 4208 79936 4216 80000
rect 4280 79936 4296 80000
rect 4360 79936 4376 80000
rect 4440 79936 4456 80000
rect 4520 79936 4528 80000
rect 4208 78912 4528 79936
rect 4208 78848 4216 78912
rect 4280 78848 4296 78912
rect 4360 78848 4376 78912
rect 4440 78848 4456 78912
rect 4520 78848 4528 78912
rect 4208 77824 4528 78848
rect 4208 77760 4216 77824
rect 4280 77760 4296 77824
rect 4360 77760 4376 77824
rect 4440 77760 4456 77824
rect 4520 77760 4528 77824
rect 4208 76736 4528 77760
rect 4208 76672 4216 76736
rect 4280 76672 4296 76736
rect 4360 76672 4376 76736
rect 4440 76672 4456 76736
rect 4520 76672 4528 76736
rect 4208 75648 4528 76672
rect 4208 75584 4216 75648
rect 4280 75584 4296 75648
rect 4360 75584 4376 75648
rect 4440 75584 4456 75648
rect 4520 75584 4528 75648
rect 4208 74560 4528 75584
rect 4208 74496 4216 74560
rect 4280 74496 4296 74560
rect 4360 74496 4376 74560
rect 4440 74496 4456 74560
rect 4520 74496 4528 74560
rect 4208 73472 4528 74496
rect 4208 73408 4216 73472
rect 4280 73408 4296 73472
rect 4360 73408 4376 73472
rect 4440 73408 4456 73472
rect 4520 73408 4528 73472
rect 4208 72384 4528 73408
rect 4208 72320 4216 72384
rect 4280 72320 4296 72384
rect 4360 72320 4376 72384
rect 4440 72320 4456 72384
rect 4520 72320 4528 72384
rect 4208 71296 4528 72320
rect 4208 71232 4216 71296
rect 4280 71232 4296 71296
rect 4360 71232 4376 71296
rect 4440 71232 4456 71296
rect 4520 71232 4528 71296
rect 4208 70208 4528 71232
rect 4208 70144 4216 70208
rect 4280 70144 4296 70208
rect 4360 70144 4376 70208
rect 4440 70144 4456 70208
rect 4520 70144 4528 70208
rect 4208 69120 4528 70144
rect 4208 69056 4216 69120
rect 4280 69056 4296 69120
rect 4360 69056 4376 69120
rect 4440 69056 4456 69120
rect 4520 69056 4528 69120
rect 4208 68032 4528 69056
rect 4208 67968 4216 68032
rect 4280 67968 4296 68032
rect 4360 67968 4376 68032
rect 4440 67968 4456 68032
rect 4520 67968 4528 68032
rect 4208 66944 4528 67968
rect 4208 66880 4216 66944
rect 4280 66896 4296 66944
rect 4360 66896 4376 66944
rect 4440 66896 4456 66944
rect 4520 66880 4528 66944
rect 4208 66660 4250 66880
rect 4486 66660 4528 66880
rect 4208 65856 4528 66660
rect 4208 65792 4216 65856
rect 4280 65792 4296 65856
rect 4360 65792 4376 65856
rect 4440 65792 4456 65856
rect 4520 65792 4528 65856
rect 4208 64768 4528 65792
rect 4208 64704 4216 64768
rect 4280 64704 4296 64768
rect 4360 64704 4376 64768
rect 4440 64704 4456 64768
rect 4520 64704 4528 64768
rect 4208 63680 4528 64704
rect 4208 63616 4216 63680
rect 4280 63616 4296 63680
rect 4360 63616 4376 63680
rect 4440 63616 4456 63680
rect 4520 63616 4528 63680
rect 4208 62592 4528 63616
rect 4208 62528 4216 62592
rect 4280 62528 4296 62592
rect 4360 62528 4376 62592
rect 4440 62528 4456 62592
rect 4520 62528 4528 62592
rect 4208 61504 4528 62528
rect 4208 61440 4216 61504
rect 4280 61440 4296 61504
rect 4360 61440 4376 61504
rect 4440 61440 4456 61504
rect 4520 61440 4528 61504
rect 4208 60416 4528 61440
rect 4208 60352 4216 60416
rect 4280 60352 4296 60416
rect 4360 60352 4376 60416
rect 4440 60352 4456 60416
rect 4520 60352 4528 60416
rect 4208 59328 4528 60352
rect 4208 59264 4216 59328
rect 4280 59264 4296 59328
rect 4360 59264 4376 59328
rect 4440 59264 4456 59328
rect 4520 59264 4528 59328
rect 4208 58240 4528 59264
rect 4208 58176 4216 58240
rect 4280 58176 4296 58240
rect 4360 58176 4376 58240
rect 4440 58176 4456 58240
rect 4520 58176 4528 58240
rect 4208 57152 4528 58176
rect 4208 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4528 57152
rect 4208 56064 4528 57088
rect 4208 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4528 56064
rect 4208 54976 4528 56000
rect 4208 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4528 54976
rect 4208 53888 4528 54912
rect 4208 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4528 53888
rect 4208 52800 4528 53824
rect 4208 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4528 52800
rect 4208 51712 4528 52736
rect 4208 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4528 51712
rect 4208 50624 4528 51648
rect 4208 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4528 50624
rect 4208 49536 4528 50560
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 48448 4528 49472
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 47360 4528 48384
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36260 4528 36416
rect 4208 36024 4250 36260
rect 4486 36024 4528 36260
rect 4208 35392 4528 36024
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5624 4528 5952
rect 4208 5388 4250 5624
rect 4486 5388 4528 5624
rect 4208 4928 4528 5388
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 934 4528 2688
rect 4208 698 4250 934
rect 4486 698 4528 934
rect -1076 38 -1034 274
rect -798 38 -756 274
rect -1076 -4 -756 38
rect 4208 -4 4528 698
rect 4868 97882 5188 97924
rect 4868 97646 4910 97882
rect 5146 97646 5188 97882
rect 4868 95776 5188 97646
rect 4868 95712 4876 95776
rect 4940 95712 4956 95776
rect 5020 95712 5036 95776
rect 5100 95712 5116 95776
rect 5180 95712 5188 95776
rect 4868 94688 5188 95712
rect 4868 94624 4876 94688
rect 4940 94624 4956 94688
rect 5020 94624 5036 94688
rect 5100 94624 5116 94688
rect 5180 94624 5188 94688
rect 4868 93600 5188 94624
rect 4868 93536 4876 93600
rect 4940 93536 4956 93600
rect 5020 93536 5036 93600
rect 5100 93536 5116 93600
rect 5180 93536 5188 93600
rect 4868 92512 5188 93536
rect 4868 92448 4876 92512
rect 4940 92448 4956 92512
rect 5020 92448 5036 92512
rect 5100 92448 5116 92512
rect 5180 92448 5188 92512
rect 4868 91424 5188 92448
rect 4868 91360 4876 91424
rect 4940 91360 4956 91424
rect 5020 91360 5036 91424
rect 5100 91360 5116 91424
rect 5180 91360 5188 91424
rect 4868 90336 5188 91360
rect 34928 97222 35248 97924
rect 34928 96986 34970 97222
rect 35206 96986 35248 97222
rect 34928 95232 35248 96986
rect 34928 95168 34936 95232
rect 35000 95168 35016 95232
rect 35080 95168 35096 95232
rect 35160 95168 35176 95232
rect 35240 95168 35248 95232
rect 34928 94144 35248 95168
rect 34928 94080 34936 94144
rect 35000 94080 35016 94144
rect 35080 94080 35096 94144
rect 35160 94080 35176 94144
rect 35240 94080 35248 94144
rect 34928 93056 35248 94080
rect 34928 92992 34936 93056
rect 35000 92992 35016 93056
rect 35080 92992 35096 93056
rect 35160 92992 35176 93056
rect 35240 92992 35248 93056
rect 34928 91057 35248 92992
rect 35588 97882 35908 97924
rect 35588 97646 35630 97882
rect 35866 97646 35908 97882
rect 35588 95776 35908 97646
rect 35588 95712 35596 95776
rect 35660 95712 35676 95776
rect 35740 95712 35756 95776
rect 35820 95712 35836 95776
rect 35900 95712 35908 95776
rect 35588 94688 35908 95712
rect 35588 94624 35596 94688
rect 35660 94624 35676 94688
rect 35740 94624 35756 94688
rect 35820 94624 35836 94688
rect 35900 94624 35908 94688
rect 35588 93600 35908 94624
rect 35588 93536 35596 93600
rect 35660 93536 35676 93600
rect 35740 93536 35756 93600
rect 35820 93536 35836 93600
rect 35900 93536 35908 93600
rect 35588 91057 35908 93536
rect 65648 97222 65968 97924
rect 65648 96986 65690 97222
rect 65926 96986 65968 97222
rect 65648 95232 65968 96986
rect 65648 95168 65656 95232
rect 65720 95168 65736 95232
rect 65800 95168 65816 95232
rect 65880 95168 65896 95232
rect 65960 95168 65968 95232
rect 65648 94144 65968 95168
rect 65648 94080 65656 94144
rect 65720 94080 65736 94144
rect 65800 94080 65816 94144
rect 65880 94080 65896 94144
rect 65960 94080 65968 94144
rect 65648 93056 65968 94080
rect 65648 92992 65656 93056
rect 65720 92992 65736 93056
rect 65800 92992 65816 93056
rect 65880 92992 65896 93056
rect 65960 92992 65968 93056
rect 65648 91057 65968 92992
rect 66308 97882 66628 97924
rect 66308 97646 66350 97882
rect 66586 97646 66628 97882
rect 66308 95776 66628 97646
rect 66308 95712 66316 95776
rect 66380 95712 66396 95776
rect 66460 95712 66476 95776
rect 66540 95712 66556 95776
rect 66620 95712 66628 95776
rect 66308 94688 66628 95712
rect 66308 94624 66316 94688
rect 66380 94624 66396 94688
rect 66460 94624 66476 94688
rect 66540 94624 66556 94688
rect 66620 94624 66628 94688
rect 66308 93600 66628 94624
rect 66308 93536 66316 93600
rect 66380 93536 66396 93600
rect 66460 93536 66476 93600
rect 66540 93536 66556 93600
rect 66620 93536 66628 93600
rect 66308 91057 66628 93536
rect 96368 97222 96688 97924
rect 96368 96986 96410 97222
rect 96646 96986 96688 97222
rect 96368 95232 96688 96986
rect 96368 95168 96376 95232
rect 96440 95168 96456 95232
rect 96520 95168 96536 95232
rect 96600 95168 96616 95232
rect 96680 95168 96688 95232
rect 96368 94144 96688 95168
rect 96368 94080 96376 94144
rect 96440 94080 96456 94144
rect 96520 94080 96536 94144
rect 96600 94080 96616 94144
rect 96680 94080 96688 94144
rect 96368 93056 96688 94080
rect 96368 92992 96376 93056
rect 96440 92992 96456 93056
rect 96520 92992 96536 93056
rect 96600 92992 96616 93056
rect 96680 92992 96688 93056
rect 96368 91968 96688 92992
rect 96368 91904 96376 91968
rect 96440 91904 96456 91968
rect 96520 91904 96536 91968
rect 96600 91904 96616 91968
rect 96680 91904 96688 91968
rect 96368 90880 96688 91904
rect 96368 90816 96376 90880
rect 96440 90816 96456 90880
rect 96520 90816 96536 90880
rect 96600 90816 96616 90880
rect 96680 90816 96688 90880
rect 50843 90540 50909 90541
rect 50843 90476 50844 90540
rect 50908 90476 50909 90540
rect 50843 90475 50909 90476
rect 4868 90272 4876 90336
rect 4940 90272 4956 90336
rect 5020 90272 5036 90336
rect 5100 90272 5116 90336
rect 5180 90272 5188 90336
rect 4868 89248 5188 90272
rect 4868 89184 4876 89248
rect 4940 89184 4956 89248
rect 5020 89184 5036 89248
rect 5100 89184 5116 89248
rect 5180 89184 5188 89248
rect 4868 88160 5188 89184
rect 4868 88096 4876 88160
rect 4940 88096 4956 88160
rect 5020 88096 5036 88160
rect 5100 88096 5116 88160
rect 5180 88096 5188 88160
rect 4868 87072 5188 88096
rect 4868 87008 4876 87072
rect 4940 87008 4956 87072
rect 5020 87008 5036 87072
rect 5100 87008 5116 87072
rect 5180 87008 5188 87072
rect 4868 85984 5188 87008
rect 12868 86684 12910 86920
rect 13146 86684 13188 86920
rect 43588 86684 43630 86920
rect 43866 86684 43908 86920
rect 12208 86024 12250 86260
rect 12486 86024 12528 86260
rect 42928 86024 42970 86260
rect 43206 86024 43248 86260
rect 4868 85920 4876 85984
rect 4940 85920 4956 85984
rect 5020 85920 5036 85984
rect 5100 85920 5116 85984
rect 5180 85920 5188 85984
rect 4868 84896 5188 85920
rect 4868 84832 4876 84896
rect 4940 84832 4956 84896
rect 5020 84832 5036 84896
rect 5100 84832 5116 84896
rect 5180 84832 5188 84896
rect 4868 83808 5188 84832
rect 4868 83744 4876 83808
rect 4940 83744 4956 83808
rect 5020 83744 5036 83808
rect 5100 83744 5116 83808
rect 5180 83744 5188 83808
rect 4868 82720 5188 83744
rect 4868 82656 4876 82720
rect 4940 82656 4956 82720
rect 5020 82656 5036 82720
rect 5100 82656 5116 82720
rect 5180 82656 5188 82720
rect 4868 81632 5188 82656
rect 4868 81568 4876 81632
rect 4940 81568 4956 81632
rect 5020 81568 5036 81632
rect 5100 81568 5116 81632
rect 5180 81568 5188 81632
rect 4868 80544 5188 81568
rect 4868 80480 4876 80544
rect 4940 80480 4956 80544
rect 5020 80480 5036 80544
rect 5100 80480 5116 80544
rect 5180 80480 5188 80544
rect 4868 79456 5188 80480
rect 4868 79392 4876 79456
rect 4940 79392 4956 79456
rect 5020 79392 5036 79456
rect 5100 79392 5116 79456
rect 5180 79392 5188 79456
rect 4868 78368 5188 79392
rect 4868 78304 4876 78368
rect 4940 78304 4956 78368
rect 5020 78304 5036 78368
rect 5100 78304 5116 78368
rect 5180 78304 5188 78368
rect 4868 77280 5188 78304
rect 4868 77216 4876 77280
rect 4940 77216 4956 77280
rect 5020 77216 5036 77280
rect 5100 77216 5116 77280
rect 5180 77216 5188 77280
rect 4868 76192 5188 77216
rect 4868 76128 4876 76192
rect 4940 76128 4956 76192
rect 5020 76128 5036 76192
rect 5100 76128 5116 76192
rect 5180 76128 5188 76192
rect 4868 75104 5188 76128
rect 4868 75040 4876 75104
rect 4940 75040 4956 75104
rect 5020 75040 5036 75104
rect 5100 75040 5116 75104
rect 5180 75040 5188 75104
rect 4868 74016 5188 75040
rect 4868 73952 4876 74016
rect 4940 73952 4956 74016
rect 5020 73952 5036 74016
rect 5100 73952 5116 74016
rect 5180 73952 5188 74016
rect 4868 72928 5188 73952
rect 4868 72864 4876 72928
rect 4940 72864 4956 72928
rect 5020 72864 5036 72928
rect 5100 72864 5116 72928
rect 5180 72864 5188 72928
rect 4868 71840 5188 72864
rect 4868 71776 4876 71840
rect 4940 71776 4956 71840
rect 5020 71776 5036 71840
rect 5100 71776 5116 71840
rect 5180 71776 5188 71840
rect 4868 70752 5188 71776
rect 4868 70688 4876 70752
rect 4940 70688 4956 70752
rect 5020 70688 5036 70752
rect 5100 70688 5116 70752
rect 5180 70688 5188 70752
rect 4868 69664 5188 70688
rect 4868 69600 4876 69664
rect 4940 69600 4956 69664
rect 5020 69600 5036 69664
rect 5100 69600 5116 69664
rect 5180 69600 5188 69664
rect 4868 68576 5188 69600
rect 4868 68512 4876 68576
rect 4940 68512 4956 68576
rect 5020 68512 5036 68576
rect 5100 68512 5116 68576
rect 5180 68512 5188 68576
rect 4868 67556 5188 68512
rect 4868 67488 4910 67556
rect 5146 67488 5188 67556
rect 4868 67424 4876 67488
rect 5180 67424 5188 67488
rect 4868 67320 4910 67424
rect 5146 67320 5188 67424
rect 12868 67320 12910 67556
rect 13146 67320 13188 67556
rect 43588 67320 43630 67556
rect 43866 67320 43908 67556
rect 4868 66400 5188 67320
rect 12208 66660 12250 66896
rect 12486 66660 12528 66896
rect 42928 66660 42970 66896
rect 43206 66660 43248 66896
rect 4868 66336 4876 66400
rect 4940 66336 4956 66400
rect 5020 66336 5036 66400
rect 5100 66336 5116 66400
rect 5180 66336 5188 66400
rect 4868 65312 5188 66336
rect 4868 65248 4876 65312
rect 4940 65248 4956 65312
rect 5020 65248 5036 65312
rect 5100 65248 5116 65312
rect 5180 65248 5188 65312
rect 4868 64224 5188 65248
rect 4868 64160 4876 64224
rect 4940 64160 4956 64224
rect 5020 64160 5036 64224
rect 5100 64160 5116 64224
rect 5180 64160 5188 64224
rect 4868 63136 5188 64160
rect 4868 63072 4876 63136
rect 4940 63072 4956 63136
rect 5020 63072 5036 63136
rect 5100 63072 5116 63136
rect 5180 63072 5188 63136
rect 4868 62048 5188 63072
rect 4868 61984 4876 62048
rect 4940 61984 4956 62048
rect 5020 61984 5036 62048
rect 5100 61984 5116 62048
rect 5180 61984 5188 62048
rect 4868 60960 5188 61984
rect 4868 60896 4876 60960
rect 4940 60896 4956 60960
rect 5020 60896 5036 60960
rect 5100 60896 5116 60960
rect 5180 60896 5188 60960
rect 4868 59872 5188 60896
rect 4868 59808 4876 59872
rect 4940 59808 4956 59872
rect 5020 59808 5036 59872
rect 5100 59808 5116 59872
rect 5180 59808 5188 59872
rect 4868 58784 5188 59808
rect 4868 58720 4876 58784
rect 4940 58720 4956 58784
rect 5020 58720 5036 58784
rect 5100 58720 5116 58784
rect 5180 58720 5188 58784
rect 4868 57696 5188 58720
rect 4868 57632 4876 57696
rect 4940 57632 4956 57696
rect 5020 57632 5036 57696
rect 5100 57632 5116 57696
rect 5180 57632 5188 57696
rect 4868 56608 5188 57632
rect 4868 56544 4876 56608
rect 4940 56544 4956 56608
rect 5020 56544 5036 56608
rect 5100 56544 5116 56608
rect 5180 56544 5188 56608
rect 4868 55520 5188 56544
rect 12868 56048 12910 56284
rect 13146 56048 13188 56284
rect 43588 56048 43630 56284
rect 43866 56048 43908 56284
rect 4868 55456 4876 55520
rect 4940 55456 4956 55520
rect 5020 55456 5036 55520
rect 5100 55456 5116 55520
rect 5180 55456 5188 55520
rect 4868 54432 5188 55456
rect 12208 55388 12250 55624
rect 12486 55388 12528 55624
rect 42928 55388 42970 55624
rect 43206 55388 43248 55624
rect 4868 54368 4876 54432
rect 4940 54368 4956 54432
rect 5020 54368 5036 54432
rect 5100 54368 5116 54432
rect 5180 54368 5188 54432
rect 4868 53344 5188 54368
rect 4868 53280 4876 53344
rect 4940 53280 4956 53344
rect 5020 53280 5036 53344
rect 5100 53280 5116 53344
rect 5180 53280 5188 53344
rect 4868 52256 5188 53280
rect 4868 52192 4876 52256
rect 4940 52192 4956 52256
rect 5020 52192 5036 52256
rect 5100 52192 5116 52256
rect 5180 52192 5188 52256
rect 4868 51168 5188 52192
rect 4868 51104 4876 51168
rect 4940 51104 4956 51168
rect 5020 51104 5036 51168
rect 5100 51104 5116 51168
rect 5180 51104 5188 51168
rect 4868 50080 5188 51104
rect 4868 50016 4876 50080
rect 4940 50016 4956 50080
rect 5020 50016 5036 50080
rect 5100 50016 5116 50080
rect 5180 50016 5188 50080
rect 4868 48992 5188 50016
rect 4868 48928 4876 48992
rect 4940 48928 4956 48992
rect 5020 48928 5036 48992
rect 5100 48928 5116 48992
rect 5180 48928 5188 48992
rect 4868 47904 5188 48928
rect 4868 47840 4876 47904
rect 4940 47840 4956 47904
rect 5020 47840 5036 47904
rect 5100 47840 5116 47904
rect 5180 47840 5188 47904
rect 4868 46816 5188 47840
rect 4868 46752 4876 46816
rect 4940 46752 4956 46816
rect 5020 46752 5036 46816
rect 5100 46752 5116 46816
rect 5180 46752 5188 46816
rect 4868 45728 5188 46752
rect 4868 45664 4876 45728
rect 4940 45664 4956 45728
rect 5020 45664 5036 45728
rect 5100 45664 5116 45728
rect 5180 45664 5188 45728
rect 4868 44640 5188 45664
rect 12868 44684 12910 44920
rect 13146 44684 13188 44920
rect 43588 44684 43630 44920
rect 43866 44684 43908 44920
rect 4868 44576 4876 44640
rect 4940 44576 4956 44640
rect 5020 44576 5036 44640
rect 5100 44576 5116 44640
rect 5180 44576 5188 44640
rect 4868 43552 5188 44576
rect 12208 44024 12250 44260
rect 12486 44024 12528 44260
rect 42928 44024 42970 44260
rect 43206 44024 43248 44260
rect 4868 43488 4876 43552
rect 4940 43488 4956 43552
rect 5020 43488 5036 43552
rect 5100 43488 5116 43552
rect 5180 43488 5188 43552
rect 4868 42464 5188 43488
rect 4868 42400 4876 42464
rect 4940 42400 4956 42464
rect 5020 42400 5036 42464
rect 5100 42400 5116 42464
rect 5180 42400 5188 42464
rect 4868 41376 5188 42400
rect 4868 41312 4876 41376
rect 4940 41312 4956 41376
rect 5020 41312 5036 41376
rect 5100 41312 5116 41376
rect 5180 41312 5188 41376
rect 4868 40288 5188 41312
rect 4868 40224 4876 40288
rect 4940 40224 4956 40288
rect 5020 40224 5036 40288
rect 5100 40224 5116 40288
rect 5180 40224 5188 40288
rect 4868 39200 5188 40224
rect 4868 39136 4876 39200
rect 4940 39136 4956 39200
rect 5020 39136 5036 39200
rect 5100 39136 5116 39200
rect 5180 39136 5188 39200
rect 4868 38112 5188 39136
rect 4868 38048 4876 38112
rect 4940 38048 4956 38112
rect 5020 38048 5036 38112
rect 5100 38048 5116 38112
rect 5180 38048 5188 38112
rect 4868 37024 5188 38048
rect 4868 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5188 37024
rect 4868 36920 5188 36960
rect 4868 36684 4910 36920
rect 5146 36684 5188 36920
rect 12868 36684 12910 36920
rect 13146 36684 13188 36920
rect 43588 36684 43630 36920
rect 43866 36684 43908 36920
rect 4868 35936 5188 36684
rect 12208 36024 12250 36260
rect 12486 36024 12528 36260
rect 42928 36024 42970 36260
rect 43206 36024 43248 36260
rect 4868 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5188 35936
rect 4868 34848 5188 35872
rect 4868 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5188 34848
rect 4868 33760 5188 34784
rect 4868 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5188 33760
rect 4868 32672 5188 33696
rect 4868 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5188 32672
rect 4868 31584 5188 32608
rect 4868 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5188 31584
rect 4868 30496 5188 31520
rect 4868 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5188 30496
rect 4868 29408 5188 30432
rect 4868 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5188 29408
rect 4868 28320 5188 29344
rect 4868 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5188 28320
rect 4868 27232 5188 28256
rect 4868 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5188 27232
rect 4868 26144 5188 27168
rect 4868 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5188 26144
rect 4868 25056 5188 26080
rect 4868 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5188 25056
rect 4868 23968 5188 24992
rect 4868 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5188 23968
rect 4868 22880 5188 23904
rect 4868 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5188 22880
rect 4868 21792 5188 22816
rect 4868 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5188 21792
rect 4868 20704 5188 21728
rect 4868 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5188 20704
rect 4868 19616 5188 20640
rect 4868 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5188 19616
rect 4868 18528 5188 19552
rect 4868 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5188 18528
rect 4868 17440 5188 18464
rect 4868 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5188 17440
rect 4868 16352 5188 17376
rect 4868 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5188 16352
rect 4868 15264 5188 16288
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4868 13088 5188 14112
rect 12868 14048 12910 14284
rect 13146 14048 13188 14284
rect 43588 14048 43630 14284
rect 43866 14048 43908 14284
rect 12208 13388 12250 13624
rect 12486 13388 12528 13624
rect 42928 13388 42970 13624
rect 43206 13388 43248 13624
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4868 10912 5188 11936
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 50846 8669 50906 90475
rect 96368 89792 96688 90816
rect 96368 89728 96376 89792
rect 96440 89728 96456 89792
rect 96520 89728 96536 89792
rect 96600 89728 96616 89792
rect 96680 89728 96688 89792
rect 96368 88704 96688 89728
rect 96368 88640 96376 88704
rect 96440 88640 96456 88704
rect 96520 88640 96536 88704
rect 96600 88640 96616 88704
rect 96680 88640 96688 88704
rect 96368 87616 96688 88640
rect 96368 87552 96376 87616
rect 96440 87552 96456 87616
rect 96520 87552 96536 87616
rect 96600 87552 96616 87616
rect 96680 87552 96688 87616
rect 54868 86684 54910 86920
rect 55146 86684 55188 86920
rect 85588 86684 85630 86920
rect 85866 86684 85908 86920
rect 96368 86528 96688 87552
rect 96368 86464 96376 86528
rect 96440 86464 96456 86528
rect 96520 86464 96536 86528
rect 96600 86464 96616 86528
rect 96680 86464 96688 86528
rect 54208 86024 54250 86260
rect 54486 86024 54528 86260
rect 84928 86024 84970 86260
rect 85206 86024 85248 86260
rect 96368 85440 96688 86464
rect 96368 85376 96376 85440
rect 96440 85376 96456 85440
rect 96520 85376 96536 85440
rect 96600 85376 96616 85440
rect 96680 85376 96688 85440
rect 96368 84352 96688 85376
rect 96368 84288 96376 84352
rect 96440 84288 96456 84352
rect 96520 84288 96536 84352
rect 96600 84288 96616 84352
rect 96680 84288 96688 84352
rect 96368 83264 96688 84288
rect 96368 83200 96376 83264
rect 96440 83200 96456 83264
rect 96520 83200 96536 83264
rect 96600 83200 96616 83264
rect 96680 83200 96688 83264
rect 96368 82176 96688 83200
rect 96368 82112 96376 82176
rect 96440 82112 96456 82176
rect 96520 82112 96536 82176
rect 96600 82112 96616 82176
rect 96680 82112 96688 82176
rect 96368 81088 96688 82112
rect 96368 81024 96376 81088
rect 96440 81024 96456 81088
rect 96520 81024 96536 81088
rect 96600 81024 96616 81088
rect 96680 81024 96688 81088
rect 96368 80000 96688 81024
rect 96368 79936 96376 80000
rect 96440 79936 96456 80000
rect 96520 79936 96536 80000
rect 96600 79936 96616 80000
rect 96680 79936 96688 80000
rect 96368 78912 96688 79936
rect 96368 78848 96376 78912
rect 96440 78848 96456 78912
rect 96520 78848 96536 78912
rect 96600 78848 96616 78912
rect 96680 78848 96688 78912
rect 96368 77824 96688 78848
rect 96368 77760 96376 77824
rect 96440 77760 96456 77824
rect 96520 77760 96536 77824
rect 96600 77760 96616 77824
rect 96680 77760 96688 77824
rect 96368 76736 96688 77760
rect 96368 76672 96376 76736
rect 96440 76672 96456 76736
rect 96520 76672 96536 76736
rect 96600 76672 96616 76736
rect 96680 76672 96688 76736
rect 96368 75648 96688 76672
rect 96368 75584 96376 75648
rect 96440 75584 96456 75648
rect 96520 75584 96536 75648
rect 96600 75584 96616 75648
rect 96680 75584 96688 75648
rect 96368 74560 96688 75584
rect 96368 74496 96376 74560
rect 96440 74496 96456 74560
rect 96520 74496 96536 74560
rect 96600 74496 96616 74560
rect 96680 74496 96688 74560
rect 96368 73472 96688 74496
rect 96368 73408 96376 73472
rect 96440 73408 96456 73472
rect 96520 73408 96536 73472
rect 96600 73408 96616 73472
rect 96680 73408 96688 73472
rect 96368 72384 96688 73408
rect 96368 72320 96376 72384
rect 96440 72320 96456 72384
rect 96520 72320 96536 72384
rect 96600 72320 96616 72384
rect 96680 72320 96688 72384
rect 96368 71296 96688 72320
rect 96368 71232 96376 71296
rect 96440 71232 96456 71296
rect 96520 71232 96536 71296
rect 96600 71232 96616 71296
rect 96680 71232 96688 71296
rect 96368 70208 96688 71232
rect 96368 70144 96376 70208
rect 96440 70144 96456 70208
rect 96520 70144 96536 70208
rect 96600 70144 96616 70208
rect 96680 70144 96688 70208
rect 96368 69120 96688 70144
rect 96368 69056 96376 69120
rect 96440 69056 96456 69120
rect 96520 69056 96536 69120
rect 96600 69056 96616 69120
rect 96680 69056 96688 69120
rect 96368 68032 96688 69056
rect 96368 67968 96376 68032
rect 96440 67968 96456 68032
rect 96520 67968 96536 68032
rect 96600 67968 96616 68032
rect 96680 67968 96688 68032
rect 54868 67320 54910 67556
rect 55146 67320 55188 67556
rect 85588 67320 85630 67556
rect 85866 67320 85908 67556
rect 96368 66944 96688 67968
rect 54208 66660 54250 66896
rect 54486 66660 54528 66896
rect 84928 66660 84970 66896
rect 85206 66660 85248 66896
rect 96368 66880 96376 66944
rect 96440 66896 96456 66944
rect 96520 66896 96536 66944
rect 96600 66896 96616 66944
rect 96680 66880 96688 66944
rect 96368 66660 96410 66880
rect 96646 66660 96688 66880
rect 96368 65856 96688 66660
rect 96368 65792 96376 65856
rect 96440 65792 96456 65856
rect 96520 65792 96536 65856
rect 96600 65792 96616 65856
rect 96680 65792 96688 65856
rect 96368 64768 96688 65792
rect 96368 64704 96376 64768
rect 96440 64704 96456 64768
rect 96520 64704 96536 64768
rect 96600 64704 96616 64768
rect 96680 64704 96688 64768
rect 96368 63680 96688 64704
rect 96368 63616 96376 63680
rect 96440 63616 96456 63680
rect 96520 63616 96536 63680
rect 96600 63616 96616 63680
rect 96680 63616 96688 63680
rect 96368 62592 96688 63616
rect 96368 62528 96376 62592
rect 96440 62528 96456 62592
rect 96520 62528 96536 62592
rect 96600 62528 96616 62592
rect 96680 62528 96688 62592
rect 96368 61504 96688 62528
rect 96368 61440 96376 61504
rect 96440 61440 96456 61504
rect 96520 61440 96536 61504
rect 96600 61440 96616 61504
rect 96680 61440 96688 61504
rect 96368 60416 96688 61440
rect 96368 60352 96376 60416
rect 96440 60352 96456 60416
rect 96520 60352 96536 60416
rect 96600 60352 96616 60416
rect 96680 60352 96688 60416
rect 96368 59328 96688 60352
rect 96368 59264 96376 59328
rect 96440 59264 96456 59328
rect 96520 59264 96536 59328
rect 96600 59264 96616 59328
rect 96680 59264 96688 59328
rect 96368 58240 96688 59264
rect 96368 58176 96376 58240
rect 96440 58176 96456 58240
rect 96520 58176 96536 58240
rect 96600 58176 96616 58240
rect 96680 58176 96688 58240
rect 96368 57152 96688 58176
rect 96368 57088 96376 57152
rect 96440 57088 96456 57152
rect 96520 57088 96536 57152
rect 96600 57088 96616 57152
rect 96680 57088 96688 57152
rect 54868 56048 54910 56284
rect 55146 56048 55188 56284
rect 85588 56048 85630 56284
rect 85866 56048 85908 56284
rect 96368 56064 96688 57088
rect 96368 56000 96376 56064
rect 96440 56000 96456 56064
rect 96520 56000 96536 56064
rect 96600 56000 96616 56064
rect 96680 56000 96688 56064
rect 54208 55388 54250 55624
rect 54486 55388 54528 55624
rect 84928 55388 84970 55624
rect 85206 55388 85248 55624
rect 96368 54976 96688 56000
rect 96368 54912 96376 54976
rect 96440 54912 96456 54976
rect 96520 54912 96536 54976
rect 96600 54912 96616 54976
rect 96680 54912 96688 54976
rect 96368 53888 96688 54912
rect 96368 53824 96376 53888
rect 96440 53824 96456 53888
rect 96520 53824 96536 53888
rect 96600 53824 96616 53888
rect 96680 53824 96688 53888
rect 96368 52800 96688 53824
rect 96368 52736 96376 52800
rect 96440 52736 96456 52800
rect 96520 52736 96536 52800
rect 96600 52736 96616 52800
rect 96680 52736 96688 52800
rect 96368 51712 96688 52736
rect 96368 51648 96376 51712
rect 96440 51648 96456 51712
rect 96520 51648 96536 51712
rect 96600 51648 96616 51712
rect 96680 51648 96688 51712
rect 96368 50624 96688 51648
rect 96368 50560 96376 50624
rect 96440 50560 96456 50624
rect 96520 50560 96536 50624
rect 96600 50560 96616 50624
rect 96680 50560 96688 50624
rect 96368 49536 96688 50560
rect 96368 49472 96376 49536
rect 96440 49472 96456 49536
rect 96520 49472 96536 49536
rect 96600 49472 96616 49536
rect 96680 49472 96688 49536
rect 96368 48448 96688 49472
rect 96368 48384 96376 48448
rect 96440 48384 96456 48448
rect 96520 48384 96536 48448
rect 96600 48384 96616 48448
rect 96680 48384 96688 48448
rect 96368 47360 96688 48384
rect 96368 47296 96376 47360
rect 96440 47296 96456 47360
rect 96520 47296 96536 47360
rect 96600 47296 96616 47360
rect 96680 47296 96688 47360
rect 96368 46272 96688 47296
rect 96368 46208 96376 46272
rect 96440 46208 96456 46272
rect 96520 46208 96536 46272
rect 96600 46208 96616 46272
rect 96680 46208 96688 46272
rect 96368 45184 96688 46208
rect 96368 45120 96376 45184
rect 96440 45120 96456 45184
rect 96520 45120 96536 45184
rect 96600 45120 96616 45184
rect 96680 45120 96688 45184
rect 54868 44684 54910 44920
rect 55146 44684 55188 44920
rect 85588 44684 85630 44920
rect 85866 44684 85908 44920
rect 54208 44024 54250 44260
rect 54486 44024 54528 44260
rect 84928 44024 84970 44260
rect 85206 44024 85248 44260
rect 96368 44096 96688 45120
rect 96368 44032 96376 44096
rect 96440 44032 96456 44096
rect 96520 44032 96536 44096
rect 96600 44032 96616 44096
rect 96680 44032 96688 44096
rect 96368 43008 96688 44032
rect 96368 42944 96376 43008
rect 96440 42944 96456 43008
rect 96520 42944 96536 43008
rect 96600 42944 96616 43008
rect 96680 42944 96688 43008
rect 96368 41920 96688 42944
rect 96368 41856 96376 41920
rect 96440 41856 96456 41920
rect 96520 41856 96536 41920
rect 96600 41856 96616 41920
rect 96680 41856 96688 41920
rect 96368 40832 96688 41856
rect 96368 40768 96376 40832
rect 96440 40768 96456 40832
rect 96520 40768 96536 40832
rect 96600 40768 96616 40832
rect 96680 40768 96688 40832
rect 96368 39744 96688 40768
rect 96368 39680 96376 39744
rect 96440 39680 96456 39744
rect 96520 39680 96536 39744
rect 96600 39680 96616 39744
rect 96680 39680 96688 39744
rect 96368 38656 96688 39680
rect 96368 38592 96376 38656
rect 96440 38592 96456 38656
rect 96520 38592 96536 38656
rect 96600 38592 96616 38656
rect 96680 38592 96688 38656
rect 96368 37568 96688 38592
rect 96368 37504 96376 37568
rect 96440 37504 96456 37568
rect 96520 37504 96536 37568
rect 96600 37504 96616 37568
rect 96680 37504 96688 37568
rect 54868 36684 54910 36920
rect 55146 36684 55188 36920
rect 85588 36684 85630 36920
rect 85866 36684 85908 36920
rect 96368 36480 96688 37504
rect 96368 36416 96376 36480
rect 96440 36416 96456 36480
rect 96520 36416 96536 36480
rect 96600 36416 96616 36480
rect 96680 36416 96688 36480
rect 96368 36260 96688 36416
rect 54208 36024 54250 36260
rect 54486 36024 54528 36260
rect 84928 36024 84970 36260
rect 85206 36024 85248 36260
rect 96368 36024 96410 36260
rect 96646 36024 96688 36260
rect 96368 35392 96688 36024
rect 96368 35328 96376 35392
rect 96440 35328 96456 35392
rect 96520 35328 96536 35392
rect 96600 35328 96616 35392
rect 96680 35328 96688 35392
rect 96368 34304 96688 35328
rect 96368 34240 96376 34304
rect 96440 34240 96456 34304
rect 96520 34240 96536 34304
rect 96600 34240 96616 34304
rect 96680 34240 96688 34304
rect 96368 33216 96688 34240
rect 96368 33152 96376 33216
rect 96440 33152 96456 33216
rect 96520 33152 96536 33216
rect 96600 33152 96616 33216
rect 96680 33152 96688 33216
rect 96368 32128 96688 33152
rect 96368 32064 96376 32128
rect 96440 32064 96456 32128
rect 96520 32064 96536 32128
rect 96600 32064 96616 32128
rect 96680 32064 96688 32128
rect 96368 31040 96688 32064
rect 96368 30976 96376 31040
rect 96440 30976 96456 31040
rect 96520 30976 96536 31040
rect 96600 30976 96616 31040
rect 96680 30976 96688 31040
rect 96368 29952 96688 30976
rect 96368 29888 96376 29952
rect 96440 29888 96456 29952
rect 96520 29888 96536 29952
rect 96600 29888 96616 29952
rect 96680 29888 96688 29952
rect 96368 28864 96688 29888
rect 96368 28800 96376 28864
rect 96440 28800 96456 28864
rect 96520 28800 96536 28864
rect 96600 28800 96616 28864
rect 96680 28800 96688 28864
rect 96368 27776 96688 28800
rect 96368 27712 96376 27776
rect 96440 27712 96456 27776
rect 96520 27712 96536 27776
rect 96600 27712 96616 27776
rect 96680 27712 96688 27776
rect 96368 26688 96688 27712
rect 96368 26624 96376 26688
rect 96440 26624 96456 26688
rect 96520 26624 96536 26688
rect 96600 26624 96616 26688
rect 96680 26624 96688 26688
rect 96368 25600 96688 26624
rect 96368 25536 96376 25600
rect 96440 25536 96456 25600
rect 96520 25536 96536 25600
rect 96600 25536 96616 25600
rect 96680 25536 96688 25600
rect 96368 24512 96688 25536
rect 96368 24448 96376 24512
rect 96440 24448 96456 24512
rect 96520 24448 96536 24512
rect 96600 24448 96616 24512
rect 96680 24448 96688 24512
rect 96368 23424 96688 24448
rect 96368 23360 96376 23424
rect 96440 23360 96456 23424
rect 96520 23360 96536 23424
rect 96600 23360 96616 23424
rect 96680 23360 96688 23424
rect 96368 22336 96688 23360
rect 96368 22272 96376 22336
rect 96440 22272 96456 22336
rect 96520 22272 96536 22336
rect 96600 22272 96616 22336
rect 96680 22272 96688 22336
rect 96368 21248 96688 22272
rect 96368 21184 96376 21248
rect 96440 21184 96456 21248
rect 96520 21184 96536 21248
rect 96600 21184 96616 21248
rect 96680 21184 96688 21248
rect 96368 20160 96688 21184
rect 96368 20096 96376 20160
rect 96440 20096 96456 20160
rect 96520 20096 96536 20160
rect 96600 20096 96616 20160
rect 96680 20096 96688 20160
rect 96368 19072 96688 20096
rect 96368 19008 96376 19072
rect 96440 19008 96456 19072
rect 96520 19008 96536 19072
rect 96600 19008 96616 19072
rect 96680 19008 96688 19072
rect 96368 17984 96688 19008
rect 96368 17920 96376 17984
rect 96440 17920 96456 17984
rect 96520 17920 96536 17984
rect 96600 17920 96616 17984
rect 96680 17920 96688 17984
rect 96368 16896 96688 17920
rect 96368 16832 96376 16896
rect 96440 16832 96456 16896
rect 96520 16832 96536 16896
rect 96600 16832 96616 16896
rect 96680 16832 96688 16896
rect 96368 15808 96688 16832
rect 96368 15744 96376 15808
rect 96440 15744 96456 15808
rect 96520 15744 96536 15808
rect 96600 15744 96616 15808
rect 96680 15744 96688 15808
rect 96368 14720 96688 15744
rect 96368 14656 96376 14720
rect 96440 14656 96456 14720
rect 96520 14656 96536 14720
rect 96600 14656 96616 14720
rect 96680 14656 96688 14720
rect 54868 14048 54910 14284
rect 55146 14048 55188 14284
rect 85588 14048 85630 14284
rect 85866 14048 85908 14284
rect 96368 13632 96688 14656
rect 54208 13388 54250 13624
rect 54486 13388 54528 13624
rect 84928 13388 84970 13624
rect 85206 13388 85248 13624
rect 96368 13568 96376 13632
rect 96440 13568 96456 13632
rect 96520 13568 96536 13632
rect 96600 13568 96616 13632
rect 96680 13568 96688 13632
rect 96368 12544 96688 13568
rect 96368 12480 96376 12544
rect 96440 12480 96456 12544
rect 96520 12480 96536 12544
rect 96600 12480 96616 12544
rect 96680 12480 96688 12544
rect 96368 11456 96688 12480
rect 96368 11392 96376 11456
rect 96440 11392 96456 11456
rect 96520 11392 96536 11456
rect 96600 11392 96616 11456
rect 96680 11392 96688 11456
rect 96368 10368 96688 11392
rect 96368 10304 96376 10368
rect 96440 10304 96456 10368
rect 96520 10304 96536 10368
rect 96600 10304 96616 10368
rect 96680 10304 96688 10368
rect 96368 9280 96688 10304
rect 96368 9216 96376 9280
rect 96440 9216 96456 9280
rect 96520 9216 96536 9280
rect 96600 9216 96616 9280
rect 96680 9216 96688 9280
rect 50843 8668 50909 8669
rect 50843 8604 50844 8668
rect 50908 8604 50909 8668
rect 50843 8603 50909 8604
rect 96368 8192 96688 9216
rect 96368 8128 96376 8192
rect 96440 8128 96456 8192
rect 96520 8128 96536 8192
rect 96600 8128 96616 8192
rect 96680 8128 96688 8192
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 6284 5188 6496
rect 4868 6048 4910 6284
rect 5146 6048 5188 6284
rect 4868 5472 5188 6048
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 274 5188 2144
rect 4868 38 4910 274
rect 5146 38 5188 274
rect 4868 -4 5188 38
rect 34928 6016 35248 8015
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5624 35248 5952
rect 34928 5388 34970 5624
rect 35206 5388 35248 5624
rect 34928 4928 35248 5388
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 934 35248 2688
rect 34928 698 34970 934
rect 35206 698 35248 934
rect 34928 -4 35248 698
rect 35588 6284 35908 8015
rect 35588 6048 35630 6284
rect 35866 6048 35908 6284
rect 35588 5472 35908 6048
rect 35588 5408 35596 5472
rect 35660 5408 35676 5472
rect 35740 5408 35756 5472
rect 35820 5408 35836 5472
rect 35900 5408 35908 5472
rect 35588 4384 35908 5408
rect 35588 4320 35596 4384
rect 35660 4320 35676 4384
rect 35740 4320 35756 4384
rect 35820 4320 35836 4384
rect 35900 4320 35908 4384
rect 35588 3296 35908 4320
rect 35588 3232 35596 3296
rect 35660 3232 35676 3296
rect 35740 3232 35756 3296
rect 35820 3232 35836 3296
rect 35900 3232 35908 3296
rect 35588 2208 35908 3232
rect 35588 2144 35596 2208
rect 35660 2144 35676 2208
rect 35740 2144 35756 2208
rect 35820 2144 35836 2208
rect 35900 2144 35908 2208
rect 35588 274 35908 2144
rect 35588 38 35630 274
rect 35866 38 35908 274
rect 35588 -4 35908 38
rect 65648 6016 65968 8015
rect 65648 5952 65656 6016
rect 65720 5952 65736 6016
rect 65800 5952 65816 6016
rect 65880 5952 65896 6016
rect 65960 5952 65968 6016
rect 65648 5624 65968 5952
rect 65648 5388 65690 5624
rect 65926 5388 65968 5624
rect 65648 4928 65968 5388
rect 65648 4864 65656 4928
rect 65720 4864 65736 4928
rect 65800 4864 65816 4928
rect 65880 4864 65896 4928
rect 65960 4864 65968 4928
rect 65648 3840 65968 4864
rect 65648 3776 65656 3840
rect 65720 3776 65736 3840
rect 65800 3776 65816 3840
rect 65880 3776 65896 3840
rect 65960 3776 65968 3840
rect 65648 2752 65968 3776
rect 65648 2688 65656 2752
rect 65720 2688 65736 2752
rect 65800 2688 65816 2752
rect 65880 2688 65896 2752
rect 65960 2688 65968 2752
rect 65648 934 65968 2688
rect 65648 698 65690 934
rect 65926 698 65968 934
rect 65648 -4 65968 698
rect 66308 6284 66628 8015
rect 66308 6048 66350 6284
rect 66586 6048 66628 6284
rect 66308 5472 66628 6048
rect 66308 5408 66316 5472
rect 66380 5408 66396 5472
rect 66460 5408 66476 5472
rect 66540 5408 66556 5472
rect 66620 5408 66628 5472
rect 66308 4384 66628 5408
rect 66308 4320 66316 4384
rect 66380 4320 66396 4384
rect 66460 4320 66476 4384
rect 66540 4320 66556 4384
rect 66620 4320 66628 4384
rect 66308 3296 66628 4320
rect 66308 3232 66316 3296
rect 66380 3232 66396 3296
rect 66460 3232 66476 3296
rect 66540 3232 66556 3296
rect 66620 3232 66628 3296
rect 66308 2208 66628 3232
rect 66308 2144 66316 2208
rect 66380 2144 66396 2208
rect 66460 2144 66476 2208
rect 66540 2144 66556 2208
rect 66620 2144 66628 2208
rect 66308 274 66628 2144
rect 66308 38 66350 274
rect 66586 38 66628 274
rect 66308 -4 66628 38
rect 96368 7104 96688 8128
rect 96368 7040 96376 7104
rect 96440 7040 96456 7104
rect 96520 7040 96536 7104
rect 96600 7040 96616 7104
rect 96680 7040 96688 7104
rect 96368 6016 96688 7040
rect 96368 5952 96376 6016
rect 96440 5952 96456 6016
rect 96520 5952 96536 6016
rect 96600 5952 96616 6016
rect 96680 5952 96688 6016
rect 96368 5624 96688 5952
rect 96368 5388 96410 5624
rect 96646 5388 96688 5624
rect 96368 4928 96688 5388
rect 96368 4864 96376 4928
rect 96440 4864 96456 4928
rect 96520 4864 96536 4928
rect 96600 4864 96616 4928
rect 96680 4864 96688 4928
rect 96368 3840 96688 4864
rect 96368 3776 96376 3840
rect 96440 3776 96456 3840
rect 96520 3776 96536 3840
rect 96600 3776 96616 3840
rect 96680 3776 96688 3840
rect 96368 2752 96688 3776
rect 96368 2688 96376 2752
rect 96440 2688 96456 2752
rect 96520 2688 96536 2752
rect 96600 2688 96616 2752
rect 96680 2688 96688 2752
rect 96368 934 96688 2688
rect 96368 698 96410 934
rect 96646 698 96688 934
rect 96368 -4 96688 698
rect 97028 97882 97348 97924
rect 97028 97646 97070 97882
rect 97306 97646 97348 97882
rect 97028 95776 97348 97646
rect 99748 97882 100068 97924
rect 99748 97646 99790 97882
rect 100026 97646 100068 97882
rect 97028 95712 97036 95776
rect 97100 95712 97116 95776
rect 97180 95712 97196 95776
rect 97260 95712 97276 95776
rect 97340 95712 97348 95776
rect 97028 94688 97348 95712
rect 97028 94624 97036 94688
rect 97100 94624 97116 94688
rect 97180 94624 97196 94688
rect 97260 94624 97276 94688
rect 97340 94624 97348 94688
rect 97028 93600 97348 94624
rect 97028 93536 97036 93600
rect 97100 93536 97116 93600
rect 97180 93536 97196 93600
rect 97260 93536 97276 93600
rect 97340 93536 97348 93600
rect 97028 92512 97348 93536
rect 97028 92448 97036 92512
rect 97100 92448 97116 92512
rect 97180 92448 97196 92512
rect 97260 92448 97276 92512
rect 97340 92448 97348 92512
rect 97028 91424 97348 92448
rect 97028 91360 97036 91424
rect 97100 91360 97116 91424
rect 97180 91360 97196 91424
rect 97260 91360 97276 91424
rect 97340 91360 97348 91424
rect 97028 90336 97348 91360
rect 97028 90272 97036 90336
rect 97100 90272 97116 90336
rect 97180 90272 97196 90336
rect 97260 90272 97276 90336
rect 97340 90272 97348 90336
rect 97028 89248 97348 90272
rect 97028 89184 97036 89248
rect 97100 89184 97116 89248
rect 97180 89184 97196 89248
rect 97260 89184 97276 89248
rect 97340 89184 97348 89248
rect 97028 88160 97348 89184
rect 97028 88096 97036 88160
rect 97100 88096 97116 88160
rect 97180 88096 97196 88160
rect 97260 88096 97276 88160
rect 97340 88096 97348 88160
rect 97028 87072 97348 88096
rect 97028 87008 97036 87072
rect 97100 87008 97116 87072
rect 97180 87008 97196 87072
rect 97260 87008 97276 87072
rect 97340 87008 97348 87072
rect 97028 85984 97348 87008
rect 97028 85920 97036 85984
rect 97100 85920 97116 85984
rect 97180 85920 97196 85984
rect 97260 85920 97276 85984
rect 97340 85920 97348 85984
rect 97028 84896 97348 85920
rect 97028 84832 97036 84896
rect 97100 84832 97116 84896
rect 97180 84832 97196 84896
rect 97260 84832 97276 84896
rect 97340 84832 97348 84896
rect 97028 83808 97348 84832
rect 97028 83744 97036 83808
rect 97100 83744 97116 83808
rect 97180 83744 97196 83808
rect 97260 83744 97276 83808
rect 97340 83744 97348 83808
rect 97028 82720 97348 83744
rect 97028 82656 97036 82720
rect 97100 82656 97116 82720
rect 97180 82656 97196 82720
rect 97260 82656 97276 82720
rect 97340 82656 97348 82720
rect 97028 81632 97348 82656
rect 97028 81568 97036 81632
rect 97100 81568 97116 81632
rect 97180 81568 97196 81632
rect 97260 81568 97276 81632
rect 97340 81568 97348 81632
rect 97028 80544 97348 81568
rect 97028 80480 97036 80544
rect 97100 80480 97116 80544
rect 97180 80480 97196 80544
rect 97260 80480 97276 80544
rect 97340 80480 97348 80544
rect 97028 79456 97348 80480
rect 97028 79392 97036 79456
rect 97100 79392 97116 79456
rect 97180 79392 97196 79456
rect 97260 79392 97276 79456
rect 97340 79392 97348 79456
rect 97028 78368 97348 79392
rect 97028 78304 97036 78368
rect 97100 78304 97116 78368
rect 97180 78304 97196 78368
rect 97260 78304 97276 78368
rect 97340 78304 97348 78368
rect 97028 77280 97348 78304
rect 97028 77216 97036 77280
rect 97100 77216 97116 77280
rect 97180 77216 97196 77280
rect 97260 77216 97276 77280
rect 97340 77216 97348 77280
rect 97028 76192 97348 77216
rect 97028 76128 97036 76192
rect 97100 76128 97116 76192
rect 97180 76128 97196 76192
rect 97260 76128 97276 76192
rect 97340 76128 97348 76192
rect 97028 75104 97348 76128
rect 97028 75040 97036 75104
rect 97100 75040 97116 75104
rect 97180 75040 97196 75104
rect 97260 75040 97276 75104
rect 97340 75040 97348 75104
rect 97028 74016 97348 75040
rect 97028 73952 97036 74016
rect 97100 73952 97116 74016
rect 97180 73952 97196 74016
rect 97260 73952 97276 74016
rect 97340 73952 97348 74016
rect 97028 72928 97348 73952
rect 97028 72864 97036 72928
rect 97100 72864 97116 72928
rect 97180 72864 97196 72928
rect 97260 72864 97276 72928
rect 97340 72864 97348 72928
rect 97028 71840 97348 72864
rect 97028 71776 97036 71840
rect 97100 71776 97116 71840
rect 97180 71776 97196 71840
rect 97260 71776 97276 71840
rect 97340 71776 97348 71840
rect 97028 70752 97348 71776
rect 97028 70688 97036 70752
rect 97100 70688 97116 70752
rect 97180 70688 97196 70752
rect 97260 70688 97276 70752
rect 97340 70688 97348 70752
rect 97028 69664 97348 70688
rect 97028 69600 97036 69664
rect 97100 69600 97116 69664
rect 97180 69600 97196 69664
rect 97260 69600 97276 69664
rect 97340 69600 97348 69664
rect 97028 68576 97348 69600
rect 97028 68512 97036 68576
rect 97100 68512 97116 68576
rect 97180 68512 97196 68576
rect 97260 68512 97276 68576
rect 97340 68512 97348 68576
rect 97028 67556 97348 68512
rect 97028 67488 97070 67556
rect 97306 67488 97348 67556
rect 97028 67424 97036 67488
rect 97340 67424 97348 67488
rect 97028 67320 97070 67424
rect 97306 67320 97348 67424
rect 97028 66400 97348 67320
rect 97028 66336 97036 66400
rect 97100 66336 97116 66400
rect 97180 66336 97196 66400
rect 97260 66336 97276 66400
rect 97340 66336 97348 66400
rect 97028 65312 97348 66336
rect 97028 65248 97036 65312
rect 97100 65248 97116 65312
rect 97180 65248 97196 65312
rect 97260 65248 97276 65312
rect 97340 65248 97348 65312
rect 97028 64224 97348 65248
rect 97028 64160 97036 64224
rect 97100 64160 97116 64224
rect 97180 64160 97196 64224
rect 97260 64160 97276 64224
rect 97340 64160 97348 64224
rect 97028 63136 97348 64160
rect 97028 63072 97036 63136
rect 97100 63072 97116 63136
rect 97180 63072 97196 63136
rect 97260 63072 97276 63136
rect 97340 63072 97348 63136
rect 97028 62048 97348 63072
rect 97028 61984 97036 62048
rect 97100 61984 97116 62048
rect 97180 61984 97196 62048
rect 97260 61984 97276 62048
rect 97340 61984 97348 62048
rect 97028 60960 97348 61984
rect 97028 60896 97036 60960
rect 97100 60896 97116 60960
rect 97180 60896 97196 60960
rect 97260 60896 97276 60960
rect 97340 60896 97348 60960
rect 97028 59872 97348 60896
rect 97028 59808 97036 59872
rect 97100 59808 97116 59872
rect 97180 59808 97196 59872
rect 97260 59808 97276 59872
rect 97340 59808 97348 59872
rect 97028 58784 97348 59808
rect 97028 58720 97036 58784
rect 97100 58720 97116 58784
rect 97180 58720 97196 58784
rect 97260 58720 97276 58784
rect 97340 58720 97348 58784
rect 97028 57696 97348 58720
rect 97028 57632 97036 57696
rect 97100 57632 97116 57696
rect 97180 57632 97196 57696
rect 97260 57632 97276 57696
rect 97340 57632 97348 57696
rect 97028 56608 97348 57632
rect 97028 56544 97036 56608
rect 97100 56544 97116 56608
rect 97180 56544 97196 56608
rect 97260 56544 97276 56608
rect 97340 56544 97348 56608
rect 97028 55520 97348 56544
rect 97028 55456 97036 55520
rect 97100 55456 97116 55520
rect 97180 55456 97196 55520
rect 97260 55456 97276 55520
rect 97340 55456 97348 55520
rect 97028 54432 97348 55456
rect 97028 54368 97036 54432
rect 97100 54368 97116 54432
rect 97180 54368 97196 54432
rect 97260 54368 97276 54432
rect 97340 54368 97348 54432
rect 97028 53344 97348 54368
rect 97028 53280 97036 53344
rect 97100 53280 97116 53344
rect 97180 53280 97196 53344
rect 97260 53280 97276 53344
rect 97340 53280 97348 53344
rect 97028 52256 97348 53280
rect 97028 52192 97036 52256
rect 97100 52192 97116 52256
rect 97180 52192 97196 52256
rect 97260 52192 97276 52256
rect 97340 52192 97348 52256
rect 97028 51168 97348 52192
rect 97028 51104 97036 51168
rect 97100 51104 97116 51168
rect 97180 51104 97196 51168
rect 97260 51104 97276 51168
rect 97340 51104 97348 51168
rect 97028 50080 97348 51104
rect 97028 50016 97036 50080
rect 97100 50016 97116 50080
rect 97180 50016 97196 50080
rect 97260 50016 97276 50080
rect 97340 50016 97348 50080
rect 97028 48992 97348 50016
rect 97028 48928 97036 48992
rect 97100 48928 97116 48992
rect 97180 48928 97196 48992
rect 97260 48928 97276 48992
rect 97340 48928 97348 48992
rect 97028 47904 97348 48928
rect 97028 47840 97036 47904
rect 97100 47840 97116 47904
rect 97180 47840 97196 47904
rect 97260 47840 97276 47904
rect 97340 47840 97348 47904
rect 97028 46816 97348 47840
rect 97028 46752 97036 46816
rect 97100 46752 97116 46816
rect 97180 46752 97196 46816
rect 97260 46752 97276 46816
rect 97340 46752 97348 46816
rect 97028 45728 97348 46752
rect 97028 45664 97036 45728
rect 97100 45664 97116 45728
rect 97180 45664 97196 45728
rect 97260 45664 97276 45728
rect 97340 45664 97348 45728
rect 97028 44640 97348 45664
rect 97028 44576 97036 44640
rect 97100 44576 97116 44640
rect 97180 44576 97196 44640
rect 97260 44576 97276 44640
rect 97340 44576 97348 44640
rect 97028 43552 97348 44576
rect 97028 43488 97036 43552
rect 97100 43488 97116 43552
rect 97180 43488 97196 43552
rect 97260 43488 97276 43552
rect 97340 43488 97348 43552
rect 97028 42464 97348 43488
rect 97028 42400 97036 42464
rect 97100 42400 97116 42464
rect 97180 42400 97196 42464
rect 97260 42400 97276 42464
rect 97340 42400 97348 42464
rect 97028 41376 97348 42400
rect 97028 41312 97036 41376
rect 97100 41312 97116 41376
rect 97180 41312 97196 41376
rect 97260 41312 97276 41376
rect 97340 41312 97348 41376
rect 97028 40288 97348 41312
rect 97028 40224 97036 40288
rect 97100 40224 97116 40288
rect 97180 40224 97196 40288
rect 97260 40224 97276 40288
rect 97340 40224 97348 40288
rect 97028 39200 97348 40224
rect 97028 39136 97036 39200
rect 97100 39136 97116 39200
rect 97180 39136 97196 39200
rect 97260 39136 97276 39200
rect 97340 39136 97348 39200
rect 97028 38112 97348 39136
rect 97028 38048 97036 38112
rect 97100 38048 97116 38112
rect 97180 38048 97196 38112
rect 97260 38048 97276 38112
rect 97340 38048 97348 38112
rect 97028 37024 97348 38048
rect 97028 36960 97036 37024
rect 97100 36960 97116 37024
rect 97180 36960 97196 37024
rect 97260 36960 97276 37024
rect 97340 36960 97348 37024
rect 97028 36920 97348 36960
rect 97028 36684 97070 36920
rect 97306 36684 97348 36920
rect 97028 35936 97348 36684
rect 97028 35872 97036 35936
rect 97100 35872 97116 35936
rect 97180 35872 97196 35936
rect 97260 35872 97276 35936
rect 97340 35872 97348 35936
rect 97028 34848 97348 35872
rect 97028 34784 97036 34848
rect 97100 34784 97116 34848
rect 97180 34784 97196 34848
rect 97260 34784 97276 34848
rect 97340 34784 97348 34848
rect 97028 33760 97348 34784
rect 97028 33696 97036 33760
rect 97100 33696 97116 33760
rect 97180 33696 97196 33760
rect 97260 33696 97276 33760
rect 97340 33696 97348 33760
rect 97028 32672 97348 33696
rect 97028 32608 97036 32672
rect 97100 32608 97116 32672
rect 97180 32608 97196 32672
rect 97260 32608 97276 32672
rect 97340 32608 97348 32672
rect 97028 31584 97348 32608
rect 97028 31520 97036 31584
rect 97100 31520 97116 31584
rect 97180 31520 97196 31584
rect 97260 31520 97276 31584
rect 97340 31520 97348 31584
rect 97028 30496 97348 31520
rect 97028 30432 97036 30496
rect 97100 30432 97116 30496
rect 97180 30432 97196 30496
rect 97260 30432 97276 30496
rect 97340 30432 97348 30496
rect 97028 29408 97348 30432
rect 97028 29344 97036 29408
rect 97100 29344 97116 29408
rect 97180 29344 97196 29408
rect 97260 29344 97276 29408
rect 97340 29344 97348 29408
rect 97028 28320 97348 29344
rect 97028 28256 97036 28320
rect 97100 28256 97116 28320
rect 97180 28256 97196 28320
rect 97260 28256 97276 28320
rect 97340 28256 97348 28320
rect 97028 27232 97348 28256
rect 97028 27168 97036 27232
rect 97100 27168 97116 27232
rect 97180 27168 97196 27232
rect 97260 27168 97276 27232
rect 97340 27168 97348 27232
rect 97028 26144 97348 27168
rect 97028 26080 97036 26144
rect 97100 26080 97116 26144
rect 97180 26080 97196 26144
rect 97260 26080 97276 26144
rect 97340 26080 97348 26144
rect 97028 25056 97348 26080
rect 97028 24992 97036 25056
rect 97100 24992 97116 25056
rect 97180 24992 97196 25056
rect 97260 24992 97276 25056
rect 97340 24992 97348 25056
rect 97028 23968 97348 24992
rect 97028 23904 97036 23968
rect 97100 23904 97116 23968
rect 97180 23904 97196 23968
rect 97260 23904 97276 23968
rect 97340 23904 97348 23968
rect 97028 22880 97348 23904
rect 97028 22816 97036 22880
rect 97100 22816 97116 22880
rect 97180 22816 97196 22880
rect 97260 22816 97276 22880
rect 97340 22816 97348 22880
rect 97028 21792 97348 22816
rect 97028 21728 97036 21792
rect 97100 21728 97116 21792
rect 97180 21728 97196 21792
rect 97260 21728 97276 21792
rect 97340 21728 97348 21792
rect 97028 20704 97348 21728
rect 97028 20640 97036 20704
rect 97100 20640 97116 20704
rect 97180 20640 97196 20704
rect 97260 20640 97276 20704
rect 97340 20640 97348 20704
rect 97028 19616 97348 20640
rect 97028 19552 97036 19616
rect 97100 19552 97116 19616
rect 97180 19552 97196 19616
rect 97260 19552 97276 19616
rect 97340 19552 97348 19616
rect 97028 18528 97348 19552
rect 97028 18464 97036 18528
rect 97100 18464 97116 18528
rect 97180 18464 97196 18528
rect 97260 18464 97276 18528
rect 97340 18464 97348 18528
rect 97028 17440 97348 18464
rect 97028 17376 97036 17440
rect 97100 17376 97116 17440
rect 97180 17376 97196 17440
rect 97260 17376 97276 17440
rect 97340 17376 97348 17440
rect 97028 16352 97348 17376
rect 97028 16288 97036 16352
rect 97100 16288 97116 16352
rect 97180 16288 97196 16352
rect 97260 16288 97276 16352
rect 97340 16288 97348 16352
rect 97028 15264 97348 16288
rect 97028 15200 97036 15264
rect 97100 15200 97116 15264
rect 97180 15200 97196 15264
rect 97260 15200 97276 15264
rect 97340 15200 97348 15264
rect 97028 14176 97348 15200
rect 97028 14112 97036 14176
rect 97100 14112 97116 14176
rect 97180 14112 97196 14176
rect 97260 14112 97276 14176
rect 97340 14112 97348 14176
rect 97028 13088 97348 14112
rect 97028 13024 97036 13088
rect 97100 13024 97116 13088
rect 97180 13024 97196 13088
rect 97260 13024 97276 13088
rect 97340 13024 97348 13088
rect 97028 12000 97348 13024
rect 97028 11936 97036 12000
rect 97100 11936 97116 12000
rect 97180 11936 97196 12000
rect 97260 11936 97276 12000
rect 97340 11936 97348 12000
rect 97028 10912 97348 11936
rect 97028 10848 97036 10912
rect 97100 10848 97116 10912
rect 97180 10848 97196 10912
rect 97260 10848 97276 10912
rect 97340 10848 97348 10912
rect 97028 9824 97348 10848
rect 97028 9760 97036 9824
rect 97100 9760 97116 9824
rect 97180 9760 97196 9824
rect 97260 9760 97276 9824
rect 97340 9760 97348 9824
rect 97028 8736 97348 9760
rect 97028 8672 97036 8736
rect 97100 8672 97116 8736
rect 97180 8672 97196 8736
rect 97260 8672 97276 8736
rect 97340 8672 97348 8736
rect 97028 7648 97348 8672
rect 97028 7584 97036 7648
rect 97100 7584 97116 7648
rect 97180 7584 97196 7648
rect 97260 7584 97276 7648
rect 97340 7584 97348 7648
rect 97028 6560 97348 7584
rect 97028 6496 97036 6560
rect 97100 6496 97116 6560
rect 97180 6496 97196 6560
rect 97260 6496 97276 6560
rect 97340 6496 97348 6560
rect 97028 6284 97348 6496
rect 97028 6048 97070 6284
rect 97306 6048 97348 6284
rect 97028 5472 97348 6048
rect 97028 5408 97036 5472
rect 97100 5408 97116 5472
rect 97180 5408 97196 5472
rect 97260 5408 97276 5472
rect 97340 5408 97348 5472
rect 97028 4384 97348 5408
rect 97028 4320 97036 4384
rect 97100 4320 97116 4384
rect 97180 4320 97196 4384
rect 97260 4320 97276 4384
rect 97340 4320 97348 4384
rect 97028 3296 97348 4320
rect 97028 3232 97036 3296
rect 97100 3232 97116 3296
rect 97180 3232 97196 3296
rect 97260 3232 97276 3296
rect 97340 3232 97348 3296
rect 97028 2208 97348 3232
rect 97028 2144 97036 2208
rect 97100 2144 97116 2208
rect 97180 2144 97196 2208
rect 97260 2144 97276 2208
rect 97340 2144 97348 2208
rect 97028 274 97348 2144
rect 99088 97222 99408 97264
rect 99088 96986 99130 97222
rect 99366 96986 99408 97222
rect 99088 66896 99408 96986
rect 99088 66660 99130 66896
rect 99366 66660 99408 66896
rect 99088 36260 99408 66660
rect 99088 36024 99130 36260
rect 99366 36024 99408 36260
rect 99088 5624 99408 36024
rect 99088 5388 99130 5624
rect 99366 5388 99408 5624
rect 99088 934 99408 5388
rect 99088 698 99130 934
rect 99366 698 99408 934
rect 99088 656 99408 698
rect 99748 67556 100068 97646
rect 99748 67320 99790 67556
rect 100026 67320 100068 67556
rect 99748 36920 100068 67320
rect 99748 36684 99790 36920
rect 100026 36684 100068 36920
rect 99748 6284 100068 36684
rect 99748 6048 99790 6284
rect 100026 6048 100068 6284
rect 97028 38 97070 274
rect 97306 38 97348 274
rect 97028 -4 97348 38
rect 99748 274 100068 6048
rect 99748 38 99790 274
rect 100026 38 100068 274
rect 99748 -4 100068 38
<< via4 >>
rect -1034 97646 -798 97882
rect -1034 67320 -798 67556
rect -1034 36684 -798 36920
rect -1034 6048 -798 6284
rect -374 96986 -138 97222
rect -374 66660 -138 66896
rect -374 36024 -138 36260
rect -374 5388 -138 5624
rect -374 698 -138 934
rect 4250 96986 4486 97222
rect 4250 66880 4280 66896
rect 4280 66880 4296 66896
rect 4296 66880 4360 66896
rect 4360 66880 4376 66896
rect 4376 66880 4440 66896
rect 4440 66880 4456 66896
rect 4456 66880 4486 66896
rect 4250 66660 4486 66880
rect 4250 36024 4486 36260
rect 4250 5388 4486 5624
rect 4250 698 4486 934
rect -1034 38 -798 274
rect 4910 97646 5146 97882
rect 34970 96986 35206 97222
rect 35630 97646 35866 97882
rect 65690 96986 65926 97222
rect 66350 97646 66586 97882
rect 96410 96986 96646 97222
rect 12910 86684 13146 86920
rect 43630 86684 43866 86920
rect 12250 86024 12486 86260
rect 42970 86024 43206 86260
rect 4910 67488 5146 67556
rect 4910 67424 4940 67488
rect 4940 67424 4956 67488
rect 4956 67424 5020 67488
rect 5020 67424 5036 67488
rect 5036 67424 5100 67488
rect 5100 67424 5116 67488
rect 5116 67424 5146 67488
rect 4910 67320 5146 67424
rect 12910 67320 13146 67556
rect 43630 67320 43866 67556
rect 12250 66660 12486 66896
rect 42970 66660 43206 66896
rect 12910 56048 13146 56284
rect 43630 56048 43866 56284
rect 12250 55388 12486 55624
rect 42970 55388 43206 55624
rect 12910 44684 13146 44920
rect 43630 44684 43866 44920
rect 12250 44024 12486 44260
rect 42970 44024 43206 44260
rect 4910 36684 5146 36920
rect 12910 36684 13146 36920
rect 43630 36684 43866 36920
rect 12250 36024 12486 36260
rect 42970 36024 43206 36260
rect 12910 14048 13146 14284
rect 43630 14048 43866 14284
rect 12250 13388 12486 13624
rect 42970 13388 43206 13624
rect 54910 86684 55146 86920
rect 85630 86684 85866 86920
rect 54250 86024 54486 86260
rect 84970 86024 85206 86260
rect 54910 67320 55146 67556
rect 85630 67320 85866 67556
rect 54250 66660 54486 66896
rect 84970 66660 85206 66896
rect 96410 66880 96440 66896
rect 96440 66880 96456 66896
rect 96456 66880 96520 66896
rect 96520 66880 96536 66896
rect 96536 66880 96600 66896
rect 96600 66880 96616 66896
rect 96616 66880 96646 66896
rect 96410 66660 96646 66880
rect 54910 56048 55146 56284
rect 85630 56048 85866 56284
rect 54250 55388 54486 55624
rect 84970 55388 85206 55624
rect 54910 44684 55146 44920
rect 85630 44684 85866 44920
rect 54250 44024 54486 44260
rect 84970 44024 85206 44260
rect 54910 36684 55146 36920
rect 85630 36684 85866 36920
rect 54250 36024 54486 36260
rect 84970 36024 85206 36260
rect 96410 36024 96646 36260
rect 54910 14048 55146 14284
rect 85630 14048 85866 14284
rect 54250 13388 54486 13624
rect 84970 13388 85206 13624
rect 4910 6048 5146 6284
rect 4910 38 5146 274
rect 34970 5388 35206 5624
rect 34970 698 35206 934
rect 35630 6048 35866 6284
rect 35630 38 35866 274
rect 65690 5388 65926 5624
rect 65690 698 65926 934
rect 66350 6048 66586 6284
rect 66350 38 66586 274
rect 96410 5388 96646 5624
rect 96410 698 96646 934
rect 97070 97646 97306 97882
rect 99790 97646 100026 97882
rect 97070 67488 97306 67556
rect 97070 67424 97100 67488
rect 97100 67424 97116 67488
rect 97116 67424 97180 67488
rect 97180 67424 97196 67488
rect 97196 67424 97260 67488
rect 97260 67424 97276 67488
rect 97276 67424 97306 67488
rect 97070 67320 97306 67424
rect 97070 36684 97306 36920
rect 97070 6048 97306 6284
rect 99130 96986 99366 97222
rect 99130 66660 99366 66896
rect 99130 36024 99366 36260
rect 99130 5388 99366 5624
rect 99130 698 99366 934
rect 99790 67320 100026 67556
rect 99790 36684 100026 36920
rect 99790 6048 100026 6284
rect 97070 38 97306 274
rect 99790 38 100026 274
<< metal5 >>
rect -1076 97882 100068 97924
rect -1076 97646 -1034 97882
rect -798 97646 4910 97882
rect 5146 97646 35630 97882
rect 35866 97646 66350 97882
rect 66586 97646 97070 97882
rect 97306 97646 99790 97882
rect 100026 97646 100068 97882
rect -1076 97604 100068 97646
rect -416 97222 99408 97264
rect -416 96986 -374 97222
rect -138 96986 4250 97222
rect 4486 96986 34970 97222
rect 35206 96986 65690 97222
rect 65926 96986 96410 97222
rect 96646 96986 99130 97222
rect 99366 96986 99408 97222
rect -416 96944 99408 96986
rect 12886 86920 13170 86962
rect 12886 86684 12910 86920
rect 13146 86684 13170 86920
rect 12886 86642 13170 86684
rect 43606 86920 43890 86962
rect 43606 86684 43630 86920
rect 43866 86684 43890 86920
rect 43606 86642 43890 86684
rect 54886 86920 55170 86962
rect 54886 86684 54910 86920
rect 55146 86684 55170 86920
rect 54886 86642 55170 86684
rect 85606 86920 85890 86962
rect 85606 86684 85630 86920
rect 85866 86684 85890 86920
rect 85606 86642 85890 86684
rect 12226 86260 12510 86302
rect 12226 86024 12250 86260
rect 12486 86024 12510 86260
rect 12226 85982 12510 86024
rect 42946 86260 43230 86302
rect 42946 86024 42970 86260
rect 43206 86024 43230 86260
rect 42946 85982 43230 86024
rect 54226 86260 54510 86302
rect 54226 86024 54250 86260
rect 54486 86024 54510 86260
rect 54226 85982 54510 86024
rect 84946 86260 85230 86302
rect 84946 86024 84970 86260
rect 85206 86024 85230 86260
rect 84946 85982 85230 86024
rect -1076 67556 100068 67598
rect -1076 67320 -1034 67556
rect -798 67320 4910 67556
rect 5146 67320 12910 67556
rect 13146 67320 43630 67556
rect 43866 67320 54910 67556
rect 55146 67320 85630 67556
rect 85866 67320 97070 67556
rect 97306 67320 99790 67556
rect 100026 67320 100068 67556
rect -1076 67278 100068 67320
rect -1076 66896 100068 66938
rect -1076 66660 -374 66896
rect -138 66660 4250 66896
rect 4486 66660 12250 66896
rect 12486 66660 42970 66896
rect 43206 66660 54250 66896
rect 54486 66660 84970 66896
rect 85206 66660 96410 66896
rect 96646 66660 99130 66896
rect 99366 66660 100068 66896
rect -1076 66618 100068 66660
rect 12886 56284 13170 56326
rect 12886 56048 12910 56284
rect 13146 56048 13170 56284
rect 12886 56006 13170 56048
rect 43606 56284 43890 56326
rect 43606 56048 43630 56284
rect 43866 56048 43890 56284
rect 43606 56006 43890 56048
rect 54886 56284 55170 56326
rect 54886 56048 54910 56284
rect 55146 56048 55170 56284
rect 54886 56006 55170 56048
rect 85606 56284 85890 56326
rect 85606 56048 85630 56284
rect 85866 56048 85890 56284
rect 85606 56006 85890 56048
rect 12226 55624 12510 55666
rect 12226 55388 12250 55624
rect 12486 55388 12510 55624
rect 12226 55346 12510 55388
rect 42946 55624 43230 55666
rect 42946 55388 42970 55624
rect 43206 55388 43230 55624
rect 42946 55346 43230 55388
rect 54226 55624 54510 55666
rect 54226 55388 54250 55624
rect 54486 55388 54510 55624
rect 54226 55346 54510 55388
rect 84946 55624 85230 55666
rect 84946 55388 84970 55624
rect 85206 55388 85230 55624
rect 84946 55346 85230 55388
rect 12886 44920 13170 44962
rect 12886 44684 12910 44920
rect 13146 44684 13170 44920
rect 12886 44642 13170 44684
rect 43606 44920 43890 44962
rect 43606 44684 43630 44920
rect 43866 44684 43890 44920
rect 43606 44642 43890 44684
rect 54886 44920 55170 44962
rect 54886 44684 54910 44920
rect 55146 44684 55170 44920
rect 54886 44642 55170 44684
rect 85606 44920 85890 44962
rect 85606 44684 85630 44920
rect 85866 44684 85890 44920
rect 85606 44642 85890 44684
rect 12226 44260 12510 44302
rect 12226 44024 12250 44260
rect 12486 44024 12510 44260
rect 12226 43982 12510 44024
rect 42946 44260 43230 44302
rect 42946 44024 42970 44260
rect 43206 44024 43230 44260
rect 42946 43982 43230 44024
rect 54226 44260 54510 44302
rect 54226 44024 54250 44260
rect 54486 44024 54510 44260
rect 54226 43982 54510 44024
rect 84946 44260 85230 44302
rect 84946 44024 84970 44260
rect 85206 44024 85230 44260
rect 84946 43982 85230 44024
rect -1076 36920 100068 36962
rect -1076 36684 -1034 36920
rect -798 36684 4910 36920
rect 5146 36684 12910 36920
rect 13146 36684 43630 36920
rect 43866 36684 54910 36920
rect 55146 36684 85630 36920
rect 85866 36684 97070 36920
rect 97306 36684 99790 36920
rect 100026 36684 100068 36920
rect -1076 36642 100068 36684
rect -1076 36260 100068 36302
rect -1076 36024 -374 36260
rect -138 36024 4250 36260
rect 4486 36024 12250 36260
rect 12486 36024 42970 36260
rect 43206 36024 54250 36260
rect 54486 36024 84970 36260
rect 85206 36024 96410 36260
rect 96646 36024 99130 36260
rect 99366 36024 100068 36260
rect -1076 35982 100068 36024
rect 12886 14284 13170 14326
rect 12886 14048 12910 14284
rect 13146 14048 13170 14284
rect 12886 14006 13170 14048
rect 43606 14284 43890 14326
rect 43606 14048 43630 14284
rect 43866 14048 43890 14284
rect 43606 14006 43890 14048
rect 54886 14284 55170 14326
rect 54886 14048 54910 14284
rect 55146 14048 55170 14284
rect 54886 14006 55170 14048
rect 85606 14284 85890 14326
rect 85606 14048 85630 14284
rect 85866 14048 85890 14284
rect 85606 14006 85890 14048
rect 12226 13624 12510 13666
rect 12226 13388 12250 13624
rect 12486 13388 12510 13624
rect 12226 13346 12510 13388
rect 42946 13624 43230 13666
rect 42946 13388 42970 13624
rect 43206 13388 43230 13624
rect 42946 13346 43230 13388
rect 54226 13624 54510 13666
rect 54226 13388 54250 13624
rect 54486 13388 54510 13624
rect 54226 13346 54510 13388
rect 84946 13624 85230 13666
rect 84946 13388 84970 13624
rect 85206 13388 85230 13624
rect 84946 13346 85230 13388
rect -1076 6284 100068 6326
rect -1076 6048 -1034 6284
rect -798 6048 4910 6284
rect 5146 6048 35630 6284
rect 35866 6048 66350 6284
rect 66586 6048 97070 6284
rect 97306 6048 99790 6284
rect 100026 6048 100068 6284
rect -1076 6006 100068 6048
rect -1076 5624 100068 5666
rect -1076 5388 -374 5624
rect -138 5388 4250 5624
rect 4486 5388 34970 5624
rect 35206 5388 65690 5624
rect 65926 5388 96410 5624
rect 96646 5388 99130 5624
rect 99366 5388 100068 5624
rect -1076 5346 100068 5388
rect -416 934 99408 976
rect -416 698 -374 934
rect -138 698 4250 934
rect 4486 698 34970 934
rect 35206 698 65690 934
rect 65926 698 96410 934
rect 96646 698 99130 934
rect 99366 698 99408 934
rect -416 656 99408 698
rect -1076 274 100068 316
rect -1076 38 -1034 274
rect -798 38 4910 274
rect 5146 38 35630 274
rect 35866 38 66350 274
rect 66586 38 97070 274
rect 97306 38 99790 274
rect 100026 38 100068 274
rect -1076 -4 100068 38
use sky130_fd_sc_hd__diode_2  ANTENNA_cell0_clk
timestamp 18001
transform 1 0 5520 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell0_config_data_out
timestamp 18001
transform -1 0 9108 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell0_config_en
timestamp 18001
transform -1 0 5520 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell0_en
timestamp 18001
transform -1 0 5336 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell0_le_clk
timestamp 18001
transform 1 0 9936 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell0_le_en
timestamp 18001
transform 1 0 11040 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell0_le_nrst
timestamp 18001
transform 1 0 12144 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell0_nrst
timestamp 18001
transform -1 0 5704 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell1_clk
timestamp 18001
transform -1 0 51060 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell1_config_data_in
timestamp 18001
transform -1 0 94484 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell1_config_data_out
timestamp 18001
transform -1 0 51244 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell1_config_en
timestamp 18001
transform -1 0 94668 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell1_en
timestamp 18001
transform -1 0 94852 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell1_le_clk
timestamp 18001
transform 1 0 51980 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell1_le_en
timestamp 18001
transform 1 0 53084 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell1_le_nrst
timestamp 18001
transform 1 0 54188 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell1_nrst
timestamp 18001
transform -1 0 95036 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell2_clk
timestamp 18001
transform -1 0 9108 0 -1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell2_config_data_in
timestamp 18001
transform -1 0 13432 0 -1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell2_config_data_out
timestamp 18001
transform -1 0 5704 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell2_config_en
timestamp 18001
transform 1 0 12144 0 -1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell2_en
timestamp 18001
transform 1 0 9936 0 -1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell2_le_clk
timestamp 18001
transform -1 0 5520 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell2_le_en
timestamp 18001
transform -1 0 5336 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell2_le_nrst
timestamp 18001
transform -1 0 5704 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell2_nrst
timestamp 18001
transform 1 0 11040 0 -1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell3_clk
timestamp 18001
transform -1 0 51060 0 -1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell3_config_data_in
timestamp 18001
transform -1 0 55200 0 -1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell3_config_data_out
timestamp 18001
transform 1 0 51060 0 -1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell3_config_en
timestamp 18001
transform 1 0 54188 0 -1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell3_en
timestamp 18001
transform 1 0 51980 0 -1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell3_le_clk
timestamp 18001
transform -1 0 94484 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell3_le_en
timestamp 18001
transform -1 0 94668 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell3_le_nrst
timestamp 18001
transform -1 0 94852 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell3_nrst
timestamp 18001
transform 1 0 52256 0 -1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 18001
transform -1 0 31924 0 -1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_X
timestamp 18001
transform 1 0 32108 0 -1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0__f_clk_A
timestamp 18001
transform 1 0 5520 0 -1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0__f_clk_X
timestamp 18001
transform 1 0 5520 0 -1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1__f_clk_A
timestamp 18001
transform 1 0 40296 0 -1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1__f_clk_X
timestamp 18001
transform 1 0 42412 0 -1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 18001
transform -1 0 1932 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 18001
transform -1 0 55200 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_X
timestamp 18001
transform -1 0 56948 0 1 94656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 18001
transform -1 0 52900 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_X
timestamp 18001
transform -1 0 53084 0 1 94656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 18001
transform -1 0 97336 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 18001
transform -1 0 97336 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 18001
transform -1 0 97336 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 18001
transform -1 0 97336 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 18001
transform -1 0 97336 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 18001
transform -1 0 97336 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 18001
transform -1 0 97336 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 18001
transform -1 0 97336 0 1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 18001
transform -1 0 97612 0 1 71808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 18001
transform -1 0 97336 0 -1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 18001
transform -1 0 97244 0 1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 18001
transform -1 0 97612 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 18001
transform -1 0 97336 0 -1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 18001
transform -1 0 97336 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 18001
transform -1 0 97336 0 -1 78336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 18001
transform -1 0 97244 0 -1 79424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 18001
transform -1 0 97336 0 1 79424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 18001
transform -1 0 97336 0 -1 81600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 18001
transform -1 0 97336 0 1 81600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 18001
transform -1 0 97336 0 -1 83776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 18001
transform -1 0 97336 0 -1 84864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 18001
transform -1 0 97336 0 1 84864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 18001
transform -1 0 97336 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 18001
transform -1 0 97336 0 -1 87040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 18001
transform -1 0 97336 0 1 87040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 18001
transform -1 0 97244 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 18001
transform -1 0 97336 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 18001
transform -1 0 97336 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 18001
transform -1 0 97336 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 18001
transform -1 0 97244 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 18001
transform -1 0 97336 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 18001
transform -1 0 97336 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 18001
transform -1 0 14260 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 18001
transform -1 0 25208 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 18001
transform -1 0 26496 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 18001
transform -1 0 27784 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 18001
transform -1 0 29072 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 18001
transform -1 0 29716 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 18001
transform -1 0 31004 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 18001
transform -1 0 57316 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 18001
transform -1 0 58052 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 18001
transform -1 0 58696 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 18001
transform -1 0 59984 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 18001
transform -1 0 15548 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 18001
transform -1 0 60628 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 18001
transform -1 0 61916 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 18001
transform -1 0 63204 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 18001
transform -1 0 63848 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 18001
transform -1 0 65136 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 18001
transform -1 0 66424 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 18001
transform -1 0 68080 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 18001
transform -1 0 69552 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 18001
transform -1 0 70104 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 18001
transform -1 0 70932 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 18001
transform -1 0 16836 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 18001
transform -1 0 71576 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 18001
transform -1 0 72864 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 18001
transform -1 0 17480 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 18001
transform -1 0 18768 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 18001
transform -1 0 20056 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 18001
transform -1 0 21344 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 18001
transform -1 0 21988 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 18001
transform -1 0 23276 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 18001
transform -1 0 24564 0 1 94656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 18001
transform -1 0 32292 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 18001
transform -1 0 43240 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 18001
transform -1 0 44528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 18001
transform -1 0 45172 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 18001
transform -1 0 46460 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 18001
transform -1 0 47748 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 18001
transform -1 0 49220 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 18001
transform -1 0 74152 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 18001
transform -1 0 75440 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input77_A
timestamp 18001
transform -1 0 76084 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input78_A
timestamp 18001
transform -1 0 77372 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 18001
transform -1 0 32936 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 18001
transform -1 0 78660 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input81_A
timestamp 18001
transform -1 0 79304 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input82_A
timestamp 18001
transform -1 0 80592 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input83_A
timestamp 18001
transform -1 0 81880 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input84_A
timestamp 18001
transform -1 0 83168 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input85_A
timestamp 18001
transform -1 0 83812 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input86_A
timestamp 18001
transform -1 0 85100 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input87_A
timestamp 18001
transform -1 0 86388 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input88_A
timestamp 18001
transform -1 0 87032 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input89_A
timestamp 18001
transform -1 0 88688 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input90_A
timestamp 18001
transform -1 0 34224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input91_A
timestamp 18001
transform -1 0 89700 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input92_A
timestamp 18001
transform -1 0 97244 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input93_A
timestamp 18001
transform -1 0 35512 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input94_A
timestamp 18001
transform -1 0 36800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input95_A
timestamp 18001
transform -1 0 37444 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input96_A
timestamp 18001
transform -1 0 38732 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input97_A
timestamp 18001
transform -1 0 40020 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input98_A
timestamp 18001
transform -1 0 40664 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input99_A
timestamp 18001
transform -1 0 41952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input100_A
timestamp 18001
transform -1 0 1932 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input101_A
timestamp 18001
transform -1 0 1932 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input102_A
timestamp 18001
transform -1 0 1932 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input103_A
timestamp 18001
transform -1 0 1932 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input104_A
timestamp 18001
transform -1 0 1932 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input105_A
timestamp 18001
transform -1 0 1932 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input106_A
timestamp 18001
transform -1 0 1840 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input107_A
timestamp 18001
transform -1 0 1932 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input108_A
timestamp 18001
transform -1 0 1932 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input109_A
timestamp 18001
transform -1 0 2116 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input110_A
timestamp 18001
transform -1 0 2116 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input111_A
timestamp 18001
transform -1 0 1932 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input112_A
timestamp 18001
transform -1 0 1932 0 1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input113_A
timestamp 18001
transform -1 0 1932 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input114_A
timestamp 18001
transform -1 0 2116 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input115_A
timestamp 18001
transform -1 0 1932 0 -1 62016
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input116_A
timestamp 18001
transform -1 0 2116 0 -1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input117_A
timestamp 18001
transform -1 0 1932 0 1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input118_A
timestamp 18001
transform -1 0 1932 0 -1 65280
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input119_A
timestamp 18001
transform -1 0 1932 0 1 65280
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input120_A
timestamp 18001
transform -1 0 1932 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input121_A
timestamp 18001
transform -1 0 1932 0 -1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input122_A
timestamp 18001
transform -1 0 2116 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input123_A
timestamp 18001
transform -1 0 1932 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input124_A
timestamp 18001
transform -1 0 1840 0 -1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input125_A
timestamp 18001
transform -1 0 2116 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input126_A
timestamp 18001
transform -1 0 1932 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input127_A
timestamp 18001
transform -1 0 1932 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input128_A
timestamp 18001
transform -1 0 2116 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input129_A
timestamp 18001
transform -1 0 1932 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input130_A
timestamp 18001
transform -1 0 2116 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input131_A
timestamp 18001
transform -1 0 1932 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input132_A
timestamp 18001
transform -1 0 11960 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input132_X
timestamp 18001
transform 1 0 11592 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input133_A
timestamp 18001
transform -1 0 11684 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input133_X
timestamp 18001
transform -1 0 13340 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input134_A
timestamp 18001
transform -1 0 12328 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input134_X
timestamp 18001
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input135_A
timestamp 18001
transform -1 0 52900 0 1 94656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input135_X
timestamp 18001
transform 1 0 54372 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_max_cap265_A
timestamp 18001
transform 1 0 52440 0 -1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_max_cap265_X
timestamp 18001
transform 1 0 54372 0 -1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_max_cap266_A
timestamp 18001
transform -1 0 56948 0 -1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_max_cap266_X
timestamp 18001
transform 1 0 56948 0 -1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_max_cap267_A
timestamp 18001
transform -1 0 54740 0 1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_max_cap267_X
timestamp 18001
transform -1 0 54924 0 1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output136_A
timestamp 18001
transform -1 0 51336 0 1 94656
box -38 -48 222 592
use fpgacell  cell0
timestamp 0
transform 1 0 8000 0 1 8000
box 0 0 42000 41000
use fpgacell  cell1
timestamp 0
transform 1 0 50000 0 1 8000
box 0 0 42000 41000
use fpgacell  cell2
timestamp 0
transform 1 0 8000 0 1 50000
box 0 0 42000 41000
use fpgacell  cell3
timestamp 0
transform 1 0 50000 0 1 50000
box 0 0 42000 41000
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 18001
transform -1 0 31740 0 -1 93568
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 18001
transform -1 0 5704 0 1 69632
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 18001
transform 1 0 40480 0 -1 93568
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3
timestamp 1636986456
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1636986456
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp 18001
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1636986456
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1636986456
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp 18001
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1636986456
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1636986456
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 18001
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85
timestamp 18001
transform 1 0 8924 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_93
timestamp 18001
transform 1 0 9660 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113
timestamp 18001
transform 1 0 11500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_118
timestamp 18001
transform 1 0 11960 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 18001
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_147
timestamp 18001
transform 1 0 14628 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_155
timestamp 18001
transform 1 0 15364 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_161
timestamp 18001
transform 1 0 15916 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 18001
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 18001
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_175
timestamp 18001
transform 1 0 17204 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_182
timestamp 18001
transform 1 0 17848 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_190
timestamp 18001
transform 1 0 18584 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_197
timestamp 18001
transform 1 0 19228 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_205
timestamp 18001
transform 1 0 19964 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_210
timestamp 18001
transform 1 0 20424 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_218
timestamp 18001
transform 1 0 21160 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 18001
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_231
timestamp 18001
transform 1 0 22356 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_239
timestamp 18001
transform 1 0 23092 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_245
timestamp 18001
transform 1 0 23644 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 18001
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 18001
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_259
timestamp 18001
transform 1 0 24932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_266
timestamp 18001
transform 1 0 25576 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_274
timestamp 18001
transform 1 0 26312 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_281
timestamp 18001
transform 1 0 26956 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_289
timestamp 18001
transform 1 0 27692 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_294
timestamp 18001
transform 1 0 28152 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_302
timestamp 18001
transform 1 0 28888 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 18001
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_315
timestamp 18001
transform 1 0 30084 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_323
timestamp 18001
transform 1 0 30820 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_329
timestamp 18001
transform 1 0 31372 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_335
timestamp 18001
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_342
timestamp 18001
transform 1 0 32568 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_349
timestamp 18001
transform 1 0 33212 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_357
timestamp 18001
transform 1 0 33948 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 18001
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_365
timestamp 18001
transform 1 0 34684 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_371
timestamp 18001
transform 1 0 35236 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_377
timestamp 18001
transform 1 0 35788 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_385
timestamp 18001
transform 1 0 36524 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_391
timestamp 18001
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_398
timestamp 18001
transform 1 0 37720 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_406
timestamp 18001
transform 1 0 38456 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_412
timestamp 18001
transform 1 0 39008 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_426
timestamp 18001
transform 1 0 40296 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_433
timestamp 18001
transform 1 0 40940 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_441
timestamp 18001
transform 1 0 41676 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_447
timestamp 18001
transform 1 0 42228 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_449
timestamp 18001
transform 1 0 42412 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_455
timestamp 18001
transform 1 0 42964 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_461
timestamp 18001
transform 1 0 43516 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_469
timestamp 18001
transform 1 0 44252 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_489
timestamp 18001
transform 1 0 46092 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_503
timestamp 18001
transform 1 0 47380 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_523
timestamp 18001
transform 1 0 49220 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_531
timestamp 18001
transform 1 0 49956 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_533
timestamp 1636986456
transform 1 0 50140 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_545
timestamp 1636986456
transform 1 0 51244 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_557
timestamp 18001
transform 1 0 52348 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_561
timestamp 1636986456
transform 1 0 52716 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_573
timestamp 1636986456
transform 1 0 53820 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_585
timestamp 18001
transform 1 0 54924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_589
timestamp 18001
transform 1 0 55292 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_597
timestamp 18001
transform 1 0 56028 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_602
timestamp 18001
transform 1 0 56488 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_610
timestamp 18001
transform 1 0 57224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_617
timestamp 18001
transform 1 0 57868 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_625
timestamp 18001
transform 1 0 58604 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_630
timestamp 18001
transform 1 0 59064 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_638
timestamp 18001
transform 1 0 59800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_645
timestamp 18001
transform 1 0 60444 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_651
timestamp 18001
transform 1 0 60996 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_659
timestamp 18001
transform 1 0 61732 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_665
timestamp 18001
transform 1 0 62284 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_671
timestamp 18001
transform 1 0 62836 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_673
timestamp 18001
transform 1 0 63020 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_679
timestamp 18001
transform 1 0 63572 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_686
timestamp 18001
transform 1 0 64216 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_694
timestamp 18001
transform 1 0 64952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_701
timestamp 18001
transform 1 0 65596 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_709
timestamp 18001
transform 1 0 66332 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_714
timestamp 18001
transform 1 0 66792 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_722
timestamp 18001
transform 1 0 67528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_729
timestamp 18001
transform 1 0 68172 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_735
timestamp 18001
transform 1 0 68724 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_743
timestamp 18001
transform 1 0 69460 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_749
timestamp 18001
transform 1 0 70012 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_755
timestamp 18001
transform 1 0 70564 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_757
timestamp 18001
transform 1 0 70748 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_763
timestamp 18001
transform 1 0 71300 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_770
timestamp 18001
transform 1 0 71944 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_778
timestamp 18001
transform 1 0 72680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_785
timestamp 18001
transform 1 0 73324 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_791
timestamp 18001
transform 1 0 73876 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_797
timestamp 18001
transform 1 0 74428 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_805
timestamp 18001
transform 1 0 75164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_811
timestamp 18001
transform 1 0 75716 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_818
timestamp 18001
transform 1 0 76360 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_826
timestamp 18001
transform 1 0 77096 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_832
timestamp 18001
transform 1 0 77648 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_846
timestamp 18001
transform 1 0 78936 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_853
timestamp 18001
transform 1 0 79580 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_861
timestamp 18001
transform 1 0 80316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_867
timestamp 18001
transform 1 0 80868 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_869
timestamp 18001
transform 1 0 81052 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_875
timestamp 18001
transform 1 0 81604 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_881
timestamp 18001
transform 1 0 82156 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_889
timestamp 18001
transform 1 0 82892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_895
timestamp 18001
transform 1 0 83444 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_902
timestamp 18001
transform 1 0 84088 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_910
timestamp 18001
transform 1 0 84824 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_916
timestamp 18001
transform 1 0 85376 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_931
timestamp 18001
transform 1 0 86756 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_944
timestamp 18001
transform 1 0 87952 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_973
timestamp 18001
transform 1 0 90620 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_979
timestamp 18001
transform 1 0 91172 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_981
timestamp 1636986456
transform 1 0 91356 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_993
timestamp 1636986456
transform 1 0 92460 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1005
timestamp 18001
transform 1 0 93564 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1009
timestamp 1636986456
transform 1 0 93932 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1021
timestamp 1636986456
transform 1 0 95036 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1033
timestamp 18001
transform 1 0 96140 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1037
timestamp 1636986456
transform 1 0 96508 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1636986456
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1636986456
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1636986456
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1636986456
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 18001
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 18001
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1636986456
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1636986456
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1636986456
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1636986456
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 18001
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 18001
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_133
timestamp 1636986456
transform 1 0 13340 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_145
timestamp 1636986456
transform 1 0 14444 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_157
timestamp 18001
transform 1 0 15548 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_165
timestamp 18001
transform 1 0 16284 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1636986456
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1636986456
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1636986456
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1636986456
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 18001
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 18001
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1636986456
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1636986456
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1636986456
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1636986456
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 18001
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 18001
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1636986456
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1636986456
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1636986456
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1636986456
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 18001
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 18001
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1636986456
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1636986456
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1636986456
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1636986456
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 18001
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 18001
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1636986456
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_405
timestamp 1636986456
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_417
timestamp 1636986456
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_429
timestamp 1636986456
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 18001
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 18001
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_449
timestamp 1636986456
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_461
timestamp 1636986456
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_473
timestamp 1636986456
transform 1 0 44620 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_485
timestamp 1636986456
transform 1 0 45724 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_497
timestamp 18001
transform 1 0 46828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 18001
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_505
timestamp 1636986456
transform 1 0 47564 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_517
timestamp 1636986456
transform 1 0 48668 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_529
timestamp 1636986456
transform 1 0 49772 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_541
timestamp 1636986456
transform 1 0 50876 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_553
timestamp 18001
transform 1 0 51980 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_559
timestamp 18001
transform 1 0 52532 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_561
timestamp 1636986456
transform 1 0 52716 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_573
timestamp 1636986456
transform 1 0 53820 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_585
timestamp 1636986456
transform 1 0 54924 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_597
timestamp 1636986456
transform 1 0 56028 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_609
timestamp 18001
transform 1 0 57132 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_615
timestamp 18001
transform 1 0 57684 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_617
timestamp 1636986456
transform 1 0 57868 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_629
timestamp 1636986456
transform 1 0 58972 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_641
timestamp 1636986456
transform 1 0 60076 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_653
timestamp 1636986456
transform 1 0 61180 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_665
timestamp 18001
transform 1 0 62284 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_671
timestamp 18001
transform 1 0 62836 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_673
timestamp 1636986456
transform 1 0 63020 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_685
timestamp 1636986456
transform 1 0 64124 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_697
timestamp 1636986456
transform 1 0 65228 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_709
timestamp 1636986456
transform 1 0 66332 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_721
timestamp 18001
transform 1 0 67436 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_727
timestamp 18001
transform 1 0 67988 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_729
timestamp 1636986456
transform 1 0 68172 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_741
timestamp 1636986456
transform 1 0 69276 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_753
timestamp 1636986456
transform 1 0 70380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_765
timestamp 1636986456
transform 1 0 71484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_777
timestamp 18001
transform 1 0 72588 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_783
timestamp 18001
transform 1 0 73140 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_785
timestamp 1636986456
transform 1 0 73324 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_797
timestamp 1636986456
transform 1 0 74428 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_809
timestamp 1636986456
transform 1 0 75532 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_821
timestamp 1636986456
transform 1 0 76636 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_833
timestamp 18001
transform 1 0 77740 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_839
timestamp 18001
transform 1 0 78292 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_841
timestamp 1636986456
transform 1 0 78476 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_853
timestamp 1636986456
transform 1 0 79580 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_865
timestamp 1636986456
transform 1 0 80684 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_877
timestamp 1636986456
transform 1 0 81788 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_889
timestamp 18001
transform 1 0 82892 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_895
timestamp 18001
transform 1 0 83444 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_897
timestamp 1636986456
transform 1 0 83628 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_909
timestamp 1636986456
transform 1 0 84732 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_921
timestamp 1636986456
transform 1 0 85836 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_933
timestamp 1636986456
transform 1 0 86940 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_945
timestamp 18001
transform 1 0 88044 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_951
timestamp 18001
transform 1 0 88596 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_953
timestamp 18001
transform 1 0 88780 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_963
timestamp 1636986456
transform 1 0 89700 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_975
timestamp 1636986456
transform 1 0 90804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_987
timestamp 1636986456
transform 1 0 91908 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_999
timestamp 18001
transform 1 0 93012 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1007
timestamp 18001
transform 1 0 93748 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1009
timestamp 1636986456
transform 1 0 93932 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1021
timestamp 1636986456
transform 1 0 95036 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1033
timestamp 1636986456
transform 1 0 96140 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1045
timestamp 18001
transform 1 0 97244 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1636986456
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1636986456
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 18001
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1636986456
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1636986456
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1636986456
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1636986456
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 18001
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 18001
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1636986456
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1636986456
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1636986456
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1636986456
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 18001
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 18001
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1636986456
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1636986456
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1636986456
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1636986456
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 18001
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 18001
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1636986456
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1636986456
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1636986456
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1636986456
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 18001
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 18001
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1636986456
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1636986456
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1636986456
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1636986456
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 18001
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 18001
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1636986456
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1636986456
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1636986456
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1636986456
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 18001
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 18001
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1636986456
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1636986456
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1636986456
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1636986456
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 18001
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 18001
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1636986456
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1636986456
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 1636986456
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_457
timestamp 1636986456
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 18001
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 18001
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_477
timestamp 1636986456
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_489
timestamp 1636986456
transform 1 0 46092 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_501
timestamp 1636986456
transform 1 0 47196 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_513
timestamp 1636986456
transform 1 0 48300 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_525
timestamp 18001
transform 1 0 49404 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 18001
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_533
timestamp 1636986456
transform 1 0 50140 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_545
timestamp 1636986456
transform 1 0 51244 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_557
timestamp 1636986456
transform 1 0 52348 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_569
timestamp 1636986456
transform 1 0 53452 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_581
timestamp 18001
transform 1 0 54556 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 18001
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_589
timestamp 1636986456
transform 1 0 55292 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_601
timestamp 1636986456
transform 1 0 56396 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_613
timestamp 1636986456
transform 1 0 57500 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_625
timestamp 1636986456
transform 1 0 58604 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_637
timestamp 18001
transform 1 0 59708 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_643
timestamp 18001
transform 1 0 60260 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_645
timestamp 1636986456
transform 1 0 60444 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_657
timestamp 1636986456
transform 1 0 61548 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_669
timestamp 1636986456
transform 1 0 62652 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_681
timestamp 1636986456
transform 1 0 63756 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_693
timestamp 18001
transform 1 0 64860 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_699
timestamp 18001
transform 1 0 65412 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_701
timestamp 1636986456
transform 1 0 65596 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_713
timestamp 1636986456
transform 1 0 66700 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_725
timestamp 1636986456
transform 1 0 67804 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_737
timestamp 1636986456
transform 1 0 68908 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_749
timestamp 18001
transform 1 0 70012 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_755
timestamp 18001
transform 1 0 70564 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_757
timestamp 1636986456
transform 1 0 70748 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_769
timestamp 1636986456
transform 1 0 71852 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_781
timestamp 1636986456
transform 1 0 72956 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_793
timestamp 1636986456
transform 1 0 74060 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_805
timestamp 18001
transform 1 0 75164 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_811
timestamp 18001
transform 1 0 75716 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_813
timestamp 1636986456
transform 1 0 75900 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_825
timestamp 1636986456
transform 1 0 77004 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_837
timestamp 1636986456
transform 1 0 78108 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_849
timestamp 1636986456
transform 1 0 79212 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_861
timestamp 18001
transform 1 0 80316 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_867
timestamp 18001
transform 1 0 80868 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_869
timestamp 1636986456
transform 1 0 81052 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_881
timestamp 1636986456
transform 1 0 82156 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_893
timestamp 1636986456
transform 1 0 83260 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_905
timestamp 1636986456
transform 1 0 84364 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_917
timestamp 18001
transform 1 0 85468 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_923
timestamp 18001
transform 1 0 86020 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_925
timestamp 1636986456
transform 1 0 86204 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_937
timestamp 1636986456
transform 1 0 87308 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_949
timestamp 1636986456
transform 1 0 88412 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_961
timestamp 1636986456
transform 1 0 89516 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_973
timestamp 18001
transform 1 0 90620 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_979
timestamp 18001
transform 1 0 91172 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_981
timestamp 1636986456
transform 1 0 91356 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_993
timestamp 1636986456
transform 1 0 92460 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1005
timestamp 1636986456
transform 1 0 93564 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1017
timestamp 1636986456
transform 1 0 94668 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1029
timestamp 18001
transform 1 0 95772 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1035
timestamp 18001
transform 1 0 96324 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1037
timestamp 1636986456
transform 1 0 96508 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1636986456
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1636986456
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1636986456
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1636986456
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 18001
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 18001
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1636986456
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1636986456
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1636986456
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1636986456
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 18001
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 18001
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1636986456
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1636986456
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1636986456
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1636986456
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 18001
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 18001
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1636986456
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1636986456
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1636986456
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1636986456
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 18001
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 18001
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1636986456
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1636986456
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1636986456
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1636986456
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 18001
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 18001
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1636986456
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1636986456
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1636986456
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1636986456
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 18001
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 18001
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1636986456
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1636986456
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1636986456
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1636986456
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 18001
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 18001
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1636986456
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1636986456
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1636986456
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1636986456
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 18001
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 18001
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1636986456
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1636986456
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1636986456
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1636986456
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 18001
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 18001
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_505
timestamp 1636986456
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_517
timestamp 1636986456
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_529
timestamp 1636986456
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_541
timestamp 1636986456
transform 1 0 50876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_553
timestamp 18001
transform 1 0 51980 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 18001
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_561
timestamp 1636986456
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_573
timestamp 1636986456
transform 1 0 53820 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_585
timestamp 1636986456
transform 1 0 54924 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_597
timestamp 1636986456
transform 1 0 56028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_609
timestamp 18001
transform 1 0 57132 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 18001
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_617
timestamp 1636986456
transform 1 0 57868 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_629
timestamp 1636986456
transform 1 0 58972 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_641
timestamp 1636986456
transform 1 0 60076 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_653
timestamp 1636986456
transform 1 0 61180 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_665
timestamp 18001
transform 1 0 62284 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_671
timestamp 18001
transform 1 0 62836 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_673
timestamp 1636986456
transform 1 0 63020 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_685
timestamp 1636986456
transform 1 0 64124 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_697
timestamp 1636986456
transform 1 0 65228 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_709
timestamp 1636986456
transform 1 0 66332 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_721
timestamp 18001
transform 1 0 67436 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_727
timestamp 18001
transform 1 0 67988 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_729
timestamp 1636986456
transform 1 0 68172 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_741
timestamp 1636986456
transform 1 0 69276 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_753
timestamp 1636986456
transform 1 0 70380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_765
timestamp 1636986456
transform 1 0 71484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_777
timestamp 18001
transform 1 0 72588 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_783
timestamp 18001
transform 1 0 73140 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_785
timestamp 1636986456
transform 1 0 73324 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_797
timestamp 1636986456
transform 1 0 74428 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_809
timestamp 1636986456
transform 1 0 75532 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_821
timestamp 1636986456
transform 1 0 76636 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_833
timestamp 18001
transform 1 0 77740 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_839
timestamp 18001
transform 1 0 78292 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_841
timestamp 1636986456
transform 1 0 78476 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_853
timestamp 1636986456
transform 1 0 79580 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_865
timestamp 1636986456
transform 1 0 80684 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_877
timestamp 1636986456
transform 1 0 81788 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_889
timestamp 18001
transform 1 0 82892 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_895
timestamp 18001
transform 1 0 83444 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_897
timestamp 1636986456
transform 1 0 83628 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_909
timestamp 1636986456
transform 1 0 84732 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_921
timestamp 1636986456
transform 1 0 85836 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_933
timestamp 1636986456
transform 1 0 86940 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_945
timestamp 18001
transform 1 0 88044 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_951
timestamp 18001
transform 1 0 88596 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_953
timestamp 1636986456
transform 1 0 88780 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_965
timestamp 1636986456
transform 1 0 89884 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_977
timestamp 1636986456
transform 1 0 90988 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_989
timestamp 1636986456
transform 1 0 92092 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1001
timestamp 18001
transform 1 0 93196 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1007
timestamp 18001
transform 1 0 93748 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1009
timestamp 1636986456
transform 1 0 93932 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1021
timestamp 1636986456
transform 1 0 95036 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1033
timestamp 1636986456
transform 1 0 96140 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1045
timestamp 18001
transform 1 0 97244 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1636986456
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1636986456
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 18001
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1636986456
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1636986456
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1636986456
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1636986456
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 18001
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 18001
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1636986456
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1636986456
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1636986456
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1636986456
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 18001
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 18001
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1636986456
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1636986456
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1636986456
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1636986456
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 18001
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 18001
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1636986456
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1636986456
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1636986456
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1636986456
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 18001
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 18001
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1636986456
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1636986456
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1636986456
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1636986456
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 18001
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 18001
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1636986456
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1636986456
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1636986456
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1636986456
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 18001
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 18001
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1636986456
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1636986456
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1636986456
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1636986456
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 18001
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 18001
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1636986456
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1636986456
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1636986456
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1636986456
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 18001
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 18001
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1636986456
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1636986456
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_501
timestamp 1636986456
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_513
timestamp 1636986456
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_525
timestamp 18001
transform 1 0 49404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 18001
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_533
timestamp 1636986456
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_545
timestamp 1636986456
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_557
timestamp 1636986456
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_569
timestamp 1636986456
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_581
timestamp 18001
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 18001
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_589
timestamp 1636986456
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_601
timestamp 1636986456
transform 1 0 56396 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_613
timestamp 1636986456
transform 1 0 57500 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_625
timestamp 1636986456
transform 1 0 58604 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_637
timestamp 18001
transform 1 0 59708 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_643
timestamp 18001
transform 1 0 60260 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_645
timestamp 1636986456
transform 1 0 60444 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_657
timestamp 1636986456
transform 1 0 61548 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_669
timestamp 1636986456
transform 1 0 62652 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_681
timestamp 1636986456
transform 1 0 63756 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_693
timestamp 18001
transform 1 0 64860 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_699
timestamp 18001
transform 1 0 65412 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_701
timestamp 1636986456
transform 1 0 65596 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_713
timestamp 1636986456
transform 1 0 66700 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_725
timestamp 1636986456
transform 1 0 67804 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_737
timestamp 1636986456
transform 1 0 68908 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_749
timestamp 18001
transform 1 0 70012 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_755
timestamp 18001
transform 1 0 70564 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_757
timestamp 1636986456
transform 1 0 70748 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_769
timestamp 1636986456
transform 1 0 71852 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_781
timestamp 1636986456
transform 1 0 72956 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_793
timestamp 1636986456
transform 1 0 74060 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_805
timestamp 18001
transform 1 0 75164 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_811
timestamp 18001
transform 1 0 75716 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_813
timestamp 1636986456
transform 1 0 75900 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_825
timestamp 1636986456
transform 1 0 77004 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_837
timestamp 1636986456
transform 1 0 78108 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_849
timestamp 1636986456
transform 1 0 79212 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_861
timestamp 18001
transform 1 0 80316 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_867
timestamp 18001
transform 1 0 80868 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_869
timestamp 1636986456
transform 1 0 81052 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_881
timestamp 1636986456
transform 1 0 82156 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_893
timestamp 1636986456
transform 1 0 83260 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_905
timestamp 1636986456
transform 1 0 84364 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_917
timestamp 18001
transform 1 0 85468 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_923
timestamp 18001
transform 1 0 86020 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_925
timestamp 1636986456
transform 1 0 86204 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_937
timestamp 1636986456
transform 1 0 87308 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_949
timestamp 1636986456
transform 1 0 88412 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_961
timestamp 1636986456
transform 1 0 89516 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_973
timestamp 18001
transform 1 0 90620 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_979
timestamp 18001
transform 1 0 91172 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_981
timestamp 1636986456
transform 1 0 91356 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_993
timestamp 1636986456
transform 1 0 92460 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1005
timestamp 1636986456
transform 1 0 93564 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1017
timestamp 1636986456
transform 1 0 94668 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1029
timestamp 18001
transform 1 0 95772 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1035
timestamp 18001
transform 1 0 96324 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1037
timestamp 1636986456
transform 1 0 96508 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1636986456
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1636986456
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1636986456
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1636986456
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 18001
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 18001
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1636986456
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1636986456
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1636986456
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1636986456
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 18001
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 18001
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1636986456
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1636986456
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1636986456
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1636986456
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 18001
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 18001
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1636986456
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1636986456
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1636986456
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1636986456
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 18001
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 18001
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1636986456
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1636986456
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1636986456
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1636986456
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 18001
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 18001
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1636986456
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1636986456
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1636986456
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1636986456
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 18001
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 18001
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1636986456
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1636986456
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1636986456
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1636986456
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 18001
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 18001
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1636986456
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1636986456
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1636986456
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1636986456
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 18001
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 18001
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1636986456
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1636986456
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1636986456
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1636986456
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 18001
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 18001
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1636986456
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_517
timestamp 1636986456
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_529
timestamp 1636986456
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_541
timestamp 1636986456
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 18001
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 18001
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_561
timestamp 1636986456
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_573
timestamp 1636986456
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_585
timestamp 1636986456
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_597
timestamp 1636986456
transform 1 0 56028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_609
timestamp 18001
transform 1 0 57132 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_615
timestamp 18001
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_617
timestamp 1636986456
transform 1 0 57868 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_629
timestamp 1636986456
transform 1 0 58972 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_641
timestamp 1636986456
transform 1 0 60076 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_653
timestamp 1636986456
transform 1 0 61180 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_665
timestamp 18001
transform 1 0 62284 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_671
timestamp 18001
transform 1 0 62836 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_673
timestamp 1636986456
transform 1 0 63020 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_685
timestamp 1636986456
transform 1 0 64124 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_697
timestamp 1636986456
transform 1 0 65228 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_709
timestamp 1636986456
transform 1 0 66332 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_721
timestamp 18001
transform 1 0 67436 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_727
timestamp 18001
transform 1 0 67988 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_729
timestamp 1636986456
transform 1 0 68172 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_741
timestamp 1636986456
transform 1 0 69276 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_753
timestamp 1636986456
transform 1 0 70380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_765
timestamp 1636986456
transform 1 0 71484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_777
timestamp 18001
transform 1 0 72588 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_783
timestamp 18001
transform 1 0 73140 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_785
timestamp 1636986456
transform 1 0 73324 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_797
timestamp 1636986456
transform 1 0 74428 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_809
timestamp 1636986456
transform 1 0 75532 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_821
timestamp 1636986456
transform 1 0 76636 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_833
timestamp 18001
transform 1 0 77740 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_839
timestamp 18001
transform 1 0 78292 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_841
timestamp 1636986456
transform 1 0 78476 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_853
timestamp 1636986456
transform 1 0 79580 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_865
timestamp 1636986456
transform 1 0 80684 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_877
timestamp 1636986456
transform 1 0 81788 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_889
timestamp 18001
transform 1 0 82892 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_895
timestamp 18001
transform 1 0 83444 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_897
timestamp 1636986456
transform 1 0 83628 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_909
timestamp 1636986456
transform 1 0 84732 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_921
timestamp 1636986456
transform 1 0 85836 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_933
timestamp 1636986456
transform 1 0 86940 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_945
timestamp 18001
transform 1 0 88044 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_951
timestamp 18001
transform 1 0 88596 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_953
timestamp 1636986456
transform 1 0 88780 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_965
timestamp 1636986456
transform 1 0 89884 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_977
timestamp 1636986456
transform 1 0 90988 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_989
timestamp 1636986456
transform 1 0 92092 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1001
timestamp 18001
transform 1 0 93196 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1007
timestamp 18001
transform 1 0 93748 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1009
timestamp 1636986456
transform 1 0 93932 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1021
timestamp 1636986456
transform 1 0 95036 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1033
timestamp 1636986456
transform 1 0 96140 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1045
timestamp 18001
transform 1 0 97244 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1636986456
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1636986456
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 18001
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1636986456
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1636986456
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_53
timestamp 18001
transform 1 0 5980 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_57
timestamp 1636986456
transform 1 0 6348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_69
timestamp 1636986456
transform 1 0 7452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_81
timestamp 18001
transform 1 0 8556 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_87
timestamp 18001
transform 1 0 9108 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_95
timestamp 18001
transform 1 0 9844 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_98
timestamp 18001
transform 1 0 10120 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_106
timestamp 18001
transform 1 0 10856 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_110
timestamp 18001
transform 1 0 11224 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_113
timestamp 18001
transform 1 0 11500 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_119
timestamp 18001
transform 1 0 12052 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_122
timestamp 1636986456
transform 1 0 12328 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_134
timestamp 18001
transform 1 0 13432 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1636986456
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1636986456
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_165
timestamp 18001
transform 1 0 16284 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_169
timestamp 1636986456
transform 1 0 16652 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_181
timestamp 1636986456
transform 1 0 17756 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_193
timestamp 18001
transform 1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1636986456
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1636986456
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_221
timestamp 18001
transform 1 0 21436 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_225
timestamp 1636986456
transform 1 0 21804 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_237
timestamp 1636986456
transform 1 0 22908 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_249
timestamp 18001
transform 1 0 24012 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1636986456
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1636986456
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_277
timestamp 18001
transform 1 0 26588 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_281
timestamp 1636986456
transform 1 0 26956 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_293
timestamp 1636986456
transform 1 0 28060 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_305
timestamp 18001
transform 1 0 29164 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1636986456
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1636986456
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_333
timestamp 18001
transform 1 0 31740 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_337
timestamp 1636986456
transform 1 0 32108 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_349
timestamp 1636986456
transform 1 0 33212 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_361
timestamp 18001
transform 1 0 34316 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1636986456
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1636986456
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_389
timestamp 18001
transform 1 0 36892 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_393
timestamp 1636986456
transform 1 0 37260 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_405
timestamp 1636986456
transform 1 0 38364 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_417
timestamp 18001
transform 1 0 39468 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1636986456
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1636986456
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_445
timestamp 18001
transform 1 0 42044 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_449
timestamp 1636986456
transform 1 0 42412 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_461
timestamp 1636986456
transform 1 0 43516 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_473
timestamp 18001
transform 1 0 44620 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1636986456
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1636986456
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_501
timestamp 18001
transform 1 0 47196 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_505
timestamp 1636986456
transform 1 0 47564 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_517
timestamp 1636986456
transform 1 0 48668 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_529
timestamp 18001
transform 1 0 49772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_533
timestamp 18001
transform 1 0 50140 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_545
timestamp 18001
transform 1 0 51244 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_555
timestamp 18001
transform 1 0 52164 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_559
timestamp 18001
transform 1 0 52532 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_561
timestamp 18001
transform 1 0 52716 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_567
timestamp 18001
transform 1 0 53268 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_575
timestamp 18001
transform 1 0 54004 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_579
timestamp 18001
transform 1 0 54372 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 18001
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_589
timestamp 1636986456
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_601
timestamp 1636986456
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_613
timestamp 18001
transform 1 0 57500 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_617
timestamp 1636986456
transform 1 0 57868 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_629
timestamp 1636986456
transform 1 0 58972 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_641
timestamp 18001
transform 1 0 60076 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_645
timestamp 1636986456
transform 1 0 60444 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_657
timestamp 1636986456
transform 1 0 61548 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_669
timestamp 18001
transform 1 0 62652 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_673
timestamp 1636986456
transform 1 0 63020 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_685
timestamp 1636986456
transform 1 0 64124 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_697
timestamp 18001
transform 1 0 65228 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_701
timestamp 1636986456
transform 1 0 65596 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_713
timestamp 1636986456
transform 1 0 66700 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_725
timestamp 18001
transform 1 0 67804 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_729
timestamp 1636986456
transform 1 0 68172 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_741
timestamp 1636986456
transform 1 0 69276 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_753
timestamp 18001
transform 1 0 70380 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_757
timestamp 1636986456
transform 1 0 70748 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_769
timestamp 1636986456
transform 1 0 71852 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_781
timestamp 18001
transform 1 0 72956 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_785
timestamp 1636986456
transform 1 0 73324 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_797
timestamp 1636986456
transform 1 0 74428 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_809
timestamp 18001
transform 1 0 75532 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_813
timestamp 1636986456
transform 1 0 75900 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_825
timestamp 1636986456
transform 1 0 77004 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_837
timestamp 18001
transform 1 0 78108 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_841
timestamp 1636986456
transform 1 0 78476 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_853
timestamp 1636986456
transform 1 0 79580 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_865
timestamp 18001
transform 1 0 80684 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_869
timestamp 1636986456
transform 1 0 81052 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_881
timestamp 1636986456
transform 1 0 82156 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_893
timestamp 18001
transform 1 0 83260 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_897
timestamp 1636986456
transform 1 0 83628 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_909
timestamp 1636986456
transform 1 0 84732 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_921
timestamp 18001
transform 1 0 85836 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_925
timestamp 1636986456
transform 1 0 86204 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_937
timestamp 1636986456
transform 1 0 87308 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_949
timestamp 18001
transform 1 0 88412 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_953
timestamp 1636986456
transform 1 0 88780 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_965
timestamp 1636986456
transform 1 0 89884 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_977
timestamp 18001
transform 1 0 90988 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_981
timestamp 1636986456
transform 1 0 91356 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_993
timestamp 1636986456
transform 1 0 92460 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_1005
timestamp 18001
transform 1 0 93564 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1009
timestamp 1636986456
transform 1 0 93932 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1021
timestamp 1636986456
transform 1 0 95036 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_1033
timestamp 18001
transform 1 0 96140 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1037
timestamp 1636986456
transform 1 0 96508 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1636986456
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1636986456
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1636986456
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_39
timestamp 18001
transform 1 0 4692 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_47
timestamp 18001
transform 1 0 5428 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1013
timestamp 1636986456
transform 1 0 94300 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1025
timestamp 1636986456
transform 1 0 95404 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1037
timestamp 1636986456
transform 1 0 96508 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1636986456
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1636986456
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 18001
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1636986456
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_41
timestamp 18001
transform 1 0 4876 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_49
timestamp 18001
transform 1 0 5612 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1013
timestamp 1636986456
transform 1 0 94300 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1025
timestamp 1636986456
transform 1 0 95404 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1037
timestamp 18001
transform 1 0 96508 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_1039
timestamp 18001
transform 1 0 96692 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_1047
timestamp 18001
transform 1 0 97428 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1636986456
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1636986456
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1636986456
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_39
timestamp 18001
transform 1 0 4692 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_47
timestamp 18001
transform 1 0 5428 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1013
timestamp 1636986456
transform 1 0 94300 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1025
timestamp 1636986456
transform 1 0 95404 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1037
timestamp 1636986456
transform 1 0 96508 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1636986456
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1636986456
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 18001
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1636986456
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_41
timestamp 18001
transform 1 0 4876 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_49
timestamp 18001
transform 1 0 5612 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1013
timestamp 1636986456
transform 1 0 94300 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1025
timestamp 1636986456
transform 1 0 95404 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1037
timestamp 18001
transform 1 0 96508 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_1039
timestamp 18001
transform 1 0 96692 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_1047
timestamp 18001
transform 1 0 97428 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1636986456
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1636986456
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1636986456
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_39
timestamp 18001
transform 1 0 4692 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_47
timestamp 18001
transform 1 0 5428 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1013
timestamp 1636986456
transform 1 0 94300 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1025
timestamp 1636986456
transform 1 0 95404 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1037
timestamp 18001
transform 1 0 96508 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1636986456
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1636986456
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 18001
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1636986456
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_41
timestamp 18001
transform 1 0 4876 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_49
timestamp 18001
transform 1 0 5612 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1013
timestamp 1636986456
transform 1 0 94300 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1025
timestamp 1636986456
transform 1 0 95404 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1037
timestamp 18001
transform 1 0 96508 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1039
timestamp 18001
transform 1 0 96692 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_1047
timestamp 18001
transform 1 0 97428 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1636986456
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1636986456
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1636986456
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_39
timestamp 18001
transform 1 0 4692 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_47
timestamp 18001
transform 1 0 5428 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1013
timestamp 1636986456
transform 1 0 94300 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1025
timestamp 1636986456
transform 1 0 95404 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1037
timestamp 1636986456
transform 1 0 96508 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1636986456
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1636986456
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 18001
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1636986456
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_41
timestamp 18001
transform 1 0 4876 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_49
timestamp 18001
transform 1 0 5612 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1013
timestamp 1636986456
transform 1 0 94300 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1025
timestamp 1636986456
transform 1 0 95404 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1037
timestamp 18001
transform 1 0 96508 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1039
timestamp 18001
transform 1 0 96692 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_1047
timestamp 18001
transform 1 0 97428 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1636986456
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1636986456
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1636986456
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_39
timestamp 18001
transform 1 0 4692 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_47
timestamp 18001
transform 1 0 5428 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1013
timestamp 1636986456
transform 1 0 94300 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1025
timestamp 1636986456
transform 1 0 95404 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1037
timestamp 1636986456
transform 1 0 96508 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1636986456
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1636986456
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 18001
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1636986456
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_41
timestamp 18001
transform 1 0 4876 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_49
timestamp 18001
transform 1 0 5612 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1013
timestamp 1636986456
transform 1 0 94300 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1025
timestamp 1636986456
transform 1 0 95404 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1037
timestamp 18001
transform 1 0 96508 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_1039
timestamp 18001
transform 1 0 96692 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_1047
timestamp 18001
transform 1 0 97428 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_9
timestamp 1636986456
transform 1 0 1932 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_21
timestamp 1636986456
transform 1 0 3036 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_33
timestamp 1636986456
transform 1 0 4140 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_45
timestamp 18001
transform 1 0 5244 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_49
timestamp 18001
transform 1 0 5612 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1013
timestamp 1636986456
transform 1 0 94300 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1025
timestamp 1636986456
transform 1 0 95404 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_1037
timestamp 18001
transform 1 0 96508 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1636986456
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1636986456
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 18001
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1636986456
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_41
timestamp 18001
transform 1 0 4876 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_49
timestamp 18001
transform 1 0 5612 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1013
timestamp 1636986456
transform 1 0 94300 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1025
timestamp 1636986456
transform 1 0 95404 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1037
timestamp 18001
transform 1 0 96508 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_1039
timestamp 18001
transform 1 0 96692 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_1047
timestamp 18001
transform 1 0 97428 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1636986456
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1636986456
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1636986456
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_39
timestamp 18001
transform 1 0 4692 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_47
timestamp 18001
transform 1 0 5428 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1013
timestamp 1636986456
transform 1 0 94300 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1025
timestamp 1636986456
transform 1 0 95404 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1037
timestamp 1636986456
transform 1 0 96508 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_9
timestamp 1636986456
transform 1 0 1932 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_21
timestamp 18001
transform 1 0 3036 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 18001
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1636986456
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_41
timestamp 18001
transform 1 0 4876 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_49
timestamp 18001
transform 1 0 5612 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1013
timestamp 1636986456
transform 1 0 94300 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1025
timestamp 1636986456
transform 1 0 95404 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1037
timestamp 18001
transform 1 0 96508 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1039
timestamp 18001
transform 1 0 96692 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_11
timestamp 1636986456
transform 1 0 2116 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_23
timestamp 1636986456
transform 1 0 3220 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_35
timestamp 1636986456
transform 1 0 4324 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_47
timestamp 18001
transform 1 0 5428 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1013
timestamp 1636986456
transform 1 0 94300 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1025
timestamp 1636986456
transform 1 0 95404 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_1037
timestamp 18001
transform 1 0 96508 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1636986456
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1636986456
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 18001
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1636986456
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_41
timestamp 18001
transform 1 0 4876 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_49
timestamp 18001
transform 1 0 5612 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1013
timestamp 1636986456
transform 1 0 94300 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1025
timestamp 1636986456
transform 1 0 95404 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_1037
timestamp 18001
transform 1 0 96508 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_1039
timestamp 18001
transform 1 0 96692 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_1047
timestamp 18001
transform 1 0 97428 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1636986456
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1636986456
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1636986456
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_39
timestamp 18001
transform 1 0 4692 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_47
timestamp 18001
transform 1 0 5428 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1013
timestamp 1636986456
transform 1 0 94300 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1025
timestamp 1636986456
transform 1 0 95404 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1037
timestamp 1636986456
transform 1 0 96508 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_11
timestamp 1636986456
transform 1 0 2116 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_23
timestamp 18001
transform 1 0 3220 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 18001
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1636986456
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_41
timestamp 18001
transform 1 0 4876 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_49
timestamp 18001
transform 1 0 5612 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1013
timestamp 1636986456
transform 1 0 94300 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1025
timestamp 1636986456
transform 1 0 95404 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_1037
timestamp 18001
transform 1 0 96508 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_1039
timestamp 18001
transform 1 0 96692 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_9
timestamp 1636986456
transform 1 0 1932 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_21
timestamp 1636986456
transform 1 0 3036 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_33
timestamp 1636986456
transform 1 0 4140 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_45
timestamp 18001
transform 1 0 5244 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_49
timestamp 18001
transform 1 0 5612 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1013
timestamp 1636986456
transform 1 0 94300 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1025
timestamp 1636986456
transform 1 0 95404 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_1037
timestamp 18001
transform 1 0 96508 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1636986456
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1636986456
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 18001
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1636986456
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_41
timestamp 18001
transform 1 0 4876 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_49
timestamp 18001
transform 1 0 5612 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1013
timestamp 1636986456
transform 1 0 94300 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1025
timestamp 1636986456
transform 1 0 95404 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_1037
timestamp 18001
transform 1 0 96508 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_1039
timestamp 18001
transform 1 0 96692 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_1047
timestamp 18001
transform 1 0 97428 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_9
timestamp 1636986456
transform 1 0 1932 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_21
timestamp 1636986456
transform 1 0 3036 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_33
timestamp 1636986456
transform 1 0 4140 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_45
timestamp 18001
transform 1 0 5244 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_49
timestamp 18001
transform 1 0 5612 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1013
timestamp 1636986456
transform 1 0 94300 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1025
timestamp 1636986456
transform 1 0 95404 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_1037
timestamp 18001
transform 1 0 96508 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1636986456
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1636986456
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 18001
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1636986456
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_41
timestamp 18001
transform 1 0 4876 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_49
timestamp 18001
transform 1 0 5612 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1013
timestamp 1636986456
transform 1 0 94300 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1025
timestamp 1636986456
transform 1 0 95404 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_1037
timestamp 18001
transform 1 0 96508 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_1039
timestamp 18001
transform 1 0 96692 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_1047
timestamp 18001
transform 1 0 97428 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1636986456
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1636986456
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1636986456
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_39
timestamp 18001
transform 1 0 4692 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_47
timestamp 18001
transform 1 0 5428 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1013
timestamp 1636986456
transform 1 0 94300 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1025
timestamp 1636986456
transform 1 0 95404 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1037
timestamp 1636986456
transform 1 0 96508 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_11
timestamp 1636986456
transform 1 0 2116 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_23
timestamp 18001
transform 1 0 3220 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 18001
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1636986456
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_41
timestamp 18001
transform 1 0 4876 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_49
timestamp 18001
transform 1 0 5612 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1013
timestamp 1636986456
transform 1 0 94300 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1025
timestamp 1636986456
transform 1 0 95404 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_1037
timestamp 18001
transform 1 0 96508 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_1039
timestamp 18001
transform 1 0 96692 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_9
timestamp 1636986456
transform 1 0 1932 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_21
timestamp 1636986456
transform 1 0 3036 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_33
timestamp 1636986456
transform 1 0 4140 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_45
timestamp 18001
transform 1 0 5244 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_49
timestamp 18001
transform 1 0 5612 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1013
timestamp 1636986456
transform 1 0 94300 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1025
timestamp 1636986456
transform 1 0 95404 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_1037
timestamp 18001
transform 1 0 96508 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1636986456
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1636986456
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 18001
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1636986456
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_41
timestamp 18001
transform 1 0 4876 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_49
timestamp 18001
transform 1 0 5612 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1013
timestamp 1636986456
transform 1 0 94300 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1025
timestamp 1636986456
transform 1 0 95404 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_1037
timestamp 18001
transform 1 0 96508 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_1039
timestamp 18001
transform 1 0 96692 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_1047
timestamp 18001
transform 1 0 97428 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1636986456
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1636986456
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1636986456
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_39
timestamp 18001
transform 1 0 4692 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_47
timestamp 18001
transform 1 0 5428 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1013
timestamp 1636986456
transform 1 0 94300 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1025
timestamp 1636986456
transform 1 0 95404 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1037
timestamp 1636986456
transform 1 0 96508 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_11
timestamp 1636986456
transform 1 0 2116 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_23
timestamp 18001
transform 1 0 3220 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 18001
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1636986456
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_41
timestamp 18001
transform 1 0 4876 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_49
timestamp 18001
transform 1 0 5612 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1013
timestamp 1636986456
transform 1 0 94300 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1025
timestamp 1636986456
transform 1 0 95404 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_1037
timestamp 18001
transform 1 0 96508 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_1039
timestamp 18001
transform 1 0 96692 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_9
timestamp 1636986456
transform 1 0 1932 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_21
timestamp 1636986456
transform 1 0 3036 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_33
timestamp 1636986456
transform 1 0 4140 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_45
timestamp 18001
transform 1 0 5244 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_49
timestamp 18001
transform 1 0 5612 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1013
timestamp 1636986456
transform 1 0 94300 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1025
timestamp 1636986456
transform 1 0 95404 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_1037
timestamp 18001
transform 1 0 96508 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1636986456
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1636986456
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 18001
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1636986456
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_41
timestamp 18001
transform 1 0 4876 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_49
timestamp 18001
transform 1 0 5612 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1013
timestamp 1636986456
transform 1 0 94300 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1025
timestamp 1636986456
transform 1 0 95404 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_1037
timestamp 18001
transform 1 0 96508 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_1039
timestamp 18001
transform 1 0 96692 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_1047
timestamp 18001
transform 1 0 97428 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_9
timestamp 1636986456
transform 1 0 1932 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_21
timestamp 1636986456
transform 1 0 3036 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_33
timestamp 1636986456
transform 1 0 4140 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_45
timestamp 18001
transform 1 0 5244 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_49
timestamp 18001
transform 1 0 5612 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1013
timestamp 1636986456
transform 1 0 94300 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1025
timestamp 1636986456
transform 1 0 95404 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_1037
timestamp 18001
transform 1 0 96508 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1636986456
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1636986456
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 18001
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1636986456
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_41
timestamp 18001
transform 1 0 4876 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_49
timestamp 18001
transform 1 0 5612 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1013
timestamp 1636986456
transform 1 0 94300 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1025
timestamp 1636986456
transform 1 0 95404 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_1037
timestamp 18001
transform 1 0 96508 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_1039
timestamp 18001
transform 1 0 96692 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_1047
timestamp 18001
transform 1 0 97428 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1636986456
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1636986456
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1636986456
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_39
timestamp 18001
transform 1 0 4692 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_47
timestamp 18001
transform 1 0 5428 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1013
timestamp 1636986456
transform 1 0 94300 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1025
timestamp 1636986456
transform 1 0 95404 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1037
timestamp 1636986456
transform 1 0 96508 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_9
timestamp 1636986456
transform 1 0 1932 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_21
timestamp 18001
transform 1 0 3036 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 18001
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1636986456
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_41
timestamp 18001
transform 1 0 4876 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_49
timestamp 18001
transform 1 0 5612 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1013
timestamp 1636986456
transform 1 0 94300 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1025
timestamp 1636986456
transform 1 0 95404 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_1037
timestamp 18001
transform 1 0 96508 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_1039
timestamp 18001
transform 1 0 96692 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_9
timestamp 1636986456
transform 1 0 1932 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_21
timestamp 1636986456
transform 1 0 3036 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_33
timestamp 1636986456
transform 1 0 4140 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_45
timestamp 18001
transform 1 0 5244 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_49
timestamp 18001
transform 1 0 5612 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1013
timestamp 1636986456
transform 1 0 94300 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1025
timestamp 1636986456
transform 1 0 95404 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_1037
timestamp 18001
transform 1 0 96508 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1636986456
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1636986456
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 18001
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1636986456
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_41
timestamp 18001
transform 1 0 4876 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_49
timestamp 18001
transform 1 0 5612 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1013
timestamp 1636986456
transform 1 0 94300 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1025
timestamp 1636986456
transform 1 0 95404 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_1037
timestamp 18001
transform 1 0 96508 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_1039
timestamp 18001
transform 1 0 96692 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_1047
timestamp 18001
transform 1 0 97428 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1636986456
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1636986456
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1636986456
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_39
timestamp 18001
transform 1 0 4692 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_47
timestamp 18001
transform 1 0 5428 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1013
timestamp 1636986456
transform 1 0 94300 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1025
timestamp 1636986456
transform 1 0 95404 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1037
timestamp 1636986456
transform 1 0 96508 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_9
timestamp 1636986456
transform 1 0 1932 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_21
timestamp 18001
transform 1 0 3036 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 18001
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1636986456
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_41
timestamp 18001
transform 1 0 4876 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_49
timestamp 18001
transform 1 0 5612 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1013
timestamp 1636986456
transform 1 0 94300 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1025
timestamp 1636986456
transform 1 0 95404 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_1037
timestamp 18001
transform 1 0 96508 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_1039
timestamp 18001
transform 1 0 96692 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_9
timestamp 1636986456
transform 1 0 1932 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_21
timestamp 1636986456
transform 1 0 3036 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_33
timestamp 1636986456
transform 1 0 4140 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_45
timestamp 18001
transform 1 0 5244 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_49
timestamp 18001
transform 1 0 5612 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1013
timestamp 1636986456
transform 1 0 94300 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1025
timestamp 1636986456
transform 1 0 95404 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_1037
timestamp 18001
transform 1 0 96508 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1636986456
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1636986456
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 18001
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1636986456
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_41
timestamp 18001
transform 1 0 4876 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_49
timestamp 18001
transform 1 0 5612 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1013
timestamp 1636986456
transform 1 0 94300 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1025
timestamp 1636986456
transform 1 0 95404 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_1037
timestamp 18001
transform 1 0 96508 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_1039
timestamp 18001
transform 1 0 96692 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_1047
timestamp 18001
transform 1 0 97428 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_8
timestamp 1636986456
transform 1 0 1840 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_20
timestamp 1636986456
transform 1 0 2944 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_32
timestamp 1636986456
transform 1 0 4048 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_44
timestamp 18001
transform 1 0 5152 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1013
timestamp 1636986456
transform 1 0 94300 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1025
timestamp 1636986456
transform 1 0 95404 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_1037
timestamp 18001
transform 1 0 96508 0 -1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1636986456
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1636986456
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 18001
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1636986456
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_41
timestamp 18001
transform 1 0 4876 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_49
timestamp 18001
transform 1 0 5612 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1013
timestamp 1636986456
transform 1 0 94300 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1025
timestamp 1636986456
transform 1 0 95404 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_1037
timestamp 18001
transform 1 0 96508 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_1039
timestamp 18001
transform 1 0 96692 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_1047
timestamp 18001
transform 1 0 97428 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1636986456
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1636986456
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1636986456
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_39
timestamp 18001
transform 1 0 4692 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_47
timestamp 18001
transform 1 0 5428 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1013
timestamp 1636986456
transform 1 0 94300 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1025
timestamp 1636986456
transform 1 0 95404 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1037
timestamp 1636986456
transform 1 0 96508 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_7
timestamp 1636986456
transform 1 0 1748 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_19
timestamp 18001
transform 1 0 2852 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 18001
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1636986456
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_41
timestamp 18001
transform 1 0 4876 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_49
timestamp 18001
transform 1 0 5612 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1013
timestamp 1636986456
transform 1 0 94300 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1025
timestamp 1636986456
transform 1 0 95404 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_1037
timestamp 18001
transform 1 0 96508 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_1039
timestamp 18001
transform 1 0 96692 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_1043
timestamp 18001
transform 1 0 97060 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_7
timestamp 1636986456
transform 1 0 1748 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_19
timestamp 1636986456
transform 1 0 2852 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_31
timestamp 1636986456
transform 1 0 3956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_43
timestamp 18001
transform 1 0 5060 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_49
timestamp 18001
transform 1 0 5612 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1013
timestamp 1636986456
transform 1 0 94300 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1025
timestamp 1636986456
transform 1 0 95404 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_1037
timestamp 18001
transform 1 0 96508 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1636986456
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1636986456
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 18001
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1636986456
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_41
timestamp 18001
transform 1 0 4876 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_49
timestamp 18001
transform 1 0 5612 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1013
timestamp 1636986456
transform 1 0 94300 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1025
timestamp 1636986456
transform 1 0 95404 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_1037
timestamp 18001
transform 1 0 96508 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_1039
timestamp 18001
transform 1 0 96692 0 1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1636986456
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1636986456
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1636986456
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_39
timestamp 18001
transform 1 0 4692 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_47
timestamp 18001
transform 1 0 5428 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1013
timestamp 1636986456
transform 1 0 94300 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1025
timestamp 1636986456
transform 1 0 95404 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1037
timestamp 1636986456
transform 1 0 96508 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_7
timestamp 1636986456
transform 1 0 1748 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_19
timestamp 18001
transform 1 0 2852 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 18001
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1636986456
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_41
timestamp 18001
transform 1 0 4876 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_49
timestamp 18001
transform 1 0 5612 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1013
timestamp 1636986456
transform 1 0 94300 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1025
timestamp 1636986456
transform 1 0 95404 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_1037
timestamp 18001
transform 1 0 96508 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_1039
timestamp 18001
transform 1 0 96692 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_1043
timestamp 18001
transform 1 0 97060 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_7
timestamp 1636986456
transform 1 0 1748 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_19
timestamp 1636986456
transform 1 0 2852 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_31
timestamp 1636986456
transform 1 0 3956 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_43
timestamp 18001
transform 1 0 5060 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_49
timestamp 18001
transform 1 0 5612 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1013
timestamp 1636986456
transform 1 0 94300 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1025
timestamp 1636986456
transform 1 0 95404 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_1037
timestamp 18001
transform 1 0 96508 0 -1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1636986456
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1636986456
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 18001
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1636986456
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_41
timestamp 18001
transform 1 0 4876 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_49
timestamp 18001
transform 1 0 5612 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1013
timestamp 1636986456
transform 1 0 94300 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1025
timestamp 1636986456
transform 1 0 95404 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_1037
timestamp 18001
transform 1 0 96508 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_1039
timestamp 18001
transform 1 0 96692 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_1047
timestamp 18001
transform 1 0 97428 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_7
timestamp 1636986456
transform 1 0 1748 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_19
timestamp 1636986456
transform 1 0 2852 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_31
timestamp 1636986456
transform 1 0 3956 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_43
timestamp 18001
transform 1 0 5060 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_49
timestamp 18001
transform 1 0 5612 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1013
timestamp 1636986456
transform 1 0 94300 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1025
timestamp 1636986456
transform 1 0 95404 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_1037
timestamp 18001
transform 1 0 96508 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_1043
timestamp 18001
transform 1 0 97060 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1636986456
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1636986456
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 18001
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1636986456
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_41
timestamp 18001
transform 1 0 4876 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_49
timestamp 18001
transform 1 0 5612 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1013
timestamp 1636986456
transform 1 0 94300 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1025
timestamp 1636986456
transform 1 0 95404 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_1037
timestamp 18001
transform 1 0 96508 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_1039
timestamp 18001
transform 1 0 96692 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_1047
timestamp 18001
transform 1 0 97428 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1636986456
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1636986456
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1636986456
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_39
timestamp 18001
transform 1 0 4692 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_47
timestamp 18001
transform 1 0 5428 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1013
timestamp 1636986456
transform 1 0 94300 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1025
timestamp 1636986456
transform 1 0 95404 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1037
timestamp 1636986456
transform 1 0 96508 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_7
timestamp 1636986456
transform 1 0 1748 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_19
timestamp 18001
transform 1 0 2852 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 18001
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1636986456
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_41
timestamp 18001
transform 1 0 4876 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_49
timestamp 18001
transform 1 0 5612 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1013
timestamp 1636986456
transform 1 0 94300 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1025
timestamp 1636986456
transform 1 0 95404 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_1037
timestamp 18001
transform 1 0 96508 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_1039
timestamp 18001
transform 1 0 96692 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_1043
timestamp 18001
transform 1 0 97060 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_7
timestamp 1636986456
transform 1 0 1748 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_19
timestamp 1636986456
transform 1 0 2852 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_31
timestamp 1636986456
transform 1 0 3956 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_43
timestamp 18001
transform 1 0 5060 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_49
timestamp 18001
transform 1 0 5612 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1013
timestamp 1636986456
transform 1 0 94300 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1025
timestamp 1636986456
transform 1 0 95404 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_1037
timestamp 18001
transform 1 0 96508 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_1043
timestamp 18001
transform 1 0 97060 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1636986456
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1636986456
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 18001
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1636986456
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_41
timestamp 18001
transform 1 0 4876 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_49
timestamp 18001
transform 1 0 5612 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_1013
timestamp 1636986456
transform 1 0 94300 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_1025
timestamp 1636986456
transform 1 0 95404 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_1037
timestamp 18001
transform 1 0 96508 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_1039
timestamp 18001
transform 1 0 96692 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_1047
timestamp 18001
transform 1 0 97428 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1636986456
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1636986456
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1636986456
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_39
timestamp 18001
transform 1 0 4692 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_47
timestamp 18001
transform 1 0 5428 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_1013
timestamp 1636986456
transform 1 0 94300 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_1025
timestamp 1636986456
transform 1 0 95404 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_1037
timestamp 1636986456
transform 1 0 96508 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_7
timestamp 1636986456
transform 1 0 1748 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_19
timestamp 18001
transform 1 0 2852 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 18001
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1636986456
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_41
timestamp 18001
transform 1 0 4876 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_49
timestamp 18001
transform 1 0 5612 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_1013
timestamp 1636986456
transform 1 0 94300 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_1025
timestamp 1636986456
transform 1 0 95404 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_1037
timestamp 18001
transform 1 0 96508 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1039
timestamp 18001
transform 1 0 96692 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_7
timestamp 1636986456
transform 1 0 1748 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_19
timestamp 1636986456
transform 1 0 2852 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_31
timestamp 1636986456
transform 1 0 3956 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_43
timestamp 18001
transform 1 0 5060 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_49
timestamp 18001
transform 1 0 5612 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_1013
timestamp 1636986456
transform 1 0 94300 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_1025
timestamp 1636986456
transform 1 0 95404 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_1037
timestamp 18001
transform 1 0 96508 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_1043
timestamp 18001
transform 1 0 97060 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1636986456
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 1636986456
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 18001
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1636986456
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_41
timestamp 18001
transform 1 0 4876 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_49
timestamp 18001
transform 1 0 5612 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_1013
timestamp 1636986456
transform 1 0 94300 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_1025
timestamp 1636986456
transform 1 0 95404 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_1037
timestamp 18001
transform 1 0 96508 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_1039
timestamp 18001
transform 1 0 96692 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_1047
timestamp 18001
transform 1 0 97428 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_7
timestamp 1636986456
transform 1 0 1748 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_19
timestamp 1636986456
transform 1 0 2852 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_31
timestamp 1636986456
transform 1 0 3956 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_43
timestamp 18001
transform 1 0 5060 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_49
timestamp 18001
transform 1 0 5612 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_1013
timestamp 1636986456
transform 1 0 94300 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_1025
timestamp 1636986456
transform 1 0 95404 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_1037
timestamp 18001
transform 1 0 96508 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_1043
timestamp 18001
transform 1 0 97060 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1636986456
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1636986456
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 18001
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1636986456
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_41
timestamp 18001
transform 1 0 4876 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_49
timestamp 18001
transform 1 0 5612 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_1013
timestamp 1636986456
transform 1 0 94300 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_1025
timestamp 1636986456
transform 1 0 95404 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_1037
timestamp 18001
transform 1 0 96508 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_1039
timestamp 18001
transform 1 0 96692 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_1047
timestamp 18001
transform 1 0 97428 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1636986456
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1636986456
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1636986456
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_39
timestamp 18001
transform 1 0 4692 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_69_47
timestamp 18001
transform 1 0 5428 0 -1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_69_1013
timestamp 1636986456
transform 1 0 94300 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_1025
timestamp 1636986456
transform 1 0 95404 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_1037
timestamp 1636986456
transform 1 0 96508 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_7
timestamp 1636986456
transform 1 0 1748 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_19
timestamp 18001
transform 1 0 2852 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 18001
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1636986456
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_41
timestamp 18001
transform 1 0 4876 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_49
timestamp 18001
transform 1 0 5612 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_1013
timestamp 1636986456
transform 1 0 94300 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_1025
timestamp 1636986456
transform 1 0 95404 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_1037
timestamp 18001
transform 1 0 96508 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_1039
timestamp 18001
transform 1 0 96692 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_1043
timestamp 18001
transform 1 0 97060 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_7
timestamp 1636986456
transform 1 0 1748 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_19
timestamp 1636986456
transform 1 0 2852 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_31
timestamp 1636986456
transform 1 0 3956 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_43
timestamp 18001
transform 1 0 5060 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_49
timestamp 18001
transform 1 0 5612 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_1013
timestamp 1636986456
transform 1 0 94300 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_1025
timestamp 1636986456
transform 1 0 95404 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_1037
timestamp 18001
transform 1 0 96508 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_1043
timestamp 18001
transform 1 0 97060 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1636986456
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1636986456
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 18001
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1636986456
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_41
timestamp 18001
transform 1 0 4876 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_49
timestamp 18001
transform 1 0 5612 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_1013
timestamp 1636986456
transform 1 0 94300 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_1025
timestamp 1636986456
transform 1 0 95404 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_1037
timestamp 18001
transform 1 0 96508 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_1039
timestamp 18001
transform 1 0 96692 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_1047
timestamp 18001
transform 1 0 97428 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1636986456
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1636986456
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1636986456
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_39
timestamp 18001
transform 1 0 4692 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_73_47
timestamp 18001
transform 1 0 5428 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_73_1013
timestamp 1636986456
transform 1 0 94300 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_1025
timestamp 1636986456
transform 1 0 95404 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_1037
timestamp 1636986456
transform 1 0 96508 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_7
timestamp 1636986456
transform 1 0 1748 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_19
timestamp 18001
transform 1 0 2852 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 18001
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1636986456
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_41
timestamp 18001
transform 1 0 4876 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_49
timestamp 18001
transform 1 0 5612 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_1013
timestamp 1636986456
transform 1 0 94300 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_1025
timestamp 1636986456
transform 1 0 95404 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_1037
timestamp 18001
transform 1 0 96508 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_1039
timestamp 18001
transform 1 0 96692 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_1043
timestamp 18001
transform 1 0 97060 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_7
timestamp 1636986456
transform 1 0 1748 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_19
timestamp 1636986456
transform 1 0 2852 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_31
timestamp 1636986456
transform 1 0 3956 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_43
timestamp 18001
transform 1 0 5060 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_49
timestamp 18001
transform 1 0 5612 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_1013
timestamp 1636986456
transform 1 0 94300 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_1025
timestamp 1636986456
transform 1 0 95404 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_1037
timestamp 18001
transform 1 0 96508 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_1043
timestamp 18001
transform 1 0 97060 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1636986456
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1636986456
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 18001
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1636986456
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_41
timestamp 18001
transform 1 0 4876 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_76_49
timestamp 18001
transform 1 0 5612 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_1013
timestamp 1636986456
transform 1 0 94300 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_1025
timestamp 1636986456
transform 1 0 95404 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_1037
timestamp 18001
transform 1 0 96508 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_1039
timestamp 18001
transform 1 0 96692 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_1047
timestamp 18001
transform 1 0 97428 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_77_7
timestamp 1636986456
transform 1 0 1748 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_19
timestamp 1636986456
transform 1 0 2852 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_31
timestamp 1636986456
transform 1 0 3956 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_43
timestamp 18001
transform 1 0 5060 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_49
timestamp 18001
transform 1 0 5612 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_1013
timestamp 1636986456
transform 1 0 94300 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_1025
timestamp 1636986456
transform 1 0 95404 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_1037
timestamp 18001
transform 1 0 96508 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_1043
timestamp 18001
transform 1 0 97060 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1636986456
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1636986456
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 18001
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1636986456
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_41
timestamp 18001
transform 1 0 4876 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_78_49
timestamp 18001
transform 1 0 5612 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_1013
timestamp 1636986456
transform 1 0 94300 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_1025
timestamp 1636986456
transform 1 0 95404 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_1037
timestamp 18001
transform 1 0 96508 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_1039
timestamp 18001
transform 1 0 96692 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_1047
timestamp 18001
transform 1 0 97428 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1636986456
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1636986456
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 1636986456
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_39
timestamp 18001
transform 1 0 4692 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_79_47
timestamp 18001
transform 1 0 5428 0 -1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_79_1013
timestamp 1636986456
transform 1 0 94300 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_1025
timestamp 1636986456
transform 1 0 95404 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_1037
timestamp 1636986456
transform 1 0 96508 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_7
timestamp 1636986456
transform 1 0 1748 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_19
timestamp 18001
transform 1 0 2852 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 18001
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1636986456
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_41
timestamp 18001
transform 1 0 4876 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_49
timestamp 18001
transform 1 0 5612 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_1013
timestamp 1636986456
transform 1 0 94300 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_1025
timestamp 1636986456
transform 1 0 95404 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_1037
timestamp 18001
transform 1 0 96508 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_1039
timestamp 18001
transform 1 0 96692 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_1043
timestamp 18001
transform 1 0 97060 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1636986456
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1636986456
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_27
timestamp 1636986456
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_39
timestamp 18001
transform 1 0 4692 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_47
timestamp 18001
transform 1 0 5428 0 -1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_81_1013
timestamp 1636986456
transform 1 0 94300 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_1025
timestamp 1636986456
transform 1 0 95404 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_1037
timestamp 1636986456
transform 1 0 96508 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_3
timestamp 1636986456
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_15
timestamp 1636986456
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 18001
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1636986456
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_41
timestamp 18001
transform 1 0 4876 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_49
timestamp 18001
transform 1 0 5612 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_1013
timestamp 1636986456
transform 1 0 94300 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_1025
timestamp 1636986456
transform 1 0 95404 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_1037
timestamp 18001
transform 1 0 96508 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_1039
timestamp 18001
transform 1 0 96692 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_1047
timestamp 18001
transform 1 0 97428 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_83_3
timestamp 1636986456
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_15
timestamp 1636986456
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_27
timestamp 1636986456
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_39
timestamp 18001
transform 1 0 4692 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_83_47
timestamp 18001
transform 1 0 5428 0 -1 47872
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_83_1013
timestamp 1636986456
transform 1 0 94300 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_1025
timestamp 1636986456
transform 1 0 95404 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_1037
timestamp 1636986456
transform 1 0 96508 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_3
timestamp 1636986456
transform 1 0 1380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_15
timestamp 1636986456
transform 1 0 2484 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 18001
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1636986456
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_41
timestamp 18001
transform 1 0 4876 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_47
timestamp 18001
transform 1 0 5428 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_1013
timestamp 1636986456
transform 1 0 94300 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_1025
timestamp 1636986456
transform 1 0 95404 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_1037
timestamp 18001
transform 1 0 96508 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_1039
timestamp 18001
transform 1 0 96692 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_84_1047
timestamp 18001
transform 1 0 97428 0 1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_85_9
timestamp 1636986456
transform 1 0 1932 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_21
timestamp 1636986456
transform 1 0 3036 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_33
timestamp 18001
transform 1 0 4140 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_85_41
timestamp 18001
transform 1 0 4876 0 -1 48960
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_85_1021
timestamp 1636986456
transform 1 0 95036 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_1033
timestamp 1636986456
transform 1 0 96140 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_1045
timestamp 18001
transform 1 0 97244 0 -1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_86_3
timestamp 1636986456
transform 1 0 1380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_15
timestamp 1636986456
transform 1 0 2484 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 18001
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_29
timestamp 1636986456
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_41
timestamp 18001
transform 1 0 4876 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_86_49
timestamp 18001
transform 1 0 5612 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_1013
timestamp 1636986456
transform 1 0 94300 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_1025
timestamp 1636986456
transform 1 0 95404 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_1037
timestamp 18001
transform 1 0 96508 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_86_1039
timestamp 18001
transform 1 0 96692 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_86_1047
timestamp 18001
transform 1 0 97428 0 1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_87_3
timestamp 1636986456
transform 1 0 1380 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_15
timestamp 1636986456
transform 1 0 2484 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_27
timestamp 1636986456
transform 1 0 3588 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_39
timestamp 18001
transform 1 0 4692 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_87_47
timestamp 18001
transform 1 0 5428 0 -1 50048
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_87_1013
timestamp 1636986456
transform 1 0 94300 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_1025
timestamp 1636986456
transform 1 0 95404 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_1037
timestamp 1636986456
transform 1 0 96508 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_3
timestamp 1636986456
transform 1 0 1380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_15
timestamp 1636986456
transform 1 0 2484 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_27
timestamp 18001
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_29
timestamp 1636986456
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_41
timestamp 18001
transform 1 0 4876 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_47
timestamp 18001
transform 1 0 5428 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_1013
timestamp 1636986456
transform 1 0 94300 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_1025
timestamp 1636986456
transform 1 0 95404 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_1037
timestamp 18001
transform 1 0 96508 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_88_1039
timestamp 18001
transform 1 0 96692 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_88_1047
timestamp 18001
transform 1 0 97428 0 1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_89_3
timestamp 1636986456
transform 1 0 1380 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_15
timestamp 1636986456
transform 1 0 2484 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_27
timestamp 1636986456
transform 1 0 3588 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_39
timestamp 18001
transform 1 0 4692 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_43
timestamp 18001
transform 1 0 5060 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_1019
timestamp 1636986456
transform 1 0 94852 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_1031
timestamp 1636986456
transform 1 0 95956 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_1043
timestamp 18001
transform 1 0 97060 0 -1 51136
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_90_3
timestamp 1636986456
transform 1 0 1380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_15
timestamp 1636986456
transform 1 0 2484 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 18001
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_29
timestamp 1636986456
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_90_41
timestamp 18001
transform 1 0 4876 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_90_49
timestamp 18001
transform 1 0 5612 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_1013
timestamp 1636986456
transform 1 0 94300 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_1025
timestamp 1636986456
transform 1 0 95404 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_1037
timestamp 18001
transform 1 0 96508 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_90_1039
timestamp 18001
transform 1 0 96692 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_90_1047
timestamp 18001
transform 1 0 97428 0 1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_91_3
timestamp 1636986456
transform 1 0 1380 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_15
timestamp 1636986456
transform 1 0 2484 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_27
timestamp 1636986456
transform 1 0 3588 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_39
timestamp 18001
transform 1 0 4692 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_91_47
timestamp 18001
transform 1 0 5428 0 -1 52224
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_91_1013
timestamp 1636986456
transform 1 0 94300 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_1025
timestamp 1636986456
transform 1 0 95404 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_1037
timestamp 1636986456
transform 1 0 96508 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_3
timestamp 1636986456
transform 1 0 1380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_15
timestamp 1636986456
transform 1 0 2484 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_27
timestamp 18001
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_29
timestamp 1636986456
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_41
timestamp 18001
transform 1 0 4876 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_92_49
timestamp 18001
transform 1 0 5612 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_1013
timestamp 1636986456
transform 1 0 94300 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_1025
timestamp 1636986456
transform 1 0 95404 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_1037
timestamp 18001
transform 1 0 96508 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_92_1039
timestamp 18001
transform 1 0 96692 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_92_1047
timestamp 18001
transform 1 0 97428 0 1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_93_3
timestamp 1636986456
transform 1 0 1380 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_15
timestamp 1636986456
transform 1 0 2484 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_27
timestamp 1636986456
transform 1 0 3588 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_39
timestamp 18001
transform 1 0 4692 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_93_47
timestamp 18001
transform 1 0 5428 0 -1 53312
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_93_1013
timestamp 1636986456
transform 1 0 94300 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_1025
timestamp 1636986456
transform 1 0 95404 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_1037
timestamp 1636986456
transform 1 0 96508 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_3
timestamp 1636986456
transform 1 0 1380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_15
timestamp 1636986456
transform 1 0 2484 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_27
timestamp 18001
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_29
timestamp 1636986456
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_41
timestamp 18001
transform 1 0 4876 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_94_49
timestamp 18001
transform 1 0 5612 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_1013
timestamp 1636986456
transform 1 0 94300 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_1025
timestamp 1636986456
transform 1 0 95404 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_1037
timestamp 18001
transform 1 0 96508 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_94_1039
timestamp 18001
transform 1 0 96692 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_94_1047
timestamp 18001
transform 1 0 97428 0 1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_95_9
timestamp 1636986456
transform 1 0 1932 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_21
timestamp 1636986456
transform 1 0 3036 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_33
timestamp 1636986456
transform 1 0 4140 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_45
timestamp 18001
transform 1 0 5244 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_49
timestamp 18001
transform 1 0 5612 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_1013
timestamp 1636986456
transform 1 0 94300 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_1025
timestamp 1636986456
transform 1 0 95404 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_1037
timestamp 18001
transform 1 0 96508 0 -1 54400
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_96_9
timestamp 1636986456
transform 1 0 1932 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_21
timestamp 18001
transform 1 0 3036 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_27
timestamp 18001
transform 1 0 3588 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_29
timestamp 1636986456
transform 1 0 3772 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_96_41
timestamp 18001
transform 1 0 4876 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_96_49
timestamp 18001
transform 1 0 5612 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_1013
timestamp 1636986456
transform 1 0 94300 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_1025
timestamp 1636986456
transform 1 0 95404 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_1037
timestamp 18001
transform 1 0 96508 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_96_1039
timestamp 18001
transform 1 0 96692 0 1 54400
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_97_3
timestamp 1636986456
transform 1 0 1380 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_15
timestamp 1636986456
transform 1 0 2484 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_27
timestamp 1636986456
transform 1 0 3588 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_39
timestamp 18001
transform 1 0 4692 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_97_47
timestamp 18001
transform 1 0 5428 0 -1 55488
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_97_1013
timestamp 1636986456
transform 1 0 94300 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_1025
timestamp 1636986456
transform 1 0 95404 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_1037
timestamp 1636986456
transform 1 0 96508 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_3
timestamp 1636986456
transform 1 0 1380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_15
timestamp 1636986456
transform 1 0 2484 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_27
timestamp 18001
transform 1 0 3588 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_29
timestamp 1636986456
transform 1 0 3772 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_41
timestamp 18001
transform 1 0 4876 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_98_49
timestamp 18001
transform 1 0 5612 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_1013
timestamp 1636986456
transform 1 0 94300 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_1025
timestamp 1636986456
transform 1 0 95404 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_1037
timestamp 18001
transform 1 0 96508 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_98_1039
timestamp 18001
transform 1 0 96692 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_98_1047
timestamp 18001
transform 1 0 97428 0 1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_99_11
timestamp 1636986456
transform 1 0 2116 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_23
timestamp 1636986456
transform 1 0 3220 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_35
timestamp 1636986456
transform 1 0 4324 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_99_47
timestamp 18001
transform 1 0 5428 0 -1 56576
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_99_1013
timestamp 1636986456
transform 1 0 94300 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_1025
timestamp 1636986456
transform 1 0 95404 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_1037
timestamp 18001
transform 1 0 96508 0 -1 56576
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_100_3
timestamp 1636986456
transform 1 0 1380 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_15
timestamp 1636986456
transform 1 0 2484 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_27
timestamp 18001
transform 1 0 3588 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_29
timestamp 1636986456
transform 1 0 3772 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_41
timestamp 18001
transform 1 0 4876 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_100_49
timestamp 18001
transform 1 0 5612 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_1013
timestamp 1636986456
transform 1 0 94300 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_1025
timestamp 1636986456
transform 1 0 95404 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_1037
timestamp 18001
transform 1 0 96508 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_100_1039
timestamp 18001
transform 1 0 96692 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_100_1047
timestamp 18001
transform 1 0 97428 0 1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_101_11
timestamp 1636986456
transform 1 0 2116 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_23
timestamp 1636986456
transform 1 0 3220 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_35
timestamp 1636986456
transform 1 0 4324 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_47
timestamp 18001
transform 1 0 5428 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_1013
timestamp 1636986456
transform 1 0 94300 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_1025
timestamp 1636986456
transform 1 0 95404 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_1037
timestamp 18001
transform 1 0 96508 0 -1 57664
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_102_9
timestamp 1636986456
transform 1 0 1932 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_21
timestamp 18001
transform 1 0 3036 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_27
timestamp 18001
transform 1 0 3588 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_29
timestamp 1636986456
transform 1 0 3772 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_102_41
timestamp 18001
transform 1 0 4876 0 1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_102_49
timestamp 18001
transform 1 0 5612 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_1013
timestamp 1636986456
transform 1 0 94300 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_1025
timestamp 1636986456
transform 1 0 95404 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_102_1037
timestamp 18001
transform 1 0 96508 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_102_1039
timestamp 18001
transform 1 0 96692 0 1 57664
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_103_3
timestamp 1636986456
transform 1 0 1380 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_15
timestamp 1636986456
transform 1 0 2484 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_27
timestamp 1636986456
transform 1 0 3588 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_103_39
timestamp 18001
transform 1 0 4692 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_103_47
timestamp 18001
transform 1 0 5428 0 -1 58752
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_103_1013
timestamp 1636986456
transform 1 0 94300 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_1025
timestamp 1636986456
transform 1 0 95404 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_1037
timestamp 1636986456
transform 1 0 96508 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_3
timestamp 1636986456
transform 1 0 1380 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_15
timestamp 1636986456
transform 1 0 2484 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_104_27
timestamp 18001
transform 1 0 3588 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_29
timestamp 1636986456
transform 1 0 3772 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_104_41
timestamp 18001
transform 1 0 4876 0 1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_104_49
timestamp 18001
transform 1 0 5612 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_1013
timestamp 1636986456
transform 1 0 94300 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_1025
timestamp 1636986456
transform 1 0 95404 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_104_1037
timestamp 18001
transform 1 0 96508 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_104_1039
timestamp 18001
transform 1 0 96692 0 1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_104_1047
timestamp 18001
transform 1 0 97428 0 1 58752
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_105_9
timestamp 1636986456
transform 1 0 1932 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_21
timestamp 1636986456
transform 1 0 3036 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_33
timestamp 1636986456
transform 1 0 4140 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_105_45
timestamp 18001
transform 1 0 5244 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_105_49
timestamp 18001
transform 1 0 5612 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_1013
timestamp 1636986456
transform 1 0 94300 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_1025
timestamp 1636986456
transform 1 0 95404 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_105_1037
timestamp 18001
transform 1 0 96508 0 -1 59840
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_106_11
timestamp 1636986456
transform 1 0 2116 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_106_23
timestamp 18001
transform 1 0 3220 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_106_27
timestamp 18001
transform 1 0 3588 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_29
timestamp 1636986456
transform 1 0 3772 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_106_41
timestamp 18001
transform 1 0 4876 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_106_49
timestamp 18001
transform 1 0 5612 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_1013
timestamp 1636986456
transform 1 0 94300 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_1025
timestamp 1636986456
transform 1 0 95404 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_106_1037
timestamp 18001
transform 1 0 96508 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_106_1039
timestamp 18001
transform 1 0 96692 0 1 59840
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_107_3
timestamp 1636986456
transform 1 0 1380 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_15
timestamp 1636986456
transform 1 0 2484 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_27
timestamp 1636986456
transform 1 0 3588 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_39
timestamp 18001
transform 1 0 4692 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_107_47
timestamp 18001
transform 1 0 5428 0 -1 60928
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_107_1013
timestamp 1636986456
transform 1 0 94300 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_1025
timestamp 1636986456
transform 1 0 95404 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_1037
timestamp 1636986456
transform 1 0 96508 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_3
timestamp 1636986456
transform 1 0 1380 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_15
timestamp 1636986456
transform 1 0 2484 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_108_27
timestamp 18001
transform 1 0 3588 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_29
timestamp 1636986456
transform 1 0 3772 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_108_41
timestamp 18001
transform 1 0 4876 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_108_49
timestamp 18001
transform 1 0 5612 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_1013
timestamp 1636986456
transform 1 0 94300 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_1025
timestamp 1636986456
transform 1 0 95404 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_108_1037
timestamp 18001
transform 1 0 96508 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_108_1039
timestamp 18001
transform 1 0 96692 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_108_1047
timestamp 18001
transform 1 0 97428 0 1 60928
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_109_9
timestamp 1636986456
transform 1 0 1932 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_21
timestamp 1636986456
transform 1 0 3036 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_33
timestamp 1636986456
transform 1 0 4140 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_109_45
timestamp 18001
transform 1 0 5244 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_109_49
timestamp 18001
transform 1 0 5612 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_1013
timestamp 1636986456
transform 1 0 94300 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_1025
timestamp 1636986456
transform 1 0 95404 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_109_1037
timestamp 18001
transform 1 0 96508 0 -1 62016
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_110_3
timestamp 1636986456
transform 1 0 1380 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_15
timestamp 1636986456
transform 1 0 2484 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_110_27
timestamp 18001
transform 1 0 3588 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_29
timestamp 1636986456
transform 1 0 3772 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_110_41
timestamp 18001
transform 1 0 4876 0 1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_110_49
timestamp 18001
transform 1 0 5612 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_1013
timestamp 1636986456
transform 1 0 94300 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_1025
timestamp 1636986456
transform 1 0 95404 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_110_1037
timestamp 18001
transform 1 0 96508 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_110_1039
timestamp 18001
transform 1 0 96692 0 1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_110_1047
timestamp 18001
transform 1 0 97428 0 1 62016
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_111_11
timestamp 1636986456
transform 1 0 2116 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_23
timestamp 1636986456
transform 1 0 3220 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_35
timestamp 1636986456
transform 1 0 4324 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_111_47
timestamp 18001
transform 1 0 5428 0 -1 63104
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_111_1013
timestamp 1636986456
transform 1 0 94300 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_1025
timestamp 1636986456
transform 1 0 95404 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_111_1037
timestamp 18001
transform 1 0 96508 0 -1 63104
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_112_9
timestamp 1636986456
transform 1 0 1932 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_21
timestamp 18001
transform 1 0 3036 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_27
timestamp 18001
transform 1 0 3588 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_29
timestamp 1636986456
transform 1 0 3772 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_112_41
timestamp 18001
transform 1 0 4876 0 1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_112_49
timestamp 18001
transform 1 0 5612 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_1013
timestamp 1636986456
transform 1 0 94300 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_1025
timestamp 1636986456
transform 1 0 95404 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_112_1037
timestamp 18001
transform 1 0 96508 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_112_1039
timestamp 18001
transform 1 0 96692 0 1 63104
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_113_3
timestamp 1636986456
transform 1 0 1380 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_15
timestamp 1636986456
transform 1 0 2484 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_27
timestamp 1636986456
transform 1 0 3588 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_113_39
timestamp 18001
transform 1 0 4692 0 -1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_113_47
timestamp 18001
transform 1 0 5428 0 -1 64192
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_113_1013
timestamp 1636986456
transform 1 0 94300 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_1025
timestamp 1636986456
transform 1 0 95404 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_1037
timestamp 1636986456
transform 1 0 96508 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_3
timestamp 1636986456
transform 1 0 1380 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_15
timestamp 1636986456
transform 1 0 2484 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_114_27
timestamp 18001
transform 1 0 3588 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_29
timestamp 1636986456
transform 1 0 3772 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_114_41
timestamp 18001
transform 1 0 4876 0 1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_114_49
timestamp 18001
transform 1 0 5612 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_1013
timestamp 1636986456
transform 1 0 94300 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_1025
timestamp 1636986456
transform 1 0 95404 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_114_1037
timestamp 18001
transform 1 0 96508 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_114_1039
timestamp 18001
transform 1 0 96692 0 1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_114_1047
timestamp 18001
transform 1 0 97428 0 1 64192
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_115_9
timestamp 1636986456
transform 1 0 1932 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_21
timestamp 1636986456
transform 1 0 3036 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_33
timestamp 1636986456
transform 1 0 4140 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_115_45
timestamp 18001
transform 1 0 5244 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_115_49
timestamp 18001
transform 1 0 5612 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_1013
timestamp 1636986456
transform 1 0 94300 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_1025
timestamp 1636986456
transform 1 0 95404 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_115_1037
timestamp 18001
transform 1 0 96508 0 -1 65280
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_116_9
timestamp 1636986456
transform 1 0 1932 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_21
timestamp 18001
transform 1 0 3036 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_27
timestamp 18001
transform 1 0 3588 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_29
timestamp 1636986456
transform 1 0 3772 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_116_41
timestamp 18001
transform 1 0 4876 0 1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_116_49
timestamp 18001
transform 1 0 5612 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_1013
timestamp 1636986456
transform 1 0 94300 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_1025
timestamp 1636986456
transform 1 0 95404 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_116_1037
timestamp 18001
transform 1 0 96508 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_116_1039
timestamp 18001
transform 1 0 96692 0 1 65280
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_117_3
timestamp 1636986456
transform 1 0 1380 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_15
timestamp 1636986456
transform 1 0 2484 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_27
timestamp 1636986456
transform 1 0 3588 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_117_39
timestamp 18001
transform 1 0 4692 0 -1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_117_47
timestamp 18001
transform 1 0 5428 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_1013
timestamp 1636986456
transform 1 0 94300 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_1025
timestamp 1636986456
transform 1 0 95404 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_1037
timestamp 1636986456
transform 1 0 96508 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_3
timestamp 1636986456
transform 1 0 1380 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_15
timestamp 1636986456
transform 1 0 2484 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_118_27
timestamp 18001
transform 1 0 3588 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_29
timestamp 1636986456
transform 1 0 3772 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_118_41
timestamp 18001
transform 1 0 4876 0 1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_118_49
timestamp 18001
transform 1 0 5612 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_1013
timestamp 1636986456
transform 1 0 94300 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_1025
timestamp 1636986456
transform 1 0 95404 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_118_1037
timestamp 18001
transform 1 0 96508 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_118_1039
timestamp 18001
transform 1 0 96692 0 1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_118_1047
timestamp 18001
transform 1 0 97428 0 1 66368
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_119_9
timestamp 1636986456
transform 1 0 1932 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_21
timestamp 1636986456
transform 1 0 3036 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_33
timestamp 1636986456
transform 1 0 4140 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_119_45
timestamp 18001
transform 1 0 5244 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_119_49
timestamp 18001
transform 1 0 5612 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_1013
timestamp 1636986456
transform 1 0 94300 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_1025
timestamp 1636986456
transform 1 0 95404 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_119_1037
timestamp 18001
transform 1 0 96508 0 -1 67456
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_120_3
timestamp 1636986456
transform 1 0 1380 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_15
timestamp 1636986456
transform 1 0 2484 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_120_27
timestamp 18001
transform 1 0 3588 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_29
timestamp 1636986456
transform 1 0 3772 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_120_41
timestamp 18001
transform 1 0 4876 0 1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_120_49
timestamp 18001
transform 1 0 5612 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_1013
timestamp 1636986456
transform 1 0 94300 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_1025
timestamp 1636986456
transform 1 0 95404 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_120_1037
timestamp 18001
transform 1 0 96508 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_120_1039
timestamp 18001
transform 1 0 96692 0 1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_120_1047
timestamp 18001
transform 1 0 97428 0 1 67456
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_121_9
timestamp 1636986456
transform 1 0 1932 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_21
timestamp 1636986456
transform 1 0 3036 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_33
timestamp 1636986456
transform 1 0 4140 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_121_45
timestamp 18001
transform 1 0 5244 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_121_49
timestamp 18001
transform 1 0 5612 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_1013
timestamp 1636986456
transform 1 0 94300 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_1025
timestamp 1636986456
transform 1 0 95404 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_121_1037
timestamp 18001
transform 1 0 96508 0 -1 68544
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_122_9
timestamp 1636986456
transform 1 0 1932 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_21
timestamp 18001
transform 1 0 3036 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_27
timestamp 18001
transform 1 0 3588 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_29
timestamp 1636986456
transform 1 0 3772 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_122_41
timestamp 18001
transform 1 0 4876 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_122_49
timestamp 18001
transform 1 0 5612 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_1013
timestamp 1636986456
transform 1 0 94300 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_1025
timestamp 1636986456
transform 1 0 95404 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_122_1037
timestamp 18001
transform 1 0 96508 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_122_1039
timestamp 18001
transform 1 0 96692 0 1 68544
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_123_3
timestamp 1636986456
transform 1 0 1380 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_15
timestamp 1636986456
transform 1 0 2484 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_27
timestamp 1636986456
transform 1 0 3588 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_123_39
timestamp 18001
transform 1 0 4692 0 -1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_123_47
timestamp 18001
transform 1 0 5428 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_1013
timestamp 1636986456
transform 1 0 94300 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_1025
timestamp 1636986456
transform 1 0 95404 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_1037
timestamp 1636986456
transform 1 0 96508 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_3
timestamp 1636986456
transform 1 0 1380 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_15
timestamp 1636986456
transform 1 0 2484 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_124_27
timestamp 18001
transform 1 0 3588 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_124_29
timestamp 18001
transform 1 0 3772 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_1013
timestamp 1636986456
transform 1 0 94300 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_1025
timestamp 1636986456
transform 1 0 95404 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_124_1037
timestamp 18001
transform 1 0 96508 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_124_1039
timestamp 18001
transform 1 0 96692 0 1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_124_1047
timestamp 18001
transform 1 0 97428 0 1 69632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_125_8
timestamp 1636986456
transform 1 0 1840 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_20
timestamp 1636986456
transform 1 0 2944 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_32
timestamp 1636986456
transform 1 0 4048 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_125_44
timestamp 18001
transform 1 0 5152 0 -1 70720
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_125_1013
timestamp 1636986456
transform 1 0 94300 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_1025
timestamp 1636986456
transform 1 0 95404 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_125_1037
timestamp 18001
transform 1 0 96508 0 -1 70720
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_126_7
timestamp 1636986456
transform 1 0 1748 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_126_19
timestamp 18001
transform 1 0 2852 0 1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_126_27
timestamp 18001
transform 1 0 3588 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_29
timestamp 1636986456
transform 1 0 3772 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_126_41
timestamp 18001
transform 1 0 4876 0 1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_126_49
timestamp 18001
transform 1 0 5612 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_1013
timestamp 1636986456
transform 1 0 94300 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_1025
timestamp 1636986456
transform 1 0 95404 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_126_1037
timestamp 18001
transform 1 0 96508 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_126_1039
timestamp 18001
transform 1 0 96692 0 1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_126_1043
timestamp 18001
transform 1 0 97060 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_3
timestamp 1636986456
transform 1 0 1380 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_15
timestamp 1636986456
transform 1 0 2484 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_27
timestamp 1636986456
transform 1 0 3588 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_127_39
timestamp 18001
transform 1 0 4692 0 -1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_127_47
timestamp 18001
transform 1 0 5428 0 -1 71808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_127_1013
timestamp 1636986456
transform 1 0 94300 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_1025
timestamp 1636986456
transform 1 0 95404 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_1037
timestamp 1636986456
transform 1 0 96508 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_3
timestamp 1636986456
transform 1 0 1380 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_15
timestamp 1636986456
transform 1 0 2484 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_128_27
timestamp 18001
transform 1 0 3588 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_29
timestamp 1636986456
transform 1 0 3772 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_128_41
timestamp 18001
transform 1 0 4876 0 1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_128_49
timestamp 18001
transform 1 0 5612 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_1013
timestamp 1636986456
transform 1 0 94300 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_1025
timestamp 1636986456
transform 1 0 95404 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_128_1037
timestamp 18001
transform 1 0 96508 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_128_1039
timestamp 18001
transform 1 0 96692 0 1 71808
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_129_7
timestamp 1636986456
transform 1 0 1748 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_19
timestamp 1636986456
transform 1 0 2852 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_31
timestamp 1636986456
transform 1 0 3956 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_43
timestamp 18001
transform 1 0 5060 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_49
timestamp 18001
transform 1 0 5612 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_1013
timestamp 1636986456
transform 1 0 94300 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_1025
timestamp 1636986456
transform 1 0 95404 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_129_1037
timestamp 18001
transform 1 0 96508 0 -1 72896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_130_3
timestamp 1636986456
transform 1 0 1380 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_15
timestamp 1636986456
transform 1 0 2484 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_130_27
timestamp 18001
transform 1 0 3588 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_29
timestamp 1636986456
transform 1 0 3772 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_130_41
timestamp 18001
transform 1 0 4876 0 1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_130_49
timestamp 18001
transform 1 0 5612 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_1013
timestamp 1636986456
transform 1 0 94300 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_1025
timestamp 1636986456
transform 1 0 95404 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_130_1037
timestamp 18001
transform 1 0 96508 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_130_1039
timestamp 18001
transform 1 0 96692 0 1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_130_1047
timestamp 18001
transform 1 0 97428 0 1 72896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_131_7
timestamp 1636986456
transform 1 0 1748 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_19
timestamp 1636986456
transform 1 0 2852 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_31
timestamp 1636986456
transform 1 0 3956 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_43
timestamp 18001
transform 1 0 5060 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_49
timestamp 18001
transform 1 0 5612 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_1013
timestamp 1636986456
transform 1 0 94300 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_1025
timestamp 1636986456
transform 1 0 95404 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_1037
timestamp 18001
transform 1 0 96508 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_1043
timestamp 18001
transform 1 0 97060 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_7
timestamp 1636986456
transform 1 0 1748 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_132_19
timestamp 18001
transform 1 0 2852 0 1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_132_27
timestamp 18001
transform 1 0 3588 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_29
timestamp 1636986456
transform 1 0 3772 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_132_41
timestamp 18001
transform 1 0 4876 0 1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_132_49
timestamp 18001
transform 1 0 5612 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_1013
timestamp 1636986456
transform 1 0 94300 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_1025
timestamp 1636986456
transform 1 0 95404 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_132_1037
timestamp 18001
transform 1 0 96508 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_132_1039
timestamp 18001
transform 1 0 96692 0 1 73984
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_133_3
timestamp 1636986456
transform 1 0 1380 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_15
timestamp 1636986456
transform 1 0 2484 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_27
timestamp 1636986456
transform 1 0 3588 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_133_39
timestamp 18001
transform 1 0 4692 0 -1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_133_47
timestamp 18001
transform 1 0 5428 0 -1 75072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_133_1013
timestamp 1636986456
transform 1 0 94300 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_1025
timestamp 1636986456
transform 1 0 95404 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_1037
timestamp 1636986456
transform 1 0 96508 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_3
timestamp 1636986456
transform 1 0 1380 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_15
timestamp 1636986456
transform 1 0 2484 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_134_27
timestamp 18001
transform 1 0 3588 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_29
timestamp 1636986456
transform 1 0 3772 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_134_41
timestamp 18001
transform 1 0 4876 0 1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_134_49
timestamp 18001
transform 1 0 5612 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_1013
timestamp 1636986456
transform 1 0 94300 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_1025
timestamp 1636986456
transform 1 0 95404 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_134_1037
timestamp 18001
transform 1 0 96508 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_134_1039
timestamp 18001
transform 1 0 96692 0 1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_134_1047
timestamp 18001
transform 1 0 97428 0 1 75072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_135_7
timestamp 1636986456
transform 1 0 1748 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_19
timestamp 1636986456
transform 1 0 2852 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_31
timestamp 1636986456
transform 1 0 3956 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_43
timestamp 18001
transform 1 0 5060 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_49
timestamp 18001
transform 1 0 5612 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_1013
timestamp 1636986456
transform 1 0 94300 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_1025
timestamp 1636986456
transform 1 0 95404 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_1037
timestamp 18001
transform 1 0 96508 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_1043
timestamp 18001
transform 1 0 97060 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_7
timestamp 1636986456
transform 1 0 1748 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_136_19
timestamp 18001
transform 1 0 2852 0 1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_136_27
timestamp 18001
transform 1 0 3588 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_29
timestamp 1636986456
transform 1 0 3772 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_136_41
timestamp 18001
transform 1 0 4876 0 1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_136_49
timestamp 18001
transform 1 0 5612 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_1013
timestamp 1636986456
transform 1 0 94300 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_1025
timestamp 1636986456
transform 1 0 95404 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_136_1037
timestamp 18001
transform 1 0 96508 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_136_1039
timestamp 18001
transform 1 0 96692 0 1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_136_1043
timestamp 18001
transform 1 0 97060 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_3
timestamp 1636986456
transform 1 0 1380 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_15
timestamp 1636986456
transform 1 0 2484 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_27
timestamp 1636986456
transform 1 0 3588 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_137_39
timestamp 18001
transform 1 0 4692 0 -1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_137_47
timestamp 18001
transform 1 0 5428 0 -1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_137_1013
timestamp 1636986456
transform 1 0 94300 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_1025
timestamp 1636986456
transform 1 0 95404 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_1037
timestamp 1636986456
transform 1 0 96508 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_3
timestamp 1636986456
transform 1 0 1380 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_15
timestamp 1636986456
transform 1 0 2484 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_138_27
timestamp 18001
transform 1 0 3588 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_138_29
timestamp 1636986456
transform 1 0 3772 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_138_41
timestamp 18001
transform 1 0 4876 0 1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_138_49
timestamp 18001
transform 1 0 5612 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_138_1013
timestamp 1636986456
transform 1 0 94300 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_1025
timestamp 1636986456
transform 1 0 95404 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_138_1037
timestamp 18001
transform 1 0 96508 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_138_1039
timestamp 18001
transform 1 0 96692 0 1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_138_1047
timestamp 18001
transform 1 0 97428 0 1 77248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_139_7
timestamp 1636986456
transform 1 0 1748 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_19
timestamp 1636986456
transform 1 0 2852 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_31
timestamp 1636986456
transform 1 0 3956 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_139_43
timestamp 18001
transform 1 0 5060 0 -1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_139_49
timestamp 18001
transform 1 0 5612 0 -1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_139_1013
timestamp 1636986456
transform 1 0 94300 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_1025
timestamp 1636986456
transform 1 0 95404 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_139_1037
timestamp 18001
transform 1 0 96508 0 -1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_139_1043
timestamp 18001
transform 1 0 97060 0 -1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_140_3
timestamp 1636986456
transform 1 0 1380 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_15
timestamp 1636986456
transform 1 0 2484 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_140_27
timestamp 18001
transform 1 0 3588 0 1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_140_29
timestamp 1636986456
transform 1 0 3772 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_140_41
timestamp 18001
transform 1 0 4876 0 1 78336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_140_49
timestamp 18001
transform 1 0 5612 0 1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_140_1013
timestamp 1636986456
transform 1 0 94300 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_1025
timestamp 1636986456
transform 1 0 95404 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_140_1037
timestamp 18001
transform 1 0 96508 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_140_1039
timestamp 18001
transform 1 0 96692 0 1 78336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_140_1047
timestamp 18001
transform 1 0 97428 0 1 78336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_141_7
timestamp 1636986456
transform 1 0 1748 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_19
timestamp 1636986456
transform 1 0 2852 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_31
timestamp 1636986456
transform 1 0 3956 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_141_43
timestamp 18001
transform 1 0 5060 0 -1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_141_49
timestamp 18001
transform 1 0 5612 0 -1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_141_1013
timestamp 1636986456
transform 1 0 94300 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_1025
timestamp 1636986456
transform 1 0 95404 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_141_1037
timestamp 18001
transform 1 0 96508 0 -1 79424
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_142_7
timestamp 1636986456
transform 1 0 1748 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_142_19
timestamp 18001
transform 1 0 2852 0 1 79424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_142_27
timestamp 18001
transform 1 0 3588 0 1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_142_29
timestamp 1636986456
transform 1 0 3772 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_142_41
timestamp 18001
transform 1 0 4876 0 1 79424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_142_49
timestamp 18001
transform 1 0 5612 0 1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_142_1013
timestamp 1636986456
transform 1 0 94300 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_1025
timestamp 1636986456
transform 1 0 95404 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_142_1037
timestamp 18001
transform 1 0 96508 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_142_1039
timestamp 18001
transform 1 0 96692 0 1 79424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_142_1043
timestamp 18001
transform 1 0 97060 0 1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_143_3
timestamp 1636986456
transform 1 0 1380 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_15
timestamp 1636986456
transform 1 0 2484 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_27
timestamp 1636986456
transform 1 0 3588 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_143_39
timestamp 18001
transform 1 0 4692 0 -1 80512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_143_47
timestamp 18001
transform 1 0 5428 0 -1 80512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_143_1013
timestamp 1636986456
transform 1 0 94300 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_1025
timestamp 1636986456
transform 1 0 95404 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_1037
timestamp 1636986456
transform 1 0 96508 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_3
timestamp 1636986456
transform 1 0 1380 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_15
timestamp 1636986456
transform 1 0 2484 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_144_27
timestamp 18001
transform 1 0 3588 0 1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_144_29
timestamp 1636986456
transform 1 0 3772 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_144_41
timestamp 18001
transform 1 0 4876 0 1 80512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_144_49
timestamp 18001
transform 1 0 5612 0 1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_144_1013
timestamp 1636986456
transform 1 0 94300 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_1025
timestamp 1636986456
transform 1 0 95404 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_144_1037
timestamp 18001
transform 1 0 96508 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_144_1039
timestamp 18001
transform 1 0 96692 0 1 80512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_144_1047
timestamp 18001
transform 1 0 97428 0 1 80512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_145_7
timestamp 1636986456
transform 1 0 1748 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_19
timestamp 1636986456
transform 1 0 2852 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_31
timestamp 1636986456
transform 1 0 3956 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_145_43
timestamp 18001
transform 1 0 5060 0 -1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_145_49
timestamp 18001
transform 1 0 5612 0 -1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_145_1013
timestamp 1636986456
transform 1 0 94300 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_1025
timestamp 1636986456
transform 1 0 95404 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_145_1037
timestamp 18001
transform 1 0 96508 0 -1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_145_1043
timestamp 18001
transform 1 0 97060 0 -1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_146_7
timestamp 1636986456
transform 1 0 1748 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_146_19
timestamp 18001
transform 1 0 2852 0 1 81600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_146_27
timestamp 18001
transform 1 0 3588 0 1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_146_29
timestamp 1636986456
transform 1 0 3772 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_146_41
timestamp 18001
transform 1 0 4876 0 1 81600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_146_49
timestamp 18001
transform 1 0 5612 0 1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_146_1013
timestamp 1636986456
transform 1 0 94300 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_1025
timestamp 1636986456
transform 1 0 95404 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_146_1037
timestamp 18001
transform 1 0 96508 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_146_1039
timestamp 18001
transform 1 0 96692 0 1 81600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_146_1043
timestamp 18001
transform 1 0 97060 0 1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_3
timestamp 1636986456
transform 1 0 1380 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_15
timestamp 1636986456
transform 1 0 2484 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_27
timestamp 1636986456
transform 1 0 3588 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_147_39
timestamp 18001
transform 1 0 4692 0 -1 82688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_147_47
timestamp 18001
transform 1 0 5428 0 -1 82688
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_147_1013
timestamp 1636986456
transform 1 0 94300 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_1025
timestamp 1636986456
transform 1 0 95404 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_1037
timestamp 1636986456
transform 1 0 96508 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_3
timestamp 1636986456
transform 1 0 1380 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_15
timestamp 1636986456
transform 1 0 2484 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_148_27
timestamp 18001
transform 1 0 3588 0 1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_29
timestamp 1636986456
transform 1 0 3772 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_148_41
timestamp 18001
transform 1 0 4876 0 1 82688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_148_49
timestamp 18001
transform 1 0 5612 0 1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_1013
timestamp 1636986456
transform 1 0 94300 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_1025
timestamp 1636986456
transform 1 0 95404 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_148_1037
timestamp 18001
transform 1 0 96508 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_148_1039
timestamp 18001
transform 1 0 96692 0 1 82688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_148_1047
timestamp 18001
transform 1 0 97428 0 1 82688
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_149_7
timestamp 1636986456
transform 1 0 1748 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_19
timestamp 1636986456
transform 1 0 2852 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_31
timestamp 1636986456
transform 1 0 3956 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_43
timestamp 18001
transform 1 0 5060 0 -1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_49
timestamp 18001
transform 1 0 5612 0 -1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_1013
timestamp 1636986456
transform 1 0 94300 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_1025
timestamp 1636986456
transform 1 0 95404 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_1037
timestamp 18001
transform 1 0 96508 0 -1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_1043
timestamp 18001
transform 1 0 97060 0 -1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_3
timestamp 1636986456
transform 1 0 1380 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_15
timestamp 1636986456
transform 1 0 2484 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_150_27
timestamp 18001
transform 1 0 3588 0 1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_29
timestamp 1636986456
transform 1 0 3772 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_150_41
timestamp 18001
transform 1 0 4876 0 1 83776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_150_49
timestamp 18001
transform 1 0 5612 0 1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_1013
timestamp 1636986456
transform 1 0 94300 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_1025
timestamp 1636986456
transform 1 0 95404 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_150_1037
timestamp 18001
transform 1 0 96508 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_150_1039
timestamp 18001
transform 1 0 96692 0 1 83776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_150_1047
timestamp 18001
transform 1 0 97428 0 1 83776
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_151_7
timestamp 1636986456
transform 1 0 1748 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_19
timestamp 1636986456
transform 1 0 2852 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_31
timestamp 1636986456
transform 1 0 3956 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_151_43
timestamp 18001
transform 1 0 5060 0 -1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_49
timestamp 18001
transform 1 0 5612 0 -1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_151_1013
timestamp 1636986456
transform 1 0 94300 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_1025
timestamp 1636986456
transform 1 0 95404 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_151_1037
timestamp 18001
transform 1 0 96508 0 -1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_1043
timestamp 18001
transform 1 0 97060 0 -1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_152_7
timestamp 1636986456
transform 1 0 1748 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_152_19
timestamp 18001
transform 1 0 2852 0 1 84864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_152_27
timestamp 18001
transform 1 0 3588 0 1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_152_29
timestamp 1636986456
transform 1 0 3772 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_152_41
timestamp 18001
transform 1 0 4876 0 1 84864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_152_49
timestamp 18001
transform 1 0 5612 0 1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_152_1013
timestamp 1636986456
transform 1 0 94300 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_1025
timestamp 1636986456
transform 1 0 95404 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_152_1037
timestamp 18001
transform 1 0 96508 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_152_1039
timestamp 18001
transform 1 0 96692 0 1 84864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_152_1043
timestamp 18001
transform 1 0 97060 0 1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_153_3
timestamp 1636986456
transform 1 0 1380 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_15
timestamp 1636986456
transform 1 0 2484 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_27
timestamp 1636986456
transform 1 0 3588 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_153_39
timestamp 18001
transform 1 0 4692 0 -1 85952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_153_47
timestamp 18001
transform 1 0 5428 0 -1 85952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_153_1013
timestamp 1636986456
transform 1 0 94300 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_1025
timestamp 1636986456
transform 1 0 95404 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_1037
timestamp 1636986456
transform 1 0 96508 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_3
timestamp 1636986456
transform 1 0 1380 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_15
timestamp 1636986456
transform 1 0 2484 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_154_27
timestamp 18001
transform 1 0 3588 0 1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_154_29
timestamp 1636986456
transform 1 0 3772 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_154_41
timestamp 18001
transform 1 0 4876 0 1 85952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_154_49
timestamp 18001
transform 1 0 5612 0 1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_154_1013
timestamp 1636986456
transform 1 0 94300 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_1025
timestamp 1636986456
transform 1 0 95404 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_154_1037
timestamp 18001
transform 1 0 96508 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_154_1039
timestamp 18001
transform 1 0 96692 0 1 85952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_154_1047
timestamp 18001
transform 1 0 97428 0 1 85952
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_155_7
timestamp 1636986456
transform 1 0 1748 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_19
timestamp 1636986456
transform 1 0 2852 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_31
timestamp 1636986456
transform 1 0 3956 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_155_43
timestamp 18001
transform 1 0 5060 0 -1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_155_49
timestamp 18001
transform 1 0 5612 0 -1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_155_1013
timestamp 1636986456
transform 1 0 94300 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_1025
timestamp 1636986456
transform 1 0 95404 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_155_1037
timestamp 18001
transform 1 0 96508 0 -1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_155_1043
timestamp 18001
transform 1 0 97060 0 -1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_156_7
timestamp 1636986456
transform 1 0 1748 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_156_19
timestamp 18001
transform 1 0 2852 0 1 87040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_156_27
timestamp 18001
transform 1 0 3588 0 1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_156_29
timestamp 1636986456
transform 1 0 3772 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_156_41
timestamp 18001
transform 1 0 4876 0 1 87040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_156_49
timestamp 18001
transform 1 0 5612 0 1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_156_1013
timestamp 1636986456
transform 1 0 94300 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_1025
timestamp 1636986456
transform 1 0 95404 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_156_1037
timestamp 18001
transform 1 0 96508 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_156_1039
timestamp 18001
transform 1 0 96692 0 1 87040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_156_1043
timestamp 18001
transform 1 0 97060 0 1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_157_3
timestamp 1636986456
transform 1 0 1380 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_15
timestamp 1636986456
transform 1 0 2484 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_27
timestamp 1636986456
transform 1 0 3588 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_157_39
timestamp 18001
transform 1 0 4692 0 -1 88128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_157_47
timestamp 18001
transform 1 0 5428 0 -1 88128
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_157_1013
timestamp 1636986456
transform 1 0 94300 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_1025
timestamp 1636986456
transform 1 0 95404 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_1037
timestamp 1636986456
transform 1 0 96508 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_3
timestamp 1636986456
transform 1 0 1380 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_15
timestamp 1636986456
transform 1 0 2484 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_158_27
timestamp 18001
transform 1 0 3588 0 1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_158_29
timestamp 1636986456
transform 1 0 3772 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_158_41
timestamp 18001
transform 1 0 4876 0 1 88128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_158_49
timestamp 18001
transform 1 0 5612 0 1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_158_1013
timestamp 1636986456
transform 1 0 94300 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_1025
timestamp 1636986456
transform 1 0 95404 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_158_1037
timestamp 18001
transform 1 0 96508 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_158_1039
timestamp 18001
transform 1 0 96692 0 1 88128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_158_1047
timestamp 18001
transform 1 0 97428 0 1 88128
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_159_3
timestamp 1636986456
transform 1 0 1380 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_15
timestamp 1636986456
transform 1 0 2484 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_27
timestamp 1636986456
transform 1 0 3588 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_159_39
timestamp 18001
transform 1 0 4692 0 -1 89216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_159_47
timestamp 18001
transform 1 0 5428 0 -1 89216
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_159_1013
timestamp 1636986456
transform 1 0 94300 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_1025
timestamp 1636986456
transform 1 0 95404 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_1037
timestamp 1636986456
transform 1 0 96508 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_3
timestamp 1636986456
transform 1 0 1380 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_15
timestamp 1636986456
transform 1 0 2484 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_160_27
timestamp 18001
transform 1 0 3588 0 1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_160_29
timestamp 1636986456
transform 1 0 3772 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_160_41
timestamp 18001
transform 1 0 4876 0 1 89216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_160_49
timestamp 18001
transform 1 0 5612 0 1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_160_1013
timestamp 1636986456
transform 1 0 94300 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_1025
timestamp 1636986456
transform 1 0 95404 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_160_1037
timestamp 18001
transform 1 0 96508 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_160_1039
timestamp 18001
transform 1 0 96692 0 1 89216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_160_1047
timestamp 18001
transform 1 0 97428 0 1 89216
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_161_3
timestamp 1636986456
transform 1 0 1380 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_15
timestamp 1636986456
transform 1 0 2484 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_27
timestamp 1636986456
transform 1 0 3588 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_161_39
timestamp 18001
transform 1 0 4692 0 -1 90304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_161_47
timestamp 18001
transform 1 0 5428 0 -1 90304
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_161_1013
timestamp 1636986456
transform 1 0 94300 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_1025
timestamp 1636986456
transform 1 0 95404 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_1037
timestamp 1636986456
transform 1 0 96508 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_3
timestamp 1636986456
transform 1 0 1380 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_15
timestamp 1636986456
transform 1 0 2484 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_162_27
timestamp 18001
transform 1 0 3588 0 1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_162_29
timestamp 1636986456
transform 1 0 3772 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_162_41
timestamp 18001
transform 1 0 4876 0 1 90304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_162_49
timestamp 18001
transform 1 0 5612 0 1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_162_1013
timestamp 1636986456
transform 1 0 94300 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_1025
timestamp 1636986456
transform 1 0 95404 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_162_1037
timestamp 18001
transform 1 0 96508 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_162_1039
timestamp 18001
transform 1 0 96692 0 1 90304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_162_1047
timestamp 18001
transform 1 0 97428 0 1 90304
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_163_3
timestamp 1636986456
transform 1 0 1380 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_15
timestamp 1636986456
transform 1 0 2484 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_27
timestamp 1636986456
transform 1 0 3588 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_163_39
timestamp 18001
transform 1 0 4692 0 -1 91392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_163_47
timestamp 18001
transform 1 0 5428 0 -1 91392
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_163_1013
timestamp 1636986456
transform 1 0 94300 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_1025
timestamp 1636986456
transform 1 0 95404 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_1037
timestamp 1636986456
transform 1 0 96508 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_3
timestamp 1636986456
transform 1 0 1380 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_15
timestamp 1636986456
transform 1 0 2484 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_164_27
timestamp 18001
transform 1 0 3588 0 1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_164_29
timestamp 1636986456
transform 1 0 3772 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_164_41
timestamp 18001
transform 1 0 4876 0 1 91392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_164_49
timestamp 18001
transform 1 0 5612 0 1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_164_1013
timestamp 1636986456
transform 1 0 94300 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_1025
timestamp 1636986456
transform 1 0 95404 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_164_1037
timestamp 18001
transform 1 0 96508 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_164_1039
timestamp 18001
transform 1 0 96692 0 1 91392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_164_1047
timestamp 18001
transform 1 0 97428 0 1 91392
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_165_3
timestamp 1636986456
transform 1 0 1380 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_15
timestamp 1636986456
transform 1 0 2484 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_27
timestamp 1636986456
transform 1 0 3588 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_165_39
timestamp 18001
transform 1 0 4692 0 -1 92480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_165_47
timestamp 18001
transform 1 0 5428 0 -1 92480
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_165_1013
timestamp 1636986456
transform 1 0 94300 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_1025
timestamp 1636986456
transform 1 0 95404 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_1037
timestamp 1636986456
transform 1 0 96508 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_3
timestamp 1636986456
transform 1 0 1380 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_15
timestamp 1636986456
transform 1 0 2484 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_166_27
timestamp 18001
transform 1 0 3588 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_29
timestamp 1636986456
transform 1 0 3772 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_166_41
timestamp 18001
transform 1 0 4876 0 1 92480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_166_49
timestamp 18001
transform 1 0 5612 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_1013
timestamp 1636986456
transform 1 0 94300 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_1025
timestamp 1636986456
transform 1 0 95404 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_166_1037
timestamp 18001
transform 1 0 96508 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_166_1039
timestamp 18001
transform 1 0 96692 0 1 92480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_166_1047
timestamp 18001
transform 1 0 97428 0 1 92480
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_167_3
timestamp 1636986456
transform 1 0 1380 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_15
timestamp 1636986456
transform 1 0 2484 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_167_27
timestamp 18001
transform 1 0 3588 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_29
timestamp 1636986456
transform 1 0 3772 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_41
timestamp 1636986456
transform 1 0 4876 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_167_53
timestamp 18001
transform 1 0 5980 0 -1 93568
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_167_57
timestamp 1636986456
transform 1 0 6348 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_69
timestamp 1636986456
transform 1 0 7452 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_167_81
timestamp 18001
transform 1 0 8556 0 -1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_167_87
timestamp 18001
transform 1 0 9108 0 -1 93568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_167_95
timestamp 18001
transform 1 0 9844 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_167_98
timestamp 18001
transform 1 0 10120 0 -1 93568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_167_106
timestamp 18001
transform 1 0 10856 0 -1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_167_110
timestamp 18001
transform 1 0 11224 0 -1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_167_113
timestamp 18001
transform 1 0 11500 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_119
timestamp 18001
transform 1 0 12052 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_167_122
timestamp 18001
transform 1 0 12328 0 -1 93568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_167_130
timestamp 18001
transform 1 0 13064 0 -1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_167_134
timestamp 18001
transform 1 0 13432 0 -1 93568
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_167_141
timestamp 1636986456
transform 1 0 14076 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_153
timestamp 1636986456
transform 1 0 15180 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_167_165
timestamp 18001
transform 1 0 16284 0 -1 93568
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_167_169
timestamp 1636986456
transform 1 0 16652 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_181
timestamp 1636986456
transform 1 0 17756 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_167_193
timestamp 18001
transform 1 0 18860 0 -1 93568
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_167_197
timestamp 1636986456
transform 1 0 19228 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_209
timestamp 1636986456
transform 1 0 20332 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_167_221
timestamp 18001
transform 1 0 21436 0 -1 93568
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_167_225
timestamp 1636986456
transform 1 0 21804 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_237
timestamp 1636986456
transform 1 0 22908 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_167_249
timestamp 18001
transform 1 0 24012 0 -1 93568
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_167_253
timestamp 1636986456
transform 1 0 24380 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_265
timestamp 1636986456
transform 1 0 25484 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_167_277
timestamp 18001
transform 1 0 26588 0 -1 93568
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_167_281
timestamp 1636986456
transform 1 0 26956 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_293
timestamp 1636986456
transform 1 0 28060 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_167_305
timestamp 18001
transform 1 0 29164 0 -1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_167_309
timestamp 18001
transform 1 0 29532 0 -1 93568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_167_335
timestamp 18001
transform 1 0 31924 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_339
timestamp 1636986456
transform 1 0 32292 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_351
timestamp 1636986456
transform 1 0 33396 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_167_363
timestamp 18001
transform 1 0 34500 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_365
timestamp 1636986456
transform 1 0 34684 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_377
timestamp 1636986456
transform 1 0 35788 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_167_389
timestamp 18001
transform 1 0 36892 0 -1 93568
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_167_393
timestamp 1636986456
transform 1 0 37260 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_405
timestamp 1636986456
transform 1 0 38364 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_167_417
timestamp 18001
transform 1 0 39468 0 -1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_167_421
timestamp 18001
transform 1 0 39836 0 -1 93568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_167_425
timestamp 18001
transform 1 0 40204 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_451
timestamp 1636986456
transform 1 0 42596 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_463
timestamp 1636986456
transform 1 0 43700 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_167_475
timestamp 18001
transform 1 0 44804 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_477
timestamp 1636986456
transform 1 0 44988 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_489
timestamp 1636986456
transform 1 0 46092 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_167_501
timestamp 18001
transform 1 0 47196 0 -1 93568
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_167_505
timestamp 1636986456
transform 1 0 47564 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_517
timestamp 1636986456
transform 1 0 48668 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_167_529
timestamp 18001
transform 1 0 49772 0 -1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_167_533
timestamp 18001
transform 1 0 50140 0 -1 93568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_167_545
timestamp 18001
transform 1 0 51244 0 -1 93568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_167_555
timestamp 18001
transform 1 0 52164 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_167_581
timestamp 18001
transform 1 0 54556 0 -1 93568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_167_585
timestamp 18001
transform 1 0 54924 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_167_609
timestamp 18001
transform 1 0 57132 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_615
timestamp 18001
transform 1 0 57684 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_617
timestamp 1636986456
transform 1 0 57868 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_629
timestamp 1636986456
transform 1 0 58972 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_167_641
timestamp 18001
transform 1 0 60076 0 -1 93568
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_167_645
timestamp 1636986456
transform 1 0 60444 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_657
timestamp 1636986456
transform 1 0 61548 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_167_669
timestamp 18001
transform 1 0 62652 0 -1 93568
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_167_673
timestamp 1636986456
transform 1 0 63020 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_685
timestamp 1636986456
transform 1 0 64124 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_167_697
timestamp 18001
transform 1 0 65228 0 -1 93568
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_167_701
timestamp 1636986456
transform 1 0 65596 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_713
timestamp 1636986456
transform 1 0 66700 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_167_725
timestamp 18001
transform 1 0 67804 0 -1 93568
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_167_729
timestamp 1636986456
transform 1 0 68172 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_741
timestamp 1636986456
transform 1 0 69276 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_167_753
timestamp 18001
transform 1 0 70380 0 -1 93568
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_167_757
timestamp 1636986456
transform 1 0 70748 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_769
timestamp 1636986456
transform 1 0 71852 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_167_781
timestamp 18001
transform 1 0 72956 0 -1 93568
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_167_785
timestamp 1636986456
transform 1 0 73324 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_797
timestamp 1636986456
transform 1 0 74428 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_167_809
timestamp 18001
transform 1 0 75532 0 -1 93568
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_167_813
timestamp 1636986456
transform 1 0 75900 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_825
timestamp 1636986456
transform 1 0 77004 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_167_837
timestamp 18001
transform 1 0 78108 0 -1 93568
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_167_841
timestamp 1636986456
transform 1 0 78476 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_853
timestamp 1636986456
transform 1 0 79580 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_167_865
timestamp 18001
transform 1 0 80684 0 -1 93568
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_167_869
timestamp 1636986456
transform 1 0 81052 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_881
timestamp 1636986456
transform 1 0 82156 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_167_893
timestamp 18001
transform 1 0 83260 0 -1 93568
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_167_897
timestamp 1636986456
transform 1 0 83628 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_909
timestamp 1636986456
transform 1 0 84732 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_167_921
timestamp 18001
transform 1 0 85836 0 -1 93568
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_167_925
timestamp 1636986456
transform 1 0 86204 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_937
timestamp 1636986456
transform 1 0 87308 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_167_949
timestamp 18001
transform 1 0 88412 0 -1 93568
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_167_953
timestamp 1636986456
transform 1 0 88780 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_965
timestamp 1636986456
transform 1 0 89884 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_167_977
timestamp 18001
transform 1 0 90988 0 -1 93568
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_167_981
timestamp 1636986456
transform 1 0 91356 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_993
timestamp 1636986456
transform 1 0 92460 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_167_1005
timestamp 18001
transform 1 0 93564 0 -1 93568
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_167_1009
timestamp 1636986456
transform 1 0 93932 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_1021
timestamp 1636986456
transform 1 0 95036 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_167_1033
timestamp 18001
transform 1 0 96140 0 -1 93568
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_167_1037
timestamp 1636986456
transform 1 0 96508 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_3
timestamp 1636986456
transform 1 0 1380 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_15
timestamp 1636986456
transform 1 0 2484 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_168_27
timestamp 18001
transform 1 0 3588 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_29
timestamp 1636986456
transform 1 0 3772 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_41
timestamp 1636986456
transform 1 0 4876 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_53
timestamp 1636986456
transform 1 0 5980 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_65
timestamp 1636986456
transform 1 0 7084 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_77
timestamp 18001
transform 1 0 8188 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_83
timestamp 18001
transform 1 0 8740 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_85
timestamp 1636986456
transform 1 0 8924 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_97
timestamp 1636986456
transform 1 0 10028 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_109
timestamp 1636986456
transform 1 0 11132 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_121
timestamp 1636986456
transform 1 0 12236 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_133
timestamp 18001
transform 1 0 13340 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_139
timestamp 18001
transform 1 0 13892 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_141
timestamp 1636986456
transform 1 0 14076 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_153
timestamp 1636986456
transform 1 0 15180 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_165
timestamp 1636986456
transform 1 0 16284 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_177
timestamp 1636986456
transform 1 0 17388 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_189
timestamp 18001
transform 1 0 18492 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_195
timestamp 18001
transform 1 0 19044 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_197
timestamp 1636986456
transform 1 0 19228 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_209
timestamp 1636986456
transform 1 0 20332 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_221
timestamp 1636986456
transform 1 0 21436 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_233
timestamp 1636986456
transform 1 0 22540 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_245
timestamp 18001
transform 1 0 23644 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_251
timestamp 18001
transform 1 0 24196 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_253
timestamp 1636986456
transform 1 0 24380 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_265
timestamp 1636986456
transform 1 0 25484 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_277
timestamp 1636986456
transform 1 0 26588 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_289
timestamp 1636986456
transform 1 0 27692 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_301
timestamp 18001
transform 1 0 28796 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_307
timestamp 18001
transform 1 0 29348 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_309
timestamp 1636986456
transform 1 0 29532 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_321
timestamp 1636986456
transform 1 0 30636 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_333
timestamp 1636986456
transform 1 0 31740 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_345
timestamp 1636986456
transform 1 0 32844 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_357
timestamp 18001
transform 1 0 33948 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_363
timestamp 18001
transform 1 0 34500 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_365
timestamp 1636986456
transform 1 0 34684 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_377
timestamp 1636986456
transform 1 0 35788 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_389
timestamp 1636986456
transform 1 0 36892 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_401
timestamp 1636986456
transform 1 0 37996 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_413
timestamp 18001
transform 1 0 39100 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_419
timestamp 18001
transform 1 0 39652 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_421
timestamp 1636986456
transform 1 0 39836 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_433
timestamp 1636986456
transform 1 0 40940 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_445
timestamp 1636986456
transform 1 0 42044 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_457
timestamp 1636986456
transform 1 0 43148 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_469
timestamp 18001
transform 1 0 44252 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_475
timestamp 18001
transform 1 0 44804 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_477
timestamp 1636986456
transform 1 0 44988 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_489
timestamp 1636986456
transform 1 0 46092 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_501
timestamp 1636986456
transform 1 0 47196 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_513
timestamp 1636986456
transform 1 0 48300 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_525
timestamp 18001
transform 1 0 49404 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_531
timestamp 18001
transform 1 0 49956 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_533
timestamp 1636986456
transform 1 0 50140 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_545
timestamp 1636986456
transform 1 0 51244 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_168_557
timestamp 18001
transform 1 0 52348 0 1 93568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_168_585
timestamp 18001
transform 1 0 54924 0 1 93568
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_168_589
timestamp 1636986456
transform 1 0 55292 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_601
timestamp 1636986456
transform 1 0 56396 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_613
timestamp 1636986456
transform 1 0 57500 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_625
timestamp 1636986456
transform 1 0 58604 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_637
timestamp 18001
transform 1 0 59708 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_643
timestamp 18001
transform 1 0 60260 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_645
timestamp 1636986456
transform 1 0 60444 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_657
timestamp 1636986456
transform 1 0 61548 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_669
timestamp 1636986456
transform 1 0 62652 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_681
timestamp 1636986456
transform 1 0 63756 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_693
timestamp 18001
transform 1 0 64860 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_699
timestamp 18001
transform 1 0 65412 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_701
timestamp 1636986456
transform 1 0 65596 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_713
timestamp 1636986456
transform 1 0 66700 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_725
timestamp 1636986456
transform 1 0 67804 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_737
timestamp 1636986456
transform 1 0 68908 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_749
timestamp 18001
transform 1 0 70012 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_755
timestamp 18001
transform 1 0 70564 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_757
timestamp 1636986456
transform 1 0 70748 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_769
timestamp 1636986456
transform 1 0 71852 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_781
timestamp 1636986456
transform 1 0 72956 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_793
timestamp 1636986456
transform 1 0 74060 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_805
timestamp 18001
transform 1 0 75164 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_811
timestamp 18001
transform 1 0 75716 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_813
timestamp 1636986456
transform 1 0 75900 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_825
timestamp 1636986456
transform 1 0 77004 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_837
timestamp 1636986456
transform 1 0 78108 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_849
timestamp 1636986456
transform 1 0 79212 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_861
timestamp 18001
transform 1 0 80316 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_867
timestamp 18001
transform 1 0 80868 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_869
timestamp 1636986456
transform 1 0 81052 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_881
timestamp 1636986456
transform 1 0 82156 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_893
timestamp 1636986456
transform 1 0 83260 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_905
timestamp 1636986456
transform 1 0 84364 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_917
timestamp 18001
transform 1 0 85468 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_923
timestamp 18001
transform 1 0 86020 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_925
timestamp 1636986456
transform 1 0 86204 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_937
timestamp 1636986456
transform 1 0 87308 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_949
timestamp 1636986456
transform 1 0 88412 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_961
timestamp 1636986456
transform 1 0 89516 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_973
timestamp 18001
transform 1 0 90620 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_979
timestamp 18001
transform 1 0 91172 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_981
timestamp 1636986456
transform 1 0 91356 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_993
timestamp 1636986456
transform 1 0 92460 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_1005
timestamp 1636986456
transform 1 0 93564 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_1017
timestamp 1636986456
transform 1 0 94668 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_1029
timestamp 18001
transform 1 0 95772 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_1035
timestamp 18001
transform 1 0 96324 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_1037
timestamp 1636986456
transform 1 0 96508 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_3
timestamp 1636986456
transform 1 0 1380 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_15
timestamp 1636986456
transform 1 0 2484 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_27
timestamp 1636986456
transform 1 0 3588 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_39
timestamp 1636986456
transform 1 0 4692 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_169_51
timestamp 18001
transform 1 0 5796 0 -1 94656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_169_55
timestamp 18001
transform 1 0 6164 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_57
timestamp 1636986456
transform 1 0 6348 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_69
timestamp 1636986456
transform 1 0 7452 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_81
timestamp 1636986456
transform 1 0 8556 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_93
timestamp 1636986456
transform 1 0 9660 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_105
timestamp 18001
transform 1 0 10764 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_111
timestamp 18001
transform 1 0 11316 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_113
timestamp 1636986456
transform 1 0 11500 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_125
timestamp 1636986456
transform 1 0 12604 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_137
timestamp 1636986456
transform 1 0 13708 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_149
timestamp 1636986456
transform 1 0 14812 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_161
timestamp 18001
transform 1 0 15916 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_167
timestamp 18001
transform 1 0 16468 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_169
timestamp 1636986456
transform 1 0 16652 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_181
timestamp 1636986456
transform 1 0 17756 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_193
timestamp 1636986456
transform 1 0 18860 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_205
timestamp 1636986456
transform 1 0 19964 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_217
timestamp 18001
transform 1 0 21068 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_223
timestamp 18001
transform 1 0 21620 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_225
timestamp 1636986456
transform 1 0 21804 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_237
timestamp 1636986456
transform 1 0 22908 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_249
timestamp 1636986456
transform 1 0 24012 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_261
timestamp 1636986456
transform 1 0 25116 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_273
timestamp 18001
transform 1 0 26220 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_279
timestamp 18001
transform 1 0 26772 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_281
timestamp 1636986456
transform 1 0 26956 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_293
timestamp 1636986456
transform 1 0 28060 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_305
timestamp 1636986456
transform 1 0 29164 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_317
timestamp 1636986456
transform 1 0 30268 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_329
timestamp 18001
transform 1 0 31372 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_335
timestamp 18001
transform 1 0 31924 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_337
timestamp 1636986456
transform 1 0 32108 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_349
timestamp 1636986456
transform 1 0 33212 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_361
timestamp 1636986456
transform 1 0 34316 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_373
timestamp 1636986456
transform 1 0 35420 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_385
timestamp 18001
transform 1 0 36524 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_391
timestamp 18001
transform 1 0 37076 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_393
timestamp 1636986456
transform 1 0 37260 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_405
timestamp 1636986456
transform 1 0 38364 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_417
timestamp 1636986456
transform 1 0 39468 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_429
timestamp 1636986456
transform 1 0 40572 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_441
timestamp 18001
transform 1 0 41676 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_447
timestamp 18001
transform 1 0 42228 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_449
timestamp 1636986456
transform 1 0 42412 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_461
timestamp 1636986456
transform 1 0 43516 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_473
timestamp 1636986456
transform 1 0 44620 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_485
timestamp 1636986456
transform 1 0 45724 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_497
timestamp 18001
transform 1 0 46828 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_503
timestamp 18001
transform 1 0 47380 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_505
timestamp 1636986456
transform 1 0 47564 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_517
timestamp 1636986456
transform 1 0 48668 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_529
timestamp 1636986456
transform 1 0 49772 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_541
timestamp 1636986456
transform 1 0 50876 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_553
timestamp 18001
transform 1 0 51980 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_559
timestamp 18001
transform 1 0 52532 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_561
timestamp 1636986456
transform 1 0 52716 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_573
timestamp 1636986456
transform 1 0 53820 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_585
timestamp 1636986456
transform 1 0 54924 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_597
timestamp 1636986456
transform 1 0 56028 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_609
timestamp 18001
transform 1 0 57132 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_615
timestamp 18001
transform 1 0 57684 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_617
timestamp 1636986456
transform 1 0 57868 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_629
timestamp 1636986456
transform 1 0 58972 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_641
timestamp 1636986456
transform 1 0 60076 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_653
timestamp 1636986456
transform 1 0 61180 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_665
timestamp 18001
transform 1 0 62284 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_671
timestamp 18001
transform 1 0 62836 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_673
timestamp 1636986456
transform 1 0 63020 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_685
timestamp 1636986456
transform 1 0 64124 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_697
timestamp 1636986456
transform 1 0 65228 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_709
timestamp 1636986456
transform 1 0 66332 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_721
timestamp 18001
transform 1 0 67436 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_727
timestamp 18001
transform 1 0 67988 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_729
timestamp 1636986456
transform 1 0 68172 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_741
timestamp 1636986456
transform 1 0 69276 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_753
timestamp 1636986456
transform 1 0 70380 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_765
timestamp 1636986456
transform 1 0 71484 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_777
timestamp 18001
transform 1 0 72588 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_783
timestamp 18001
transform 1 0 73140 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_785
timestamp 1636986456
transform 1 0 73324 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_797
timestamp 1636986456
transform 1 0 74428 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_809
timestamp 1636986456
transform 1 0 75532 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_821
timestamp 1636986456
transform 1 0 76636 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_833
timestamp 18001
transform 1 0 77740 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_839
timestamp 18001
transform 1 0 78292 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_841
timestamp 1636986456
transform 1 0 78476 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_853
timestamp 1636986456
transform 1 0 79580 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_865
timestamp 1636986456
transform 1 0 80684 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_877
timestamp 1636986456
transform 1 0 81788 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_889
timestamp 18001
transform 1 0 82892 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_895
timestamp 18001
transform 1 0 83444 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_897
timestamp 1636986456
transform 1 0 83628 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_909
timestamp 1636986456
transform 1 0 84732 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_921
timestamp 1636986456
transform 1 0 85836 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_933
timestamp 1636986456
transform 1 0 86940 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_945
timestamp 18001
transform 1 0 88044 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_951
timestamp 18001
transform 1 0 88596 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_953
timestamp 1636986456
transform 1 0 88780 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_965
timestamp 1636986456
transform 1 0 89884 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_977
timestamp 1636986456
transform 1 0 90988 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_989
timestamp 1636986456
transform 1 0 92092 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_1001
timestamp 18001
transform 1 0 93196 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_1007
timestamp 18001
transform 1 0 93748 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_1009
timestamp 1636986456
transform 1 0 93932 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_1021
timestamp 1636986456
transform 1 0 95036 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_1033
timestamp 1636986456
transform 1 0 96140 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_169_1045
timestamp 18001
transform 1 0 97244 0 -1 94656
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_170_3
timestamp 1636986456
transform 1 0 1380 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_15
timestamp 1636986456
transform 1 0 2484 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_170_27
timestamp 18001
transform 1 0 3588 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_29
timestamp 1636986456
transform 1 0 3772 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_41
timestamp 1636986456
transform 1 0 4876 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_53
timestamp 1636986456
transform 1 0 5980 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_65
timestamp 1636986456
transform 1 0 7084 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_77
timestamp 18001
transform 1 0 8188 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_83
timestamp 18001
transform 1 0 8740 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_85
timestamp 1636986456
transform 1 0 8924 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_97
timestamp 1636986456
transform 1 0 10028 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_109
timestamp 1636986456
transform 1 0 11132 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_121
timestamp 1636986456
transform 1 0 12236 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_133
timestamp 18001
transform 1 0 13340 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_139
timestamp 18001
transform 1 0 13892 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_141
timestamp 1636986456
transform 1 0 14076 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_153
timestamp 1636986456
transform 1 0 15180 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_165
timestamp 1636986456
transform 1 0 16284 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_177
timestamp 1636986456
transform 1 0 17388 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_189
timestamp 18001
transform 1 0 18492 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_195
timestamp 18001
transform 1 0 19044 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_197
timestamp 1636986456
transform 1 0 19228 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_209
timestamp 1636986456
transform 1 0 20332 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_221
timestamp 1636986456
transform 1 0 21436 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_233
timestamp 1636986456
transform 1 0 22540 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_245
timestamp 18001
transform 1 0 23644 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_251
timestamp 18001
transform 1 0 24196 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_265
timestamp 1636986456
transform 1 0 25484 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_277
timestamp 1636986456
transform 1 0 26588 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_289
timestamp 1636986456
transform 1 0 27692 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_301
timestamp 18001
transform 1 0 28796 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_307
timestamp 18001
transform 1 0 29348 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_309
timestamp 1636986456
transform 1 0 29532 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_321
timestamp 1636986456
transform 1 0 30636 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_333
timestamp 1636986456
transform 1 0 31740 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_345
timestamp 1636986456
transform 1 0 32844 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_357
timestamp 18001
transform 1 0 33948 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_363
timestamp 18001
transform 1 0 34500 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_365
timestamp 1636986456
transform 1 0 34684 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_377
timestamp 1636986456
transform 1 0 35788 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_389
timestamp 1636986456
transform 1 0 36892 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_401
timestamp 1636986456
transform 1 0 37996 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_413
timestamp 18001
transform 1 0 39100 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_419
timestamp 18001
transform 1 0 39652 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_421
timestamp 1636986456
transform 1 0 39836 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_433
timestamp 1636986456
transform 1 0 40940 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_445
timestamp 1636986456
transform 1 0 42044 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_457
timestamp 1636986456
transform 1 0 43148 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_469
timestamp 18001
transform 1 0 44252 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_475
timestamp 18001
transform 1 0 44804 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_477
timestamp 1636986456
transform 1 0 44988 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_489
timestamp 1636986456
transform 1 0 46092 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_501
timestamp 1636986456
transform 1 0 47196 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_513
timestamp 1636986456
transform 1 0 48300 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_525
timestamp 18001
transform 1 0 49404 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_531
timestamp 18001
transform 1 0 49956 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_170_533
timestamp 18001
transform 1 0 50140 0 1 94656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_170_541
timestamp 18001
transform 1 0 50876 0 1 94656
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_170_546
timestamp 1636986456
transform 1 0 51336 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_170_558
timestamp 18001
transform 1 0 52440 0 1 94656
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_170_565
timestamp 1636986456
transform 1 0 53084 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_170_577
timestamp 18001
transform 1 0 54188 0 1 94656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_170_585
timestamp 18001
transform 1 0 54924 0 1 94656
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_170_589
timestamp 1636986456
transform 1 0 55292 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_170_601
timestamp 18001
transform 1 0 56396 0 1 94656
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_170_607
timestamp 1636986456
transform 1 0 56948 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_619
timestamp 1636986456
transform 1 0 58052 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_631
timestamp 1636986456
transform 1 0 59156 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_170_643
timestamp 18001
transform 1 0 60260 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_645
timestamp 1636986456
transform 1 0 60444 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_657
timestamp 1636986456
transform 1 0 61548 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_669
timestamp 1636986456
transform 1 0 62652 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_681
timestamp 1636986456
transform 1 0 63756 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_693
timestamp 18001
transform 1 0 64860 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_699
timestamp 18001
transform 1 0 65412 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_701
timestamp 1636986456
transform 1 0 65596 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_713
timestamp 1636986456
transform 1 0 66700 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_725
timestamp 1636986456
transform 1 0 67804 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_737
timestamp 1636986456
transform 1 0 68908 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_749
timestamp 18001
transform 1 0 70012 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_755
timestamp 18001
transform 1 0 70564 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_757
timestamp 1636986456
transform 1 0 70748 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_769
timestamp 1636986456
transform 1 0 71852 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_781
timestamp 1636986456
transform 1 0 72956 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_793
timestamp 1636986456
transform 1 0 74060 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_805
timestamp 18001
transform 1 0 75164 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_811
timestamp 18001
transform 1 0 75716 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_813
timestamp 1636986456
transform 1 0 75900 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_825
timestamp 1636986456
transform 1 0 77004 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_837
timestamp 1636986456
transform 1 0 78108 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_849
timestamp 1636986456
transform 1 0 79212 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_861
timestamp 18001
transform 1 0 80316 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_867
timestamp 18001
transform 1 0 80868 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_869
timestamp 1636986456
transform 1 0 81052 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_881
timestamp 1636986456
transform 1 0 82156 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_893
timestamp 1636986456
transform 1 0 83260 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_905
timestamp 1636986456
transform 1 0 84364 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_917
timestamp 18001
transform 1 0 85468 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_923
timestamp 18001
transform 1 0 86020 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_925
timestamp 1636986456
transform 1 0 86204 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_937
timestamp 1636986456
transform 1 0 87308 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_949
timestamp 1636986456
transform 1 0 88412 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_961
timestamp 1636986456
transform 1 0 89516 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_973
timestamp 18001
transform 1 0 90620 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_979
timestamp 18001
transform 1 0 91172 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_981
timestamp 1636986456
transform 1 0 91356 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_993
timestamp 1636986456
transform 1 0 92460 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_1005
timestamp 1636986456
transform 1 0 93564 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_1017
timestamp 1636986456
transform 1 0 94668 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_1029
timestamp 18001
transform 1 0 95772 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_1035
timestamp 18001
transform 1 0 96324 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_1037
timestamp 1636986456
transform 1 0 96508 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_3
timestamp 1636986456
transform 1 0 1380 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_15
timestamp 1636986456
transform 1 0 2484 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_171_27
timestamp 18001
transform 1 0 3588 0 -1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_171_29
timestamp 1636986456
transform 1 0 3772 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_41
timestamp 1636986456
transform 1 0 4876 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_171_53
timestamp 18001
transform 1 0 5980 0 -1 95744
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_171_57
timestamp 1636986456
transform 1 0 6348 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_69
timestamp 1636986456
transform 1 0 7452 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_171_81
timestamp 18001
transform 1 0 8556 0 -1 95744
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_171_85
timestamp 1636986456
transform 1 0 8924 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_97
timestamp 1636986456
transform 1 0 10028 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_171_109
timestamp 18001
transform 1 0 11132 0 -1 95744
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_171_113
timestamp 1636986456
transform 1 0 11500 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_125
timestamp 1636986456
transform 1 0 12604 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_171_137
timestamp 18001
transform 1 0 13708 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_171_147
timestamp 18001
transform 1 0 14628 0 -1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_171_161
timestamp 18001
transform 1 0 15916 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_167
timestamp 18001
transform 1 0 16468 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_171_175
timestamp 18001
transform 1 0 17204 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_171_182
timestamp 18001
transform 1 0 17848 0 -1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_171_197
timestamp 18001
transform 1 0 19228 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_203
timestamp 18001
transform 1 0 19780 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_171_210
timestamp 18001
transform 1 0 20424 0 -1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_171_230
timestamp 18001
transform 1 0 22264 0 -1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_171_238
timestamp 18001
transform 1 0 23000 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_171_245
timestamp 18001
transform 1 0 23644 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_251
timestamp 18001
transform 1 0 24196 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_171_253
timestamp 18001
transform 1 0 24380 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_259
timestamp 18001
transform 1 0 24932 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_171_272
timestamp 18001
transform 1 0 26128 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_171_279
timestamp 18001
transform 1 0 26772 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_171_281
timestamp 18001
transform 1 0 26956 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_287
timestamp 18001
transform 1 0 27508 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_171_293
timestamp 18001
transform 1 0 28060 0 -1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_171_301
timestamp 18001
transform 1 0 28796 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_171_307
timestamp 18001
transform 1 0 29348 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_171_314
timestamp 18001
transform 1 0 29992 0 -1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_171_322
timestamp 18001
transform 1 0 30728 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_171_328
timestamp 18001
transform 1 0 31280 0 -1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_171_337
timestamp 18001
transform 1 0 32108 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_171_343
timestamp 18001
transform 1 0 32660 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_171_350
timestamp 18001
transform 1 0 33304 0 -1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_171_358
timestamp 18001
transform 1 0 34040 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_171_365
timestamp 18001
transform 1 0 34684 0 -1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_171_373
timestamp 18001
transform 1 0 35420 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_171_378
timestamp 18001
transform 1 0 35880 0 -1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_171_386
timestamp 18001
transform 1 0 36616 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_171_393
timestamp 18001
transform 1 0 37260 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_171_399
timestamp 18001
transform 1 0 37812 0 -1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_171_407
timestamp 18001
transform 1 0 38548 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_171_413
timestamp 18001
transform 1 0 39100 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_419
timestamp 18001
transform 1 0 39652 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_171_421
timestamp 18001
transform 1 0 39836 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_171_427
timestamp 18001
transform 1 0 40388 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_171_434
timestamp 18001
transform 1 0 41032 0 -1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_171_442
timestamp 18001
transform 1 0 41768 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_171_449
timestamp 18001
transform 1 0 42412 0 -1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_171_457
timestamp 18001
transform 1 0 43148 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_171_462
timestamp 18001
transform 1 0 43608 0 -1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_171_470
timestamp 18001
transform 1 0 44344 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_171_477
timestamp 18001
transform 1 0 44988 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_171_483
timestamp 18001
transform 1 0 45540 0 -1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_171_491
timestamp 18001
transform 1 0 46276 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_171_497
timestamp 18001
transform 1 0 46828 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_503
timestamp 18001
transform 1 0 47380 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_171_505
timestamp 18001
transform 1 0 47564 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_171_511
timestamp 18001
transform 1 0 48116 0 -1 95744
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_171_518
timestamp 1636986456
transform 1 0 48760 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_171_530
timestamp 18001
transform 1 0 49864 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_171_533
timestamp 18001
transform 1 0 50140 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_539
timestamp 18001
transform 1 0 50692 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_171_581
timestamp 18001
transform 1 0 54556 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_171_585
timestamp 18001
transform 1 0 54924 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_171_611
timestamp 18001
transform 1 0 57316 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_171_619
timestamp 18001
transform 1 0 58052 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_171_623
timestamp 18001
transform 1 0 58420 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_171_630
timestamp 18001
transform 1 0 59064 0 -1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_171_651
timestamp 18001
transform 1 0 60996 0 -1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_171_665
timestamp 18001
transform 1 0 62284 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_671
timestamp 18001
transform 1 0 62836 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_171_679
timestamp 18001
transform 1 0 63572 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_171_685
timestamp 18001
transform 1 0 64124 0 -1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_171_693
timestamp 18001
transform 1 0 64860 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_171_701
timestamp 18001
transform 1 0 65596 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_707
timestamp 18001
transform 1 0 66148 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_171_720
timestamp 18001
transform 1 0 67344 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_744
timestamp 18001
transform 1 0 69552 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_171_750
timestamp 18001
transform 1 0 70104 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_171_762
timestamp 18001
transform 1 0 71208 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_171_769
timestamp 18001
transform 1 0 71852 0 -1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_171_777
timestamp 18001
transform 1 0 72588 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_171_783
timestamp 18001
transform 1 0 73140 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_171_785
timestamp 18001
transform 1 0 73324 0 -1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_171_793
timestamp 18001
transform 1 0 74060 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_171_798
timestamp 18001
transform 1 0 74520 0 -1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_171_806
timestamp 18001
transform 1 0 75256 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_171_813
timestamp 18001
transform 1 0 75900 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_171_819
timestamp 18001
transform 1 0 76452 0 -1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_171_827
timestamp 18001
transform 1 0 77188 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_171_833
timestamp 18001
transform 1 0 77740 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_839
timestamp 18001
transform 1 0 78292 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_171_841
timestamp 18001
transform 1 0 78476 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_171_847
timestamp 18001
transform 1 0 79028 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_171_854
timestamp 18001
transform 1 0 79672 0 -1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_171_862
timestamp 18001
transform 1 0 80408 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_171_869
timestamp 18001
transform 1 0 81052 0 -1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_171_877
timestamp 18001
transform 1 0 81788 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_171_882
timestamp 18001
transform 1 0 82248 0 -1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_171_890
timestamp 18001
transform 1 0 82984 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_171_897
timestamp 18001
transform 1 0 83628 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_171_903
timestamp 18001
transform 1 0 84180 0 -1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_171_911
timestamp 18001
transform 1 0 84916 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_171_917
timestamp 18001
transform 1 0 85468 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_923
timestamp 18001
transform 1 0 86020 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_171_925
timestamp 18001
transform 1 0 86204 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_171_931
timestamp 18001
transform 1 0 86756 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_171_938
timestamp 18001
transform 1 0 87400 0 -1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_171_946
timestamp 18001
transform 1 0 88136 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_171_953
timestamp 18001
transform 1 0 88780 0 -1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_171_961
timestamp 18001
transform 1 0 89516 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_171_966
timestamp 18001
transform 1 0 89976 0 -1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_171_974
timestamp 18001
transform 1 0 90712 0 -1 95744
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_171_981
timestamp 1636986456
transform 1 0 91356 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_993
timestamp 1636986456
transform 1 0 92460 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_171_1005
timestamp 18001
transform 1 0 93564 0 -1 95744
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_171_1009
timestamp 1636986456
transform 1 0 93932 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_1021
timestamp 1636986456
transform 1 0 95036 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_171_1033
timestamp 18001
transform 1 0 96140 0 -1 95744
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_171_1037
timestamp 1636986456
transform 1 0 96508 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  input1
timestamp 18001
transform 1 0 1380 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_12  input2
timestamp 18001
transform 1 0 55292 0 -1 95744
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  input3
timestamp 18001
transform -1 0 52624 0 -1 95744
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 18001
transform -1 0 97612 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 18001
transform -1 0 97612 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 18001
transform -1 0 97612 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 18001
transform -1 0 97612 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 18001
transform -1 0 97612 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 18001
transform -1 0 97612 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 18001
transform -1 0 97612 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input11
timestamp 18001
transform -1 0 97612 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input12
timestamp 18001
transform -1 0 97612 0 -1 72896
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 18001
transform -1 0 97612 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 18001
transform -1 0 97612 0 1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 18001
transform -1 0 97612 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 18001
transform -1 0 97612 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 18001
transform -1 0 97612 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input18
timestamp 18001
transform -1 0 97612 0 -1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 18001
transform -1 0 97612 0 -1 79424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input20
timestamp 18001
transform -1 0 97612 0 1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input21
timestamp 18001
transform -1 0 97612 0 -1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 18001
transform -1 0 97612 0 1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input23
timestamp 18001
transform -1 0 97612 0 -1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input24
timestamp 18001
transform -1 0 97612 0 -1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input25
timestamp 18001
transform -1 0 97612 0 1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input26
timestamp 18001
transform -1 0 97612 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input27
timestamp 18001
transform -1 0 97612 0 -1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input28
timestamp 18001
transform -1 0 97612 0 1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp 18001
transform -1 0 97612 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input30
timestamp 18001
transform -1 0 97612 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input31
timestamp 18001
transform -1 0 97612 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input32
timestamp 18001
transform -1 0 97612 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input33
timestamp 18001
transform -1 0 97612 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input34
timestamp 18001
transform -1 0 97612 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input35
timestamp 18001
transform -1 0 97612 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input36
timestamp 18001
transform 1 0 14260 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input37
timestamp 18001
transform 1 0 25208 0 -1 95744
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input38
timestamp 18001
transform -1 0 26772 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input39
timestamp 18001
transform -1 0 28060 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input40
timestamp 18001
transform -1 0 29348 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input41
timestamp 18001
transform 1 0 29716 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input42
timestamp 18001
transform -1 0 31280 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input43
timestamp 18001
transform -1 0 57132 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input44
timestamp 18001
transform -1 0 57776 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input45
timestamp 18001
transform 1 0 58696 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input46
timestamp 18001
transform -1 0 60352 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input47
timestamp 18001
transform 1 0 15548 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input48
timestamp 18001
transform 1 0 60628 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input49
timestamp 18001
transform -1 0 62284 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 18001
transform -1 0 63572 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input51
timestamp 18001
transform 1 0 63848 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input52
timestamp 18001
transform -1 0 65504 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input53
timestamp 18001
transform 1 0 66424 0 -1 95744
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input54
timestamp 18001
transform 1 0 68172 0 -1 95744
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input55
timestamp 18001
transform -1 0 69368 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input56
timestamp 18001
transform -1 0 69920 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input57
timestamp 18001
transform -1 0 71208 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input58
timestamp 18001
transform 1 0 16836 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input59
timestamp 18001
transform 1 0 71576 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input60
timestamp 18001
transform 1 0 72864 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input61
timestamp 18001
transform 1 0 17480 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input62
timestamp 18001
transform -1 0 19136 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input63
timestamp 18001
transform -1 0 20424 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input64
timestamp 18001
transform -1 0 21712 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input65
timestamp 18001
transform 1 0 21988 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input66
timestamp 18001
transform -1 0 23644 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input67
timestamp 18001
transform 1 0 24564 0 1 94656
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input68
timestamp 18001
transform -1 0 32568 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input69
timestamp 18001
transform -1 0 43516 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input70
timestamp 18001
transform -1 0 44896 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input71
timestamp 18001
transform 1 0 45172 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input72
timestamp 18001
transform 1 0 46460 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input73
timestamp 18001
transform 1 0 47748 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input74
timestamp 18001
transform -1 0 49036 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input75
timestamp 18001
transform -1 0 74428 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input76
timestamp 18001
transform -1 0 75716 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input77
timestamp 18001
transform -1 0 76360 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input78
timestamp 18001
transform 1 0 77372 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input79
timestamp 18001
transform 1 0 32936 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input80
timestamp 18001
transform -1 0 78936 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input81
timestamp 18001
transform 1 0 79304 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input82
timestamp 18001
transform 1 0 80592 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input83
timestamp 18001
transform -1 0 82156 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input84
timestamp 18001
transform -1 0 83444 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input85
timestamp 18001
transform 1 0 83812 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input86
timestamp 18001
transform -1 0 85376 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input87
timestamp 18001
transform -1 0 86756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input88
timestamp 18001
transform 1 0 87032 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input89
timestamp 18001
transform 1 0 88780 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input90
timestamp 18001
transform 1 0 34224 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input91
timestamp 18001
transform 1 0 89700 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input92
timestamp 18001
transform -1 0 97612 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input93
timestamp 18001
transform 1 0 35512 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input94
timestamp 18001
transform -1 0 37076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input95
timestamp 18001
transform -1 0 37720 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input96
timestamp 18001
transform -1 0 39008 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input97
timestamp 18001
transform -1 0 40296 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input98
timestamp 18001
transform 1 0 40664 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input99
timestamp 18001
transform -1 0 42228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input100
timestamp 18001
transform 1 0 1380 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input101
timestamp 18001
transform 1 0 1380 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input102
timestamp 18001
transform 1 0 1380 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input103
timestamp 18001
transform 1 0 1380 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input104
timestamp 18001
transform 1 0 1380 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input105
timestamp 18001
transform 1 0 1380 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input106
timestamp 18001
transform 1 0 1380 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input107
timestamp 18001
transform 1 0 1380 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input108
timestamp 18001
transform 1 0 1380 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input109
timestamp 18001
transform 1 0 1380 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input110
timestamp 18001
transform 1 0 1380 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input111
timestamp 18001
transform 1 0 1380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input112
timestamp 18001
transform 1 0 1380 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input113
timestamp 18001
transform 1 0 1380 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input114
timestamp 18001
transform 1 0 1380 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input115
timestamp 18001
transform 1 0 1380 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input116
timestamp 18001
transform 1 0 1380 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input117
timestamp 18001
transform 1 0 1380 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input118
timestamp 18001
transform 1 0 1380 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input119
timestamp 18001
transform 1 0 1380 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input120
timestamp 18001
transform 1 0 1380 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input121
timestamp 18001
transform 1 0 1380 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input122
timestamp 18001
transform 1 0 1380 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input123
timestamp 18001
transform 1 0 1380 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input124
timestamp 18001
transform 1 0 1380 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input125
timestamp 18001
transform 1 0 1380 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input126
timestamp 18001
transform 1 0 1380 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input127
timestamp 18001
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input128
timestamp 18001
transform 1 0 1380 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input129
timestamp 18001
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input130
timestamp 18001
transform 1 0 1380 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input131
timestamp 18001
transform 1 0 1380 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_12  input132
timestamp 18001
transform -1 0 11408 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  input133
timestamp 18001
transform 1 0 11684 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  input134
timestamp 18001
transform 1 0 12328 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  input135
timestamp 18001
transform 1 0 52900 0 -1 95744
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  max_cap265
timestamp 18001
transform 1 0 52716 0 -1 93568
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  max_cap266
timestamp 18001
transform -1 0 56764 0 -1 93568
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  max_cap267
timestamp 18001
transform 1 0 53084 0 1 93568
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  output136
timestamp 18001
transform -1 0 51152 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output137
timestamp 18001
transform 1 0 97244 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output138
timestamp 18001
transform 1 0 97244 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp 18001
transform 1 0 97244 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output140
timestamp 18001
transform 1 0 97244 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output141
timestamp 18001
transform 1 0 97244 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output142
timestamp 18001
transform 1 0 97244 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output143
timestamp 18001
transform 1 0 97244 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output144
timestamp 18001
transform 1 0 97244 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output145
timestamp 18001
transform 1 0 97244 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output146
timestamp 18001
transform 1 0 97244 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output147
timestamp 18001
transform 1 0 97244 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output148
timestamp 18001
transform 1 0 97244 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output149
timestamp 18001
transform 1 0 97244 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output150
timestamp 18001
transform 1 0 97244 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output151
timestamp 18001
transform 1 0 97244 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output152
timestamp 18001
transform 1 0 97244 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output153
timestamp 18001
transform 1 0 97244 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output154
timestamp 18001
transform 1 0 97244 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output155
timestamp 18001
transform 1 0 97244 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output156
timestamp 18001
transform 1 0 97244 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output157
timestamp 18001
transform 1 0 97244 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output158
timestamp 18001
transform 1 0 97244 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output159
timestamp 18001
transform 1 0 97244 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output160
timestamp 18001
transform 1 0 97244 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output161
timestamp 18001
transform 1 0 97244 0 -1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output162
timestamp 18001
transform 1 0 97244 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output163
timestamp 18001
transform 1 0 97244 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output164
timestamp 18001
transform 1 0 97244 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output165
timestamp 18001
transform 1 0 97244 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output166
timestamp 18001
transform 1 0 97244 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output167
timestamp 18001
transform 1 0 97244 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output168
timestamp 18001
transform 1 0 97244 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output169
timestamp 18001
transform 1 0 32292 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output170
timestamp 18001
transform 1 0 43240 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output171
timestamp 18001
transform 1 0 44528 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output172
timestamp 18001
transform -1 0 45540 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output173
timestamp 18001
transform 1 0 46460 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output174
timestamp 18001
transform 1 0 47748 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output175
timestamp 18001
transform -1 0 48760 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output176
timestamp 18001
transform 1 0 74152 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output177
timestamp 18001
transform 1 0 75440 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output178
timestamp 18001
transform -1 0 76452 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output179
timestamp 18001
transform 1 0 77372 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output180
timestamp 18001
transform -1 0 33304 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output181
timestamp 18001
transform 1 0 78660 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output182
timestamp 18001
transform -1 0 79672 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output183
timestamp 18001
transform 1 0 80592 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output184
timestamp 18001
transform 1 0 81880 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output185
timestamp 18001
transform 1 0 83168 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output186
timestamp 18001
transform -1 0 84180 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output187
timestamp 18001
transform 1 0 85100 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output188
timestamp 18001
transform 1 0 86388 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output189
timestamp 18001
transform -1 0 87400 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output190
timestamp 18001
transform 1 0 88320 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output191
timestamp 18001
transform 1 0 34224 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output192
timestamp 18001
transform 1 0 89608 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output193
timestamp 18001
transform 1 0 90896 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output194
timestamp 18001
transform 1 0 35512 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output195
timestamp 18001
transform 1 0 36800 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output196
timestamp 18001
transform -1 0 37812 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output197
timestamp 18001
transform 1 0 38732 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output198
timestamp 18001
transform 1 0 40020 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output199
timestamp 18001
transform -1 0 41032 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output200
timestamp 18001
transform 1 0 41952 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output201
timestamp 18001
transform -1 0 14628 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output202
timestamp 18001
transform -1 0 25576 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output203
timestamp 18001
transform 1 0 26496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output204
timestamp 18001
transform 1 0 27784 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output205
timestamp 18001
transform 1 0 29072 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output206
timestamp 18001
transform -1 0 30084 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output207
timestamp 18001
transform 1 0 31004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output208
timestamp 18001
transform -1 0 56488 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output209
timestamp 18001
transform 1 0 57408 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output210
timestamp 18001
transform 1 0 58696 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output211
timestamp 18001
transform 1 0 59984 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output212
timestamp 18001
transform 1 0 15548 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output213
timestamp 18001
transform -1 0 60996 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output214
timestamp 18001
transform 1 0 61916 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output215
timestamp 18001
transform 1 0 63204 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output216
timestamp 18001
transform -1 0 64216 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output217
timestamp 18001
transform 1 0 65136 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output218
timestamp 18001
transform 1 0 66424 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output219
timestamp 18001
transform 1 0 67712 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output220
timestamp 18001
transform -1 0 68724 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output221
timestamp 18001
transform 1 0 69644 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output222
timestamp 18001
transform 1 0 70932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output223
timestamp 18001
transform 1 0 16836 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output224
timestamp 18001
transform -1 0 71944 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output225
timestamp 18001
transform 1 0 72864 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output226
timestamp 18001
transform -1 0 17848 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output227
timestamp 18001
transform 1 0 18768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output228
timestamp 18001
transform 1 0 20056 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output229
timestamp 18001
transform 1 0 21344 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output230
timestamp 18001
transform -1 0 22356 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output231
timestamp 18001
transform 1 0 23276 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output232
timestamp 18001
transform 1 0 24564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output233
timestamp 18001
transform -1 0 1748 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output234
timestamp 18001
transform -1 0 1748 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output235
timestamp 18001
transform -1 0 1748 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output236
timestamp 18001
transform -1 0 1748 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output237
timestamp 18001
transform -1 0 1748 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output238
timestamp 18001
transform -1 0 1748 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output239
timestamp 18001
transform -1 0 1748 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output240
timestamp 18001
transform -1 0 1748 0 1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output241
timestamp 18001
transform -1 0 1748 0 -1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output242
timestamp 18001
transform -1 0 1748 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output243
timestamp 18001
transform -1 0 1748 0 1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output244
timestamp 18001
transform -1 0 1748 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output245
timestamp 18001
transform -1 0 1748 0 -1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output246
timestamp 18001
transform -1 0 1748 0 1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output247
timestamp 18001
transform -1 0 1748 0 -1 78336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output248
timestamp 18001
transform -1 0 1748 0 -1 79424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output249
timestamp 18001
transform -1 0 1748 0 1 79424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output250
timestamp 18001
transform -1 0 1748 0 -1 81600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output251
timestamp 18001
transform -1 0 1748 0 1 81600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output252
timestamp 18001
transform -1 0 1748 0 -1 83776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output253
timestamp 18001
transform -1 0 1748 0 -1 84864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output254
timestamp 18001
transform -1 0 1748 0 1 84864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output255
timestamp 18001
transform -1 0 1748 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output256
timestamp 18001
transform -1 0 1748 0 -1 87040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output257
timestamp 18001
transform -1 0 1748 0 1 87040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output258
timestamp 18001
transform -1 0 1748 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output259
timestamp 18001
transform -1 0 1748 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output260
timestamp 18001
transform -1 0 1748 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output261
timestamp 18001
transform -1 0 1748 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output262
timestamp 18001
transform -1 0 1748 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output263
timestamp 18001
transform -1 0 1748 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output264
timestamp 18001
transform -1 0 1748 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_172
timestamp 18001
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 18001
transform -1 0 97888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_173
timestamp 18001
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 18001
transform -1 0 97888 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_174
timestamp 18001
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 18001
transform -1 0 97888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_175
timestamp 18001
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 18001
transform -1 0 97888 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_176
timestamp 18001
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 18001
transform -1 0 97888 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_177
timestamp 18001
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 18001
transform -1 0 97888 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_178
timestamp 18001
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 18001
transform -1 0 97888 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_1_Left_343
timestamp 18001
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_1_Right_663
timestamp 18001
transform -1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_3_Left_344
timestamp 18001
transform 1 0 94024 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_3_Right_12
timestamp 18001
transform -1 0 97888 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_1_Left_179
timestamp 18001
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_1_Right_504
timestamp 18001
transform -1 0 5980 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_3_Left_345
timestamp 18001
transform 1 0 94024 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_3_Right_13
timestamp 18001
transform -1 0 97888 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_1_Left_180
timestamp 18001
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_1_Right_505
timestamp 18001
transform -1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_3_Left_346
timestamp 18001
transform 1 0 94024 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_3_Right_14
timestamp 18001
transform -1 0 97888 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_1_Left_181
timestamp 18001
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_1_Right_506
timestamp 18001
transform -1 0 5980 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_3_Left_347
timestamp 18001
transform 1 0 94024 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_3_Right_15
timestamp 18001
transform -1 0 97888 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_1_Left_182
timestamp 18001
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_1_Right_507
timestamp 18001
transform -1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_3_Left_348
timestamp 18001
transform 1 0 94024 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_3_Right_16
timestamp 18001
transform -1 0 97888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_1_Left_183
timestamp 18001
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_1_Right_508
timestamp 18001
transform -1 0 5980 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_3_Left_349
timestamp 18001
transform 1 0 94024 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_3_Right_17
timestamp 18001
transform -1 0 97888 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_1_Left_184
timestamp 18001
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_1_Right_509
timestamp 18001
transform -1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_3_Left_350
timestamp 18001
transform 1 0 94024 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_3_Right_18
timestamp 18001
transform -1 0 97888 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_1_Left_185
timestamp 18001
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_1_Right_510
timestamp 18001
transform -1 0 5980 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_3_Left_351
timestamp 18001
transform 1 0 94024 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_3_Right_19
timestamp 18001
transform -1 0 97888 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_1_Left_186
timestamp 18001
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_1_Right_511
timestamp 18001
transform -1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_3_Left_352
timestamp 18001
transform 1 0 94024 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_3_Right_20
timestamp 18001
transform -1 0 97888 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_1_Left_187
timestamp 18001
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_1_Right_512
timestamp 18001
transform -1 0 5980 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_3_Left_353
timestamp 18001
transform 1 0 94024 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_3_Right_21
timestamp 18001
transform -1 0 97888 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_1_Left_188
timestamp 18001
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_1_Right_513
timestamp 18001
transform -1 0 5980 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_3_Left_354
timestamp 18001
transform 1 0 94024 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_3_Right_22
timestamp 18001
transform -1 0 97888 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_1_Left_189
timestamp 18001
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_1_Right_514
timestamp 18001
transform -1 0 5980 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_3_Left_355
timestamp 18001
transform 1 0 94024 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_3_Right_23
timestamp 18001
transform -1 0 97888 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_1_Left_190
timestamp 18001
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_1_Right_515
timestamp 18001
transform -1 0 5980 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_3_Left_356
timestamp 18001
transform 1 0 94024 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_3_Right_24
timestamp 18001
transform -1 0 97888 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_1_Left_191
timestamp 18001
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_1_Right_516
timestamp 18001
transform -1 0 5980 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_3_Left_357
timestamp 18001
transform 1 0 94024 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_3_Right_25
timestamp 18001
transform -1 0 97888 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_1_Left_192
timestamp 18001
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_1_Right_517
timestamp 18001
transform -1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_3_Left_358
timestamp 18001
transform 1 0 94024 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_3_Right_26
timestamp 18001
transform -1 0 97888 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_1_Left_193
timestamp 18001
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_1_Right_518
timestamp 18001
transform -1 0 5980 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_3_Left_359
timestamp 18001
transform 1 0 94024 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_3_Right_27
timestamp 18001
transform -1 0 97888 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_1_Left_194
timestamp 18001
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_1_Right_519
timestamp 18001
transform -1 0 5980 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_3_Left_360
timestamp 18001
transform 1 0 94024 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_3_Right_28
timestamp 18001
transform -1 0 97888 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_1_Left_195
timestamp 18001
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_1_Right_520
timestamp 18001
transform -1 0 5980 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_3_Left_361
timestamp 18001
transform 1 0 94024 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_3_Right_29
timestamp 18001
transform -1 0 97888 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_1_Left_196
timestamp 18001
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_1_Right_521
timestamp 18001
transform -1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_3_Left_362
timestamp 18001
transform 1 0 94024 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_3_Right_30
timestamp 18001
transform -1 0 97888 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_1_Left_197
timestamp 18001
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_1_Right_522
timestamp 18001
transform -1 0 5980 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_3_Left_363
timestamp 18001
transform 1 0 94024 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_3_Right_31
timestamp 18001
transform -1 0 97888 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_1_Left_198
timestamp 18001
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_1_Right_523
timestamp 18001
transform -1 0 5980 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_3_Left_364
timestamp 18001
transform 1 0 94024 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_3_Right_32
timestamp 18001
transform -1 0 97888 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_1_Left_199
timestamp 18001
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_1_Right_524
timestamp 18001
transform -1 0 5980 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_3_Left_365
timestamp 18001
transform 1 0 94024 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_3_Right_33
timestamp 18001
transform -1 0 97888 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_1_Left_200
timestamp 18001
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_1_Right_525
timestamp 18001
transform -1 0 5980 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_3_Left_366
timestamp 18001
transform 1 0 94024 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_3_Right_34
timestamp 18001
transform -1 0 97888 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_1_Left_201
timestamp 18001
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_1_Right_526
timestamp 18001
transform -1 0 5980 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_3_Left_367
timestamp 18001
transform 1 0 94024 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_3_Right_35
timestamp 18001
transform -1 0 97888 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_1_Left_202
timestamp 18001
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_1_Right_527
timestamp 18001
transform -1 0 5980 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_3_Left_368
timestamp 18001
transform 1 0 94024 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_3_Right_36
timestamp 18001
transform -1 0 97888 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_1_Left_203
timestamp 18001
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_1_Right_528
timestamp 18001
transform -1 0 5980 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_3_Left_369
timestamp 18001
transform 1 0 94024 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_3_Right_37
timestamp 18001
transform -1 0 97888 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_1_Left_204
timestamp 18001
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_1_Right_529
timestamp 18001
transform -1 0 5980 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_3_Left_370
timestamp 18001
transform 1 0 94024 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_3_Right_38
timestamp 18001
transform -1 0 97888 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_1_Left_205
timestamp 18001
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_1_Right_530
timestamp 18001
transform -1 0 5980 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_3_Left_371
timestamp 18001
transform 1 0 94024 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_3_Right_39
timestamp 18001
transform -1 0 97888 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_1_Left_206
timestamp 18001
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_1_Right_531
timestamp 18001
transform -1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_3_Left_372
timestamp 18001
transform 1 0 94024 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_3_Right_40
timestamp 18001
transform -1 0 97888 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_1_Left_207
timestamp 18001
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_1_Right_532
timestamp 18001
transform -1 0 5980 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_3_Left_373
timestamp 18001
transform 1 0 94024 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_3_Right_41
timestamp 18001
transform -1 0 97888 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_1_Left_208
timestamp 18001
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_1_Right_533
timestamp 18001
transform -1 0 5980 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_3_Left_374
timestamp 18001
transform 1 0 94024 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_3_Right_42
timestamp 18001
transform -1 0 97888 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_1_Left_209
timestamp 18001
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_1_Right_534
timestamp 18001
transform -1 0 5980 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_3_Left_375
timestamp 18001
transform 1 0 94024 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_3_Right_43
timestamp 18001
transform -1 0 97888 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_1_Left_210
timestamp 18001
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_1_Right_535
timestamp 18001
transform -1 0 5980 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_3_Left_376
timestamp 18001
transform 1 0 94024 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_3_Right_44
timestamp 18001
transform -1 0 97888 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_1_Left_211
timestamp 18001
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_1_Right_536
timestamp 18001
transform -1 0 5980 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_3_Left_377
timestamp 18001
transform 1 0 94024 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_3_Right_45
timestamp 18001
transform -1 0 97888 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_1_Left_212
timestamp 18001
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_1_Right_537
timestamp 18001
transform -1 0 5980 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_3_Left_378
timestamp 18001
transform 1 0 94024 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_3_Right_46
timestamp 18001
transform -1 0 97888 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_1_Left_213
timestamp 18001
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_1_Right_538
timestamp 18001
transform -1 0 5980 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_3_Left_379
timestamp 18001
transform 1 0 94024 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_3_Right_47
timestamp 18001
transform -1 0 97888 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_1_Left_214
timestamp 18001
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_1_Right_539
timestamp 18001
transform -1 0 5980 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_3_Left_380
timestamp 18001
transform 1 0 94024 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_3_Right_48
timestamp 18001
transform -1 0 97888 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_1_Left_215
timestamp 18001
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_1_Right_540
timestamp 18001
transform -1 0 5980 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_3_Left_381
timestamp 18001
transform 1 0 94024 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_3_Right_49
timestamp 18001
transform -1 0 97888 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_1_Left_216
timestamp 18001
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_1_Right_541
timestamp 18001
transform -1 0 5980 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_3_Left_382
timestamp 18001
transform 1 0 94024 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_3_Right_50
timestamp 18001
transform -1 0 97888 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_1_Left_217
timestamp 18001
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_1_Right_542
timestamp 18001
transform -1 0 5980 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_3_Left_383
timestamp 18001
transform 1 0 94024 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_3_Right_51
timestamp 18001
transform -1 0 97888 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_1_Left_218
timestamp 18001
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_1_Right_543
timestamp 18001
transform -1 0 5980 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_3_Left_384
timestamp 18001
transform 1 0 94024 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_3_Right_52
timestamp 18001
transform -1 0 97888 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_1_Left_219
timestamp 18001
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_1_Right_544
timestamp 18001
transform -1 0 5980 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_3_Left_385
timestamp 18001
transform 1 0 94024 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_3_Right_53
timestamp 18001
transform -1 0 97888 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_1_Left_220
timestamp 18001
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_1_Right_545
timestamp 18001
transform -1 0 5980 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_3_Left_386
timestamp 18001
transform 1 0 94024 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_3_Right_54
timestamp 18001
transform -1 0 97888 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_1_Left_221
timestamp 18001
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_1_Right_546
timestamp 18001
transform -1 0 5980 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_3_Left_387
timestamp 18001
transform 1 0 94024 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_3_Right_55
timestamp 18001
transform -1 0 97888 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_1_Left_222
timestamp 18001
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_1_Right_547
timestamp 18001
transform -1 0 5980 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_3_Left_388
timestamp 18001
transform 1 0 94024 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_3_Right_56
timestamp 18001
transform -1 0 97888 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_1_Left_223
timestamp 18001
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_1_Right_548
timestamp 18001
transform -1 0 5980 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_3_Left_389
timestamp 18001
transform 1 0 94024 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_3_Right_57
timestamp 18001
transform -1 0 97888 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_1_Left_224
timestamp 18001
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_1_Right_549
timestamp 18001
transform -1 0 5980 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_3_Left_390
timestamp 18001
transform 1 0 94024 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_3_Right_58
timestamp 18001
transform -1 0 97888 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_1_Left_225
timestamp 18001
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_1_Right_550
timestamp 18001
transform -1 0 5980 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_3_Left_391
timestamp 18001
transform 1 0 94024 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_3_Right_59
timestamp 18001
transform -1 0 97888 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_1_Left_226
timestamp 18001
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_1_Right_551
timestamp 18001
transform -1 0 5980 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_3_Left_392
timestamp 18001
transform 1 0 94024 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_3_Right_60
timestamp 18001
transform -1 0 97888 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_1_Left_227
timestamp 18001
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_1_Right_552
timestamp 18001
transform -1 0 5980 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_3_Left_393
timestamp 18001
transform 1 0 94024 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_3_Right_61
timestamp 18001
transform -1 0 97888 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_1_Left_228
timestamp 18001
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_1_Right_553
timestamp 18001
transform -1 0 5980 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_3_Left_394
timestamp 18001
transform 1 0 94024 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_3_Right_62
timestamp 18001
transform -1 0 97888 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_1_Left_229
timestamp 18001
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_1_Right_554
timestamp 18001
transform -1 0 5980 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_3_Left_395
timestamp 18001
transform 1 0 94024 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_3_Right_63
timestamp 18001
transform -1 0 97888 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_1_Left_230
timestamp 18001
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_1_Right_555
timestamp 18001
transform -1 0 5980 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_3_Left_396
timestamp 18001
transform 1 0 94024 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_3_Right_64
timestamp 18001
transform -1 0 97888 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_1_Left_231
timestamp 18001
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_1_Right_556
timestamp 18001
transform -1 0 5980 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_3_Left_397
timestamp 18001
transform 1 0 94024 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_3_Right_65
timestamp 18001
transform -1 0 97888 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_1_Left_232
timestamp 18001
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_1_Right_557
timestamp 18001
transform -1 0 5980 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_3_Left_398
timestamp 18001
transform 1 0 94024 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_3_Right_66
timestamp 18001
transform -1 0 97888 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_1_Left_233
timestamp 18001
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_1_Right_558
timestamp 18001
transform -1 0 5980 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_3_Left_399
timestamp 18001
transform 1 0 94024 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_3_Right_67
timestamp 18001
transform -1 0 97888 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_1_Left_234
timestamp 18001
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_1_Right_559
timestamp 18001
transform -1 0 5980 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_3_Left_400
timestamp 18001
transform 1 0 94024 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_3_Right_68
timestamp 18001
transform -1 0 97888 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_1_Left_235
timestamp 18001
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_1_Right_560
timestamp 18001
transform -1 0 5980 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_3_Left_401
timestamp 18001
transform 1 0 94024 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_3_Right_69
timestamp 18001
transform -1 0 97888 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_1_Left_236
timestamp 18001
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_1_Right_561
timestamp 18001
transform -1 0 5980 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_3_Left_402
timestamp 18001
transform 1 0 94024 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_3_Right_70
timestamp 18001
transform -1 0 97888 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_1_Left_237
timestamp 18001
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_1_Right_562
timestamp 18001
transform -1 0 5980 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_3_Left_403
timestamp 18001
transform 1 0 94024 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_3_Right_71
timestamp 18001
transform -1 0 97888 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_1_Left_238
timestamp 18001
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_1_Right_563
timestamp 18001
transform -1 0 5980 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_3_Left_404
timestamp 18001
transform 1 0 94024 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_3_Right_72
timestamp 18001
transform -1 0 97888 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_1_Left_239
timestamp 18001
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_1_Right_564
timestamp 18001
transform -1 0 5980 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_3_Left_405
timestamp 18001
transform 1 0 94024 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_3_Right_73
timestamp 18001
transform -1 0 97888 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_1_Left_240
timestamp 18001
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_1_Right_565
timestamp 18001
transform -1 0 5980 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_3_Left_406
timestamp 18001
transform 1 0 94024 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_3_Right_74
timestamp 18001
transform -1 0 97888 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_1_Left_241
timestamp 18001
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_1_Right_566
timestamp 18001
transform -1 0 5980 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_3_Left_407
timestamp 18001
transform 1 0 94024 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_3_Right_75
timestamp 18001
transform -1 0 97888 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_1_Left_242
timestamp 18001
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_1_Right_567
timestamp 18001
transform -1 0 5980 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_3_Left_408
timestamp 18001
transform 1 0 94024 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_3_Right_76
timestamp 18001
transform -1 0 97888 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_1_Left_243
timestamp 18001
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_1_Right_568
timestamp 18001
transform -1 0 5980 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_3_Left_409
timestamp 18001
transform 1 0 94024 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_3_Right_77
timestamp 18001
transform -1 0 97888 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_1_Left_244
timestamp 18001
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_1_Right_569
timestamp 18001
transform -1 0 5980 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_3_Left_410
timestamp 18001
transform 1 0 94024 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_3_Right_78
timestamp 18001
transform -1 0 97888 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_1_Left_245
timestamp 18001
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_1_Right_570
timestamp 18001
transform -1 0 5980 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_3_Left_411
timestamp 18001
transform 1 0 94024 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_3_Right_79
timestamp 18001
transform -1 0 97888 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_1_Left_246
timestamp 18001
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_1_Right_571
timestamp 18001
transform -1 0 5980 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_3_Left_412
timestamp 18001
transform 1 0 94024 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_3_Right_80
timestamp 18001
transform -1 0 97888 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_1_Left_247
timestamp 18001
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_1_Right_572
timestamp 18001
transform -1 0 5980 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_3_Left_413
timestamp 18001
transform 1 0 94024 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_3_Right_81
timestamp 18001
transform -1 0 97888 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_1_Left_248
timestamp 18001
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_1_Right_573
timestamp 18001
transform -1 0 5980 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_3_Left_414
timestamp 18001
transform 1 0 94024 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_3_Right_82
timestamp 18001
transform -1 0 97888 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_1_Left_249
timestamp 18001
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_1_Right_574
timestamp 18001
transform -1 0 5980 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_3_Left_415
timestamp 18001
transform 1 0 94024 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_3_Right_83
timestamp 18001
transform -1 0 97888 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_1_Left_250
timestamp 18001
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_1_Right_575
timestamp 18001
transform -1 0 5980 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_3_Left_416
timestamp 18001
transform 1 0 94024 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_3_Right_84
timestamp 18001
transform -1 0 97888 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_1_Left_251
timestamp 18001
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_1_Right_576
timestamp 18001
transform -1 0 5980 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_3_Left_417
timestamp 18001
transform 1 0 94024 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_3_Right_85
timestamp 18001
transform -1 0 97888 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_1_Left_252
timestamp 18001
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_1_Right_577
timestamp 18001
transform -1 0 5980 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_3_Left_418
timestamp 18001
transform 1 0 94024 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_3_Right_86
timestamp 18001
transform -1 0 97888 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_1_Left_253
timestamp 18001
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_1_Right_578
timestamp 18001
transform -1 0 5980 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_3_Left_419
timestamp 18001
transform 1 0 94024 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_3_Right_87
timestamp 18001
transform -1 0 97888 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_1_Left_254
timestamp 18001
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_1_Right_579
timestamp 18001
transform -1 0 5980 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_3_Left_420
timestamp 18001
transform 1 0 94024 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_3_Right_88
timestamp 18001
transform -1 0 97888 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_1_Left_255
timestamp 18001
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_1_Right_580
timestamp 18001
transform -1 0 5980 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_5_Left_421
timestamp 18001
transform 1 0 94024 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_5_Right_89
timestamp 18001
transform -1 0 97888 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_1_Left_256
timestamp 18001
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_1_Right_581
timestamp 18001
transform -1 0 5980 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_5_Left_422
timestamp 18001
transform 1 0 94024 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_5_Right_90
timestamp 18001
transform -1 0 97888 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_1_Left_257
timestamp 18001
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_1_Right_582
timestamp 18001
transform -1 0 5980 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_5_Left_423
timestamp 18001
transform 1 0 94024 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_5_Right_91
timestamp 18001
transform -1 0 97888 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_1_Left_258
timestamp 18001
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_1_Right_583
timestamp 18001
transform -1 0 5980 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_5_Left_424
timestamp 18001
transform 1 0 94024 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_5_Right_92
timestamp 18001
transform -1 0 97888 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_1_Left_259
timestamp 18001
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_1_Right_584
timestamp 18001
transform -1 0 5980 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_5_Left_425
timestamp 18001
transform 1 0 94024 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_5_Right_93
timestamp 18001
transform -1 0 97888 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_1_Left_260
timestamp 18001
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_1_Right_585
timestamp 18001
transform -1 0 5980 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_5_Left_426
timestamp 18001
transform 1 0 94024 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_5_Right_94
timestamp 18001
transform -1 0 97888 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_1_Left_261
timestamp 18001
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_1_Right_586
timestamp 18001
transform -1 0 5980 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_3_Left_427
timestamp 18001
transform 1 0 94024 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_3_Right_95
timestamp 18001
transform -1 0 97888 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_1_Left_262
timestamp 18001
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_1_Right_587
timestamp 18001
transform -1 0 5980 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_3_Left_428
timestamp 18001
transform 1 0 94024 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_3_Right_96
timestamp 18001
transform -1 0 97888 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_1_Left_263
timestamp 18001
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_1_Right_588
timestamp 18001
transform -1 0 5980 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_3_Left_429
timestamp 18001
transform 1 0 94024 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_3_Right_97
timestamp 18001
transform -1 0 97888 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_1_Left_264
timestamp 18001
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_1_Right_589
timestamp 18001
transform -1 0 5980 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_3_Left_430
timestamp 18001
transform 1 0 94024 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_3_Right_98
timestamp 18001
transform -1 0 97888 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_1_Left_265
timestamp 18001
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_1_Right_590
timestamp 18001
transform -1 0 5980 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_3_Left_431
timestamp 18001
transform 1 0 94024 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_3_Right_99
timestamp 18001
transform -1 0 97888 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_1_Left_266
timestamp 18001
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_1_Right_591
timestamp 18001
transform -1 0 5980 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_3_Left_432
timestamp 18001
transform 1 0 94024 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_3_Right_100
timestamp 18001
transform -1 0 97888 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_1_Left_267
timestamp 18001
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_1_Right_592
timestamp 18001
transform -1 0 5980 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_3_Left_433
timestamp 18001
transform 1 0 94024 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_3_Right_101
timestamp 18001
transform -1 0 97888 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_1_Left_268
timestamp 18001
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_1_Right_593
timestamp 18001
transform -1 0 5980 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_3_Left_434
timestamp 18001
transform 1 0 94024 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_3_Right_102
timestamp 18001
transform -1 0 97888 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_1_Left_269
timestamp 18001
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_1_Right_594
timestamp 18001
transform -1 0 5980 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_3_Left_435
timestamp 18001
transform 1 0 94024 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_3_Right_103
timestamp 18001
transform -1 0 97888 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_1_Left_270
timestamp 18001
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_1_Right_595
timestamp 18001
transform -1 0 5980 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_3_Left_436
timestamp 18001
transform 1 0 94024 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_3_Right_104
timestamp 18001
transform -1 0 97888 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_1_Left_271
timestamp 18001
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_1_Right_596
timestamp 18001
transform -1 0 5980 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_3_Left_437
timestamp 18001
transform 1 0 94024 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_3_Right_105
timestamp 18001
transform -1 0 97888 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_1_Left_272
timestamp 18001
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_1_Right_597
timestamp 18001
transform -1 0 5980 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_3_Left_438
timestamp 18001
transform 1 0 94024 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_3_Right_106
timestamp 18001
transform -1 0 97888 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_1_Left_273
timestamp 18001
transform 1 0 1104 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_1_Right_598
timestamp 18001
transform -1 0 5980 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_3_Left_439
timestamp 18001
transform 1 0 94024 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_3_Right_107
timestamp 18001
transform -1 0 97888 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_1_Left_274
timestamp 18001
transform 1 0 1104 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_1_Right_599
timestamp 18001
transform -1 0 5980 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_3_Left_440
timestamp 18001
transform 1 0 94024 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_3_Right_108
timestamp 18001
transform -1 0 97888 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_1_Left_275
timestamp 18001
transform 1 0 1104 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_1_Right_600
timestamp 18001
transform -1 0 5980 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_3_Left_441
timestamp 18001
transform 1 0 94024 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_3_Right_109
timestamp 18001
transform -1 0 97888 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_1_Left_276
timestamp 18001
transform 1 0 1104 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_1_Right_601
timestamp 18001
transform -1 0 5980 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_3_Left_442
timestamp 18001
transform 1 0 94024 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_3_Right_110
timestamp 18001
transform -1 0 97888 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_1_Left_277
timestamp 18001
transform 1 0 1104 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_1_Right_602
timestamp 18001
transform -1 0 5980 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_3_Left_443
timestamp 18001
transform 1 0 94024 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_3_Right_111
timestamp 18001
transform -1 0 97888 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_1_Left_278
timestamp 18001
transform 1 0 1104 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_1_Right_603
timestamp 18001
transform -1 0 5980 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_3_Left_444
timestamp 18001
transform 1 0 94024 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_3_Right_112
timestamp 18001
transform -1 0 97888 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_1_Left_279
timestamp 18001
transform 1 0 1104 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_1_Right_604
timestamp 18001
transform -1 0 5980 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_3_Left_445
timestamp 18001
transform 1 0 94024 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_3_Right_113
timestamp 18001
transform -1 0 97888 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_1_Left_280
timestamp 18001
transform 1 0 1104 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_1_Right_605
timestamp 18001
transform -1 0 5980 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_3_Left_446
timestamp 18001
transform 1 0 94024 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_3_Right_114
timestamp 18001
transform -1 0 97888 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_1_Left_281
timestamp 18001
transform 1 0 1104 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_1_Right_606
timestamp 18001
transform -1 0 5980 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_3_Left_447
timestamp 18001
transform 1 0 94024 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_3_Right_115
timestamp 18001
transform -1 0 97888 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_1_Left_282
timestamp 18001
transform 1 0 1104 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_1_Right_607
timestamp 18001
transform -1 0 5980 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_3_Left_448
timestamp 18001
transform 1 0 94024 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_3_Right_116
timestamp 18001
transform -1 0 97888 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_1_Left_283
timestamp 18001
transform 1 0 1104 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_1_Right_608
timestamp 18001
transform -1 0 5980 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_3_Left_449
timestamp 18001
transform 1 0 94024 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_3_Right_117
timestamp 18001
transform -1 0 97888 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_1_Left_284
timestamp 18001
transform 1 0 1104 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_1_Right_609
timestamp 18001
transform -1 0 5980 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_3_Left_450
timestamp 18001
transform 1 0 94024 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_3_Right_118
timestamp 18001
transform -1 0 97888 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_1_Left_285
timestamp 18001
transform 1 0 1104 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_1_Right_610
timestamp 18001
transform -1 0 5980 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_3_Left_451
timestamp 18001
transform 1 0 94024 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_3_Right_119
timestamp 18001
transform -1 0 97888 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_1_Left_286
timestamp 18001
transform 1 0 1104 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_1_Right_611
timestamp 18001
transform -1 0 5980 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_3_Left_452
timestamp 18001
transform 1 0 94024 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_3_Right_120
timestamp 18001
transform -1 0 97888 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_1_Left_287
timestamp 18001
transform 1 0 1104 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_1_Right_612
timestamp 18001
transform -1 0 5980 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_3_Left_453
timestamp 18001
transform 1 0 94024 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_3_Right_121
timestamp 18001
transform -1 0 97888 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_117_1_Left_288
timestamp 18001
transform 1 0 1104 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_117_1_Right_613
timestamp 18001
transform -1 0 5980 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_117_3_Left_454
timestamp 18001
transform 1 0 94024 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_117_3_Right_122
timestamp 18001
transform -1 0 97888 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_118_1_Left_289
timestamp 18001
transform 1 0 1104 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_118_1_Right_614
timestamp 18001
transform -1 0 5980 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_118_3_Left_455
timestamp 18001
transform 1 0 94024 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_118_3_Right_123
timestamp 18001
transform -1 0 97888 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_119_1_Left_290
timestamp 18001
transform 1 0 1104 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_119_1_Right_615
timestamp 18001
transform -1 0 5980 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_119_3_Left_456
timestamp 18001
transform 1 0 94024 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_119_3_Right_124
timestamp 18001
transform -1 0 97888 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_120_1_Left_291
timestamp 18001
transform 1 0 1104 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_120_1_Right_616
timestamp 18001
transform -1 0 5980 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_120_3_Left_457
timestamp 18001
transform 1 0 94024 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_120_3_Right_125
timestamp 18001
transform -1 0 97888 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_121_1_Left_292
timestamp 18001
transform 1 0 1104 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_121_1_Right_617
timestamp 18001
transform -1 0 5980 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_121_3_Left_458
timestamp 18001
transform 1 0 94024 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_121_3_Right_126
timestamp 18001
transform -1 0 97888 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_122_1_Left_293
timestamp 18001
transform 1 0 1104 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_122_1_Right_618
timestamp 18001
transform -1 0 5980 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_122_3_Left_459
timestamp 18001
transform 1 0 94024 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_122_3_Right_127
timestamp 18001
transform -1 0 97888 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_123_1_Left_294
timestamp 18001
transform 1 0 1104 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_123_1_Right_619
timestamp 18001
transform -1 0 5980 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_123_3_Left_460
timestamp 18001
transform 1 0 94024 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_123_3_Right_128
timestamp 18001
transform -1 0 97888 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_124_1_Left_295
timestamp 18001
transform 1 0 1104 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_124_1_Right_620
timestamp 18001
transform -1 0 5980 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_124_3_Left_461
timestamp 18001
transform 1 0 94024 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_124_3_Right_129
timestamp 18001
transform -1 0 97888 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_125_1_Left_296
timestamp 18001
transform 1 0 1104 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_125_1_Right_621
timestamp 18001
transform -1 0 5980 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_125_3_Left_462
timestamp 18001
transform 1 0 94024 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_125_3_Right_130
timestamp 18001
transform -1 0 97888 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_126_1_Left_297
timestamp 18001
transform 1 0 1104 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_126_1_Right_622
timestamp 18001
transform -1 0 5980 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_126_3_Left_463
timestamp 18001
transform 1 0 94024 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_126_3_Right_131
timestamp 18001
transform -1 0 97888 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_127_1_Left_298
timestamp 18001
transform 1 0 1104 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_127_1_Right_623
timestamp 18001
transform -1 0 5980 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_127_3_Left_464
timestamp 18001
transform 1 0 94024 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_127_3_Right_132
timestamp 18001
transform -1 0 97888 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_128_1_Left_299
timestamp 18001
transform 1 0 1104 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_128_1_Right_624
timestamp 18001
transform -1 0 5980 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_128_3_Left_465
timestamp 18001
transform 1 0 94024 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_128_3_Right_133
timestamp 18001
transform -1 0 97888 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_129_1_Left_300
timestamp 18001
transform 1 0 1104 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_129_1_Right_625
timestamp 18001
transform -1 0 5980 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_129_3_Left_466
timestamp 18001
transform 1 0 94024 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_129_3_Right_134
timestamp 18001
transform -1 0 97888 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_130_1_Left_301
timestamp 18001
transform 1 0 1104 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_130_1_Right_626
timestamp 18001
transform -1 0 5980 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_130_3_Left_467
timestamp 18001
transform 1 0 94024 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_130_3_Right_135
timestamp 18001
transform -1 0 97888 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_131_1_Left_302
timestamp 18001
transform 1 0 1104 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_131_1_Right_627
timestamp 18001
transform -1 0 5980 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_131_3_Left_468
timestamp 18001
transform 1 0 94024 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_131_3_Right_136
timestamp 18001
transform -1 0 97888 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_132_1_Left_303
timestamp 18001
transform 1 0 1104 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_132_1_Right_628
timestamp 18001
transform -1 0 5980 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_132_3_Left_469
timestamp 18001
transform 1 0 94024 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_132_3_Right_137
timestamp 18001
transform -1 0 97888 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_133_1_Left_304
timestamp 18001
transform 1 0 1104 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_133_1_Right_629
timestamp 18001
transform -1 0 5980 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_133_3_Left_470
timestamp 18001
transform 1 0 94024 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_133_3_Right_138
timestamp 18001
transform -1 0 97888 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_134_1_Left_305
timestamp 18001
transform 1 0 1104 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_134_1_Right_630
timestamp 18001
transform -1 0 5980 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_134_3_Left_471
timestamp 18001
transform 1 0 94024 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_134_3_Right_139
timestamp 18001
transform -1 0 97888 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_135_1_Left_306
timestamp 18001
transform 1 0 1104 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_135_1_Right_631
timestamp 18001
transform -1 0 5980 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_135_3_Left_472
timestamp 18001
transform 1 0 94024 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_135_3_Right_140
timestamp 18001
transform -1 0 97888 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_136_1_Left_307
timestamp 18001
transform 1 0 1104 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_136_1_Right_632
timestamp 18001
transform -1 0 5980 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_136_3_Left_473
timestamp 18001
transform 1 0 94024 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_136_3_Right_141
timestamp 18001
transform -1 0 97888 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_137_1_Left_308
timestamp 18001
transform 1 0 1104 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_137_1_Right_633
timestamp 18001
transform -1 0 5980 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_137_3_Left_474
timestamp 18001
transform 1 0 94024 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_137_3_Right_142
timestamp 18001
transform -1 0 97888 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_138_1_Left_309
timestamp 18001
transform 1 0 1104 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_138_1_Right_634
timestamp 18001
transform -1 0 5980 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_138_3_Left_475
timestamp 18001
transform 1 0 94024 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_138_3_Right_143
timestamp 18001
transform -1 0 97888 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_139_1_Left_310
timestamp 18001
transform 1 0 1104 0 -1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_139_1_Right_635
timestamp 18001
transform -1 0 5980 0 -1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_139_3_Left_476
timestamp 18001
transform 1 0 94024 0 -1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_139_3_Right_144
timestamp 18001
transform -1 0 97888 0 -1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_140_1_Left_311
timestamp 18001
transform 1 0 1104 0 1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_140_1_Right_636
timestamp 18001
transform -1 0 5980 0 1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_140_3_Left_477
timestamp 18001
transform 1 0 94024 0 1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_140_3_Right_145
timestamp 18001
transform -1 0 97888 0 1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_141_1_Left_312
timestamp 18001
transform 1 0 1104 0 -1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_141_1_Right_637
timestamp 18001
transform -1 0 5980 0 -1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_141_3_Left_478
timestamp 18001
transform 1 0 94024 0 -1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_141_3_Right_146
timestamp 18001
transform -1 0 97888 0 -1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_142_1_Left_313
timestamp 18001
transform 1 0 1104 0 1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_142_1_Right_638
timestamp 18001
transform -1 0 5980 0 1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_142_3_Left_479
timestamp 18001
transform 1 0 94024 0 1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_142_3_Right_147
timestamp 18001
transform -1 0 97888 0 1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_143_1_Left_314
timestamp 18001
transform 1 0 1104 0 -1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_143_1_Right_639
timestamp 18001
transform -1 0 5980 0 -1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_143_3_Left_480
timestamp 18001
transform 1 0 94024 0 -1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_143_3_Right_148
timestamp 18001
transform -1 0 97888 0 -1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_144_1_Left_315
timestamp 18001
transform 1 0 1104 0 1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_144_1_Right_640
timestamp 18001
transform -1 0 5980 0 1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_144_3_Left_481
timestamp 18001
transform 1 0 94024 0 1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_144_3_Right_149
timestamp 18001
transform -1 0 97888 0 1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_145_1_Left_316
timestamp 18001
transform 1 0 1104 0 -1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_145_1_Right_641
timestamp 18001
transform -1 0 5980 0 -1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_145_3_Left_482
timestamp 18001
transform 1 0 94024 0 -1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_145_3_Right_150
timestamp 18001
transform -1 0 97888 0 -1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_146_1_Left_317
timestamp 18001
transform 1 0 1104 0 1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_146_1_Right_642
timestamp 18001
transform -1 0 5980 0 1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_146_3_Left_483
timestamp 18001
transform 1 0 94024 0 1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_146_3_Right_151
timestamp 18001
transform -1 0 97888 0 1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_147_1_Left_318
timestamp 18001
transform 1 0 1104 0 -1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_147_1_Right_643
timestamp 18001
transform -1 0 5980 0 -1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_147_3_Left_484
timestamp 18001
transform 1 0 94024 0 -1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_147_3_Right_152
timestamp 18001
transform -1 0 97888 0 -1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_148_1_Left_319
timestamp 18001
transform 1 0 1104 0 1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_148_1_Right_644
timestamp 18001
transform -1 0 5980 0 1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_148_3_Left_485
timestamp 18001
transform 1 0 94024 0 1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_148_3_Right_153
timestamp 18001
transform -1 0 97888 0 1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_149_1_Left_320
timestamp 18001
transform 1 0 1104 0 -1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_149_1_Right_645
timestamp 18001
transform -1 0 5980 0 -1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_149_3_Left_486
timestamp 18001
transform 1 0 94024 0 -1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_149_3_Right_154
timestamp 18001
transform -1 0 97888 0 -1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_150_1_Left_321
timestamp 18001
transform 1 0 1104 0 1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_150_1_Right_646
timestamp 18001
transform -1 0 5980 0 1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_150_3_Left_487
timestamp 18001
transform 1 0 94024 0 1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_150_3_Right_155
timestamp 18001
transform -1 0 97888 0 1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_151_1_Left_322
timestamp 18001
transform 1 0 1104 0 -1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_151_1_Right_647
timestamp 18001
transform -1 0 5980 0 -1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_151_3_Left_488
timestamp 18001
transform 1 0 94024 0 -1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_151_3_Right_156
timestamp 18001
transform -1 0 97888 0 -1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_152_1_Left_323
timestamp 18001
transform 1 0 1104 0 1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_152_1_Right_648
timestamp 18001
transform -1 0 5980 0 1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_152_3_Left_489
timestamp 18001
transform 1 0 94024 0 1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_152_3_Right_157
timestamp 18001
transform -1 0 97888 0 1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_153_1_Left_324
timestamp 18001
transform 1 0 1104 0 -1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_153_1_Right_649
timestamp 18001
transform -1 0 5980 0 -1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_153_3_Left_490
timestamp 18001
transform 1 0 94024 0 -1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_153_3_Right_158
timestamp 18001
transform -1 0 97888 0 -1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_154_1_Left_325
timestamp 18001
transform 1 0 1104 0 1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_154_1_Right_650
timestamp 18001
transform -1 0 5980 0 1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_154_3_Left_491
timestamp 18001
transform 1 0 94024 0 1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_154_3_Right_159
timestamp 18001
transform -1 0 97888 0 1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_155_1_Left_326
timestamp 18001
transform 1 0 1104 0 -1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_155_1_Right_651
timestamp 18001
transform -1 0 5980 0 -1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_155_3_Left_492
timestamp 18001
transform 1 0 94024 0 -1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_155_3_Right_160
timestamp 18001
transform -1 0 97888 0 -1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_156_1_Left_327
timestamp 18001
transform 1 0 1104 0 1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_156_1_Right_652
timestamp 18001
transform -1 0 5980 0 1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_156_3_Left_493
timestamp 18001
transform 1 0 94024 0 1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_156_3_Right_161
timestamp 18001
transform -1 0 97888 0 1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_157_1_Left_328
timestamp 18001
transform 1 0 1104 0 -1 88128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_157_1_Right_653
timestamp 18001
transform -1 0 5980 0 -1 88128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_157_3_Left_494
timestamp 18001
transform 1 0 94024 0 -1 88128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_157_3_Right_162
timestamp 18001
transform -1 0 97888 0 -1 88128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_158_1_Left_329
timestamp 18001
transform 1 0 1104 0 1 88128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_158_1_Right_654
timestamp 18001
transform -1 0 5980 0 1 88128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_158_3_Left_495
timestamp 18001
transform 1 0 94024 0 1 88128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_158_3_Right_163
timestamp 18001
transform -1 0 97888 0 1 88128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_159_1_Left_330
timestamp 18001
transform 1 0 1104 0 -1 89216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_159_1_Right_655
timestamp 18001
transform -1 0 5980 0 -1 89216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_159_3_Left_496
timestamp 18001
transform 1 0 94024 0 -1 89216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_159_3_Right_164
timestamp 18001
transform -1 0 97888 0 -1 89216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_160_1_Left_331
timestamp 18001
transform 1 0 1104 0 1 89216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_160_1_Right_656
timestamp 18001
transform -1 0 5980 0 1 89216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_160_3_Left_497
timestamp 18001
transform 1 0 94024 0 1 89216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_160_3_Right_165
timestamp 18001
transform -1 0 97888 0 1 89216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_161_1_Left_332
timestamp 18001
transform 1 0 1104 0 -1 90304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_161_1_Right_657
timestamp 18001
transform -1 0 5980 0 -1 90304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_161_3_Left_498
timestamp 18001
transform 1 0 94024 0 -1 90304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_161_3_Right_166
timestamp 18001
transform -1 0 97888 0 -1 90304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_162_1_Left_333
timestamp 18001
transform 1 0 1104 0 1 90304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_162_1_Right_658
timestamp 18001
transform -1 0 5980 0 1 90304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_162_3_Left_499
timestamp 18001
transform 1 0 94024 0 1 90304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_162_3_Right_167
timestamp 18001
transform -1 0 97888 0 1 90304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_163_1_Left_334
timestamp 18001
transform 1 0 1104 0 -1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_163_1_Right_659
timestamp 18001
transform -1 0 5980 0 -1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_163_3_Left_500
timestamp 18001
transform 1 0 94024 0 -1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_163_3_Right_168
timestamp 18001
transform -1 0 97888 0 -1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_164_1_Left_335
timestamp 18001
transform 1 0 1104 0 1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_164_1_Right_660
timestamp 18001
transform -1 0 5980 0 1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_164_3_Left_501
timestamp 18001
transform 1 0 94024 0 1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_164_3_Right_169
timestamp 18001
transform -1 0 97888 0 1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_165_1_Left_336
timestamp 18001
transform 1 0 1104 0 -1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_165_1_Right_661
timestamp 18001
transform -1 0 5980 0 -1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_165_3_Left_502
timestamp 18001
transform 1 0 94024 0 -1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_165_3_Right_170
timestamp 18001
transform -1 0 97888 0 -1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_166_1_Left_337
timestamp 18001
transform 1 0 1104 0 1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_166_1_Right_662
timestamp 18001
transform -1 0 5980 0 1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_166_3_Left_503
timestamp 18001
transform 1 0 94024 0 1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_166_3_Right_171
timestamp 18001
transform -1 0 97888 0 1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_167_Left_338
timestamp 18001
transform 1 0 1104 0 -1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_167_Right_7
timestamp 18001
transform -1 0 97888 0 -1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_168_Left_339
timestamp 18001
transform 1 0 1104 0 1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_168_Right_8
timestamp 18001
transform -1 0 97888 0 1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_169_Left_340
timestamp 18001
transform 1 0 1104 0 -1 94656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_169_Right_9
timestamp 18001
transform -1 0 97888 0 -1 94656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_170_Left_341
timestamp 18001
transform 1 0 1104 0 1 94656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_170_Right_10
timestamp 18001
transform -1 0 97888 0 1 94656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_171_Left_342
timestamp 18001
transform 1 0 1104 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_171_Right_11
timestamp 18001
transform -1 0 97888 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_664
timestamp 18001
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_665
timestamp 18001
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_666
timestamp 18001
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_667
timestamp 18001
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_668
timestamp 18001
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_669
timestamp 18001
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_670
timestamp 18001
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_671
timestamp 18001
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_672
timestamp 18001
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_673
timestamp 18001
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_674
timestamp 18001
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_675
timestamp 18001
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_676
timestamp 18001
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_677
timestamp 18001
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_678
timestamp 18001
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_679
timestamp 18001
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_680
timestamp 18001
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_681
timestamp 18001
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_682
timestamp 18001
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_683
timestamp 18001
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_684
timestamp 18001
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_685
timestamp 18001
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_686
timestamp 18001
transform 1 0 60352 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_687
timestamp 18001
transform 1 0 62928 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_688
timestamp 18001
transform 1 0 65504 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_689
timestamp 18001
transform 1 0 68080 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_690
timestamp 18001
transform 1 0 70656 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_691
timestamp 18001
transform 1 0 73232 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_692
timestamp 18001
transform 1 0 75808 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_693
timestamp 18001
transform 1 0 78384 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_694
timestamp 18001
transform 1 0 80960 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_695
timestamp 18001
transform 1 0 83536 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_696
timestamp 18001
transform 1 0 86112 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_697
timestamp 18001
transform 1 0 88688 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_698
timestamp 18001
transform 1 0 91264 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_699
timestamp 18001
transform 1 0 93840 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_700
timestamp 18001
transform 1 0 96416 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_701
timestamp 18001
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_702
timestamp 18001
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_703
timestamp 18001
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_704
timestamp 18001
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_705
timestamp 18001
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_706
timestamp 18001
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_707
timestamp 18001
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_708
timestamp 18001
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_709
timestamp 18001
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_710
timestamp 18001
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_711
timestamp 18001
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_712
timestamp 18001
transform 1 0 62928 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_713
timestamp 18001
transform 1 0 68080 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_714
timestamp 18001
transform 1 0 73232 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_715
timestamp 18001
transform 1 0 78384 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_716
timestamp 18001
transform 1 0 83536 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_717
timestamp 18001
transform 1 0 88688 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_718
timestamp 18001
transform 1 0 93840 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_719
timestamp 18001
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_720
timestamp 18001
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_721
timestamp 18001
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_722
timestamp 18001
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_723
timestamp 18001
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_724
timestamp 18001
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_725
timestamp 18001
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_726
timestamp 18001
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_727
timestamp 18001
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_728
timestamp 18001
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_729
timestamp 18001
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_730
timestamp 18001
transform 1 0 60352 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_731
timestamp 18001
transform 1 0 65504 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_732
timestamp 18001
transform 1 0 70656 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_733
timestamp 18001
transform 1 0 75808 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_734
timestamp 18001
transform 1 0 80960 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_735
timestamp 18001
transform 1 0 86112 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_736
timestamp 18001
transform 1 0 91264 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_737
timestamp 18001
transform 1 0 96416 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_738
timestamp 18001
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_739
timestamp 18001
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_740
timestamp 18001
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_741
timestamp 18001
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_742
timestamp 18001
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_743
timestamp 18001
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_744
timestamp 18001
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_745
timestamp 18001
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_746
timestamp 18001
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_747
timestamp 18001
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_748
timestamp 18001
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_749
timestamp 18001
transform 1 0 62928 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_750
timestamp 18001
transform 1 0 68080 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_751
timestamp 18001
transform 1 0 73232 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_752
timestamp 18001
transform 1 0 78384 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_753
timestamp 18001
transform 1 0 83536 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_754
timestamp 18001
transform 1 0 88688 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_755
timestamp 18001
transform 1 0 93840 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_756
timestamp 18001
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_757
timestamp 18001
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_758
timestamp 18001
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_759
timestamp 18001
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_760
timestamp 18001
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_761
timestamp 18001
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_762
timestamp 18001
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_763
timestamp 18001
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_764
timestamp 18001
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_765
timestamp 18001
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_766
timestamp 18001
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_767
timestamp 18001
transform 1 0 60352 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_768
timestamp 18001
transform 1 0 65504 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_769
timestamp 18001
transform 1 0 70656 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_770
timestamp 18001
transform 1 0 75808 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_771
timestamp 18001
transform 1 0 80960 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_772
timestamp 18001
transform 1 0 86112 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_773
timestamp 18001
transform 1 0 91264 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_774
timestamp 18001
transform 1 0 96416 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_775
timestamp 18001
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_776
timestamp 18001
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_777
timestamp 18001
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_778
timestamp 18001
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_779
timestamp 18001
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_780
timestamp 18001
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_781
timestamp 18001
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_782
timestamp 18001
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_783
timestamp 18001
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_784
timestamp 18001
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_785
timestamp 18001
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_786
timestamp 18001
transform 1 0 62928 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_787
timestamp 18001
transform 1 0 68080 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_788
timestamp 18001
transform 1 0 73232 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_789
timestamp 18001
transform 1 0 78384 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_790
timestamp 18001
transform 1 0 83536 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_791
timestamp 18001
transform 1 0 88688 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_792
timestamp 18001
transform 1 0 93840 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_793
timestamp 18001
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_794
timestamp 18001
transform 1 0 6256 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_795
timestamp 18001
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_796
timestamp 18001
transform 1 0 11408 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_797
timestamp 18001
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_798
timestamp 18001
transform 1 0 16560 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_799
timestamp 18001
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_800
timestamp 18001
transform 1 0 21712 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_801
timestamp 18001
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_802
timestamp 18001
transform 1 0 26864 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_803
timestamp 18001
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_804
timestamp 18001
transform 1 0 32016 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_805
timestamp 18001
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_806
timestamp 18001
transform 1 0 37168 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_807
timestamp 18001
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_808
timestamp 18001
transform 1 0 42320 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_809
timestamp 18001
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_810
timestamp 18001
transform 1 0 47472 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_811
timestamp 18001
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_812
timestamp 18001
transform 1 0 52624 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_813
timestamp 18001
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_814
timestamp 18001
transform 1 0 57776 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_815
timestamp 18001
transform 1 0 60352 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_816
timestamp 18001
transform 1 0 62928 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_817
timestamp 18001
transform 1 0 65504 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_818
timestamp 18001
transform 1 0 68080 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_819
timestamp 18001
transform 1 0 70656 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_820
timestamp 18001
transform 1 0 73232 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_821
timestamp 18001
transform 1 0 75808 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_822
timestamp 18001
transform 1 0 78384 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_823
timestamp 18001
transform 1 0 80960 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_824
timestamp 18001
transform 1 0 83536 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_825
timestamp 18001
transform 1 0 86112 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_826
timestamp 18001
transform 1 0 88688 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_827
timestamp 18001
transform 1 0 91264 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_828
timestamp 18001
transform 1 0 93840 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_829
timestamp 18001
transform 1 0 96416 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1_830
timestamp 18001
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_3_1040
timestamp 18001
transform 1 0 96600 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_1_831
timestamp 18001
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_3_1041
timestamp 18001
transform 1 0 96600 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_1_832
timestamp 18001
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_3_1042
timestamp 18001
transform 1 0 96600 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_1_833
timestamp 18001
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_3_1043
timestamp 18001
transform 1 0 96600 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_1_834
timestamp 18001
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_3_1044
timestamp 18001
transform 1 0 96600 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_1_835
timestamp 18001
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_3_1045
timestamp 18001
transform 1 0 96600 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_1_836
timestamp 18001
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_3_1046
timestamp 18001
transform 1 0 96600 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_1_837
timestamp 18001
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_3_1047
timestamp 18001
transform 1 0 96600 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_1_838
timestamp 18001
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_3_1048
timestamp 18001
transform 1 0 96600 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_1_839
timestamp 18001
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_3_1049
timestamp 18001
transform 1 0 96600 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_1_840
timestamp 18001
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_3_1050
timestamp 18001
transform 1 0 96600 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_1_841
timestamp 18001
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_3_1051
timestamp 18001
transform 1 0 96600 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_1_842
timestamp 18001
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_3_1052
timestamp 18001
transform 1 0 96600 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_1_843
timestamp 18001
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_3_1053
timestamp 18001
transform 1 0 96600 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_1_844
timestamp 18001
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_3_1054
timestamp 18001
transform 1 0 96600 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_1_845
timestamp 18001
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_3_1055
timestamp 18001
transform 1 0 96600 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_1_846
timestamp 18001
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_3_1056
timestamp 18001
transform 1 0 96600 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_1_847
timestamp 18001
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_3_1057
timestamp 18001
transform 1 0 96600 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_1_848
timestamp 18001
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_3_1058
timestamp 18001
transform 1 0 96600 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_1_849
timestamp 18001
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_3_1059
timestamp 18001
transform 1 0 96600 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_1_850
timestamp 18001
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_3_1060
timestamp 18001
transform 1 0 96600 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_1_851
timestamp 18001
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_3_1061
timestamp 18001
transform 1 0 96600 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_1_852
timestamp 18001
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_3_1062
timestamp 18001
transform 1 0 96600 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_1_853
timestamp 18001
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_3_1063
timestamp 18001
transform 1 0 96600 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_1_854
timestamp 18001
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_3_1064
timestamp 18001
transform 1 0 96600 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_1_855
timestamp 18001
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_3_1065
timestamp 18001
transform 1 0 96600 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1_856
timestamp 18001
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_3_1066
timestamp 18001
transform 1 0 96600 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1_857
timestamp 18001
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_3_1067
timestamp 18001
transform 1 0 96600 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1_858
timestamp 18001
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_3_1068
timestamp 18001
transform 1 0 96600 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_1_859
timestamp 18001
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_3_1069
timestamp 18001
transform 1 0 96600 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_1_860
timestamp 18001
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_3_1070
timestamp 18001
transform 1 0 96600 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_1_861
timestamp 18001
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_3_1071
timestamp 18001
transform 1 0 96600 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1_862
timestamp 18001
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_3_1072
timestamp 18001
transform 1 0 96600 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1_863
timestamp 18001
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_3_1073
timestamp 18001
transform 1 0 96600 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1_864
timestamp 18001
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_3_1074
timestamp 18001
transform 1 0 96600 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1_865
timestamp 18001
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_3_1075
timestamp 18001
transform 1 0 96600 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1_866
timestamp 18001
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_3_1076
timestamp 18001
transform 1 0 96600 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1_867
timestamp 18001
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_3_1077
timestamp 18001
transform 1 0 96600 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1_868
timestamp 18001
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_5_1078
timestamp 18001
transform 1 0 96600 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1_869
timestamp 18001
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_5_1079
timestamp 18001
transform 1 0 96600 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1_870
timestamp 18001
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_5_1080
timestamp 18001
transform 1 0 96600 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1_871
timestamp 18001
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_3_1081
timestamp 18001
transform 1 0 96600 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1_872
timestamp 18001
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_3_1082
timestamp 18001
transform 1 0 96600 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1_873
timestamp 18001
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_3_1083
timestamp 18001
transform 1 0 96600 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1_874
timestamp 18001
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_3_1084
timestamp 18001
transform 1 0 96600 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1_875
timestamp 18001
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_3_1085
timestamp 18001
transform 1 0 96600 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1_876
timestamp 18001
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_3_1086
timestamp 18001
transform 1 0 96600 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_1_877
timestamp 18001
transform 1 0 3680 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_3_1087
timestamp 18001
transform 1 0 96600 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_1_878
timestamp 18001
transform 1 0 3680 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_3_1088
timestamp 18001
transform 1 0 96600 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_1_879
timestamp 18001
transform 1 0 3680 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_3_1089
timestamp 18001
transform 1 0 96600 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_1_880
timestamp 18001
transform 1 0 3680 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_3_1090
timestamp 18001
transform 1 0 96600 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_1_881
timestamp 18001
transform 1 0 3680 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_3_1091
timestamp 18001
transform 1 0 96600 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_1_882
timestamp 18001
transform 1 0 3680 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_3_1092
timestamp 18001
transform 1 0 96600 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_1_883
timestamp 18001
transform 1 0 3680 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_3_1093
timestamp 18001
transform 1 0 96600 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_1_884
timestamp 18001
transform 1 0 3680 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_3_1094
timestamp 18001
transform 1 0 96600 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1_885
timestamp 18001
transform 1 0 3680 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_3_1095
timestamp 18001
transform 1 0 96600 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1_886
timestamp 18001
transform 1 0 3680 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_3_1096
timestamp 18001
transform 1 0 96600 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1_887
timestamp 18001
transform 1 0 3680 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_3_1097
timestamp 18001
transform 1 0 96600 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1_888
timestamp 18001
transform 1 0 3680 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_3_1098
timestamp 18001
transform 1 0 96600 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1_889
timestamp 18001
transform 1 0 3680 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_3_1099
timestamp 18001
transform 1 0 96600 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1_890
timestamp 18001
transform 1 0 3680 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_3_1100
timestamp 18001
transform 1 0 96600 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1_891
timestamp 18001
transform 1 0 3680 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_3_1101
timestamp 18001
transform 1 0 96600 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1_892
timestamp 18001
transform 1 0 3680 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_3_1102
timestamp 18001
transform 1 0 96600 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1_893
timestamp 18001
transform 1 0 3680 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_3_1103
timestamp 18001
transform 1 0 96600 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1_894
timestamp 18001
transform 1 0 3680 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_3_1104
timestamp 18001
transform 1 0 96600 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1_895
timestamp 18001
transform 1 0 3680 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_3_1105
timestamp 18001
transform 1 0 96600 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_140_1_896
timestamp 18001
transform 1 0 3680 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_140_3_1106
timestamp 18001
transform 1 0 96600 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_142_1_897
timestamp 18001
transform 1 0 3680 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_142_3_1107
timestamp 18001
transform 1 0 96600 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_144_1_898
timestamp 18001
transform 1 0 3680 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_144_3_1108
timestamp 18001
transform 1 0 96600 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_1_899
timestamp 18001
transform 1 0 3680 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_3_1109
timestamp 18001
transform 1 0 96600 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_1_900
timestamp 18001
transform 1 0 3680 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_3_1110
timestamp 18001
transform 1 0 96600 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_1_901
timestamp 18001
transform 1 0 3680 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_3_1111
timestamp 18001
transform 1 0 96600 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_1_902
timestamp 18001
transform 1 0 3680 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_3_1112
timestamp 18001
transform 1 0 96600 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_1_903
timestamp 18001
transform 1 0 3680 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_3_1113
timestamp 18001
transform 1 0 96600 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_156_1_904
timestamp 18001
transform 1 0 3680 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_156_3_1114
timestamp 18001
transform 1 0 96600 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_158_1_905
timestamp 18001
transform 1 0 3680 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_158_3_1115
timestamp 18001
transform 1 0 96600 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_160_1_906
timestamp 18001
transform 1 0 3680 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_160_3_1116
timestamp 18001
transform 1 0 96600 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_162_1_907
timestamp 18001
transform 1 0 3680 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_162_3_1117
timestamp 18001
transform 1 0 96600 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_1_908
timestamp 18001
transform 1 0 3680 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_3_1118
timestamp 18001
transform 1 0 96600 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_1_909
timestamp 18001
transform 1 0 3680 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_3_1119
timestamp 18001
transform 1 0 96600 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_910
timestamp 18001
transform 1 0 3680 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_911
timestamp 18001
transform 1 0 6256 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_912
timestamp 18001
transform 1 0 8832 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_913
timestamp 18001
transform 1 0 11408 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_914
timestamp 18001
transform 1 0 13984 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_915
timestamp 18001
transform 1 0 16560 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_916
timestamp 18001
transform 1 0 19136 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_917
timestamp 18001
transform 1 0 21712 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_918
timestamp 18001
transform 1 0 24288 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_919
timestamp 18001
transform 1 0 26864 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_920
timestamp 18001
transform 1 0 29440 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_921
timestamp 18001
transform 1 0 32016 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_922
timestamp 18001
transform 1 0 34592 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_923
timestamp 18001
transform 1 0 37168 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_924
timestamp 18001
transform 1 0 39744 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_925
timestamp 18001
transform 1 0 42320 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_926
timestamp 18001
transform 1 0 44896 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_927
timestamp 18001
transform 1 0 47472 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_928
timestamp 18001
transform 1 0 50048 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_929
timestamp 18001
transform 1 0 52624 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_930
timestamp 18001
transform 1 0 55200 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_931
timestamp 18001
transform 1 0 57776 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_932
timestamp 18001
transform 1 0 60352 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_933
timestamp 18001
transform 1 0 62928 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_934
timestamp 18001
transform 1 0 65504 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_935
timestamp 18001
transform 1 0 68080 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_936
timestamp 18001
transform 1 0 70656 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_937
timestamp 18001
transform 1 0 73232 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_938
timestamp 18001
transform 1 0 75808 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_939
timestamp 18001
transform 1 0 78384 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_940
timestamp 18001
transform 1 0 80960 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_941
timestamp 18001
transform 1 0 83536 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_942
timestamp 18001
transform 1 0 86112 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_943
timestamp 18001
transform 1 0 88688 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_944
timestamp 18001
transform 1 0 91264 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_945
timestamp 18001
transform 1 0 93840 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_946
timestamp 18001
transform 1 0 96416 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_947
timestamp 18001
transform 1 0 3680 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_948
timestamp 18001
transform 1 0 8832 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_949
timestamp 18001
transform 1 0 13984 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_950
timestamp 18001
transform 1 0 19136 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_951
timestamp 18001
transform 1 0 24288 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_952
timestamp 18001
transform 1 0 29440 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_953
timestamp 18001
transform 1 0 34592 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_954
timestamp 18001
transform 1 0 39744 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_955
timestamp 18001
transform 1 0 44896 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_956
timestamp 18001
transform 1 0 50048 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_957
timestamp 18001
transform 1 0 55200 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_958
timestamp 18001
transform 1 0 60352 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_959
timestamp 18001
transform 1 0 65504 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_960
timestamp 18001
transform 1 0 70656 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_961
timestamp 18001
transform 1 0 75808 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_962
timestamp 18001
transform 1 0 80960 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_963
timestamp 18001
transform 1 0 86112 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_964
timestamp 18001
transform 1 0 91264 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_965
timestamp 18001
transform 1 0 96416 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_966
timestamp 18001
transform 1 0 6256 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_967
timestamp 18001
transform 1 0 11408 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_968
timestamp 18001
transform 1 0 16560 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_969
timestamp 18001
transform 1 0 21712 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_970
timestamp 18001
transform 1 0 26864 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_971
timestamp 18001
transform 1 0 32016 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_972
timestamp 18001
transform 1 0 37168 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_973
timestamp 18001
transform 1 0 42320 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_974
timestamp 18001
transform 1 0 47472 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_975
timestamp 18001
transform 1 0 52624 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_976
timestamp 18001
transform 1 0 57776 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_977
timestamp 18001
transform 1 0 62928 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_978
timestamp 18001
transform 1 0 68080 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_979
timestamp 18001
transform 1 0 73232 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_980
timestamp 18001
transform 1 0 78384 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_981
timestamp 18001
transform 1 0 83536 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_982
timestamp 18001
transform 1 0 88688 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_983
timestamp 18001
transform 1 0 93840 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_984
timestamp 18001
transform 1 0 3680 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_985
timestamp 18001
transform 1 0 8832 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_986
timestamp 18001
transform 1 0 13984 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_987
timestamp 18001
transform 1 0 19136 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_988
timestamp 18001
transform 1 0 24288 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_989
timestamp 18001
transform 1 0 29440 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_990
timestamp 18001
transform 1 0 34592 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_991
timestamp 18001
transform 1 0 39744 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_992
timestamp 18001
transform 1 0 44896 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_993
timestamp 18001
transform 1 0 50048 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_994
timestamp 18001
transform 1 0 55200 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_995
timestamp 18001
transform 1 0 60352 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_996
timestamp 18001
transform 1 0 65504 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_997
timestamp 18001
transform 1 0 70656 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_998
timestamp 18001
transform 1 0 75808 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_999
timestamp 18001
transform 1 0 80960 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_1000
timestamp 18001
transform 1 0 86112 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_1001
timestamp 18001
transform 1 0 91264 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_1002
timestamp 18001
transform 1 0 96416 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1003
timestamp 18001
transform 1 0 3680 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1004
timestamp 18001
transform 1 0 6256 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1005
timestamp 18001
transform 1 0 8832 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1006
timestamp 18001
transform 1 0 11408 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1007
timestamp 18001
transform 1 0 13984 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1008
timestamp 18001
transform 1 0 16560 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1009
timestamp 18001
transform 1 0 19136 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1010
timestamp 18001
transform 1 0 21712 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1011
timestamp 18001
transform 1 0 24288 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1012
timestamp 18001
transform 1 0 26864 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1013
timestamp 18001
transform 1 0 29440 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1014
timestamp 18001
transform 1 0 32016 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1015
timestamp 18001
transform 1 0 34592 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1016
timestamp 18001
transform 1 0 37168 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1017
timestamp 18001
transform 1 0 39744 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1018
timestamp 18001
transform 1 0 42320 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1019
timestamp 18001
transform 1 0 44896 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1020
timestamp 18001
transform 1 0 47472 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1021
timestamp 18001
transform 1 0 50048 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1022
timestamp 18001
transform 1 0 52624 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1023
timestamp 18001
transform 1 0 55200 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1024
timestamp 18001
transform 1 0 57776 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1025
timestamp 18001
transform 1 0 60352 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1026
timestamp 18001
transform 1 0 62928 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1027
timestamp 18001
transform 1 0 65504 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1028
timestamp 18001
transform 1 0 68080 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1029
timestamp 18001
transform 1 0 70656 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1030
timestamp 18001
transform 1 0 73232 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1031
timestamp 18001
transform 1 0 75808 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1032
timestamp 18001
transform 1 0 78384 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1033
timestamp 18001
transform 1 0 80960 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1034
timestamp 18001
transform 1 0 83536 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1035
timestamp 18001
transform 1 0 86112 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1036
timestamp 18001
transform 1 0 88688 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1037
timestamp 18001
transform 1 0 91264 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1038
timestamp 18001
transform 1 0 93840 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1039
timestamp 18001
transform 1 0 96416 0 -1 95744
box -38 -48 130 592
<< labels >>
flabel metal2 s 50250 97200 50306 98000 0 FreeSans 224 90 0 0 clk
port 0 nsew signal input
flabel metal3 s 0 48288 800 48408 0 FreeSans 480 0 0 0 config_data_in
port 1 nsew signal input
flabel metal2 s 50894 97200 50950 98000 0 FreeSans 224 90 0 0 config_data_out
port 2 nsew signal output
flabel metal2 s 54114 97200 54170 98000 0 FreeSans 224 90 0 0 config_en
port 3 nsew signal input
flabel metal2 s 51538 97200 51594 98000 0 FreeSans 224 90 0 0 en
port 4 nsew signal input
flabel metal3 s 98200 29248 99000 29368 0 FreeSans 480 0 0 0 io_east_in[0]
port 5 nsew signal input
flabel metal3 s 98200 40128 99000 40248 0 FreeSans 480 0 0 0 io_east_in[10]
port 6 nsew signal input
flabel metal3 s 98200 40808 99000 40928 0 FreeSans 480 0 0 0 io_east_in[11]
port 7 nsew signal input
flabel metal3 s 98200 42168 99000 42288 0 FreeSans 480 0 0 0 io_east_in[12]
port 8 nsew signal input
flabel metal3 s 98200 42848 99000 42968 0 FreeSans 480 0 0 0 io_east_in[13]
port 9 nsew signal input
flabel metal3 s 98200 44208 99000 44328 0 FreeSans 480 0 0 0 io_east_in[14]
port 10 nsew signal input
flabel metal3 s 98200 45568 99000 45688 0 FreeSans 480 0 0 0 io_east_in[15]
port 11 nsew signal input
flabel metal3 s 98200 70728 99000 70848 0 FreeSans 480 0 0 0 io_east_in[16]
port 12 nsew signal input
flabel metal3 s 98200 72088 99000 72208 0 FreeSans 480 0 0 0 io_east_in[17]
port 13 nsew signal input
flabel metal3 s 98200 73448 99000 73568 0 FreeSans 480 0 0 0 io_east_in[18]
port 14 nsew signal input
flabel metal3 s 98200 74128 99000 74248 0 FreeSans 480 0 0 0 io_east_in[19]
port 15 nsew signal input
flabel metal3 s 98200 29928 99000 30048 0 FreeSans 480 0 0 0 io_east_in[1]
port 16 nsew signal input
flabel metal3 s 98200 75488 99000 75608 0 FreeSans 480 0 0 0 io_east_in[20]
port 17 nsew signal input
flabel metal3 s 98200 76168 99000 76288 0 FreeSans 480 0 0 0 io_east_in[21]
port 18 nsew signal input
flabel metal3 s 98200 77528 99000 77648 0 FreeSans 480 0 0 0 io_east_in[22]
port 19 nsew signal input
flabel metal3 s 98200 78888 99000 79008 0 FreeSans 480 0 0 0 io_east_in[23]
port 20 nsew signal input
flabel metal3 s 98200 79568 99000 79688 0 FreeSans 480 0 0 0 io_east_in[24]
port 21 nsew signal input
flabel metal3 s 98200 80928 99000 81048 0 FreeSans 480 0 0 0 io_east_in[25]
port 22 nsew signal input
flabel metal3 s 98200 81608 99000 81728 0 FreeSans 480 0 0 0 io_east_in[26]
port 23 nsew signal input
flabel metal3 s 98200 82968 99000 83088 0 FreeSans 480 0 0 0 io_east_in[27]
port 24 nsew signal input
flabel metal3 s 98200 84328 99000 84448 0 FreeSans 480 0 0 0 io_east_in[28]
port 25 nsew signal input
flabel metal3 s 98200 85008 99000 85128 0 FreeSans 480 0 0 0 io_east_in[29]
port 26 nsew signal input
flabel metal3 s 98200 31288 99000 31408 0 FreeSans 480 0 0 0 io_east_in[2]
port 27 nsew signal input
flabel metal3 s 98200 86368 99000 86488 0 FreeSans 480 0 0 0 io_east_in[30]
port 28 nsew signal input
flabel metal3 s 98200 87048 99000 87168 0 FreeSans 480 0 0 0 io_east_in[31]
port 29 nsew signal input
flabel metal3 s 98200 31968 99000 32088 0 FreeSans 480 0 0 0 io_east_in[3]
port 30 nsew signal input
flabel metal3 s 98200 33328 99000 33448 0 FreeSans 480 0 0 0 io_east_in[4]
port 31 nsew signal input
flabel metal3 s 98200 34688 99000 34808 0 FreeSans 480 0 0 0 io_east_in[5]
port 32 nsew signal input
flabel metal3 s 98200 35368 99000 35488 0 FreeSans 480 0 0 0 io_east_in[6]
port 33 nsew signal input
flabel metal3 s 98200 36728 99000 36848 0 FreeSans 480 0 0 0 io_east_in[7]
port 34 nsew signal input
flabel metal3 s 98200 37408 99000 37528 0 FreeSans 480 0 0 0 io_east_in[8]
port 35 nsew signal input
flabel metal3 s 98200 38768 99000 38888 0 FreeSans 480 0 0 0 io_east_in[9]
port 36 nsew signal input
flabel metal3 s 98200 11568 99000 11688 0 FreeSans 480 0 0 0 io_east_out[0]
port 37 nsew signal output
flabel metal3 s 98200 22448 99000 22568 0 FreeSans 480 0 0 0 io_east_out[10]
port 38 nsew signal output
flabel metal3 s 98200 23808 99000 23928 0 FreeSans 480 0 0 0 io_east_out[11]
port 39 nsew signal output
flabel metal3 s 98200 24488 99000 24608 0 FreeSans 480 0 0 0 io_east_out[12]
port 40 nsew signal output
flabel metal3 s 98200 25848 99000 25968 0 FreeSans 480 0 0 0 io_east_out[13]
port 41 nsew signal output
flabel metal3 s 98200 26528 99000 26648 0 FreeSans 480 0 0 0 io_east_out[14]
port 42 nsew signal output
flabel metal3 s 98200 27888 99000 28008 0 FreeSans 480 0 0 0 io_east_out[15]
port 43 nsew signal output
flabel metal3 s 98200 53728 99000 53848 0 FreeSans 480 0 0 0 io_east_out[16]
port 44 nsew signal output
flabel metal3 s 98200 54408 99000 54528 0 FreeSans 480 0 0 0 io_east_out[17]
port 45 nsew signal output
flabel metal3 s 98200 55768 99000 55888 0 FreeSans 480 0 0 0 io_east_out[18]
port 46 nsew signal output
flabel metal3 s 98200 57128 99000 57248 0 FreeSans 480 0 0 0 io_east_out[19]
port 47 nsew signal output
flabel metal3 s 98200 12928 99000 13048 0 FreeSans 480 0 0 0 io_east_out[1]
port 48 nsew signal output
flabel metal3 s 98200 57808 99000 57928 0 FreeSans 480 0 0 0 io_east_out[20]
port 49 nsew signal output
flabel metal3 s 98200 59168 99000 59288 0 FreeSans 480 0 0 0 io_east_out[21]
port 50 nsew signal output
flabel metal3 s 98200 59848 99000 59968 0 FreeSans 480 0 0 0 io_east_out[22]
port 51 nsew signal output
flabel metal3 s 98200 61208 99000 61328 0 FreeSans 480 0 0 0 io_east_out[23]
port 52 nsew signal output
flabel metal3 s 98200 62568 99000 62688 0 FreeSans 480 0 0 0 io_east_out[24]
port 53 nsew signal output
flabel metal3 s 98200 63248 99000 63368 0 FreeSans 480 0 0 0 io_east_out[25]
port 54 nsew signal output
flabel metal3 s 98200 64608 99000 64728 0 FreeSans 480 0 0 0 io_east_out[26]
port 55 nsew signal output
flabel metal3 s 98200 65288 99000 65408 0 FreeSans 480 0 0 0 io_east_out[27]
port 56 nsew signal output
flabel metal3 s 98200 66648 99000 66768 0 FreeSans 480 0 0 0 io_east_out[28]
port 57 nsew signal output
flabel metal3 s 98200 68008 99000 68128 0 FreeSans 480 0 0 0 io_east_out[29]
port 58 nsew signal output
flabel metal3 s 98200 13608 99000 13728 0 FreeSans 480 0 0 0 io_east_out[2]
port 59 nsew signal output
flabel metal3 s 98200 68688 99000 68808 0 FreeSans 480 0 0 0 io_east_out[30]
port 60 nsew signal output
flabel metal3 s 98200 70048 99000 70168 0 FreeSans 480 0 0 0 io_east_out[31]
port 61 nsew signal output
flabel metal3 s 98200 14968 99000 15088 0 FreeSans 480 0 0 0 io_east_out[3]
port 62 nsew signal output
flabel metal3 s 98200 15648 99000 15768 0 FreeSans 480 0 0 0 io_east_out[4]
port 63 nsew signal output
flabel metal3 s 98200 17008 99000 17128 0 FreeSans 480 0 0 0 io_east_out[5]
port 64 nsew signal output
flabel metal3 s 98200 18368 99000 18488 0 FreeSans 480 0 0 0 io_east_out[6]
port 65 nsew signal output
flabel metal3 s 98200 19048 99000 19168 0 FreeSans 480 0 0 0 io_east_out[7]
port 66 nsew signal output
flabel metal3 s 98200 20408 99000 20528 0 FreeSans 480 0 0 0 io_east_out[8]
port 67 nsew signal output
flabel metal3 s 98200 21088 99000 21208 0 FreeSans 480 0 0 0 io_east_out[9]
port 68 nsew signal output
flabel metal2 s 14186 97200 14242 98000 0 FreeSans 224 90 0 0 io_north_in[0]
port 69 nsew signal input
flabel metal2 s 25134 97200 25190 98000 0 FreeSans 224 90 0 0 io_north_in[10]
port 70 nsew signal input
flabel metal2 s 26422 97200 26478 98000 0 FreeSans 224 90 0 0 io_north_in[11]
port 71 nsew signal input
flabel metal2 s 27710 97200 27766 98000 0 FreeSans 224 90 0 0 io_north_in[12]
port 72 nsew signal input
flabel metal2 s 28998 97200 29054 98000 0 FreeSans 224 90 0 0 io_north_in[13]
port 73 nsew signal input
flabel metal2 s 29642 97200 29698 98000 0 FreeSans 224 90 0 0 io_north_in[14]
port 74 nsew signal input
flabel metal2 s 30930 97200 30986 98000 0 FreeSans 224 90 0 0 io_north_in[15]
port 75 nsew signal input
flabel metal2 s 56046 97200 56102 98000 0 FreeSans 224 90 0 0 io_north_in[16]
port 76 nsew signal input
flabel metal2 s 57334 97200 57390 98000 0 FreeSans 224 90 0 0 io_north_in[17]
port 77 nsew signal input
flabel metal2 s 58622 97200 58678 98000 0 FreeSans 224 90 0 0 io_north_in[18]
port 78 nsew signal input
flabel metal2 s 59910 97200 59966 98000 0 FreeSans 224 90 0 0 io_north_in[19]
port 79 nsew signal input
flabel metal2 s 15474 97200 15530 98000 0 FreeSans 224 90 0 0 io_north_in[1]
port 80 nsew signal input
flabel metal2 s 60554 97200 60610 98000 0 FreeSans 224 90 0 0 io_north_in[20]
port 81 nsew signal input
flabel metal2 s 61842 97200 61898 98000 0 FreeSans 224 90 0 0 io_north_in[21]
port 82 nsew signal input
flabel metal2 s 63130 97200 63186 98000 0 FreeSans 224 90 0 0 io_north_in[22]
port 83 nsew signal input
flabel metal2 s 63774 97200 63830 98000 0 FreeSans 224 90 0 0 io_north_in[23]
port 84 nsew signal input
flabel metal2 s 65062 97200 65118 98000 0 FreeSans 224 90 0 0 io_north_in[24]
port 85 nsew signal input
flabel metal2 s 66350 97200 66406 98000 0 FreeSans 224 90 0 0 io_north_in[25]
port 86 nsew signal input
flabel metal2 s 67638 97200 67694 98000 0 FreeSans 224 90 0 0 io_north_in[26]
port 87 nsew signal input
flabel metal2 s 68282 97200 68338 98000 0 FreeSans 224 90 0 0 io_north_in[27]
port 88 nsew signal input
flabel metal2 s 69570 97200 69626 98000 0 FreeSans 224 90 0 0 io_north_in[28]
port 89 nsew signal input
flabel metal2 s 70858 97200 70914 98000 0 FreeSans 224 90 0 0 io_north_in[29]
port 90 nsew signal input
flabel metal2 s 16762 97200 16818 98000 0 FreeSans 224 90 0 0 io_north_in[2]
port 91 nsew signal input
flabel metal2 s 71502 97200 71558 98000 0 FreeSans 224 90 0 0 io_north_in[30]
port 92 nsew signal input
flabel metal2 s 72790 97200 72846 98000 0 FreeSans 224 90 0 0 io_north_in[31]
port 93 nsew signal input
flabel metal2 s 17406 97200 17462 98000 0 FreeSans 224 90 0 0 io_north_in[3]
port 94 nsew signal input
flabel metal2 s 18694 97200 18750 98000 0 FreeSans 224 90 0 0 io_north_in[4]
port 95 nsew signal input
flabel metal2 s 19982 97200 20038 98000 0 FreeSans 224 90 0 0 io_north_in[5]
port 96 nsew signal input
flabel metal2 s 21270 97200 21326 98000 0 FreeSans 224 90 0 0 io_north_in[6]
port 97 nsew signal input
flabel metal2 s 21914 97200 21970 98000 0 FreeSans 224 90 0 0 io_north_in[7]
port 98 nsew signal input
flabel metal2 s 23202 97200 23258 98000 0 FreeSans 224 90 0 0 io_north_in[8]
port 99 nsew signal input
flabel metal2 s 24490 97200 24546 98000 0 FreeSans 224 90 0 0 io_north_in[9]
port 100 nsew signal input
flabel metal2 s 32218 97200 32274 98000 0 FreeSans 224 90 0 0 io_north_out[0]
port 101 nsew signal output
flabel metal2 s 43166 97200 43222 98000 0 FreeSans 224 90 0 0 io_north_out[10]
port 102 nsew signal output
flabel metal2 s 44454 97200 44510 98000 0 FreeSans 224 90 0 0 io_north_out[11]
port 103 nsew signal output
flabel metal2 s 45098 97200 45154 98000 0 FreeSans 224 90 0 0 io_north_out[12]
port 104 nsew signal output
flabel metal2 s 46386 97200 46442 98000 0 FreeSans 224 90 0 0 io_north_out[13]
port 105 nsew signal output
flabel metal2 s 47674 97200 47730 98000 0 FreeSans 224 90 0 0 io_north_out[14]
port 106 nsew signal output
flabel metal2 s 48318 97200 48374 98000 0 FreeSans 224 90 0 0 io_north_out[15]
port 107 nsew signal output
flabel metal2 s 74078 97200 74134 98000 0 FreeSans 224 90 0 0 io_north_out[16]
port 108 nsew signal output
flabel metal2 s 75366 97200 75422 98000 0 FreeSans 224 90 0 0 io_north_out[17]
port 109 nsew signal output
flabel metal2 s 76010 97200 76066 98000 0 FreeSans 224 90 0 0 io_north_out[18]
port 110 nsew signal output
flabel metal2 s 77298 97200 77354 98000 0 FreeSans 224 90 0 0 io_north_out[19]
port 111 nsew signal output
flabel metal2 s 32862 97200 32918 98000 0 FreeSans 224 90 0 0 io_north_out[1]
port 112 nsew signal output
flabel metal2 s 78586 97200 78642 98000 0 FreeSans 224 90 0 0 io_north_out[20]
port 113 nsew signal output
flabel metal2 s 79230 97200 79286 98000 0 FreeSans 224 90 0 0 io_north_out[21]
port 114 nsew signal output
flabel metal2 s 80518 97200 80574 98000 0 FreeSans 224 90 0 0 io_north_out[22]
port 115 nsew signal output
flabel metal2 s 81806 97200 81862 98000 0 FreeSans 224 90 0 0 io_north_out[23]
port 116 nsew signal output
flabel metal2 s 83094 97200 83150 98000 0 FreeSans 224 90 0 0 io_north_out[24]
port 117 nsew signal output
flabel metal2 s 83738 97200 83794 98000 0 FreeSans 224 90 0 0 io_north_out[25]
port 118 nsew signal output
flabel metal2 s 85026 97200 85082 98000 0 FreeSans 224 90 0 0 io_north_out[26]
port 119 nsew signal output
flabel metal2 s 86314 97200 86370 98000 0 FreeSans 224 90 0 0 io_north_out[27]
port 120 nsew signal output
flabel metal2 s 86958 97200 87014 98000 0 FreeSans 224 90 0 0 io_north_out[28]
port 121 nsew signal output
flabel metal2 s 88246 97200 88302 98000 0 FreeSans 224 90 0 0 io_north_out[29]
port 122 nsew signal output
flabel metal2 s 34150 97200 34206 98000 0 FreeSans 224 90 0 0 io_north_out[2]
port 123 nsew signal output
flabel metal2 s 89534 97200 89590 98000 0 FreeSans 224 90 0 0 io_north_out[30]
port 124 nsew signal output
flabel metal2 s 90822 97200 90878 98000 0 FreeSans 224 90 0 0 io_north_out[31]
port 125 nsew signal output
flabel metal2 s 35438 97200 35494 98000 0 FreeSans 224 90 0 0 io_north_out[3]
port 126 nsew signal output
flabel metal2 s 36726 97200 36782 98000 0 FreeSans 224 90 0 0 io_north_out[4]
port 127 nsew signal output
flabel metal2 s 37370 97200 37426 98000 0 FreeSans 224 90 0 0 io_north_out[5]
port 128 nsew signal output
flabel metal2 s 38658 97200 38714 98000 0 FreeSans 224 90 0 0 io_north_out[6]
port 129 nsew signal output
flabel metal2 s 39946 97200 40002 98000 0 FreeSans 224 90 0 0 io_north_out[7]
port 130 nsew signal output
flabel metal2 s 40590 97200 40646 98000 0 FreeSans 224 90 0 0 io_north_out[8]
port 131 nsew signal output
flabel metal2 s 41878 97200 41934 98000 0 FreeSans 224 90 0 0 io_north_out[9]
port 132 nsew signal output
flabel metal2 s 32218 0 32274 800 0 FreeSans 224 90 0 0 io_south_in[0]
port 133 nsew signal input
flabel metal2 s 43166 0 43222 800 0 FreeSans 224 90 0 0 io_south_in[10]
port 134 nsew signal input
flabel metal2 s 44454 0 44510 800 0 FreeSans 224 90 0 0 io_south_in[11]
port 135 nsew signal input
flabel metal2 s 45098 0 45154 800 0 FreeSans 224 90 0 0 io_south_in[12]
port 136 nsew signal input
flabel metal2 s 46386 0 46442 800 0 FreeSans 224 90 0 0 io_south_in[13]
port 137 nsew signal input
flabel metal2 s 47674 0 47730 800 0 FreeSans 224 90 0 0 io_south_in[14]
port 138 nsew signal input
flabel metal2 s 48318 0 48374 800 0 FreeSans 224 90 0 0 io_south_in[15]
port 139 nsew signal input
flabel metal2 s 74078 0 74134 800 0 FreeSans 224 90 0 0 io_south_in[16]
port 140 nsew signal input
flabel metal2 s 75366 0 75422 800 0 FreeSans 224 90 0 0 io_south_in[17]
port 141 nsew signal input
flabel metal2 s 76010 0 76066 800 0 FreeSans 224 90 0 0 io_south_in[18]
port 142 nsew signal input
flabel metal2 s 77298 0 77354 800 0 FreeSans 224 90 0 0 io_south_in[19]
port 143 nsew signal input
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 io_south_in[1]
port 144 nsew signal input
flabel metal2 s 78586 0 78642 800 0 FreeSans 224 90 0 0 io_south_in[20]
port 145 nsew signal input
flabel metal2 s 79230 0 79286 800 0 FreeSans 224 90 0 0 io_south_in[21]
port 146 nsew signal input
flabel metal2 s 80518 0 80574 800 0 FreeSans 224 90 0 0 io_south_in[22]
port 147 nsew signal input
flabel metal2 s 81806 0 81862 800 0 FreeSans 224 90 0 0 io_south_in[23]
port 148 nsew signal input
flabel metal2 s 83094 0 83150 800 0 FreeSans 224 90 0 0 io_south_in[24]
port 149 nsew signal input
flabel metal2 s 83738 0 83794 800 0 FreeSans 224 90 0 0 io_south_in[25]
port 150 nsew signal input
flabel metal2 s 85026 0 85082 800 0 FreeSans 224 90 0 0 io_south_in[26]
port 151 nsew signal input
flabel metal2 s 86314 0 86370 800 0 FreeSans 224 90 0 0 io_south_in[27]
port 152 nsew signal input
flabel metal2 s 86958 0 87014 800 0 FreeSans 224 90 0 0 io_south_in[28]
port 153 nsew signal input
flabel metal2 s 88246 0 88302 800 0 FreeSans 224 90 0 0 io_south_in[29]
port 154 nsew signal input
flabel metal2 s 34150 0 34206 800 0 FreeSans 224 90 0 0 io_south_in[2]
port 155 nsew signal input
flabel metal2 s 89534 0 89590 800 0 FreeSans 224 90 0 0 io_south_in[30]
port 156 nsew signal input
flabel metal3 s 98200 8168 99000 8288 0 FreeSans 480 0 0 0 io_south_in[31]
port 157 nsew signal input
flabel metal2 s 35438 0 35494 800 0 FreeSans 224 90 0 0 io_south_in[3]
port 158 nsew signal input
flabel metal2 s 36726 0 36782 800 0 FreeSans 224 90 0 0 io_south_in[4]
port 159 nsew signal input
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 io_south_in[5]
port 160 nsew signal input
flabel metal2 s 38658 0 38714 800 0 FreeSans 224 90 0 0 io_south_in[6]
port 161 nsew signal input
flabel metal2 s 39946 0 40002 800 0 FreeSans 224 90 0 0 io_south_in[7]
port 162 nsew signal input
flabel metal2 s 40590 0 40646 800 0 FreeSans 224 90 0 0 io_south_in[8]
port 163 nsew signal input
flabel metal2 s 41878 0 41934 800 0 FreeSans 224 90 0 0 io_south_in[9]
port 164 nsew signal input
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 io_south_out[0]
port 165 nsew signal output
flabel metal2 s 25134 0 25190 800 0 FreeSans 224 90 0 0 io_south_out[10]
port 166 nsew signal output
flabel metal2 s 26422 0 26478 800 0 FreeSans 224 90 0 0 io_south_out[11]
port 167 nsew signal output
flabel metal2 s 27710 0 27766 800 0 FreeSans 224 90 0 0 io_south_out[12]
port 168 nsew signal output
flabel metal2 s 28998 0 29054 800 0 FreeSans 224 90 0 0 io_south_out[13]
port 169 nsew signal output
flabel metal2 s 29642 0 29698 800 0 FreeSans 224 90 0 0 io_south_out[14]
port 170 nsew signal output
flabel metal2 s 30930 0 30986 800 0 FreeSans 224 90 0 0 io_south_out[15]
port 171 nsew signal output
flabel metal2 s 56046 0 56102 800 0 FreeSans 224 90 0 0 io_south_out[16]
port 172 nsew signal output
flabel metal2 s 57334 0 57390 800 0 FreeSans 224 90 0 0 io_south_out[17]
port 173 nsew signal output
flabel metal2 s 58622 0 58678 800 0 FreeSans 224 90 0 0 io_south_out[18]
port 174 nsew signal output
flabel metal2 s 59910 0 59966 800 0 FreeSans 224 90 0 0 io_south_out[19]
port 175 nsew signal output
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 io_south_out[1]
port 176 nsew signal output
flabel metal2 s 60554 0 60610 800 0 FreeSans 224 90 0 0 io_south_out[20]
port 177 nsew signal output
flabel metal2 s 61842 0 61898 800 0 FreeSans 224 90 0 0 io_south_out[21]
port 178 nsew signal output
flabel metal2 s 63130 0 63186 800 0 FreeSans 224 90 0 0 io_south_out[22]
port 179 nsew signal output
flabel metal2 s 63774 0 63830 800 0 FreeSans 224 90 0 0 io_south_out[23]
port 180 nsew signal output
flabel metal2 s 65062 0 65118 800 0 FreeSans 224 90 0 0 io_south_out[24]
port 181 nsew signal output
flabel metal2 s 66350 0 66406 800 0 FreeSans 224 90 0 0 io_south_out[25]
port 182 nsew signal output
flabel metal2 s 67638 0 67694 800 0 FreeSans 224 90 0 0 io_south_out[26]
port 183 nsew signal output
flabel metal2 s 68282 0 68338 800 0 FreeSans 224 90 0 0 io_south_out[27]
port 184 nsew signal output
flabel metal2 s 69570 0 69626 800 0 FreeSans 224 90 0 0 io_south_out[28]
port 185 nsew signal output
flabel metal2 s 70858 0 70914 800 0 FreeSans 224 90 0 0 io_south_out[29]
port 186 nsew signal output
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 io_south_out[2]
port 187 nsew signal output
flabel metal2 s 71502 0 71558 800 0 FreeSans 224 90 0 0 io_south_out[30]
port 188 nsew signal output
flabel metal2 s 72790 0 72846 800 0 FreeSans 224 90 0 0 io_south_out[31]
port 189 nsew signal output
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 io_south_out[3]
port 190 nsew signal output
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 io_south_out[4]
port 191 nsew signal output
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 io_south_out[5]
port 192 nsew signal output
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 io_south_out[6]
port 193 nsew signal output
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 io_south_out[7]
port 194 nsew signal output
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 io_south_out[8]
port 195 nsew signal output
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 io_south_out[9]
port 196 nsew signal output
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 io_west_in[0]
port 197 nsew signal input
flabel metal3 s 0 22448 800 22568 0 FreeSans 480 0 0 0 io_west_in[10]
port 198 nsew signal input
flabel metal3 s 0 23808 800 23928 0 FreeSans 480 0 0 0 io_west_in[11]
port 199 nsew signal input
flabel metal3 s 0 24488 800 24608 0 FreeSans 480 0 0 0 io_west_in[12]
port 200 nsew signal input
flabel metal3 s 0 25848 800 25968 0 FreeSans 480 0 0 0 io_west_in[13]
port 201 nsew signal input
flabel metal3 s 0 26528 800 26648 0 FreeSans 480 0 0 0 io_west_in[14]
port 202 nsew signal input
flabel metal3 s 0 27888 800 28008 0 FreeSans 480 0 0 0 io_west_in[15]
port 203 nsew signal input
flabel metal3 s 0 53728 800 53848 0 FreeSans 480 0 0 0 io_west_in[16]
port 204 nsew signal input
flabel metal3 s 0 54408 800 54528 0 FreeSans 480 0 0 0 io_west_in[17]
port 205 nsew signal input
flabel metal3 s 0 55768 800 55888 0 FreeSans 480 0 0 0 io_west_in[18]
port 206 nsew signal input
flabel metal3 s 0 57128 800 57248 0 FreeSans 480 0 0 0 io_west_in[19]
port 207 nsew signal input
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 io_west_in[1]
port 208 nsew signal input
flabel metal3 s 0 57808 800 57928 0 FreeSans 480 0 0 0 io_west_in[20]
port 209 nsew signal input
flabel metal3 s 0 59168 800 59288 0 FreeSans 480 0 0 0 io_west_in[21]
port 210 nsew signal input
flabel metal3 s 0 59848 800 59968 0 FreeSans 480 0 0 0 io_west_in[22]
port 211 nsew signal input
flabel metal3 s 0 61208 800 61328 0 FreeSans 480 0 0 0 io_west_in[23]
port 212 nsew signal input
flabel metal3 s 0 62568 800 62688 0 FreeSans 480 0 0 0 io_west_in[24]
port 213 nsew signal input
flabel metal3 s 0 63248 800 63368 0 FreeSans 480 0 0 0 io_west_in[25]
port 214 nsew signal input
flabel metal3 s 0 64608 800 64728 0 FreeSans 480 0 0 0 io_west_in[26]
port 215 nsew signal input
flabel metal3 s 0 65288 800 65408 0 FreeSans 480 0 0 0 io_west_in[27]
port 216 nsew signal input
flabel metal3 s 0 66648 800 66768 0 FreeSans 480 0 0 0 io_west_in[28]
port 217 nsew signal input
flabel metal3 s 0 68008 800 68128 0 FreeSans 480 0 0 0 io_west_in[29]
port 218 nsew signal input
flabel metal3 s 0 13608 800 13728 0 FreeSans 480 0 0 0 io_west_in[2]
port 219 nsew signal input
flabel metal3 s 0 68688 800 68808 0 FreeSans 480 0 0 0 io_west_in[30]
port 220 nsew signal input
flabel metal3 s 0 70048 800 70168 0 FreeSans 480 0 0 0 io_west_in[31]
port 221 nsew signal input
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 io_west_in[3]
port 222 nsew signal input
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 io_west_in[4]
port 223 nsew signal input
flabel metal3 s 0 17008 800 17128 0 FreeSans 480 0 0 0 io_west_in[5]
port 224 nsew signal input
flabel metal3 s 0 18368 800 18488 0 FreeSans 480 0 0 0 io_west_in[6]
port 225 nsew signal input
flabel metal3 s 0 19048 800 19168 0 FreeSans 480 0 0 0 io_west_in[7]
port 226 nsew signal input
flabel metal3 s 0 20408 800 20528 0 FreeSans 480 0 0 0 io_west_in[8]
port 227 nsew signal input
flabel metal3 s 0 21088 800 21208 0 FreeSans 480 0 0 0 io_west_in[9]
port 228 nsew signal input
flabel metal3 s 0 29248 800 29368 0 FreeSans 480 0 0 0 io_west_out[0]
port 229 nsew signal output
flabel metal3 s 0 40128 800 40248 0 FreeSans 480 0 0 0 io_west_out[10]
port 230 nsew signal output
flabel metal3 s 0 40808 800 40928 0 FreeSans 480 0 0 0 io_west_out[11]
port 231 nsew signal output
flabel metal3 s 0 42168 800 42288 0 FreeSans 480 0 0 0 io_west_out[12]
port 232 nsew signal output
flabel metal3 s 0 42848 800 42968 0 FreeSans 480 0 0 0 io_west_out[13]
port 233 nsew signal output
flabel metal3 s 0 44208 800 44328 0 FreeSans 480 0 0 0 io_west_out[14]
port 234 nsew signal output
flabel metal3 s 0 45568 800 45688 0 FreeSans 480 0 0 0 io_west_out[15]
port 235 nsew signal output
flabel metal3 s 0 70728 800 70848 0 FreeSans 480 0 0 0 io_west_out[16]
port 236 nsew signal output
flabel metal3 s 0 72088 800 72208 0 FreeSans 480 0 0 0 io_west_out[17]
port 237 nsew signal output
flabel metal3 s 0 73448 800 73568 0 FreeSans 480 0 0 0 io_west_out[18]
port 238 nsew signal output
flabel metal3 s 0 74128 800 74248 0 FreeSans 480 0 0 0 io_west_out[19]
port 239 nsew signal output
flabel metal3 s 0 29928 800 30048 0 FreeSans 480 0 0 0 io_west_out[1]
port 240 nsew signal output
flabel metal3 s 0 75488 800 75608 0 FreeSans 480 0 0 0 io_west_out[20]
port 241 nsew signal output
flabel metal3 s 0 76168 800 76288 0 FreeSans 480 0 0 0 io_west_out[21]
port 242 nsew signal output
flabel metal3 s 0 77528 800 77648 0 FreeSans 480 0 0 0 io_west_out[22]
port 243 nsew signal output
flabel metal3 s 0 78888 800 79008 0 FreeSans 480 0 0 0 io_west_out[23]
port 244 nsew signal output
flabel metal3 s 0 79568 800 79688 0 FreeSans 480 0 0 0 io_west_out[24]
port 245 nsew signal output
flabel metal3 s 0 80928 800 81048 0 FreeSans 480 0 0 0 io_west_out[25]
port 246 nsew signal output
flabel metal3 s 0 81608 800 81728 0 FreeSans 480 0 0 0 io_west_out[26]
port 247 nsew signal output
flabel metal3 s 0 82968 800 83088 0 FreeSans 480 0 0 0 io_west_out[27]
port 248 nsew signal output
flabel metal3 s 0 84328 800 84448 0 FreeSans 480 0 0 0 io_west_out[28]
port 249 nsew signal output
flabel metal3 s 0 85008 800 85128 0 FreeSans 480 0 0 0 io_west_out[29]
port 250 nsew signal output
flabel metal3 s 0 31288 800 31408 0 FreeSans 480 0 0 0 io_west_out[2]
port 251 nsew signal output
flabel metal3 s 0 86368 800 86488 0 FreeSans 480 0 0 0 io_west_out[30]
port 252 nsew signal output
flabel metal3 s 0 87048 800 87168 0 FreeSans 480 0 0 0 io_west_out[31]
port 253 nsew signal output
flabel metal3 s 0 31968 800 32088 0 FreeSans 480 0 0 0 io_west_out[3]
port 254 nsew signal output
flabel metal3 s 0 33328 800 33448 0 FreeSans 480 0 0 0 io_west_out[4]
port 255 nsew signal output
flabel metal3 s 0 34688 800 34808 0 FreeSans 480 0 0 0 io_west_out[5]
port 256 nsew signal output
flabel metal3 s 0 35368 800 35488 0 FreeSans 480 0 0 0 io_west_out[6]
port 257 nsew signal output
flabel metal3 s 0 36728 800 36848 0 FreeSans 480 0 0 0 io_west_out[7]
port 258 nsew signal output
flabel metal3 s 0 37408 800 37528 0 FreeSans 480 0 0 0 io_west_out[8]
port 259 nsew signal output
flabel metal3 s 0 38768 800 38888 0 FreeSans 480 0 0 0 io_west_out[9]
port 260 nsew signal output
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 le_clk
port 261 nsew signal input
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 le_en
port 262 nsew signal input
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 le_nrst
port 263 nsew signal input
flabel metal2 s 52826 97200 52882 98000 0 FreeSans 224 90 0 0 nrst
port 264 nsew signal input
flabel metal4 s -416 656 -96 97264 0 FreeSans 1920 90 0 0 vccd1
port 265 nsew power bidirectional
flabel metal5 s -416 656 99408 976 0 FreeSans 2560 0 0 0 vccd1
port 265 nsew power bidirectional
flabel metal5 s -416 96944 99408 97264 0 FreeSans 2560 0 0 0 vccd1
port 265 nsew power bidirectional
flabel metal4 s 99088 656 99408 97264 0 FreeSans 1920 90 0 0 vccd1
port 265 nsew power bidirectional
flabel metal4 s 4208 -4 4528 97924 0 FreeSans 1920 90 0 0 vccd1
port 265 nsew power bidirectional
flabel metal4 s 34928 -4 35248 8015 0 FreeSans 1920 90 0 0 vccd1
port 265 nsew power bidirectional
flabel metal4 s 34928 91057 35248 97924 0 FreeSans 1920 90 0 0 vccd1
port 265 nsew power bidirectional
flabel metal4 s 65648 -4 65968 8015 0 FreeSans 1920 90 0 0 vccd1
port 265 nsew power bidirectional
flabel metal4 s 65648 91057 65968 97924 0 FreeSans 1920 90 0 0 vccd1
port 265 nsew power bidirectional
flabel metal4 s 96368 -4 96688 97924 0 FreeSans 1920 90 0 0 vccd1
port 265 nsew power bidirectional
flabel metal5 s -1076 5346 100068 5666 0 FreeSans 2560 0 0 0 vccd1
port 265 nsew power bidirectional
flabel metal5 s -1076 35982 100068 36302 0 FreeSans 2560 0 0 0 vccd1
port 265 nsew power bidirectional
flabel metal5 s -1076 66618 100068 66938 0 FreeSans 2560 0 0 0 vccd1
port 265 nsew power bidirectional
flabel metal4 s -1076 -4 -756 97924 0 FreeSans 1920 90 0 0 vssd1
port 266 nsew ground bidirectional
flabel metal5 s -1076 -4 100068 316 0 FreeSans 2560 0 0 0 vssd1
port 266 nsew ground bidirectional
flabel metal5 s -1076 97604 100068 97924 0 FreeSans 2560 0 0 0 vssd1
port 266 nsew ground bidirectional
flabel metal4 s 99748 -4 100068 97924 0 FreeSans 1920 90 0 0 vssd1
port 266 nsew ground bidirectional
flabel metal4 s 4868 -4 5188 97924 0 FreeSans 1920 90 0 0 vssd1
port 266 nsew ground bidirectional
flabel metal4 s 35588 -4 35908 8015 0 FreeSans 1920 90 0 0 vssd1
port 266 nsew ground bidirectional
flabel metal4 s 35588 91057 35908 97924 0 FreeSans 1920 90 0 0 vssd1
port 266 nsew ground bidirectional
flabel metal4 s 66308 -4 66628 8015 0 FreeSans 1920 90 0 0 vssd1
port 266 nsew ground bidirectional
flabel metal4 s 66308 91057 66628 97924 0 FreeSans 1920 90 0 0 vssd1
port 266 nsew ground bidirectional
flabel metal4 s 97028 -4 97348 97924 0 FreeSans 1920 90 0 0 vssd1
port 266 nsew ground bidirectional
flabel metal5 s -1076 6006 100068 6326 0 FreeSans 2560 0 0 0 vssd1
port 266 nsew ground bidirectional
flabel metal5 s -1076 36642 100068 36962 0 FreeSans 2560 0 0 0 vssd1
port 266 nsew ground bidirectional
flabel metal5 s -1076 67278 100068 67598 0 FreeSans 2560 0 0 0 vssd1
port 266 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 99000 98000
<< end >>
