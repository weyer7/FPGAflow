magic
tech sky130A
magscale 1 2
timestamp 1746142391
<< viali >>
rect 15393 25925 15427 25959
rect 17325 25925 17359 25959
rect 8125 25857 8159 25891
rect 8217 25857 8251 25891
rect 8401 25857 8435 25891
rect 9505 25857 9539 25891
rect 9597 25857 9631 25891
rect 9781 25857 9815 25891
rect 15301 25857 15335 25891
rect 15577 25857 15611 25891
rect 20085 25857 20119 25891
rect 20637 25857 20671 25891
rect 12081 25789 12115 25823
rect 16221 25789 16255 25823
rect 16773 25789 16807 25823
rect 20177 25789 20211 25823
rect 21189 25789 21223 25823
rect 23305 25789 23339 25823
rect 23581 25789 23615 25823
rect 24041 25789 24075 25823
rect 24317 25789 24351 25823
rect 15577 25721 15611 25755
rect 5549 25653 5583 25687
rect 8401 25653 8435 25687
rect 9781 25653 9815 25687
rect 11529 25653 11563 25687
rect 15669 25653 15703 25687
rect 19717 25653 19751 25687
rect 21833 25653 21867 25687
rect 25789 25653 25823 25687
rect 8585 25449 8619 25483
rect 8953 25449 8987 25483
rect 10425 25449 10459 25483
rect 12449 25449 12483 25483
rect 21005 25449 21039 25483
rect 24133 25449 24167 25483
rect 9781 25381 9815 25415
rect 12909 25381 12943 25415
rect 5181 25313 5215 25347
rect 8401 25313 8435 25347
rect 8493 25313 8527 25347
rect 10149 25313 10183 25347
rect 15485 25313 15519 25347
rect 19533 25313 19567 25347
rect 23489 25313 23523 25347
rect 23765 25313 23799 25347
rect 4905 25245 4939 25279
rect 8677 25245 8711 25279
rect 8769 25245 8803 25279
rect 9505 25245 9539 25279
rect 10701 25245 10735 25279
rect 12725 25245 12759 25279
rect 13001 25245 13035 25279
rect 13277 25245 13311 25279
rect 13829 25245 13863 25279
rect 14473 25245 14507 25279
rect 15209 25245 15243 25279
rect 19257 25245 19291 25279
rect 21281 25245 21315 25279
rect 21465 25245 21499 25279
rect 22109 25245 22143 25279
rect 22293 25245 22327 25279
rect 22385 25245 22419 25279
rect 22937 25245 22971 25279
rect 23121 25245 23155 25279
rect 23305 25245 23339 25279
rect 23857 25245 23891 25279
rect 26157 25245 26191 25279
rect 26341 25245 26375 25279
rect 26893 25245 26927 25279
rect 26985 25245 27019 25279
rect 27169 25245 27203 25279
rect 5457 25177 5491 25211
rect 10241 25177 10275 25211
rect 10977 25177 11011 25211
rect 25881 25177 25915 25211
rect 27077 25177 27111 25211
rect 6929 25109 6963 25143
rect 7757 25109 7791 25143
rect 9689 25109 9723 25143
rect 10441 25109 10475 25143
rect 10609 25109 10643 25143
rect 12541 25109 12575 25143
rect 15117 25109 15151 25143
rect 16957 25109 16991 25143
rect 21373 25109 21407 25143
rect 22201 25109 22235 25143
rect 24409 25109 24443 25143
rect 7849 24905 7883 24939
rect 10241 24905 10275 24939
rect 22937 24905 22971 24939
rect 23121 24905 23155 24939
rect 26249 24905 26283 24939
rect 4721 24837 4755 24871
rect 7297 24837 7331 24871
rect 10333 24837 10367 24871
rect 17785 24837 17819 24871
rect 22569 24837 22603 24871
rect 22769 24837 22803 24871
rect 25881 24837 25915 24871
rect 26097 24837 26131 24871
rect 7113 24769 7147 24803
rect 10057 24769 10091 24803
rect 10885 24769 10919 24803
rect 11529 24769 11563 24803
rect 11713 24769 11747 24803
rect 13645 24769 13679 24803
rect 13829 24769 13863 24803
rect 13921 24769 13955 24803
rect 14105 24769 14139 24803
rect 14197 24769 14231 24803
rect 14381 24769 14415 24803
rect 16313 24769 16347 24803
rect 16497 24769 16531 24803
rect 17693 24769 17727 24803
rect 17969 24769 18003 24803
rect 18061 24769 18095 24803
rect 19901 24769 19935 24803
rect 23029 24769 23063 24803
rect 23213 24769 23247 24803
rect 24961 24769 24995 24803
rect 25053 24769 25087 24803
rect 25145 24769 25179 24803
rect 25789 24769 25823 24803
rect 26341 24769 26375 24803
rect 26525 24769 26559 24803
rect 26617 24769 26651 24803
rect 26985 24769 27019 24803
rect 27169 24769 27203 24803
rect 27813 24769 27847 24803
rect 4445 24701 4479 24735
rect 6193 24701 6227 24735
rect 9321 24701 9355 24735
rect 9597 24701 9631 24735
rect 9781 24701 9815 24735
rect 11805 24701 11839 24735
rect 12081 24701 12115 24735
rect 14473 24701 14507 24735
rect 14749 24701 14783 24735
rect 16405 24701 16439 24735
rect 16681 24701 16715 24735
rect 17417 24701 17451 24735
rect 19165 24701 19199 24735
rect 20177 24701 20211 24735
rect 21649 24701 21683 24735
rect 22385 24701 22419 24735
rect 13645 24633 13679 24667
rect 14381 24633 14415 24667
rect 16221 24633 16255 24667
rect 17509 24633 17543 24667
rect 17785 24633 17819 24667
rect 26341 24633 26375 24667
rect 7389 24565 7423 24599
rect 9873 24565 9907 24599
rect 11529 24565 11563 24599
rect 13553 24565 13587 24599
rect 17325 24565 17359 24599
rect 17601 24565 17635 24599
rect 18613 24565 18647 24599
rect 21833 24565 21867 24599
rect 22753 24565 22787 24599
rect 26065 24565 26099 24599
rect 26985 24565 27019 24599
rect 27721 24565 27755 24599
rect 8677 24361 8711 24395
rect 10701 24361 10735 24395
rect 13001 24361 13035 24395
rect 16313 24361 16347 24395
rect 19257 24361 19291 24395
rect 21741 24361 21775 24395
rect 26433 24361 26467 24395
rect 12817 24293 12851 24327
rect 16129 24293 16163 24327
rect 16681 24293 16715 24327
rect 22431 24293 22465 24327
rect 6929 24225 6963 24259
rect 8953 24225 8987 24259
rect 10977 24225 11011 24259
rect 14289 24225 14323 24259
rect 16037 24225 16071 24259
rect 17325 24225 17359 24259
rect 19809 24225 19843 24259
rect 21281 24225 21315 24259
rect 21925 24225 21959 24259
rect 24225 24225 24259 24259
rect 25513 24225 25547 24259
rect 25973 24225 26007 24259
rect 26525 24225 26559 24259
rect 26801 24225 26835 24259
rect 20637 24157 20671 24191
rect 21005 24157 21039 24191
rect 21097 24157 21131 24191
rect 21373 24157 21407 24191
rect 21465 24157 21499 24191
rect 21557 24157 21591 24191
rect 21741 24157 21775 24191
rect 22017 24157 22051 24191
rect 22293 24157 22327 24191
rect 23857 24157 23891 24191
rect 25697 24157 25731 24191
rect 25789 24157 25823 24191
rect 25881 24157 25915 24191
rect 26249 24157 26283 24191
rect 26433 24157 26467 24191
rect 7205 24089 7239 24123
rect 9229 24089 9263 24123
rect 11253 24089 11287 24123
rect 12985 24089 13019 24123
rect 13185 24089 13219 24123
rect 14565 24089 14599 24123
rect 16313 24089 16347 24123
rect 17601 24089 17635 24123
rect 20085 24089 20119 24123
rect 12725 24021 12759 24055
rect 19073 24021 19107 24055
rect 19625 24021 19659 24055
rect 19717 24021 19751 24055
rect 20821 24021 20855 24055
rect 22201 24021 22235 24055
rect 28273 24021 28307 24055
rect 9229 23817 9263 23851
rect 12265 23817 12299 23851
rect 15209 23817 15243 23851
rect 15945 23817 15979 23851
rect 16773 23817 16807 23851
rect 19349 23817 19383 23851
rect 20177 23817 20211 23851
rect 22569 23817 22603 23851
rect 27077 23817 27111 23851
rect 8953 23749 8987 23783
rect 17877 23749 17911 23783
rect 20269 23749 20303 23783
rect 21281 23749 21315 23783
rect 9137 23681 9171 23715
rect 9229 23681 9263 23715
rect 10977 23681 11011 23715
rect 11069 23681 11103 23715
rect 11253 23681 11287 23715
rect 11897 23681 11931 23715
rect 12173 23681 12207 23715
rect 12357 23681 12391 23715
rect 15853 23681 15887 23715
rect 16129 23681 16163 23715
rect 16313 23681 16347 23715
rect 16681 23681 16715 23715
rect 16865 23681 16899 23715
rect 19717 23681 19751 23715
rect 19809 23681 19843 23715
rect 21005 23681 21039 23715
rect 21153 23681 21187 23715
rect 21373 23681 21407 23715
rect 21511 23681 21545 23715
rect 22293 23681 22327 23715
rect 22661 23681 22695 23715
rect 25697 23681 25731 23715
rect 26433 23681 26467 23715
rect 26617 23681 26651 23715
rect 26801 23681 26835 23715
rect 28181 23681 28215 23715
rect 11161 23613 11195 23647
rect 11713 23613 11747 23647
rect 12081 23613 12115 23647
rect 17601 23613 17635 23647
rect 19533 23613 19567 23647
rect 20821 23613 20855 23647
rect 27721 23613 27755 23647
rect 28089 23613 28123 23647
rect 27813 23545 27847 23579
rect 10793 23477 10827 23511
rect 21649 23477 21683 23511
rect 22201 23477 22235 23511
rect 25605 23477 25639 23511
rect 11345 23273 11379 23307
rect 20177 23273 20211 23307
rect 28273 23273 28307 23307
rect 15301 23205 15335 23239
rect 18981 23205 19015 23239
rect 10977 23137 11011 23171
rect 16037 23137 16071 23171
rect 17233 23137 17267 23171
rect 21925 23137 21959 23171
rect 26525 23137 26559 23171
rect 26801 23137 26835 23171
rect 11161 23069 11195 23103
rect 15025 23069 15059 23103
rect 15853 23069 15887 23103
rect 16129 23069 16163 23103
rect 19533 23069 19567 23103
rect 21649 23069 21683 23103
rect 21833 23069 21867 23103
rect 22017 23069 22051 23103
rect 22201 23069 22235 23103
rect 26249 23069 26283 23103
rect 15301 23001 15335 23035
rect 17509 23001 17543 23035
rect 15117 22933 15151 22967
rect 22385 22933 22419 22967
rect 26341 22933 26375 22967
rect 15669 22729 15703 22763
rect 7849 22661 7883 22695
rect 13277 22661 13311 22695
rect 14933 22661 14967 22695
rect 24317 22661 24351 22695
rect 26249 22661 26283 22695
rect 7481 22593 7515 22627
rect 7757 22593 7791 22627
rect 8033 22593 8067 22627
rect 12173 22593 12207 22627
rect 14105 22593 14139 22627
rect 15117 22593 15151 22627
rect 15209 22593 15243 22627
rect 15301 22593 15335 22627
rect 17233 22593 17267 22627
rect 23949 22593 23983 22627
rect 24042 22593 24076 22627
rect 24225 22593 24259 22627
rect 24414 22593 24448 22627
rect 24685 22593 24719 22627
rect 24869 22593 24903 22627
rect 24961 22593 24995 22627
rect 25237 22593 25271 22627
rect 26433 22593 26467 22627
rect 26525 22593 26559 22627
rect 26801 22593 26835 22627
rect 27721 22593 27755 22627
rect 14289 22525 14323 22559
rect 16221 22525 16255 22559
rect 20361 22525 20395 22559
rect 22385 22525 22419 22559
rect 23765 22525 23799 22559
rect 25053 22525 25087 22559
rect 25605 22525 25639 22559
rect 27629 22525 27663 22559
rect 24593 22457 24627 22491
rect 25421 22457 25455 22491
rect 26709 22457 26743 22491
rect 8033 22389 8067 22423
rect 11989 22389 12023 22423
rect 14841 22389 14875 22423
rect 15209 22389 15243 22423
rect 15485 22389 15519 22423
rect 16681 22389 16715 22423
rect 19809 22389 19843 22423
rect 21833 22389 21867 22423
rect 23213 22389 23247 22423
rect 26157 22389 26191 22423
rect 26985 22389 27019 22423
rect 28365 22389 28399 22423
rect 15945 22185 15979 22219
rect 16221 22185 16255 22219
rect 19520 22185 19554 22219
rect 21360 22185 21394 22219
rect 22845 22185 22879 22219
rect 25991 22185 26025 22219
rect 26604 22185 26638 22219
rect 16405 22117 16439 22151
rect 5825 22049 5859 22083
rect 6009 22049 6043 22083
rect 9229 22049 9263 22083
rect 11253 22049 11287 22083
rect 12173 22049 12207 22083
rect 14197 22049 14231 22083
rect 14473 22049 14507 22083
rect 16589 22049 16623 22083
rect 17325 22049 17359 22083
rect 19257 22049 19291 22083
rect 21097 22049 21131 22083
rect 23949 22049 23983 22083
rect 26249 22049 26283 22083
rect 26341 22049 26375 22083
rect 9321 21981 9355 22015
rect 11161 21981 11195 22015
rect 11437 21981 11471 22015
rect 12081 21981 12115 22015
rect 16497 21981 16531 22015
rect 16681 21981 16715 22015
rect 5549 21913 5583 21947
rect 6285 21913 6319 21947
rect 7849 21913 7883 21947
rect 8677 21913 8711 21947
rect 12449 21913 12483 21947
rect 16037 21913 16071 21947
rect 17601 21913 17635 21947
rect 23765 21913 23799 21947
rect 4077 21845 4111 21879
rect 7757 21845 7791 21879
rect 8953 21845 8987 21879
rect 11621 21845 11655 21879
rect 11897 21845 11931 21879
rect 13921 21845 13955 21879
rect 16237 21845 16271 21879
rect 19073 21845 19107 21879
rect 21005 21845 21039 21879
rect 23305 21845 23339 21879
rect 23673 21845 23707 21879
rect 24501 21845 24535 21879
rect 28089 21845 28123 21879
rect 4905 21641 4939 21675
rect 6469 21641 6503 21675
rect 16497 21641 16531 21675
rect 20085 21641 20119 21675
rect 20545 21641 20579 21675
rect 21833 21641 21867 21675
rect 24501 21641 24535 21675
rect 25697 21641 25731 21675
rect 5687 21573 5721 21607
rect 5917 21573 5951 21607
rect 9137 21573 9171 21607
rect 11805 21573 11839 21607
rect 19809 21573 19843 21607
rect 22293 21573 22327 21607
rect 23029 21573 23063 21607
rect 27353 21573 27387 21607
rect 4445 21505 4479 21539
rect 5089 21505 5123 21539
rect 5181 21505 5215 21539
rect 5273 21505 5307 21539
rect 5457 21505 5491 21539
rect 5825 21505 5859 21539
rect 6009 21505 6043 21539
rect 6837 21505 6871 21539
rect 8861 21505 8895 21539
rect 9413 21505 9447 21539
rect 9597 21505 9631 21539
rect 13461 21505 13495 21539
rect 14289 21505 14323 21539
rect 19073 21505 19107 21539
rect 20453 21505 20487 21539
rect 20913 21505 20947 21539
rect 22201 21505 22235 21539
rect 25329 21505 25363 21539
rect 25789 21505 25823 21539
rect 26985 21505 27019 21539
rect 27078 21505 27112 21539
rect 27261 21505 27295 21539
rect 27450 21505 27484 21539
rect 4353 21437 4387 21471
rect 5549 21437 5583 21471
rect 6745 21437 6779 21471
rect 9137 21437 9171 21471
rect 9873 21437 9907 21471
rect 11529 21437 11563 21471
rect 14381 21437 14415 21471
rect 14749 21437 14783 21471
rect 15025 21437 15059 21471
rect 20637 21437 20671 21471
rect 21465 21437 21499 21471
rect 22477 21437 22511 21471
rect 22753 21437 22787 21471
rect 25145 21437 25179 21471
rect 25237 21437 25271 21471
rect 26341 21437 26375 21471
rect 28273 21437 28307 21471
rect 4813 21369 4847 21403
rect 11345 21369 11379 21403
rect 13277 21369 13311 21403
rect 27721 21369 27755 21403
rect 6193 21301 6227 21335
rect 6837 21301 6871 21335
rect 9321 21301 9355 21335
rect 14657 21301 14691 21335
rect 27629 21301 27663 21335
rect 4997 21097 5031 21131
rect 6745 21097 6779 21131
rect 12081 21097 12115 21131
rect 12173 21097 12207 21131
rect 15485 21097 15519 21131
rect 17509 21097 17543 21131
rect 24225 21097 24259 21131
rect 9597 20961 9631 20995
rect 11345 20961 11379 20995
rect 11437 20961 11471 20995
rect 14841 20961 14875 20995
rect 19901 20961 19935 20995
rect 21741 20961 21775 20995
rect 23489 20961 23523 20995
rect 23581 20961 23615 20995
rect 25145 20961 25179 20995
rect 26525 20961 26559 20995
rect 26801 20961 26835 20995
rect 5181 20893 5215 20927
rect 5365 20893 5399 20927
rect 5549 20893 5583 20927
rect 6193 20893 6227 20927
rect 6561 20893 6595 20927
rect 6929 20893 6963 20927
rect 8677 20893 8711 20927
rect 8953 20893 8987 20927
rect 9137 20893 9171 20927
rect 9321 20893 9355 20927
rect 12357 20893 12391 20927
rect 12541 20893 12575 20927
rect 12633 20893 12667 20927
rect 12725 20893 12759 20927
rect 12909 20893 12943 20927
rect 15577 20893 15611 20927
rect 15853 20893 15887 20927
rect 17693 20893 17727 20927
rect 17969 20893 18003 20927
rect 19349 20893 19383 20927
rect 5273 20825 5307 20859
rect 6377 20825 6411 20859
rect 6469 20825 6503 20859
rect 7665 20825 7699 20859
rect 9229 20825 9263 20859
rect 9873 20825 9907 20859
rect 12817 20825 12851 20859
rect 15669 20825 15703 20859
rect 20177 20825 20211 20859
rect 22017 20825 22051 20859
rect 24409 20825 24443 20859
rect 8125 20757 8159 20791
rect 9505 20757 9539 20791
rect 16037 20757 16071 20791
rect 17877 20757 17911 20791
rect 21649 20757 21683 20791
rect 28273 20757 28307 20791
rect 7481 20553 7515 20587
rect 9597 20553 9631 20587
rect 10333 20553 10367 20587
rect 19901 20553 19935 20587
rect 22661 20553 22695 20587
rect 25237 20553 25271 20587
rect 26985 20553 27019 20587
rect 5825 20485 5859 20519
rect 7021 20485 7055 20519
rect 10057 20485 10091 20519
rect 13461 20485 13495 20519
rect 21097 20485 21131 20519
rect 27445 20485 27479 20519
rect 28089 20485 28123 20519
rect 28181 20485 28215 20519
rect 5641 20417 5675 20451
rect 5733 20417 5767 20451
rect 6009 20417 6043 20451
rect 7205 20417 7239 20451
rect 7297 20417 7331 20451
rect 9781 20417 9815 20451
rect 9965 20417 9999 20451
rect 10149 20417 10183 20451
rect 12357 20417 12391 20451
rect 13369 20417 13403 20451
rect 17325 20417 17359 20451
rect 18153 20417 18187 20451
rect 21465 20417 21499 20451
rect 22017 20417 22051 20451
rect 26801 20417 26835 20451
rect 27353 20417 27387 20451
rect 27997 20417 28031 20451
rect 28365 20417 28399 20451
rect 3617 20349 3651 20383
rect 3893 20349 3927 20383
rect 7849 20349 7883 20383
rect 8125 20349 8159 20383
rect 14197 20349 14231 20383
rect 14657 20349 14691 20383
rect 14933 20349 14967 20383
rect 17233 20349 17267 20383
rect 18429 20349 18463 20383
rect 23489 20349 23523 20383
rect 23765 20349 23799 20383
rect 26249 20349 26283 20383
rect 27537 20349 27571 20383
rect 5457 20281 5491 20315
rect 12173 20281 12207 20315
rect 5365 20213 5399 20247
rect 7021 20213 7055 20247
rect 16405 20213 16439 20247
rect 17693 20213 17727 20247
rect 27813 20213 27847 20247
rect 7159 20009 7193 20043
rect 7389 20009 7423 20043
rect 7941 20009 7975 20043
rect 8677 20009 8711 20043
rect 13645 20009 13679 20043
rect 17417 20009 17451 20043
rect 17785 20009 17819 20043
rect 19901 20009 19935 20043
rect 26801 20009 26835 20043
rect 27813 20009 27847 20043
rect 7297 19941 7331 19975
rect 8953 19873 8987 19907
rect 12081 19873 12115 19907
rect 13829 19873 13863 19907
rect 14197 19873 14231 19907
rect 16773 19873 16807 19907
rect 20361 19873 20395 19907
rect 20821 19873 20855 19907
rect 22109 19873 22143 19907
rect 22385 19873 22419 19907
rect 27261 19873 27295 19907
rect 27353 19873 27387 19907
rect 7021 19805 7055 19839
rect 7481 19805 7515 19839
rect 8125 19805 8159 19839
rect 8217 19805 8251 19839
rect 8493 19805 8527 19839
rect 8769 19805 8803 19839
rect 9137 19805 9171 19839
rect 9413 19805 9447 19839
rect 11529 19805 11563 19839
rect 11897 19805 11931 19839
rect 12449 19805 12483 19839
rect 12541 19815 12575 19849
rect 12909 19805 12943 19839
rect 13553 19805 13587 19839
rect 14105 19805 14139 19839
rect 15853 19805 15887 19839
rect 17964 19805 17998 19839
rect 18281 19805 18315 19839
rect 18429 19805 18463 19839
rect 19257 19805 19291 19839
rect 19405 19805 19439 19839
rect 19625 19805 19659 19839
rect 19722 19805 19756 19839
rect 20453 19805 20487 19839
rect 22017 19805 22051 19839
rect 23397 19805 23431 19839
rect 23581 19805 23615 19839
rect 23674 19805 23708 19839
rect 24087 19805 24121 19839
rect 24777 19805 24811 19839
rect 25053 19805 25087 19839
rect 27997 19805 28031 19839
rect 28365 19805 28399 19839
rect 8309 19737 8343 19771
rect 13461 19737 13495 19771
rect 18061 19737 18095 19771
rect 18153 19737 18187 19771
rect 19533 19737 19567 19771
rect 23857 19737 23891 19771
rect 23949 19737 23983 19771
rect 25329 19737 25363 19771
rect 9321 19669 9355 19703
rect 11621 19669 11655 19703
rect 12725 19669 12759 19703
rect 13829 19669 13863 19703
rect 15669 19669 15703 19703
rect 24225 19669 24259 19703
rect 27445 19669 27479 19703
rect 5917 19465 5951 19499
rect 11253 19465 11287 19499
rect 11713 19465 11747 19499
rect 12035 19465 12069 19499
rect 16037 19465 16071 19499
rect 18153 19465 18187 19499
rect 18889 19465 18923 19499
rect 22477 19465 22511 19499
rect 23949 19465 23983 19499
rect 27721 19465 27755 19499
rect 4879 19397 4913 19431
rect 18521 19397 18555 19431
rect 22201 19397 22235 19431
rect 22569 19397 22603 19431
rect 24317 19397 24351 19431
rect 4997 19329 5031 19363
rect 5089 19329 5123 19363
rect 5181 19329 5215 19363
rect 5457 19329 5491 19363
rect 5641 19329 5675 19363
rect 5825 19329 5859 19363
rect 5917 19329 5951 19363
rect 6101 19329 6135 19363
rect 7573 19329 7607 19363
rect 11161 19329 11195 19363
rect 11345 19329 11379 19363
rect 11897 19329 11931 19363
rect 13461 19329 13495 19363
rect 16221 19329 16255 19363
rect 17049 19329 17083 19363
rect 18245 19329 18279 19363
rect 18338 19329 18372 19363
rect 18613 19329 18647 19363
rect 18751 19329 18785 19363
rect 21281 19329 21315 19363
rect 21833 19329 21867 19363
rect 21926 19329 21960 19363
rect 22109 19329 22143 19363
rect 22298 19329 22332 19363
rect 23305 19329 23339 19363
rect 23398 19329 23432 19363
rect 23581 19329 23615 19363
rect 23673 19329 23707 19363
rect 23770 19329 23804 19363
rect 4721 19261 4755 19295
rect 5365 19261 5399 19295
rect 7849 19261 7883 19295
rect 13829 19261 13863 19295
rect 15761 19261 15795 19295
rect 17141 19261 17175 19295
rect 17509 19261 17543 19295
rect 23213 19261 23247 19295
rect 25145 19261 25179 19295
rect 28273 19261 28307 19295
rect 17417 19193 17451 19227
rect 9321 19125 9355 19159
rect 15117 19125 15151 19159
rect 5549 18921 5583 18955
rect 6285 18921 6319 18955
rect 9045 18921 9079 18955
rect 11897 18921 11931 18955
rect 14473 18921 14507 18955
rect 14841 18921 14875 18955
rect 18429 18921 18463 18955
rect 23949 18921 23983 18955
rect 27905 18921 27939 18955
rect 5733 18853 5767 18887
rect 11437 18853 11471 18887
rect 13829 18853 13863 18887
rect 18337 18853 18371 18887
rect 12173 18785 12207 18819
rect 12541 18785 12575 18819
rect 15117 18785 15151 18819
rect 16865 18785 16899 18819
rect 17509 18785 17543 18819
rect 18061 18785 18095 18819
rect 18981 18785 19015 18819
rect 20177 18785 20211 18819
rect 20453 18785 20487 18819
rect 22201 18785 22235 18819
rect 22937 18785 22971 18819
rect 24501 18785 24535 18819
rect 4813 18717 4847 18751
rect 5365 18717 5399 18751
rect 5457 18717 5491 18751
rect 5733 18717 5767 18751
rect 6009 18717 6043 18751
rect 6101 18717 6135 18751
rect 6469 18717 6503 18751
rect 9321 18717 9355 18751
rect 9781 18717 9815 18751
rect 11253 18717 11287 18751
rect 11437 18717 11471 18751
rect 11621 18717 11655 18751
rect 12081 18717 12115 18751
rect 12817 18717 12851 18751
rect 13093 18717 13127 18751
rect 13277 18717 13311 18751
rect 13369 18717 13403 18751
rect 13553 18717 13587 18751
rect 14289 18717 14323 18751
rect 14565 18717 14599 18751
rect 14657 18717 14691 18751
rect 17969 18717 18003 18751
rect 23305 18717 23339 18751
rect 24685 18717 24719 18751
rect 24869 18717 24903 18751
rect 26157 18717 26191 18751
rect 11805 18649 11839 18683
rect 15393 18649 15427 18683
rect 19349 18649 19383 18683
rect 20729 18649 20763 18683
rect 22293 18649 22327 18683
rect 26433 18649 26467 18683
rect 4261 18581 4295 18615
rect 5825 18581 5859 18615
rect 9597 18581 9631 18615
rect 12633 18581 12667 18615
rect 13645 18581 13679 18615
rect 14105 18581 14139 18615
rect 16957 18581 16991 18615
rect 3893 18377 3927 18411
rect 7573 18377 7607 18411
rect 8217 18377 8251 18411
rect 10885 18377 10919 18411
rect 15761 18377 15795 18411
rect 16129 18377 16163 18411
rect 20561 18377 20595 18411
rect 20729 18377 20763 18411
rect 20821 18377 20855 18411
rect 21189 18377 21223 18411
rect 24501 18377 24535 18411
rect 24685 18377 24719 18411
rect 25789 18377 25823 18411
rect 4629 18309 4663 18343
rect 17141 18309 17175 18343
rect 17341 18309 17375 18343
rect 20361 18309 20395 18343
rect 22293 18309 22327 18343
rect 22753 18309 22787 18343
rect 24869 18309 24903 18343
rect 4169 18241 4203 18275
rect 4261 18241 4295 18275
rect 4537 18241 4571 18275
rect 4813 18241 4847 18275
rect 4997 18241 5031 18275
rect 5089 18241 5123 18275
rect 5457 18241 5491 18275
rect 5549 18241 5583 18275
rect 5825 18241 5859 18275
rect 7757 18241 7791 18275
rect 7849 18241 7883 18275
rect 7941 18241 7975 18275
rect 8125 18241 8159 18275
rect 8493 18241 8527 18275
rect 8953 18241 8987 18275
rect 10793 18241 10827 18275
rect 10977 18241 11011 18275
rect 11529 18241 11563 18275
rect 11897 18241 11931 18275
rect 12357 18241 12391 18275
rect 15945 18241 15979 18275
rect 16221 18241 16255 18275
rect 17877 18241 17911 18275
rect 18153 18241 18187 18275
rect 19073 18241 19107 18275
rect 19349 18241 19383 18275
rect 21005 18241 21039 18275
rect 21281 18241 21315 18275
rect 22109 18241 22143 18275
rect 22385 18241 22419 18275
rect 23673 18241 23707 18275
rect 25145 18241 25179 18275
rect 25329 18241 25363 18275
rect 25421 18241 25455 18275
rect 25513 18241 25547 18275
rect 2145 18173 2179 18207
rect 2421 18173 2455 18207
rect 3985 18173 4019 18207
rect 5181 18173 5215 18207
rect 5641 18173 5675 18207
rect 8401 18173 8435 18207
rect 8769 18173 8803 18207
rect 8861 18173 8895 18207
rect 9229 18173 9263 18207
rect 13829 18173 13863 18207
rect 14105 18173 14139 18207
rect 15577 18173 15611 18207
rect 23305 18173 23339 18207
rect 23581 18173 23615 18207
rect 24041 18173 24075 18207
rect 4445 18105 4479 18139
rect 12173 18105 12207 18139
rect 5273 18037 5307 18071
rect 5365 18037 5399 18071
rect 5641 18037 5675 18071
rect 6009 18037 6043 18071
rect 10701 18037 10735 18071
rect 17325 18037 17359 18071
rect 17509 18037 17543 18071
rect 18889 18037 18923 18071
rect 19533 18037 19567 18071
rect 20545 18037 20579 18071
rect 21925 18037 21959 18071
rect 24685 18037 24719 18071
rect 4169 17833 4203 17867
rect 4353 17833 4387 17867
rect 5641 17833 5675 17867
rect 6009 17833 6043 17867
rect 7113 17833 7147 17867
rect 8493 17833 8527 17867
rect 9413 17833 9447 17867
rect 15669 17833 15703 17867
rect 15853 17833 15887 17867
rect 18613 17833 18647 17867
rect 18889 17833 18923 17867
rect 21005 17833 21039 17867
rect 23305 17833 23339 17867
rect 23489 17833 23523 17867
rect 24869 17833 24903 17867
rect 4905 17765 4939 17799
rect 24225 17765 24259 17799
rect 1869 17697 1903 17731
rect 2145 17697 2179 17731
rect 3801 17697 3835 17731
rect 9781 17697 9815 17731
rect 10609 17697 10643 17731
rect 11161 17697 11195 17731
rect 16865 17697 16899 17731
rect 19257 17697 19291 17731
rect 21465 17697 21499 17731
rect 21741 17697 21775 17731
rect 26525 17697 26559 17731
rect 3985 17629 4019 17663
rect 4261 17629 4295 17663
rect 4537 17629 4571 17663
rect 4721 17629 4755 17663
rect 4813 17629 4847 17663
rect 5084 17629 5118 17663
rect 5456 17629 5490 17663
rect 5549 17629 5583 17663
rect 5641 17629 5675 17663
rect 5825 17629 5859 17663
rect 6561 17629 6595 17663
rect 6653 17629 6687 17663
rect 6837 17629 6871 17663
rect 6929 17629 6963 17663
rect 8769 17629 8803 17663
rect 9597 17629 9631 17663
rect 9689 17629 9723 17663
rect 9873 17629 9907 17663
rect 10977 17629 11011 17663
rect 11253 17629 11287 17663
rect 11437 17629 11471 17663
rect 23949 17629 23983 17663
rect 24133 17629 24167 17663
rect 24225 17629 24259 17663
rect 24409 17629 24443 17663
rect 24685 17629 24719 17663
rect 25145 17629 25179 17663
rect 25237 17629 25271 17663
rect 25513 17629 25547 17663
rect 25605 17629 25639 17663
rect 25881 17629 25915 17663
rect 5181 17561 5215 17595
rect 5273 17561 5307 17595
rect 8493 17561 8527 17595
rect 8677 17561 8711 17595
rect 15485 17561 15519 17595
rect 17141 17561 17175 17595
rect 18705 17561 18739 17595
rect 18921 17561 18955 17595
rect 19533 17561 19567 17595
rect 23673 17561 23707 17595
rect 24501 17561 24535 17595
rect 26801 17561 26835 17595
rect 3617 17493 3651 17527
rect 10057 17493 10091 17527
rect 10793 17493 10827 17527
rect 11345 17493 11379 17527
rect 15685 17493 15719 17527
rect 19073 17493 19107 17527
rect 23213 17493 23247 17527
rect 23463 17493 23497 17527
rect 25053 17493 25087 17527
rect 25789 17493 25823 17527
rect 28273 17493 28307 17527
rect 5273 17289 5307 17323
rect 8953 17289 8987 17323
rect 10149 17289 10183 17323
rect 17417 17289 17451 17323
rect 22411 17289 22445 17323
rect 8309 17221 8343 17255
rect 17785 17221 17819 17255
rect 18245 17221 18279 17255
rect 19073 17221 19107 17255
rect 20085 17221 20119 17255
rect 22201 17221 22235 17255
rect 22905 17221 22939 17255
rect 23121 17221 23155 17255
rect 27721 17221 27755 17255
rect 28089 17221 28123 17255
rect 5181 17153 5215 17187
rect 5365 17153 5399 17187
rect 5641 17153 5675 17187
rect 6745 17153 6779 17187
rect 6929 17153 6963 17187
rect 7021 17153 7055 17187
rect 8493 17153 8527 17187
rect 8585 17153 8619 17187
rect 8769 17153 8803 17187
rect 8861 17153 8895 17187
rect 9113 17153 9147 17187
rect 9229 17153 9263 17187
rect 9321 17153 9355 17187
rect 9505 17153 9539 17187
rect 9781 17153 9815 17187
rect 9965 17153 9999 17187
rect 10241 17153 10275 17187
rect 12357 17153 12391 17187
rect 15301 17153 15335 17187
rect 17233 17153 17267 17187
rect 17601 17153 17635 17187
rect 17877 17153 17911 17187
rect 18797 17153 18831 17187
rect 18981 17153 19015 17187
rect 19257 17153 19291 17187
rect 19441 17153 19475 17187
rect 20729 17153 20763 17187
rect 25605 17153 25639 17187
rect 5733 17085 5767 17119
rect 6561 17085 6595 17119
rect 13921 17085 13955 17119
rect 14197 17085 14231 17119
rect 15577 17085 15611 17119
rect 16681 17085 16715 17119
rect 25329 17085 25363 17119
rect 25513 17085 25547 17119
rect 6009 17017 6043 17051
rect 22753 17017 22787 17051
rect 9597 16949 9631 16983
rect 12173 16949 12207 16983
rect 12449 16949 12483 16983
rect 15117 16949 15151 16983
rect 15485 16949 15519 16983
rect 22385 16949 22419 16983
rect 22569 16949 22603 16983
rect 22937 16949 22971 16983
rect 25421 16949 25455 16983
rect 5641 16745 5675 16779
rect 25053 16745 25087 16779
rect 27169 16745 27203 16779
rect 6101 16677 6135 16711
rect 5549 16609 5583 16643
rect 9413 16609 9447 16643
rect 12725 16609 12759 16643
rect 14473 16609 14507 16643
rect 14749 16609 14783 16643
rect 23765 16609 23799 16643
rect 25145 16609 25179 16643
rect 25237 16609 25271 16643
rect 27721 16609 27755 16643
rect 5825 16541 5859 16575
rect 6280 16541 6314 16575
rect 6469 16541 6503 16575
rect 6597 16541 6631 16575
rect 6745 16541 6779 16575
rect 9243 16541 9277 16575
rect 12817 16541 12851 16575
rect 13829 16541 13863 16575
rect 18521 16541 18555 16575
rect 22385 16541 22419 16575
rect 22661 16541 22695 16575
rect 24869 16541 24903 16575
rect 27629 16541 27663 16575
rect 6377 16473 6411 16507
rect 12449 16473 12483 16507
rect 25513 16473 25547 16507
rect 6009 16405 6043 16439
rect 9045 16405 9079 16439
rect 10977 16405 11011 16439
rect 13461 16405 13495 16439
rect 13645 16405 13679 16439
rect 16221 16405 16255 16439
rect 18705 16405 18739 16439
rect 22201 16405 22235 16439
rect 22569 16405 22603 16439
rect 23121 16405 23155 16439
rect 24685 16405 24719 16439
rect 26985 16405 27019 16439
rect 27537 16405 27571 16439
rect 4445 16201 4479 16235
rect 7757 16201 7791 16235
rect 8125 16201 8159 16235
rect 9321 16201 9355 16235
rect 23581 16201 23615 16235
rect 24869 16201 24903 16235
rect 25329 16201 25363 16235
rect 25789 16201 25823 16235
rect 5917 16133 5951 16167
rect 9045 16133 9079 16167
rect 9965 16133 9999 16167
rect 13737 16133 13771 16167
rect 22109 16133 22143 16167
rect 26617 16133 26651 16167
rect 8401 16065 8435 16099
rect 8835 16065 8869 16099
rect 8953 16065 8987 16099
rect 9137 16065 9171 16099
rect 9413 16065 9447 16099
rect 9505 16065 9539 16099
rect 9689 16065 9723 16099
rect 9781 16065 9815 16099
rect 12628 16065 12662 16099
rect 12725 16065 12759 16099
rect 12817 16065 12851 16099
rect 13000 16065 13034 16099
rect 13093 16065 13127 16099
rect 13461 16065 13495 16099
rect 13554 16065 13588 16099
rect 13829 16065 13863 16099
rect 13967 16065 14001 16099
rect 14749 16065 14783 16099
rect 17877 16065 17911 16099
rect 21097 16065 21131 16099
rect 25053 16065 25087 16099
rect 25237 16065 25271 16099
rect 25697 16065 25731 16099
rect 28365 16065 28399 16099
rect 6193 15997 6227 16031
rect 7916 15997 7950 16031
rect 8033 15997 8067 16031
rect 8677 15997 8711 16031
rect 11529 15997 11563 16031
rect 15025 15997 15059 16031
rect 16497 15997 16531 16031
rect 17233 15997 17267 16031
rect 18153 15997 18187 16031
rect 19625 15997 19659 16031
rect 20269 15997 20303 16031
rect 21373 15997 21407 16031
rect 21833 15997 21867 16031
rect 25973 15997 26007 16031
rect 26157 15997 26191 16031
rect 21281 15929 21315 15963
rect 26249 15929 26283 15963
rect 12173 15861 12207 15895
rect 12449 15861 12483 15895
rect 14105 15861 14139 15895
rect 16681 15861 16715 15895
rect 19717 15861 19751 15895
rect 20913 15861 20947 15895
rect 28181 15861 28215 15895
rect 9045 15657 9079 15691
rect 12265 15657 12299 15691
rect 12909 15657 12943 15691
rect 13645 15657 13679 15691
rect 15945 15657 15979 15691
rect 16313 15657 16347 15691
rect 18245 15657 18279 15691
rect 20637 15657 20671 15691
rect 21097 15657 21131 15691
rect 21373 15657 21407 15691
rect 26157 15657 26191 15691
rect 15853 15589 15887 15623
rect 10149 15521 10183 15555
rect 11805 15521 11839 15555
rect 13185 15521 13219 15555
rect 13277 15521 13311 15555
rect 16405 15521 16439 15555
rect 18889 15521 18923 15555
rect 22109 15521 22143 15555
rect 24409 15521 24443 15555
rect 9229 15453 9263 15487
rect 9781 15453 9815 15487
rect 9873 15453 9907 15487
rect 10425 15453 10459 15487
rect 11897 15453 11931 15487
rect 12081 15453 12115 15487
rect 13461 15453 13495 15487
rect 15209 15453 15243 15487
rect 15357 15453 15391 15487
rect 15674 15453 15708 15487
rect 16129 15453 16163 15487
rect 18429 15453 18463 15487
rect 19809 15453 19843 15487
rect 19993 15453 20027 15487
rect 20086 15453 20120 15487
rect 20269 15453 20303 15487
rect 20458 15453 20492 15487
rect 21925 15453 21959 15487
rect 24133 15453 24167 15487
rect 27813 15453 27847 15487
rect 13001 15385 13035 15419
rect 15485 15385 15519 15419
rect 15577 15385 15611 15419
rect 18521 15385 18555 15419
rect 18613 15385 18647 15419
rect 18731 15385 18765 15419
rect 20361 15385 20395 15419
rect 20821 15385 20855 15419
rect 22385 15385 22419 15419
rect 24685 15385 24719 15419
rect 27905 15385 27939 15419
rect 28089 15385 28123 15419
rect 19257 15317 19291 15351
rect 27629 15317 27663 15351
rect 9597 15113 9631 15147
rect 11897 15113 11931 15147
rect 21649 15113 21683 15147
rect 22201 15113 22235 15147
rect 22569 15113 22603 15147
rect 27813 15113 27847 15147
rect 8493 15045 8527 15079
rect 13737 15045 13771 15079
rect 14105 15045 14139 15079
rect 27905 15045 27939 15079
rect 7021 14977 7055 15011
rect 7205 14977 7239 15011
rect 8401 14977 8435 15011
rect 8677 14977 8711 15011
rect 9321 14977 9355 15011
rect 9781 14977 9815 15011
rect 10057 14977 10091 15011
rect 15853 14977 15887 15011
rect 16037 14977 16071 15011
rect 17233 14977 17267 15011
rect 17877 14977 17911 15011
rect 19901 14977 19935 15011
rect 22385 14977 22419 15011
rect 22661 14977 22695 15011
rect 9229 14909 9263 14943
rect 13369 14909 13403 14943
rect 13645 14909 13679 14943
rect 16129 14909 16163 14943
rect 16681 14909 16715 14943
rect 18153 14909 18187 14943
rect 20177 14909 20211 14943
rect 8861 14841 8895 14875
rect 6837 14773 6871 14807
rect 8953 14773 8987 14807
rect 9965 14773 9999 14807
rect 15669 14773 15703 14807
rect 19625 14773 19659 14807
rect 6745 14569 6779 14603
rect 10241 14569 10275 14603
rect 13645 14569 13679 14603
rect 18245 14569 18279 14603
rect 8953 14501 8987 14535
rect 13461 14501 13495 14535
rect 18981 14501 19015 14535
rect 6469 14433 6503 14467
rect 7481 14433 7515 14467
rect 9597 14433 9631 14467
rect 11621 14433 11655 14467
rect 19533 14433 19567 14467
rect 26801 14433 26835 14467
rect 5457 14365 5491 14399
rect 5549 14365 5583 14399
rect 5825 14365 5859 14399
rect 7297 14365 7331 14399
rect 7665 14365 7699 14399
rect 7757 14365 7791 14399
rect 7941 14365 7975 14399
rect 8125 14365 8159 14399
rect 8217 14365 8251 14399
rect 8493 14365 8527 14399
rect 8585 14365 8619 14399
rect 9137 14365 9171 14399
rect 9229 14365 9263 14399
rect 9321 14365 9355 14399
rect 9689 14365 9723 14399
rect 9965 14365 9999 14399
rect 10057 14365 10091 14399
rect 10333 14365 10367 14399
rect 10517 14365 10551 14399
rect 11345 14365 11379 14399
rect 11529 14365 11563 14399
rect 18153 14365 18187 14399
rect 18337 14365 18371 14399
rect 18705 14365 18739 14399
rect 18797 14365 18831 14399
rect 19257 14365 19291 14399
rect 26525 14365 26559 14399
rect 5641 14297 5675 14331
rect 8401 14297 8435 14331
rect 9439 14297 9473 14331
rect 9873 14297 9907 14331
rect 11437 14297 11471 14331
rect 11897 14297 11931 14331
rect 13613 14297 13647 14331
rect 13829 14297 13863 14331
rect 15301 14297 15335 14331
rect 18981 14297 19015 14331
rect 5273 14229 5307 14263
rect 5917 14229 5951 14263
rect 6285 14229 6319 14263
rect 6377 14229 6411 14263
rect 7481 14229 7515 14263
rect 8033 14229 8067 14263
rect 8769 14229 8803 14263
rect 10701 14229 10735 14263
rect 13369 14229 13403 14263
rect 16589 14229 16623 14263
rect 21005 14229 21039 14263
rect 28273 14229 28307 14263
rect 6193 14025 6227 14059
rect 6377 14025 6411 14059
rect 12265 14025 12299 14059
rect 12909 14025 12943 14059
rect 16497 14025 16531 14059
rect 18981 14025 19015 14059
rect 27813 14025 27847 14059
rect 28273 14025 28307 14059
rect 4721 13957 4755 13991
rect 7021 13957 7055 13991
rect 8861 13957 8895 13991
rect 10609 13957 10643 13991
rect 12449 13957 12483 13991
rect 12633 13957 12667 13991
rect 12817 13957 12851 13991
rect 13369 13957 13403 13991
rect 19901 13957 19935 13991
rect 22109 13957 22143 13991
rect 4445 13889 4479 13923
rect 6561 13889 6595 13923
rect 6653 13889 6687 13923
rect 7573 13889 7607 13923
rect 12173 13889 12207 13923
rect 12357 13889 12391 13923
rect 13093 13889 13127 13923
rect 13277 13889 13311 13923
rect 13645 13889 13679 13923
rect 14749 13889 14783 13923
rect 17693 13889 17727 13923
rect 19257 13889 19291 13923
rect 21971 13889 22005 13923
rect 22201 13889 22235 13923
rect 22329 13889 22363 13923
rect 22477 13889 22511 13923
rect 24133 13889 24167 13923
rect 27261 13889 27295 13923
rect 27537 13889 27571 13923
rect 27997 13889 28031 13923
rect 28089 13889 28123 13923
rect 6929 13821 6963 13855
rect 7205 13821 7239 13855
rect 7665 13821 7699 13855
rect 8585 13821 8619 13855
rect 13369 13821 13403 13855
rect 15025 13821 15059 13855
rect 16681 13821 16715 13855
rect 17325 13821 17359 13855
rect 17417 13821 17451 13855
rect 17509 13821 17543 13855
rect 18981 13821 19015 13855
rect 20453 13821 20487 13855
rect 25881 13821 25915 13855
rect 27353 13821 27387 13855
rect 27721 13821 27755 13855
rect 27445 13753 27479 13787
rect 13553 13685 13587 13719
rect 17877 13685 17911 13719
rect 19165 13685 19199 13719
rect 21833 13685 21867 13719
rect 24396 13685 24430 13719
rect 6837 13481 6871 13515
rect 15945 13481 15979 13515
rect 16129 13481 16163 13515
rect 5089 13345 5123 13379
rect 17601 13345 17635 13379
rect 17877 13345 17911 13379
rect 26525 13345 26559 13379
rect 26801 13345 26835 13379
rect 15301 13277 15335 13311
rect 15394 13277 15428 13311
rect 15577 13277 15611 13311
rect 15807 13277 15841 13311
rect 21557 13277 21591 13311
rect 23949 13277 23983 13311
rect 5365 13209 5399 13243
rect 15669 13209 15703 13243
rect 21833 13209 21867 13243
rect 23305 13141 23339 13175
rect 23397 13141 23431 13175
rect 28273 13141 28307 13175
rect 13553 12937 13587 12971
rect 15577 12937 15611 12971
rect 16313 12937 16347 12971
rect 17785 12937 17819 12971
rect 21833 12937 21867 12971
rect 27905 12937 27939 12971
rect 12633 12869 12667 12903
rect 12725 12869 12759 12903
rect 15945 12869 15979 12903
rect 17417 12869 17451 12903
rect 27445 12869 27479 12903
rect 11897 12801 11931 12835
rect 12541 12801 12575 12835
rect 12909 12801 12943 12835
rect 13737 12801 13771 12835
rect 13829 12801 13863 12835
rect 15669 12801 15703 12835
rect 15762 12801 15796 12835
rect 16037 12801 16071 12835
rect 16175 12801 16209 12835
rect 17141 12801 17175 12835
rect 17234 12801 17268 12835
rect 17509 12801 17543 12835
rect 17647 12801 17681 12835
rect 19533 12801 19567 12835
rect 20729 12801 20763 12835
rect 22017 12801 22051 12835
rect 22293 12801 22327 12835
rect 23305 12801 23339 12835
rect 26433 12801 26467 12835
rect 27169 12801 27203 12835
rect 28089 12801 28123 12835
rect 28365 12801 28399 12835
rect 14105 12733 14139 12767
rect 19717 12733 19751 12767
rect 20361 12733 20395 12767
rect 20453 12733 20487 12767
rect 22201 12733 22235 12767
rect 22477 12733 22511 12767
rect 23581 12733 23615 12767
rect 23765 12733 23799 12767
rect 24317 12733 24351 12767
rect 26157 12733 26191 12767
rect 27353 12733 27387 12767
rect 20545 12665 20579 12699
rect 23121 12665 23155 12699
rect 28181 12665 28215 12699
rect 11713 12597 11747 12631
rect 12357 12597 12391 12631
rect 18981 12597 19015 12631
rect 20913 12597 20947 12631
rect 23029 12597 23063 12631
rect 23489 12597 23523 12631
rect 24685 12597 24719 12631
rect 26985 12597 27019 12631
rect 27169 12597 27203 12631
rect 5825 12393 5859 12427
rect 13737 12393 13771 12427
rect 13921 12393 13955 12427
rect 18705 12393 18739 12427
rect 19257 12393 19291 12427
rect 22385 12393 22419 12427
rect 11161 12325 11195 12359
rect 14197 12325 14231 12359
rect 12081 12257 12115 12291
rect 18613 12257 18647 12291
rect 19073 12257 19107 12291
rect 20729 12257 20763 12291
rect 22477 12257 22511 12291
rect 26249 12257 26283 12291
rect 5273 12189 5307 12223
rect 5641 12189 5675 12223
rect 5917 12189 5951 12223
rect 6101 12189 6135 12223
rect 10241 12189 10275 12223
rect 10425 12189 10459 12223
rect 10517 12189 10551 12223
rect 11340 12189 11374 12223
rect 11437 12189 11471 12223
rect 11712 12189 11746 12223
rect 11805 12189 11839 12223
rect 11989 12189 12023 12223
rect 12265 12189 12299 12223
rect 12357 12189 12391 12223
rect 12817 12189 12851 12223
rect 13093 12189 13127 12223
rect 13277 12189 13311 12223
rect 13369 12189 13403 12223
rect 14381 12189 14415 12223
rect 14473 12189 14507 12223
rect 14565 12189 14599 12223
rect 14657 12189 14691 12223
rect 18889 12189 18923 12223
rect 21005 12189 21039 12223
rect 21741 12189 21775 12223
rect 21834 12189 21868 12223
rect 22206 12189 22240 12223
rect 5457 12121 5491 12155
rect 5549 12121 5583 12155
rect 11529 12121 11563 12155
rect 12541 12121 12575 12155
rect 22017 12121 22051 12155
rect 22109 12121 22143 12155
rect 22753 12121 22787 12155
rect 26525 12121 26559 12155
rect 6009 12053 6043 12087
rect 10057 12053 10091 12087
rect 12633 12053 12667 12087
rect 13737 12053 13771 12087
rect 24225 12053 24259 12087
rect 27997 12053 28031 12087
rect 19073 11849 19107 11883
rect 19165 11849 19199 11883
rect 22661 11849 22695 11883
rect 27353 11849 27387 11883
rect 6837 11781 6871 11815
rect 11989 11781 12023 11815
rect 12817 11781 12851 11815
rect 13737 11781 13771 11815
rect 18705 11781 18739 11815
rect 18797 11781 18831 11815
rect 20637 11781 20671 11815
rect 3341 11713 3375 11747
rect 5917 11713 5951 11747
rect 6101 11713 6135 11747
rect 6193 11713 6227 11747
rect 6469 11713 6503 11747
rect 6653 11713 6687 11747
rect 7389 11713 7423 11747
rect 7573 11713 7607 11747
rect 7757 11713 7791 11747
rect 13001 11713 13035 11747
rect 13185 11713 13219 11747
rect 13277 11713 13311 11747
rect 13369 11713 13403 11747
rect 18429 11713 18463 11747
rect 18577 11713 18611 11747
rect 18935 11713 18969 11747
rect 22109 11713 22143 11747
rect 22385 11713 22419 11747
rect 24409 11713 24443 11747
rect 26801 11713 26835 11747
rect 26985 11713 27019 11747
rect 27169 11713 27203 11747
rect 28365 11713 28399 11747
rect 3617 11645 3651 11679
rect 5089 11645 5123 11679
rect 5825 11645 5859 11679
rect 9597 11645 9631 11679
rect 9873 11645 9907 11679
rect 20913 11645 20947 11679
rect 22569 11645 22603 11679
rect 24133 11645 24167 11679
rect 26525 11645 26559 11679
rect 5181 11509 5215 11543
rect 5917 11509 5951 11543
rect 6561 11509 6595 11543
rect 8309 11509 8343 11543
rect 11345 11509 11379 11543
rect 13645 11509 13679 11543
rect 22201 11509 22235 11543
rect 25053 11509 25087 11543
rect 26985 11509 27019 11543
rect 28181 11509 28215 11543
rect 4353 11305 4387 11339
rect 5365 11305 5399 11339
rect 10793 11305 10827 11339
rect 12909 11305 12943 11339
rect 13093 11305 13127 11339
rect 13369 11305 13403 11339
rect 13553 11305 13587 11339
rect 21189 11305 21223 11339
rect 22385 11305 22419 11339
rect 7941 11237 7975 11271
rect 17233 11237 17267 11271
rect 4997 11169 5031 11203
rect 5733 11169 5767 11203
rect 5917 11169 5951 11203
rect 6745 11169 6779 11203
rect 6929 11169 6963 11203
rect 8953 11169 8987 11203
rect 9229 11169 9263 11203
rect 10701 11169 10735 11203
rect 11345 11169 11379 11203
rect 12817 11169 12851 11203
rect 15485 11169 15519 11203
rect 24225 11169 24259 11203
rect 26341 11169 26375 11203
rect 26617 11169 26651 11203
rect 28089 11169 28123 11203
rect 4721 11101 4755 11135
rect 5641 11101 5675 11135
rect 6101 11101 6135 11135
rect 6285 11101 6319 11135
rect 6561 11101 6595 11135
rect 7849 11101 7883 11135
rect 8033 11101 8067 11135
rect 11667 11101 11701 11135
rect 11897 11101 11931 11135
rect 12080 11101 12114 11135
rect 12173 11101 12207 11135
rect 12265 11101 12299 11135
rect 12357 11101 12391 11135
rect 12633 11101 12667 11135
rect 12725 11101 12759 11135
rect 14289 11101 14323 11135
rect 14381 11101 14415 11135
rect 14657 11101 14691 11135
rect 19533 11101 19567 11135
rect 20545 11101 20579 11135
rect 20638 11101 20672 11135
rect 20913 11101 20947 11135
rect 21051 11101 21085 11135
rect 21741 11101 21775 11135
rect 21834 11101 21868 11135
rect 22109 11101 22143 11135
rect 22247 11101 22281 11135
rect 6377 11033 6411 11067
rect 7757 11033 7791 11067
rect 11805 11033 11839 11067
rect 12541 11033 12575 11067
rect 13277 11033 13311 11067
rect 13537 11033 13571 11067
rect 13737 11033 13771 11067
rect 14473 11033 14507 11067
rect 15761 11033 15795 11067
rect 20821 11033 20855 11067
rect 22017 11033 22051 11067
rect 23949 11033 23983 11067
rect 4813 10965 4847 10999
rect 11529 10965 11563 10999
rect 13077 10965 13111 10999
rect 14105 10965 14139 10999
rect 22477 10965 22511 10999
rect 5457 10761 5491 10795
rect 6561 10761 6595 10795
rect 12173 10761 12207 10795
rect 15485 10761 15519 10795
rect 16297 10761 16331 10795
rect 24317 10761 24351 10795
rect 7021 10693 7055 10727
rect 8309 10693 8343 10727
rect 13461 10693 13495 10727
rect 15669 10693 15703 10727
rect 16497 10693 16531 10727
rect 22661 10693 22695 10727
rect 22753 10693 22787 10727
rect 26065 10693 26099 10727
rect 27261 10693 27295 10727
rect 27813 10693 27847 10727
rect 4997 10625 5031 10659
rect 5641 10625 5675 10659
rect 5733 10625 5767 10659
rect 5825 10625 5859 10659
rect 6009 10625 6043 10659
rect 6377 10625 6411 10659
rect 6561 10625 6595 10659
rect 6929 10625 6963 10659
rect 8033 10625 8067 10659
rect 10149 10625 10183 10659
rect 11805 10625 11839 10659
rect 12541 10625 12575 10659
rect 12633 10625 12667 10659
rect 13737 10625 13771 10659
rect 18797 10625 18831 10659
rect 19809 10625 19843 10659
rect 22385 10625 22419 10659
rect 22533 10625 22567 10659
rect 22891 10625 22925 10659
rect 23121 10625 23155 10659
rect 23949 10625 23983 10659
rect 24133 10625 24167 10659
rect 25237 10625 25271 10659
rect 27445 10625 27479 10659
rect 5089 10557 5123 10591
rect 5365 10557 5399 10591
rect 7849 10557 7883 10591
rect 10333 10557 10367 10591
rect 10425 10557 10459 10591
rect 10609 10557 10643 10591
rect 11161 10557 11195 10591
rect 11897 10557 11931 10591
rect 13461 10557 13495 10591
rect 13645 10557 13679 10591
rect 17049 10557 17083 10591
rect 18521 10557 18555 10591
rect 20085 10557 20119 10591
rect 23765 10557 23799 10591
rect 23857 10557 23891 10591
rect 9781 10489 9815 10523
rect 12817 10489 12851 10523
rect 16037 10489 16071 10523
rect 16129 10489 16163 10523
rect 23029 10489 23063 10523
rect 9965 10421 9999 10455
rect 15669 10421 15703 10455
rect 16313 10421 16347 10455
rect 21557 10421 21591 10455
rect 27077 10421 27111 10455
rect 27905 10421 27939 10455
rect 5457 10217 5491 10251
rect 14105 10217 14139 10251
rect 15669 10217 15703 10251
rect 16405 10217 16439 10251
rect 18429 10217 18463 10251
rect 18613 10217 18647 10251
rect 7665 10149 7699 10183
rect 6561 10081 6595 10115
rect 7021 10081 7055 10115
rect 7113 10081 7147 10115
rect 9229 10081 9263 10115
rect 14473 10081 14507 10115
rect 15853 10081 15887 10115
rect 18153 10081 18187 10115
rect 18245 10081 18279 10115
rect 19625 10081 19659 10115
rect 26525 10081 26559 10115
rect 26801 10081 26835 10115
rect 5273 10013 5307 10047
rect 5457 10013 5491 10047
rect 6653 10013 6687 10047
rect 6745 10013 6779 10047
rect 6929 10013 6963 10047
rect 7205 10013 7239 10047
rect 7665 10013 7699 10047
rect 7849 10013 7883 10047
rect 8953 10013 8987 10047
rect 12541 10013 12575 10047
rect 14289 10013 14323 10047
rect 15945 10013 15979 10047
rect 16037 10013 16071 10047
rect 16129 10013 16163 10047
rect 18521 10013 18555 10047
rect 18613 10013 18647 10047
rect 18797 10013 18831 10047
rect 20453 10013 20487 10047
rect 24593 10013 24627 10047
rect 26433 10013 26467 10047
rect 7389 9945 7423 9979
rect 7481 9945 7515 9979
rect 11805 9945 11839 9979
rect 17877 9945 17911 9979
rect 20545 9945 20579 9979
rect 20729 9945 20763 9979
rect 25329 9945 25363 9979
rect 10701 9877 10735 9911
rect 18245 9877 18279 9911
rect 20913 9877 20947 9911
rect 26341 9877 26375 9911
rect 28273 9877 28307 9911
rect 6377 9673 6411 9707
rect 7573 9673 7607 9707
rect 20085 9673 20119 9707
rect 12725 9605 12759 9639
rect 13093 9605 13127 9639
rect 14473 9605 14507 9639
rect 17509 9605 17543 9639
rect 17693 9605 17727 9639
rect 17877 9605 17911 9639
rect 19073 9605 19107 9639
rect 19289 9605 19323 9639
rect 19901 9605 19935 9639
rect 22753 9605 22787 9639
rect 6561 9537 6595 9571
rect 6837 9537 6871 9571
rect 7021 9537 7055 9571
rect 7113 9537 7147 9571
rect 7389 9537 7423 9571
rect 11897 9537 11931 9571
rect 12909 9537 12943 9571
rect 13001 9537 13035 9571
rect 13277 9537 13311 9571
rect 13369 9537 13403 9571
rect 14197 9537 14231 9571
rect 14289 9537 14323 9571
rect 14565 9537 14599 9571
rect 14749 9537 14783 9571
rect 17601 9537 17635 9571
rect 17969 9537 18003 9571
rect 20361 9537 20395 9571
rect 20545 9537 20579 9571
rect 21465 9537 21499 9571
rect 21925 9537 21959 9571
rect 24593 9537 24627 9571
rect 26065 9537 26099 9571
rect 26249 9537 26283 9571
rect 26341 9537 26375 9571
rect 26479 9537 26513 9571
rect 26801 9537 26835 9571
rect 27537 9537 27571 9571
rect 27905 9537 27939 9571
rect 28181 9537 28215 9571
rect 7205 9469 7239 9503
rect 13093 9469 13127 9503
rect 14105 9469 14139 9503
rect 14473 9469 14507 9503
rect 16865 9469 16899 9503
rect 18245 9469 18279 9503
rect 20453 9469 20487 9503
rect 20637 9469 20671 9503
rect 26617 9469 26651 9503
rect 27261 9469 27295 9503
rect 13461 9401 13495 9435
rect 17877 9401 17911 9435
rect 18153 9401 18187 9435
rect 19441 9401 19475 9435
rect 19533 9401 19567 9435
rect 26709 9401 26743 9435
rect 27629 9401 27663 9435
rect 7297 9333 7331 9367
rect 12725 9333 12759 9367
rect 14565 9333 14599 9367
rect 18061 9333 18095 9367
rect 19257 9333 19291 9367
rect 19901 9333 19935 9367
rect 20177 9333 20211 9367
rect 26065 9333 26099 9367
rect 26985 9333 27019 9367
rect 27169 9333 27203 9367
rect 27813 9333 27847 9367
rect 6745 9129 6779 9163
rect 14657 9129 14691 9163
rect 16681 9129 16715 9163
rect 20177 9129 20211 9163
rect 20637 9129 20671 9163
rect 26433 9129 26467 9163
rect 26893 9129 26927 9163
rect 10149 9061 10183 9095
rect 20269 9061 20303 9095
rect 24409 9061 24443 9095
rect 6561 8993 6595 9027
rect 7205 8993 7239 9027
rect 12357 8993 12391 9027
rect 15117 8993 15151 9027
rect 17049 8993 17083 9027
rect 19809 8993 19843 9027
rect 20913 8993 20947 9027
rect 22661 8993 22695 9027
rect 23397 8993 23431 9027
rect 25605 8993 25639 9027
rect 25881 8993 25915 9027
rect 25973 8993 26007 9027
rect 5641 8925 5675 8959
rect 6193 8925 6227 8959
rect 6377 8925 6411 8959
rect 6469 8925 6503 8959
rect 6653 8925 6687 8959
rect 7389 8925 7423 8959
rect 9597 8925 9631 8959
rect 9781 8925 9815 8959
rect 9873 8925 9907 8959
rect 9965 8925 9999 8959
rect 10425 8925 10459 8959
rect 10517 8925 10551 8959
rect 10793 8925 10827 8959
rect 10885 8925 10919 8959
rect 11437 8925 11471 8959
rect 12081 8925 12115 8959
rect 14841 8925 14875 8959
rect 15025 8925 15059 8959
rect 15209 8925 15243 8959
rect 15393 8925 15427 8959
rect 16865 8925 16899 8959
rect 19993 8925 20027 8959
rect 24225 8925 24259 8959
rect 25053 8925 25087 8959
rect 25789 8925 25823 8959
rect 26065 8925 26099 8959
rect 26249 8925 26283 8959
rect 26617 8925 26651 8959
rect 26709 8925 26743 8959
rect 27077 8925 27111 8959
rect 27353 8925 27387 8959
rect 27537 8925 27571 8959
rect 6929 8857 6963 8891
rect 7113 8857 7147 8891
rect 10609 8857 10643 8891
rect 21189 8857 21223 8891
rect 24133 8857 24167 8891
rect 24777 8857 24811 8891
rect 24961 8857 24995 8891
rect 25145 8857 25179 8891
rect 27261 8857 27295 8891
rect 5089 8789 5123 8823
rect 6285 8789 6319 8823
rect 7573 8789 7607 8823
rect 10241 8789 10275 8823
rect 13829 8789 13863 8823
rect 15209 8789 15243 8823
rect 20637 8789 20671 8823
rect 20821 8789 20855 8823
rect 22845 8789 22879 8823
rect 24593 8789 24627 8823
rect 24685 8789 24719 8823
rect 27721 8789 27755 8823
rect 4813 8585 4847 8619
rect 5273 8585 5307 8619
rect 6745 8585 6779 8619
rect 8401 8585 8435 8619
rect 10793 8585 10827 8619
rect 14749 8585 14783 8619
rect 20545 8585 20579 8619
rect 21103 8585 21137 8619
rect 21925 8585 21959 8619
rect 23949 8585 23983 8619
rect 9321 8517 9355 8551
rect 12725 8517 12759 8551
rect 14473 8517 14507 8551
rect 15117 8517 15151 8551
rect 16957 8517 16991 8551
rect 17049 8517 17083 8551
rect 19717 8517 19751 8551
rect 20177 8517 20211 8551
rect 20377 8517 20411 8551
rect 20637 8517 20671 8551
rect 21005 8517 21039 8551
rect 21189 8517 21223 8551
rect 3065 8449 3099 8483
rect 6561 8449 6595 8483
rect 6837 8449 6871 8483
rect 6929 8449 6963 8483
rect 7021 8449 7055 8483
rect 7113 8449 7147 8483
rect 7297 8449 7331 8483
rect 8309 8449 8343 8483
rect 14289 8449 14323 8483
rect 14933 8449 14967 8483
rect 15025 8449 15059 8483
rect 15301 8449 15335 8483
rect 15393 8449 15427 8483
rect 15577 8449 15611 8483
rect 15669 8449 15703 8483
rect 15945 8449 15979 8483
rect 16865 8449 16899 8483
rect 17233 8449 17267 8483
rect 17509 8449 17543 8483
rect 17601 8449 17635 8483
rect 17693 8449 17727 8483
rect 17877 8449 17911 8483
rect 20085 8449 20119 8483
rect 20913 8449 20947 8483
rect 21281 8449 21315 8483
rect 23857 8449 23891 8483
rect 24041 8449 24075 8483
rect 24133 8449 24167 8483
rect 24593 8449 24627 8483
rect 25237 8449 25271 8483
rect 25329 8449 25363 8483
rect 25697 8449 25731 8483
rect 25789 8449 25823 8483
rect 25973 8449 26007 8483
rect 26065 8449 26099 8483
rect 3341 8381 3375 8415
rect 5365 8381 5399 8415
rect 5457 8381 5491 8415
rect 6377 8381 6411 8415
rect 9045 8381 9079 8415
rect 12449 8381 12483 8415
rect 14197 8381 14231 8415
rect 15761 8381 15795 8415
rect 20637 8381 20671 8415
rect 23397 8381 23431 8415
rect 23673 8381 23707 8415
rect 24409 8381 24443 8415
rect 24869 8381 24903 8415
rect 25053 8381 25087 8415
rect 25145 8381 25179 8415
rect 4905 8313 4939 8347
rect 20821 8313 20855 8347
rect 25513 8313 25547 8347
rect 7297 8245 7331 8279
rect 14657 8245 14691 8279
rect 16129 8245 16163 8279
rect 16681 8245 16715 8279
rect 17325 8245 17359 8279
rect 19533 8245 19567 8279
rect 19717 8245 19751 8279
rect 20361 8245 20395 8279
rect 24317 8245 24351 8279
rect 24777 8245 24811 8279
rect 5181 8041 5215 8075
rect 7205 8041 7239 8075
rect 10057 8041 10091 8075
rect 14749 8041 14783 8075
rect 15945 8041 15979 8075
rect 16313 8041 16347 8075
rect 19809 8041 19843 8075
rect 25053 8041 25087 8075
rect 26157 8041 26191 8075
rect 26341 8041 26375 8075
rect 6009 7973 6043 8007
rect 10885 7973 10919 8007
rect 24133 7973 24167 8007
rect 25789 7973 25823 8007
rect 26433 7973 26467 8007
rect 6469 7905 6503 7939
rect 9137 7905 9171 7939
rect 11345 7905 11379 7939
rect 15209 7905 15243 7939
rect 17049 7905 17083 7939
rect 24225 7905 24259 7939
rect 24593 7905 24627 7939
rect 24870 7905 24904 7939
rect 25237 7905 25271 7939
rect 26065 7905 26099 7939
rect 4629 7837 4663 7871
rect 4813 7837 4847 7871
rect 4997 7837 5031 7871
rect 5917 7837 5951 7871
rect 6377 7837 6411 7871
rect 6837 7837 6871 7871
rect 7021 7837 7055 7871
rect 7113 7837 7147 7871
rect 7573 7837 7607 7871
rect 9321 7837 9355 7871
rect 9597 7837 9631 7871
rect 9873 7837 9907 7871
rect 10333 7837 10367 7871
rect 10609 7837 10643 7871
rect 10793 7837 10827 7871
rect 11161 7837 11195 7871
rect 11253 7837 11287 7871
rect 11437 7837 11471 7871
rect 14933 7837 14967 7871
rect 15025 7837 15059 7871
rect 15301 7837 15335 7871
rect 16129 7837 16163 7871
rect 16405 7837 16439 7871
rect 16589 7837 16623 7871
rect 16773 7837 16807 7871
rect 16957 7837 16991 7871
rect 17141 7837 17175 7871
rect 17325 7837 17359 7871
rect 18061 7837 18095 7871
rect 18521 7837 18555 7871
rect 18613 7837 18647 7871
rect 18889 7837 18923 7871
rect 19349 7837 19383 7871
rect 19441 7837 19475 7871
rect 19625 7837 19659 7871
rect 23765 7837 23799 7871
rect 24685 7837 24719 7871
rect 24777 7837 24811 7871
rect 25329 7837 25363 7871
rect 26157 7837 26191 7871
rect 26525 7837 26559 7871
rect 28365 7837 28399 7871
rect 4905 7769 4939 7803
rect 7389 7769 7423 7803
rect 10885 7769 10919 7803
rect 17877 7769 17911 7803
rect 18245 7769 18279 7803
rect 18705 7769 18739 7803
rect 25053 7769 25087 7803
rect 26249 7769 26283 7803
rect 5273 7701 5307 7735
rect 6653 7701 6687 7735
rect 9505 7701 9539 7735
rect 9689 7701 9723 7735
rect 10149 7701 10183 7735
rect 11069 7701 11103 7735
rect 18337 7701 18371 7735
rect 24409 7701 24443 7735
rect 25513 7701 25547 7735
rect 28181 7701 28215 7735
rect 4997 7497 5031 7531
rect 5457 7497 5491 7531
rect 5549 7497 5583 7531
rect 6377 7497 6411 7531
rect 7205 7497 7239 7531
rect 10609 7497 10643 7531
rect 17601 7497 17635 7531
rect 21649 7497 21683 7531
rect 26525 7497 26559 7531
rect 12127 7429 12161 7463
rect 12357 7429 12391 7463
rect 18429 7429 18463 7463
rect 19165 7429 19199 7463
rect 19257 7429 19291 7463
rect 20177 7429 20211 7463
rect 25697 7429 25731 7463
rect 6561 7361 6595 7395
rect 6653 7361 6687 7395
rect 7113 7361 7147 7395
rect 7297 7361 7331 7395
rect 10977 7361 11011 7395
rect 11989 7361 12023 7395
rect 12265 7361 12299 7395
rect 12449 7361 12483 7395
rect 13093 7361 13127 7395
rect 17785 7361 17819 7395
rect 17969 7361 18003 7395
rect 18061 7361 18095 7395
rect 18291 7361 18325 7395
rect 18521 7361 18555 7395
rect 18704 7361 18738 7395
rect 18797 7361 18831 7395
rect 19073 7361 19107 7395
rect 19441 7361 19475 7395
rect 24225 7361 24259 7395
rect 24409 7361 24443 7395
rect 25881 7361 25915 7395
rect 26157 7361 26191 7395
rect 26341 7361 26375 7395
rect 26433 7361 26467 7395
rect 26617 7361 26651 7395
rect 28365 7361 28399 7395
rect 3249 7293 3283 7327
rect 3525 7293 3559 7327
rect 5641 7293 5675 7327
rect 6929 7293 6963 7327
rect 7021 7293 7055 7327
rect 8769 7293 8803 7327
rect 9045 7293 9079 7327
rect 10517 7293 10551 7327
rect 10885 7293 10919 7327
rect 12633 7293 12667 7327
rect 13001 7293 13035 7327
rect 19901 7293 19935 7327
rect 24685 7293 24719 7327
rect 26065 7293 26099 7327
rect 5089 7225 5123 7259
rect 18889 7225 18923 7259
rect 12725 7157 12759 7191
rect 18153 7157 18187 7191
rect 24409 7157 24443 7191
rect 26157 7157 26191 7191
rect 28181 7157 28215 7191
rect 9597 6953 9631 6987
rect 10517 6953 10551 6987
rect 11437 6953 11471 6987
rect 12160 6953 12194 6987
rect 14289 6953 14323 6987
rect 18429 6953 18463 6987
rect 18889 6953 18923 6987
rect 28009 6953 28043 6987
rect 11345 6885 11379 6919
rect 10149 6817 10183 6851
rect 10977 6817 11011 6851
rect 17877 6817 17911 6851
rect 9778 6749 9812 6783
rect 10241 6749 10275 6783
rect 10609 6749 10643 6783
rect 10701 6749 10735 6783
rect 11161 6749 11195 6783
rect 11437 6749 11471 6783
rect 11529 6749 11563 6783
rect 11897 6749 11931 6783
rect 14105 6749 14139 6783
rect 18061 6749 18095 6783
rect 18613 6749 18647 6783
rect 18705 6749 18739 6783
rect 18981 6749 19015 6783
rect 28273 6749 28307 6783
rect 18245 6681 18279 6715
rect 23857 6681 23891 6715
rect 9781 6613 9815 6647
rect 10333 6613 10367 6647
rect 11805 6613 11839 6647
rect 13645 6613 13679 6647
rect 23949 6613 23983 6647
rect 26525 6613 26559 6647
rect 12265 6409 12299 6443
rect 12725 6409 12759 6443
rect 17969 6409 18003 6443
rect 23581 6409 23615 6443
rect 24869 6409 24903 6443
rect 27169 6409 27203 6443
rect 13461 6341 13495 6375
rect 15301 6341 15335 6375
rect 16865 6341 16899 6375
rect 17141 6341 17175 6375
rect 17325 6341 17359 6375
rect 11897 6273 11931 6307
rect 11989 6273 12023 6307
rect 12633 6273 12667 6307
rect 16037 6273 16071 6307
rect 16129 6273 16163 6307
rect 16221 6273 16255 6307
rect 16405 6273 16439 6307
rect 17049 6273 17083 6307
rect 18153 6273 18187 6307
rect 18337 6273 18371 6307
rect 23857 6273 23891 6307
rect 24041 6273 24075 6307
rect 24133 6273 24167 6307
rect 24317 6273 24351 6307
rect 24593 6273 24627 6307
rect 24777 6273 24811 6307
rect 26157 6273 26191 6307
rect 26249 6273 26283 6307
rect 26433 6273 26467 6307
rect 27353 6273 27387 6307
rect 27629 6273 27663 6307
rect 28365 6273 28399 6307
rect 12173 6205 12207 6239
rect 12909 6205 12943 6239
rect 21833 6205 21867 6239
rect 22109 6205 22143 6239
rect 23673 6205 23707 6239
rect 27537 6205 27571 6239
rect 12081 6137 12115 6171
rect 15577 6137 15611 6171
rect 15853 6137 15887 6171
rect 16681 6137 16715 6171
rect 23949 6137 23983 6171
rect 25973 6137 26007 6171
rect 28181 6137 28215 6171
rect 13185 6069 13219 6103
rect 15761 6069 15795 6103
rect 24501 6069 24535 6103
rect 26157 6069 26191 6103
rect 27537 6069 27571 6103
rect 17049 5865 17083 5899
rect 17417 5865 17451 5899
rect 22937 5865 22971 5899
rect 25881 5865 25915 5899
rect 26433 5865 26467 5899
rect 14749 5797 14783 5831
rect 15485 5797 15519 5831
rect 23581 5797 23615 5831
rect 6745 5729 6779 5763
rect 16681 5729 16715 5763
rect 17509 5729 17543 5763
rect 21465 5729 21499 5763
rect 23305 5729 23339 5763
rect 24777 5729 24811 5763
rect 27997 5729 28031 5763
rect 6009 5661 6043 5695
rect 6193 5661 6227 5695
rect 6285 5661 6319 5695
rect 6469 5661 6503 5695
rect 6929 5661 6963 5695
rect 14933 5661 14967 5695
rect 15209 5661 15243 5695
rect 15301 5661 15335 5695
rect 16129 5661 16163 5695
rect 16589 5661 16623 5695
rect 17049 5661 17083 5695
rect 17325 5661 17359 5695
rect 17693 5661 17727 5695
rect 21189 5661 21223 5695
rect 23489 5661 23523 5695
rect 23673 5661 23707 5695
rect 23765 5661 23799 5695
rect 23949 5661 23983 5695
rect 24593 5661 24627 5695
rect 24685 5661 24719 5695
rect 24869 5661 24903 5695
rect 25053 5661 25087 5695
rect 25329 5661 25363 5695
rect 25605 5661 25639 5695
rect 25973 5661 26007 5695
rect 26065 5661 26099 5695
rect 28273 5661 28307 5695
rect 25145 5593 25179 5627
rect 25513 5593 25547 5627
rect 26249 5593 26283 5627
rect 6101 5525 6135 5559
rect 6653 5525 6687 5559
rect 7113 5525 7147 5559
rect 15117 5525 15151 5559
rect 16865 5525 16899 5559
rect 24409 5525 24443 5559
rect 26525 5525 26559 5559
rect 6469 5321 6503 5355
rect 15393 5321 15427 5355
rect 15761 5321 15795 5355
rect 17233 5321 17267 5355
rect 18429 5321 18463 5355
rect 19073 5321 19107 5355
rect 19901 5321 19935 5355
rect 21833 5321 21867 5355
rect 24317 5321 24351 5355
rect 25697 5321 25731 5355
rect 28181 5321 28215 5355
rect 7389 5253 7423 5287
rect 8217 5253 8251 5287
rect 9505 5253 9539 5287
rect 9623 5253 9657 5287
rect 16405 5253 16439 5287
rect 16865 5253 16899 5287
rect 17877 5253 17911 5287
rect 19809 5253 19843 5287
rect 23305 5253 23339 5287
rect 6009 5185 6043 5219
rect 6377 5185 6411 5219
rect 6653 5185 6687 5219
rect 6903 5185 6937 5219
rect 7021 5185 7055 5219
rect 7113 5185 7147 5219
rect 7205 5185 7239 5219
rect 7665 5185 7699 5219
rect 8033 5185 8067 5219
rect 8309 5185 8343 5219
rect 8401 5185 8435 5219
rect 8585 5185 8619 5219
rect 8861 5185 8895 5219
rect 9321 5185 9355 5219
rect 9413 5185 9447 5219
rect 12909 5185 12943 5219
rect 13093 5185 13127 5219
rect 15301 5185 15335 5219
rect 15577 5185 15611 5219
rect 16037 5185 16071 5219
rect 16313 5185 16347 5219
rect 16681 5185 16715 5219
rect 16957 5185 16991 5219
rect 17049 5185 17083 5219
rect 18061 5185 18095 5219
rect 18153 5185 18187 5219
rect 18613 5185 18647 5219
rect 18797 5185 18831 5219
rect 18889 5185 18923 5219
rect 19349 5185 19383 5219
rect 24593 5185 24627 5219
rect 24777 5185 24811 5219
rect 25053 5185 25087 5219
rect 25329 5185 25363 5219
rect 25881 5185 25915 5219
rect 26525 5185 26559 5219
rect 26617 5185 26651 5219
rect 28365 5185 28399 5219
rect 3341 5117 3375 5151
rect 3617 5117 3651 5151
rect 5825 5117 5859 5151
rect 5917 5117 5951 5151
rect 6101 5117 6135 5151
rect 6745 5117 6779 5151
rect 7941 5117 7975 5151
rect 8677 5117 8711 5151
rect 9781 5117 9815 5151
rect 15669 5117 15703 5151
rect 16221 5117 16255 5151
rect 18694 5117 18728 5151
rect 19257 5117 19291 5151
rect 19441 5117 19475 5151
rect 19533 5117 19567 5151
rect 23581 5117 23615 5151
rect 23673 5117 23707 5151
rect 24869 5117 24903 5151
rect 25605 5117 25639 5151
rect 26157 5117 26191 5151
rect 26249 5117 26283 5151
rect 26433 5117 26467 5151
rect 5641 5049 5675 5083
rect 6653 5049 6687 5083
rect 8493 5049 8527 5083
rect 9045 5049 9079 5083
rect 15577 5049 15611 5083
rect 17877 5049 17911 5083
rect 24685 5049 24719 5083
rect 25145 5049 25179 5083
rect 5089 4981 5123 5015
rect 7481 4981 7515 5015
rect 7849 4981 7883 5015
rect 8125 4981 8159 5015
rect 9137 4981 9171 5015
rect 13001 4981 13035 5015
rect 24409 4981 24443 5015
rect 25513 4981 25547 5015
rect 26065 4981 26099 5015
rect 4721 4777 4755 4811
rect 5181 4777 5215 4811
rect 6101 4777 6135 4811
rect 6285 4777 6319 4811
rect 6745 4777 6779 4811
rect 7757 4777 7791 4811
rect 9137 4777 9171 4811
rect 10425 4777 10459 4811
rect 13553 4777 13587 4811
rect 16129 4777 16163 4811
rect 16405 4777 16439 4811
rect 16681 4777 16715 4811
rect 18337 4777 18371 4811
rect 18521 4777 18555 4811
rect 23581 4777 23615 4811
rect 25973 4777 26007 4811
rect 26525 4777 26559 4811
rect 6653 4709 6687 4743
rect 7205 4709 7239 4743
rect 8217 4709 8251 4743
rect 5733 4641 5767 4675
rect 6837 4641 6871 4675
rect 8493 4641 8527 4675
rect 8585 4641 8619 4675
rect 10517 4641 10551 4675
rect 13001 4641 13035 4675
rect 15761 4641 15795 4675
rect 16497 4641 16531 4675
rect 22569 4641 22603 4675
rect 22845 4641 22879 4675
rect 27997 4641 28031 4675
rect 4905 4573 4939 4607
rect 4997 4573 5031 4607
rect 5273 4573 5307 4607
rect 5549 4573 5583 4607
rect 6377 4573 6411 4607
rect 6469 4573 6503 4607
rect 6561 4573 6595 4607
rect 7021 4573 7055 4607
rect 7481 4573 7515 4607
rect 7849 4573 7883 4607
rect 8125 4573 8159 4607
rect 8401 4573 8435 4607
rect 8677 4573 8711 4607
rect 9051 4573 9085 4607
rect 9229 4573 9263 4607
rect 9505 4573 9539 4607
rect 9597 4573 9631 4607
rect 10241 4573 10275 4607
rect 10701 4573 10735 4607
rect 10793 4573 10827 4607
rect 11989 4573 12023 4607
rect 12173 4573 12207 4607
rect 12449 4551 12483 4585
rect 12541 4573 12575 4607
rect 12633 4573 12667 4607
rect 12817 4573 12851 4607
rect 12909 4573 12943 4607
rect 13185 4573 13219 4607
rect 13461 4573 13495 4607
rect 13645 4573 13679 4607
rect 13737 4573 13771 4607
rect 13921 4573 13955 4607
rect 15853 4573 15887 4607
rect 16221 4573 16255 4607
rect 16405 4573 16439 4607
rect 16773 4573 16807 4607
rect 17049 4573 17083 4607
rect 17233 4573 17267 4607
rect 18429 4573 18463 4607
rect 18889 4573 18923 4607
rect 19625 4573 19659 4607
rect 20177 4573 20211 4607
rect 20453 4573 20487 4607
rect 22937 4573 22971 4607
rect 25973 4573 26007 4607
rect 26157 4573 26191 4607
rect 26249 4573 26283 4607
rect 26433 4573 26467 4607
rect 28273 4573 28307 4607
rect 5365 4505 5399 4539
rect 7389 4505 7423 4539
rect 9321 4505 9355 4539
rect 10057 4505 10091 4539
rect 12081 4505 12115 4539
rect 13369 4505 13403 4539
rect 18705 4505 18739 4539
rect 19257 4505 19291 4539
rect 19809 4505 19843 4539
rect 7573 4437 7607 4471
rect 9965 4437 9999 4471
rect 12265 4437 12299 4471
rect 13829 4437 13863 4471
rect 16865 4437 16899 4471
rect 19441 4437 19475 4471
rect 19533 4437 19567 4471
rect 19993 4437 20027 4471
rect 20269 4437 20303 4471
rect 21097 4437 21131 4471
rect 26341 4437 26375 4471
rect 6193 4233 6227 4267
rect 8493 4233 8527 4267
rect 9229 4233 9263 4267
rect 16497 4233 16531 4267
rect 17693 4233 17727 4267
rect 20545 4233 20579 4267
rect 26065 4233 26099 4267
rect 27445 4233 27479 4267
rect 6745 4165 6779 4199
rect 9597 4165 9631 4199
rect 9965 4165 9999 4199
rect 11989 4165 12023 4199
rect 12199 4165 12233 4199
rect 12771 4165 12805 4199
rect 12909 4165 12943 4199
rect 13001 4165 13035 4199
rect 14105 4165 14139 4199
rect 16037 4165 16071 4199
rect 18337 4165 18371 4199
rect 19257 4165 19291 4199
rect 26709 4165 26743 4199
rect 26985 4165 27019 4199
rect 6009 4097 6043 4131
rect 6377 4097 6411 4131
rect 7021 4097 7055 4131
rect 7113 4097 7147 4131
rect 7297 4097 7331 4131
rect 8493 4097 8527 4131
rect 8677 4097 8711 4131
rect 9137 4097 9171 4131
rect 9781 4097 9815 4131
rect 10701 4097 10735 4131
rect 11897 4097 11931 4131
rect 12081 4097 12115 4131
rect 13093 4097 13127 4131
rect 13737 4097 13771 4131
rect 13829 4097 13863 4131
rect 13921 4097 13955 4131
rect 14381 4097 14415 4131
rect 14565 4097 14599 4131
rect 16313 4097 16347 4131
rect 16681 4097 16715 4131
rect 16957 4097 16991 4131
rect 17325 4097 17359 4131
rect 17969 4097 18003 4131
rect 18797 4097 18831 4131
rect 19165 4097 19199 4131
rect 19993 4097 20027 4131
rect 20085 4097 20119 4131
rect 20269 4097 20303 4131
rect 20637 4097 20671 4131
rect 21005 4097 21039 4131
rect 23029 4097 23063 4131
rect 25605 4097 25639 4131
rect 25881 4097 25915 4131
rect 26249 4097 26283 4131
rect 27261 4097 27295 4131
rect 27537 4097 27571 4131
rect 27905 4097 27939 4131
rect 5825 4029 5859 4063
rect 9321 4029 9355 4063
rect 10425 4029 10459 4063
rect 10609 4029 10643 4063
rect 11713 4029 11747 4063
rect 12357 4029 12391 4063
rect 12633 4029 12667 4063
rect 13461 4029 13495 4063
rect 13553 4029 13587 4063
rect 14289 4029 14323 4063
rect 16129 4029 16163 4063
rect 16865 4029 16899 4063
rect 17049 4029 17083 4063
rect 17141 4029 17175 4063
rect 17877 4029 17911 4063
rect 18245 4029 18279 4063
rect 18613 4029 18647 4063
rect 18705 4029 18739 4063
rect 18889 4029 18923 4063
rect 20453 4029 20487 4063
rect 23305 4029 23339 4063
rect 25421 4029 25455 4063
rect 25697 4029 25731 4063
rect 25789 4029 25823 4063
rect 26433 4029 26467 4063
rect 27077 4029 27111 4063
rect 13369 3961 13403 3995
rect 14473 3961 14507 3995
rect 20269 3961 20303 3995
rect 27721 3961 27755 3995
rect 28089 3961 28123 3995
rect 6745 3893 6779 3927
rect 6929 3893 6963 3927
rect 7481 3893 7515 3927
rect 8769 3893 8803 3927
rect 11069 3893 11103 3927
rect 13277 3893 13311 3927
rect 16313 3893 16347 3927
rect 18429 3893 18463 3927
rect 20821 3893 20855 3927
rect 24777 3893 24811 3927
rect 26249 3893 26283 3927
rect 26985 3893 27019 3927
rect 4813 3689 4847 3723
rect 6303 3689 6337 3723
rect 7389 3689 7423 3723
rect 9413 3689 9447 3723
rect 13737 3689 13771 3723
rect 16957 3689 16991 3723
rect 17141 3689 17175 3723
rect 17509 3689 17543 3723
rect 18613 3689 18647 3723
rect 19257 3689 19291 3723
rect 20177 3689 20211 3723
rect 23121 3689 23155 3723
rect 23581 3689 23615 3723
rect 26433 3689 26467 3723
rect 26525 3689 26559 3723
rect 7849 3621 7883 3655
rect 16221 3621 16255 3655
rect 25697 3621 25731 3655
rect 6653 3553 6687 3587
rect 7297 3553 7331 3587
rect 10885 3553 10919 3587
rect 11161 3553 11195 3587
rect 11529 3553 11563 3587
rect 11989 3553 12023 3587
rect 14657 3553 14691 3587
rect 17785 3553 17819 3587
rect 19073 3553 19107 3587
rect 19717 3553 19751 3587
rect 19809 3553 19843 3587
rect 28273 3553 28307 3587
rect 6561 3485 6595 3519
rect 7573 3485 7607 3519
rect 7665 3485 7699 3519
rect 7941 3485 7975 3519
rect 11437 3485 11471 3519
rect 15209 3485 15243 3519
rect 15393 3485 15427 3519
rect 15485 3485 15519 3519
rect 15945 3485 15979 3519
rect 16586 3485 16620 3519
rect 17049 3485 17083 3519
rect 17325 3485 17359 3519
rect 17601 3485 17635 3519
rect 17693 3485 17727 3519
rect 17877 3485 17911 3519
rect 18797 3485 18831 3519
rect 18981 3485 19015 3519
rect 20177 3485 20211 3519
rect 20545 3485 20579 3519
rect 21281 3485 21315 3519
rect 23305 3485 23339 3519
rect 23397 3485 23431 3519
rect 25329 3485 25363 3519
rect 25513 3485 25547 3519
rect 26249 3485 26283 3519
rect 12265 3417 12299 3451
rect 15025 3417 15059 3451
rect 15669 3417 15703 3451
rect 21557 3417 21591 3451
rect 23121 3417 23155 3451
rect 24869 3417 24903 3451
rect 25421 3417 25455 3451
rect 25697 3417 25731 3451
rect 26157 3417 26191 3451
rect 27997 3417 28031 3451
rect 11805 3349 11839 3383
rect 14105 3349 14139 3383
rect 15761 3349 15795 3383
rect 16405 3349 16439 3383
rect 16589 3349 16623 3383
rect 19625 3349 19659 3383
rect 23029 3349 23063 3383
rect 24593 3349 24627 3383
rect 12449 3145 12483 3179
rect 12909 3145 12943 3179
rect 13369 3145 13403 3179
rect 16405 3145 16439 3179
rect 16773 3145 16807 3179
rect 19257 3145 19291 3179
rect 19533 3145 19567 3179
rect 23581 3145 23615 3179
rect 25421 3145 25455 3179
rect 26433 3145 26467 3179
rect 27721 3145 27755 3179
rect 8493 3077 8527 3111
rect 12817 3077 12851 3111
rect 14473 3077 14507 3111
rect 17049 3077 17083 3111
rect 28181 3077 28215 3111
rect 6561 3009 6595 3043
rect 8217 3009 8251 3043
rect 12357 3009 12391 3043
rect 13645 3009 13679 3043
rect 16681 3009 16715 3043
rect 16865 3009 16899 3043
rect 16957 3009 16991 3043
rect 17141 3009 17175 3043
rect 18981 3009 19015 3043
rect 19165 3009 19199 3043
rect 19441 3009 19475 3043
rect 19747 3009 19781 3043
rect 19901 3009 19935 3043
rect 21833 3009 21867 3043
rect 23673 3009 23707 3043
rect 25789 3009 25823 3043
rect 25881 3009 25915 3043
rect 26249 3009 26283 3043
rect 27537 3009 27571 3043
rect 6653 2941 6687 2975
rect 6929 2941 6963 2975
rect 9965 2941 9999 2975
rect 13093 2941 13127 2975
rect 14197 2941 14231 2975
rect 15945 2941 15979 2975
rect 22109 2941 22143 2975
rect 12265 2873 12299 2907
rect 16313 2873 16347 2907
rect 27905 2873 27939 2907
rect 23936 2805 23970 2839
rect 26249 2805 26283 2839
rect 21557 2601 21591 2635
rect 22201 2601 22235 2635
rect 22845 2601 22879 2635
rect 23489 2601 23523 2635
rect 21373 2397 21407 2431
rect 22017 2397 22051 2431
rect 22661 2397 22695 2431
rect 23305 2397 23339 2431
<< metal1 >>
rect 1104 29402 28704 29424
rect 1104 29350 4874 29402
rect 4926 29350 4938 29402
rect 4990 29350 5002 29402
rect 5054 29350 5066 29402
rect 5118 29350 5130 29402
rect 5182 29350 28704 29402
rect 1104 29328 28704 29350
rect 1104 28858 28704 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 28704 28858
rect 1104 28784 28704 28806
rect 1104 28314 28704 28336
rect 1104 28262 4874 28314
rect 4926 28262 4938 28314
rect 4990 28262 5002 28314
rect 5054 28262 5066 28314
rect 5118 28262 5130 28314
rect 5182 28262 28704 28314
rect 1104 28240 28704 28262
rect 1104 27770 28704 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 28704 27770
rect 1104 27696 28704 27718
rect 1104 27226 28704 27248
rect 1104 27174 4874 27226
rect 4926 27174 4938 27226
rect 4990 27174 5002 27226
rect 5054 27174 5066 27226
rect 5118 27174 5130 27226
rect 5182 27174 28704 27226
rect 1104 27152 28704 27174
rect 1104 26682 28704 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 28704 26682
rect 1104 26608 28704 26630
rect 1104 26138 28704 26160
rect 1104 26086 4874 26138
rect 4926 26086 4938 26138
rect 4990 26086 5002 26138
rect 5054 26086 5066 26138
rect 5118 26086 5130 26138
rect 5182 26086 28704 26138
rect 1104 26064 28704 26086
rect 15381 25959 15439 25965
rect 8128 25928 9536 25956
rect 7834 25848 7840 25900
rect 7892 25888 7898 25900
rect 8128 25897 8156 25928
rect 8113 25891 8171 25897
rect 8113 25888 8125 25891
rect 7892 25860 8125 25888
rect 7892 25848 7898 25860
rect 8113 25857 8125 25860
rect 8159 25857 8171 25891
rect 8113 25851 8171 25857
rect 8205 25891 8263 25897
rect 8205 25857 8217 25891
rect 8251 25857 8263 25891
rect 8205 25851 8263 25857
rect 8389 25891 8447 25897
rect 8389 25857 8401 25891
rect 8435 25888 8447 25891
rect 8570 25888 8576 25900
rect 8435 25860 8576 25888
rect 8435 25857 8447 25860
rect 8389 25851 8447 25857
rect 8220 25820 8248 25851
rect 8570 25848 8576 25860
rect 8628 25848 8634 25900
rect 9508 25897 9536 25928
rect 15381 25925 15393 25959
rect 15427 25956 15439 25959
rect 17313 25959 17371 25965
rect 17313 25956 17325 25959
rect 15427 25928 17325 25956
rect 15427 25925 15439 25928
rect 15381 25919 15439 25925
rect 17313 25925 17325 25928
rect 17359 25956 17371 25959
rect 17770 25956 17776 25968
rect 17359 25928 17776 25956
rect 17359 25925 17371 25928
rect 17313 25919 17371 25925
rect 17770 25916 17776 25928
rect 17828 25916 17834 25968
rect 22830 25916 22836 25968
rect 22888 25956 22894 25968
rect 22888 25928 24794 25956
rect 22888 25916 22894 25928
rect 9493 25891 9551 25897
rect 9493 25857 9505 25891
rect 9539 25857 9551 25891
rect 9493 25851 9551 25857
rect 9582 25848 9588 25900
rect 9640 25848 9646 25900
rect 9769 25891 9827 25897
rect 9769 25857 9781 25891
rect 9815 25888 9827 25891
rect 10318 25888 10324 25900
rect 9815 25860 10324 25888
rect 9815 25857 9827 25860
rect 9769 25851 9827 25857
rect 10318 25848 10324 25860
rect 10376 25848 10382 25900
rect 15286 25848 15292 25900
rect 15344 25848 15350 25900
rect 15565 25891 15623 25897
rect 15565 25857 15577 25891
rect 15611 25888 15623 25891
rect 17678 25888 17684 25900
rect 15611 25860 17684 25888
rect 15611 25857 15623 25860
rect 15565 25851 15623 25857
rect 17678 25848 17684 25860
rect 17736 25848 17742 25900
rect 20073 25891 20131 25897
rect 20073 25857 20085 25891
rect 20119 25888 20131 25891
rect 20625 25891 20683 25897
rect 20625 25888 20637 25891
rect 20119 25860 20637 25888
rect 20119 25857 20131 25860
rect 20073 25851 20131 25857
rect 20625 25857 20637 25860
rect 20671 25857 20683 25891
rect 20625 25851 20683 25857
rect 8938 25820 8944 25832
rect 8220 25792 8944 25820
rect 8938 25780 8944 25792
rect 8996 25780 9002 25832
rect 11974 25780 11980 25832
rect 12032 25820 12038 25832
rect 12069 25823 12127 25829
rect 12069 25820 12081 25823
rect 12032 25792 12081 25820
rect 12032 25780 12038 25792
rect 12069 25789 12081 25792
rect 12115 25789 12127 25823
rect 12069 25783 12127 25789
rect 16209 25823 16267 25829
rect 16209 25789 16221 25823
rect 16255 25789 16267 25823
rect 16209 25783 16267 25789
rect 16761 25823 16819 25829
rect 16761 25789 16773 25823
rect 16807 25820 16819 25823
rect 16942 25820 16948 25832
rect 16807 25792 16948 25820
rect 16807 25789 16819 25792
rect 16761 25783 16819 25789
rect 15565 25755 15623 25761
rect 15565 25721 15577 25755
rect 15611 25752 15623 25755
rect 16224 25752 16252 25783
rect 16942 25780 16948 25792
rect 17000 25780 17006 25832
rect 20165 25823 20223 25829
rect 20165 25789 20177 25823
rect 20211 25789 20223 25823
rect 20165 25783 20223 25789
rect 15611 25724 16252 25752
rect 20180 25752 20208 25783
rect 21174 25780 21180 25832
rect 21232 25780 21238 25832
rect 23290 25780 23296 25832
rect 23348 25780 23354 25832
rect 23569 25823 23627 25829
rect 23569 25789 23581 25823
rect 23615 25820 23627 25823
rect 24026 25820 24032 25832
rect 23615 25792 24032 25820
rect 23615 25789 23627 25792
rect 23569 25783 23627 25789
rect 24026 25780 24032 25792
rect 24084 25780 24090 25832
rect 24302 25780 24308 25832
rect 24360 25780 24366 25832
rect 21450 25752 21456 25764
rect 20180 25724 21456 25752
rect 15611 25721 15623 25724
rect 15565 25715 15623 25721
rect 21450 25712 21456 25724
rect 21508 25712 21514 25764
rect 5534 25644 5540 25696
rect 5592 25644 5598 25696
rect 8386 25644 8392 25696
rect 8444 25644 8450 25696
rect 9766 25644 9772 25696
rect 9824 25644 9830 25696
rect 11054 25644 11060 25696
rect 11112 25684 11118 25696
rect 11517 25687 11575 25693
rect 11517 25684 11529 25687
rect 11112 25656 11529 25684
rect 11112 25644 11118 25656
rect 11517 25653 11529 25656
rect 11563 25653 11575 25687
rect 11517 25647 11575 25653
rect 15470 25644 15476 25696
rect 15528 25684 15534 25696
rect 15657 25687 15715 25693
rect 15657 25684 15669 25687
rect 15528 25656 15669 25684
rect 15528 25644 15534 25656
rect 15657 25653 15669 25656
rect 15703 25653 15715 25687
rect 15657 25647 15715 25653
rect 19518 25644 19524 25696
rect 19576 25684 19582 25696
rect 19705 25687 19763 25693
rect 19705 25684 19717 25687
rect 19576 25656 19717 25684
rect 19576 25644 19582 25656
rect 19705 25653 19717 25656
rect 19751 25653 19763 25687
rect 19705 25647 19763 25653
rect 21821 25687 21879 25693
rect 21821 25653 21833 25687
rect 21867 25684 21879 25687
rect 22922 25684 22928 25696
rect 21867 25656 22928 25684
rect 21867 25653 21879 25656
rect 21821 25647 21879 25653
rect 22922 25644 22928 25656
rect 22980 25644 22986 25696
rect 25774 25644 25780 25696
rect 25832 25644 25838 25696
rect 1104 25594 28704 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 28704 25594
rect 1104 25520 28704 25542
rect 8570 25440 8576 25492
rect 8628 25440 8634 25492
rect 8938 25440 8944 25492
rect 8996 25440 9002 25492
rect 10413 25483 10471 25489
rect 10413 25480 10425 25483
rect 10152 25452 10425 25480
rect 9769 25415 9827 25421
rect 9769 25412 9781 25415
rect 8496 25384 9781 25412
rect 5169 25347 5227 25353
rect 5169 25313 5181 25347
rect 5215 25344 5227 25347
rect 5442 25344 5448 25356
rect 5215 25316 5448 25344
rect 5215 25313 5227 25316
rect 5169 25307 5227 25313
rect 5442 25304 5448 25316
rect 5500 25304 5506 25356
rect 8386 25304 8392 25356
rect 8444 25304 8450 25356
rect 8496 25353 8524 25384
rect 9769 25381 9781 25384
rect 9815 25412 9827 25415
rect 9950 25412 9956 25424
rect 9815 25384 9956 25412
rect 9815 25381 9827 25384
rect 9769 25375 9827 25381
rect 9950 25372 9956 25384
rect 10008 25372 10014 25424
rect 10152 25353 10180 25452
rect 10413 25449 10425 25452
rect 10459 25449 10471 25483
rect 10413 25443 10471 25449
rect 11974 25440 11980 25492
rect 12032 25480 12038 25492
rect 12437 25483 12495 25489
rect 12437 25480 12449 25483
rect 12032 25452 12449 25480
rect 12032 25440 12038 25452
rect 12437 25449 12449 25452
rect 12483 25449 12495 25483
rect 12437 25443 12495 25449
rect 20993 25483 21051 25489
rect 20993 25449 21005 25483
rect 21039 25480 21051 25483
rect 21174 25480 21180 25492
rect 21039 25452 21180 25480
rect 21039 25449 21051 25452
rect 20993 25443 21051 25449
rect 21174 25440 21180 25452
rect 21232 25480 21238 25492
rect 21542 25480 21548 25492
rect 21232 25452 21548 25480
rect 21232 25440 21238 25452
rect 21542 25440 21548 25452
rect 21600 25440 21606 25492
rect 24121 25483 24179 25489
rect 24121 25449 24133 25483
rect 24167 25480 24179 25483
rect 24302 25480 24308 25492
rect 24167 25452 24308 25480
rect 24167 25449 24179 25452
rect 24121 25443 24179 25449
rect 24302 25440 24308 25452
rect 24360 25440 24366 25492
rect 12897 25415 12955 25421
rect 12897 25381 12909 25415
rect 12943 25412 12955 25415
rect 12986 25412 12992 25424
rect 12943 25384 12992 25412
rect 12943 25381 12955 25384
rect 12897 25375 12955 25381
rect 12986 25372 12992 25384
rect 13044 25372 13050 25424
rect 8481 25347 8539 25353
rect 8481 25313 8493 25347
rect 8527 25313 8539 25347
rect 10137 25347 10195 25353
rect 10137 25344 10149 25347
rect 8481 25307 8539 25313
rect 8680 25316 10149 25344
rect 4706 25236 4712 25288
rect 4764 25276 4770 25288
rect 4893 25279 4951 25285
rect 4893 25276 4905 25279
rect 4764 25248 4905 25276
rect 4764 25236 4770 25248
rect 4893 25245 4905 25248
rect 4939 25245 4951 25279
rect 4893 25239 4951 25245
rect 7834 25236 7840 25288
rect 7892 25276 7898 25288
rect 8680 25285 8708 25316
rect 10137 25313 10149 25316
rect 10183 25313 10195 25347
rect 10137 25307 10195 25313
rect 15470 25304 15476 25356
rect 15528 25304 15534 25356
rect 19518 25304 19524 25356
rect 19576 25304 19582 25356
rect 23477 25347 23535 25353
rect 22112 25316 23336 25344
rect 22112 25288 22140 25316
rect 8665 25279 8723 25285
rect 8665 25276 8677 25279
rect 7892 25248 8677 25276
rect 7892 25236 7898 25248
rect 8665 25245 8677 25248
rect 8711 25245 8723 25279
rect 8665 25239 8723 25245
rect 8754 25236 8760 25288
rect 8812 25276 8818 25288
rect 9493 25279 9551 25285
rect 9493 25276 9505 25279
rect 8812 25248 9505 25276
rect 8812 25236 8818 25248
rect 9493 25245 9505 25248
rect 9539 25276 9551 25279
rect 9582 25276 9588 25288
rect 9539 25248 9588 25276
rect 9539 25245 9551 25248
rect 9493 25239 9551 25245
rect 9582 25236 9588 25248
rect 9640 25276 9646 25288
rect 9640 25248 10272 25276
rect 9640 25236 9646 25248
rect 5445 25211 5503 25217
rect 5445 25177 5457 25211
rect 5491 25208 5503 25211
rect 5534 25208 5540 25220
rect 5491 25180 5540 25208
rect 5491 25177 5503 25180
rect 5445 25171 5503 25177
rect 5534 25168 5540 25180
rect 5592 25168 5598 25220
rect 5902 25168 5908 25220
rect 5960 25168 5966 25220
rect 10244 25217 10272 25248
rect 10686 25236 10692 25288
rect 10744 25236 10750 25288
rect 12713 25279 12771 25285
rect 12713 25245 12725 25279
rect 12759 25245 12771 25279
rect 12713 25239 12771 25245
rect 12989 25279 13047 25285
rect 12989 25245 13001 25279
rect 13035 25276 13047 25279
rect 13265 25279 13323 25285
rect 13265 25276 13277 25279
rect 13035 25248 13277 25276
rect 13035 25245 13047 25248
rect 12989 25239 13047 25245
rect 13265 25245 13277 25248
rect 13311 25245 13323 25279
rect 13265 25239 13323 25245
rect 10229 25211 10287 25217
rect 10229 25177 10241 25211
rect 10275 25177 10287 25211
rect 10229 25171 10287 25177
rect 10336 25180 10640 25208
rect 6914 25100 6920 25152
rect 6972 25100 6978 25152
rect 7190 25100 7196 25152
rect 7248 25140 7254 25152
rect 7745 25143 7803 25149
rect 7745 25140 7757 25143
rect 7248 25112 7757 25140
rect 7248 25100 7254 25112
rect 7745 25109 7757 25112
rect 7791 25109 7803 25143
rect 7745 25103 7803 25109
rect 9674 25100 9680 25152
rect 9732 25100 9738 25152
rect 9858 25100 9864 25152
rect 9916 25140 9922 25152
rect 10336 25140 10364 25180
rect 9916 25112 10364 25140
rect 9916 25100 9922 25112
rect 10410 25100 10416 25152
rect 10468 25149 10474 25152
rect 10612 25149 10640 25180
rect 10962 25168 10968 25220
rect 11020 25168 11026 25220
rect 12618 25208 12624 25220
rect 12190 25180 12624 25208
rect 12618 25168 12624 25180
rect 12676 25168 12682 25220
rect 12728 25208 12756 25239
rect 13814 25236 13820 25288
rect 13872 25236 13878 25288
rect 14366 25236 14372 25288
rect 14424 25276 14430 25288
rect 14461 25279 14519 25285
rect 14461 25276 14473 25279
rect 14424 25248 14473 25276
rect 14424 25236 14430 25248
rect 14461 25245 14473 25248
rect 14507 25245 14519 25279
rect 14461 25239 14519 25245
rect 15194 25236 15200 25288
rect 15252 25236 15258 25288
rect 17586 25236 17592 25288
rect 17644 25276 17650 25288
rect 19242 25276 19248 25288
rect 17644 25248 19248 25276
rect 17644 25236 17650 25248
rect 19242 25236 19248 25248
rect 19300 25236 19306 25288
rect 21266 25236 21272 25288
rect 21324 25236 21330 25288
rect 21453 25279 21511 25285
rect 21453 25245 21465 25279
rect 21499 25276 21511 25279
rect 22094 25276 22100 25288
rect 21499 25248 22100 25276
rect 21499 25245 21511 25248
rect 21453 25239 21511 25245
rect 22094 25236 22100 25248
rect 22152 25236 22158 25288
rect 22281 25279 22339 25285
rect 22281 25245 22293 25279
rect 22327 25276 22339 25279
rect 22373 25279 22431 25285
rect 22373 25276 22385 25279
rect 22327 25248 22385 25276
rect 22327 25245 22339 25248
rect 22281 25239 22339 25245
rect 22373 25245 22385 25248
rect 22419 25245 22431 25279
rect 22373 25239 22431 25245
rect 22922 25236 22928 25288
rect 22980 25276 22986 25288
rect 23308 25285 23336 25316
rect 23477 25313 23489 25347
rect 23523 25344 23535 25347
rect 23750 25344 23756 25356
rect 23523 25316 23756 25344
rect 23523 25313 23535 25316
rect 23477 25307 23535 25313
rect 23750 25304 23756 25316
rect 23808 25304 23814 25356
rect 24854 25344 24860 25356
rect 23860 25316 24860 25344
rect 23860 25285 23888 25316
rect 24854 25304 24860 25316
rect 24912 25304 24918 25356
rect 23109 25279 23167 25285
rect 23109 25276 23121 25279
rect 22980 25248 23121 25276
rect 22980 25236 22986 25248
rect 23109 25245 23121 25248
rect 23155 25245 23167 25279
rect 23109 25239 23167 25245
rect 23293 25279 23351 25285
rect 23293 25245 23305 25279
rect 23339 25245 23351 25279
rect 23293 25239 23351 25245
rect 23845 25279 23903 25285
rect 23845 25245 23857 25279
rect 23891 25245 23903 25279
rect 23845 25239 23903 25245
rect 26142 25236 26148 25288
rect 26200 25236 26206 25288
rect 26326 25236 26332 25288
rect 26384 25236 26390 25288
rect 26881 25279 26939 25285
rect 26881 25245 26893 25279
rect 26927 25276 26939 25279
rect 26973 25279 27031 25285
rect 26973 25276 26985 25279
rect 26927 25248 26985 25276
rect 26927 25245 26939 25248
rect 26881 25239 26939 25245
rect 26973 25245 26985 25248
rect 27019 25245 27031 25279
rect 26973 25239 27031 25245
rect 27154 25236 27160 25288
rect 27212 25236 27218 25288
rect 13630 25208 13636 25220
rect 12728 25180 13636 25208
rect 13630 25168 13636 25180
rect 13688 25168 13694 25220
rect 16022 25168 16028 25220
rect 16080 25168 16086 25220
rect 20530 25168 20536 25220
rect 20588 25168 20594 25220
rect 25869 25211 25927 25217
rect 25438 25180 25544 25208
rect 10468 25143 10487 25149
rect 10475 25109 10487 25143
rect 10468 25103 10487 25109
rect 10597 25143 10655 25149
rect 10597 25109 10609 25143
rect 10643 25109 10655 25143
rect 10597 25103 10655 25109
rect 10468 25100 10474 25103
rect 12526 25100 12532 25152
rect 12584 25100 12590 25152
rect 14550 25100 14556 25152
rect 14608 25140 14614 25152
rect 15105 25143 15163 25149
rect 15105 25140 15117 25143
rect 14608 25112 15117 25140
rect 14608 25100 14614 25112
rect 15105 25109 15117 25112
rect 15151 25109 15163 25143
rect 15105 25103 15163 25109
rect 16942 25100 16948 25152
rect 17000 25100 17006 25152
rect 21358 25100 21364 25152
rect 21416 25100 21422 25152
rect 22189 25143 22247 25149
rect 22189 25109 22201 25143
rect 22235 25140 22247 25143
rect 23014 25140 23020 25152
rect 22235 25112 23020 25140
rect 22235 25109 22247 25112
rect 22189 25103 22247 25109
rect 23014 25100 23020 25112
rect 23072 25100 23078 25152
rect 24397 25143 24455 25149
rect 24397 25109 24409 25143
rect 24443 25140 24455 25143
rect 25130 25140 25136 25152
rect 24443 25112 25136 25140
rect 24443 25109 24455 25112
rect 24397 25103 24455 25109
rect 25130 25100 25136 25112
rect 25188 25100 25194 25152
rect 25516 25140 25544 25180
rect 25869 25177 25881 25211
rect 25915 25208 25927 25211
rect 27065 25211 27123 25217
rect 27065 25208 27077 25211
rect 25915 25180 27077 25208
rect 25915 25177 25927 25180
rect 25869 25171 25927 25177
rect 27065 25177 27077 25180
rect 27111 25177 27123 25211
rect 27065 25171 27123 25177
rect 27798 25140 27804 25152
rect 25516 25112 27804 25140
rect 27798 25100 27804 25112
rect 27856 25100 27862 25152
rect 1104 25050 28704 25072
rect 1104 24998 4874 25050
rect 4926 24998 4938 25050
rect 4990 24998 5002 25050
rect 5054 24998 5066 25050
rect 5118 24998 5130 25050
rect 5182 24998 28704 25050
rect 1104 24976 28704 24998
rect 7834 24896 7840 24948
rect 7892 24896 7898 24948
rect 10229 24939 10287 24945
rect 10229 24905 10241 24939
rect 10275 24936 10287 24939
rect 10962 24936 10968 24948
rect 10275 24908 10968 24936
rect 10275 24905 10287 24908
rect 10229 24899 10287 24905
rect 10962 24896 10968 24908
rect 11020 24896 11026 24948
rect 15378 24936 15384 24948
rect 14476 24908 15384 24936
rect 4706 24828 4712 24880
rect 4764 24828 4770 24880
rect 6914 24828 6920 24880
rect 6972 24868 6978 24880
rect 7285 24871 7343 24877
rect 7285 24868 7297 24871
rect 6972 24840 7297 24868
rect 6972 24828 6978 24840
rect 7285 24837 7297 24840
rect 7331 24837 7343 24871
rect 7285 24831 7343 24837
rect 10318 24828 10324 24880
rect 10376 24828 10382 24880
rect 13354 24868 13360 24880
rect 13294 24840 13360 24868
rect 13354 24828 13360 24840
rect 13412 24828 13418 24880
rect 7101 24803 7159 24809
rect 4433 24735 4491 24741
rect 4433 24701 4445 24735
rect 4479 24732 4491 24735
rect 4479 24704 4568 24732
rect 4479 24701 4491 24704
rect 4433 24695 4491 24701
rect 4540 24596 4568 24704
rect 4798 24692 4804 24744
rect 4856 24732 4862 24744
rect 5828 24732 5856 24786
rect 7101 24769 7113 24803
rect 7147 24769 7159 24803
rect 7101 24763 7159 24769
rect 5902 24732 5908 24744
rect 4856 24704 5908 24732
rect 4856 24692 4862 24704
rect 5902 24692 5908 24704
rect 5960 24692 5966 24744
rect 6181 24735 6239 24741
rect 6181 24701 6193 24735
rect 6227 24732 6239 24735
rect 7116 24732 7144 24763
rect 6227 24704 7144 24732
rect 6227 24701 6239 24704
rect 6181 24695 6239 24701
rect 5920 24664 5948 24692
rect 8220 24664 8248 24786
rect 10042 24760 10048 24812
rect 10100 24760 10106 24812
rect 10410 24760 10416 24812
rect 10468 24800 10474 24812
rect 10873 24803 10931 24809
rect 10873 24800 10885 24803
rect 10468 24772 10885 24800
rect 10468 24760 10474 24772
rect 10873 24769 10885 24772
rect 10919 24769 10931 24803
rect 10873 24763 10931 24769
rect 11514 24760 11520 24812
rect 11572 24760 11578 24812
rect 11701 24803 11759 24809
rect 11701 24769 11713 24803
rect 11747 24769 11759 24803
rect 11701 24763 11759 24769
rect 9309 24735 9367 24741
rect 9309 24701 9321 24735
rect 9355 24732 9367 24735
rect 9355 24704 9536 24732
rect 9355 24701 9367 24704
rect 9309 24695 9367 24701
rect 5920 24636 8248 24664
rect 9508 24664 9536 24704
rect 9582 24692 9588 24744
rect 9640 24692 9646 24744
rect 9769 24735 9827 24741
rect 9769 24701 9781 24735
rect 9815 24732 9827 24735
rect 11054 24732 11060 24744
rect 9815 24704 11060 24732
rect 9815 24701 9827 24704
rect 9769 24695 9827 24701
rect 11054 24692 11060 24704
rect 11112 24692 11118 24744
rect 9674 24664 9680 24676
rect 9508 24636 9680 24664
rect 9674 24624 9680 24636
rect 9732 24624 9738 24676
rect 9950 24624 9956 24676
rect 10008 24664 10014 24676
rect 10008 24636 10640 24664
rect 10008 24624 10014 24636
rect 5442 24596 5448 24608
rect 4540 24568 5448 24596
rect 5442 24556 5448 24568
rect 5500 24556 5506 24608
rect 7377 24599 7435 24605
rect 7377 24565 7389 24599
rect 7423 24596 7435 24599
rect 9122 24596 9128 24608
rect 7423 24568 9128 24596
rect 7423 24565 7435 24568
rect 7377 24559 7435 24565
rect 9122 24556 9128 24568
rect 9180 24556 9186 24608
rect 9858 24556 9864 24608
rect 9916 24556 9922 24608
rect 10612 24596 10640 24636
rect 10962 24596 10968 24608
rect 10612 24568 10968 24596
rect 10962 24556 10968 24568
rect 11020 24596 11026 24608
rect 11517 24599 11575 24605
rect 11517 24596 11529 24599
rect 11020 24568 11529 24596
rect 11020 24556 11026 24568
rect 11517 24565 11529 24568
rect 11563 24565 11575 24599
rect 11716 24596 11744 24763
rect 13446 24760 13452 24812
rect 13504 24800 13510 24812
rect 13633 24803 13691 24809
rect 13633 24800 13645 24803
rect 13504 24772 13645 24800
rect 13504 24760 13510 24772
rect 13633 24769 13645 24772
rect 13679 24769 13691 24803
rect 13633 24763 13691 24769
rect 13814 24760 13820 24812
rect 13872 24760 13878 24812
rect 13909 24803 13967 24809
rect 13909 24769 13921 24803
rect 13955 24769 13967 24803
rect 13909 24763 13967 24769
rect 11790 24692 11796 24744
rect 11848 24692 11854 24744
rect 12069 24735 12127 24741
rect 12069 24701 12081 24735
rect 12115 24732 12127 24735
rect 12526 24732 12532 24744
rect 12115 24704 12532 24732
rect 12115 24701 12127 24704
rect 12069 24695 12127 24701
rect 12526 24692 12532 24704
rect 12584 24692 12590 24744
rect 13078 24692 13084 24744
rect 13136 24732 13142 24744
rect 13924 24732 13952 24763
rect 14090 24760 14096 24812
rect 14148 24760 14154 24812
rect 14182 24760 14188 24812
rect 14240 24760 14246 24812
rect 14369 24803 14427 24809
rect 14369 24769 14381 24803
rect 14415 24800 14427 24803
rect 14476 24800 14504 24908
rect 15378 24896 15384 24908
rect 15436 24896 15442 24948
rect 17862 24936 17868 24948
rect 17696 24908 17868 24936
rect 16022 24868 16028 24880
rect 15962 24840 16028 24868
rect 16022 24828 16028 24840
rect 16080 24868 16086 24880
rect 17696 24868 17724 24908
rect 17862 24896 17868 24908
rect 17920 24896 17926 24948
rect 22094 24896 22100 24948
rect 22152 24936 22158 24948
rect 22925 24939 22983 24945
rect 22925 24936 22937 24939
rect 22152 24908 22937 24936
rect 22152 24896 22158 24908
rect 22925 24905 22937 24908
rect 22971 24905 22983 24939
rect 22925 24899 22983 24905
rect 23109 24939 23167 24945
rect 23109 24905 23121 24939
rect 23155 24936 23167 24939
rect 23290 24936 23296 24948
rect 23155 24908 23296 24936
rect 23155 24905 23167 24908
rect 23109 24899 23167 24905
rect 23290 24896 23296 24908
rect 23348 24896 23354 24948
rect 23750 24896 23756 24948
rect 23808 24936 23814 24948
rect 26237 24939 26295 24945
rect 23808 24908 26004 24936
rect 23808 24896 23814 24908
rect 16080 24840 17724 24868
rect 16080 24828 16086 24840
rect 17770 24828 17776 24880
rect 17828 24828 17834 24880
rect 22557 24871 22615 24877
rect 22557 24837 22569 24871
rect 22603 24837 22615 24871
rect 22757 24871 22815 24877
rect 22757 24868 22769 24871
rect 22557 24831 22615 24837
rect 22756 24837 22769 24868
rect 22803 24837 22815 24871
rect 22756 24831 22815 24837
rect 14415 24772 14504 24800
rect 14415 24769 14427 24772
rect 14369 24763 14427 24769
rect 16206 24760 16212 24812
rect 16264 24800 16270 24812
rect 16301 24803 16359 24809
rect 16301 24800 16313 24803
rect 16264 24772 16313 24800
rect 16264 24760 16270 24772
rect 16301 24769 16313 24772
rect 16347 24769 16359 24803
rect 16301 24763 16359 24769
rect 16485 24803 16543 24809
rect 16485 24769 16497 24803
rect 16531 24800 16543 24803
rect 16758 24800 16764 24812
rect 16531 24772 16764 24800
rect 16531 24769 16543 24772
rect 16485 24763 16543 24769
rect 16758 24760 16764 24772
rect 16816 24760 16822 24812
rect 17034 24760 17040 24812
rect 17092 24800 17098 24812
rect 17681 24803 17739 24809
rect 17681 24800 17693 24803
rect 17092 24772 17693 24800
rect 17092 24760 17098 24772
rect 17681 24769 17693 24772
rect 17727 24800 17739 24803
rect 17957 24803 18015 24809
rect 17957 24800 17969 24803
rect 17727 24772 17969 24800
rect 17727 24769 17739 24772
rect 17681 24763 17739 24769
rect 17957 24769 17969 24772
rect 18003 24769 18015 24803
rect 17957 24763 18015 24769
rect 18049 24803 18107 24809
rect 18049 24769 18061 24803
rect 18095 24769 18107 24803
rect 18049 24763 18107 24769
rect 13136 24704 13952 24732
rect 14461 24735 14519 24741
rect 13136 24692 13142 24704
rect 14461 24701 14473 24735
rect 14507 24701 14519 24735
rect 14461 24695 14519 24701
rect 14737 24735 14795 24741
rect 14737 24701 14749 24735
rect 14783 24732 14795 24735
rect 16393 24735 16451 24741
rect 16393 24732 16405 24735
rect 14783 24704 16405 24732
rect 14783 24701 14795 24704
rect 14737 24695 14795 24701
rect 16393 24701 16405 24704
rect 16439 24701 16451 24735
rect 16393 24695 16451 24701
rect 16669 24735 16727 24741
rect 16669 24701 16681 24735
rect 16715 24701 16727 24735
rect 16669 24695 16727 24701
rect 13630 24624 13636 24676
rect 13688 24624 13694 24676
rect 14366 24624 14372 24676
rect 14424 24624 14430 24676
rect 12802 24596 12808 24608
rect 11716 24568 12808 24596
rect 11517 24559 11575 24565
rect 12802 24556 12808 24568
rect 12860 24556 12866 24608
rect 13541 24599 13599 24605
rect 13541 24565 13553 24599
rect 13587 24596 13599 24599
rect 13814 24596 13820 24608
rect 13587 24568 13820 24596
rect 13587 24565 13599 24568
rect 13541 24559 13599 24565
rect 13814 24556 13820 24568
rect 13872 24556 13878 24608
rect 14476 24596 14504 24695
rect 16209 24667 16267 24673
rect 16209 24633 16221 24667
rect 16255 24664 16267 24667
rect 16298 24664 16304 24676
rect 16255 24636 16304 24664
rect 16255 24633 16267 24636
rect 16209 24627 16267 24633
rect 16298 24624 16304 24636
rect 16356 24664 16362 24676
rect 16684 24664 16712 24695
rect 17126 24692 17132 24744
rect 17184 24732 17190 24744
rect 17405 24735 17463 24741
rect 17405 24732 17417 24735
rect 17184 24704 17417 24732
rect 17184 24692 17190 24704
rect 17405 24701 17417 24704
rect 17451 24701 17463 24735
rect 18064 24732 18092 24763
rect 19242 24760 19248 24812
rect 19300 24800 19306 24812
rect 19889 24803 19947 24809
rect 19889 24800 19901 24803
rect 19300 24772 19901 24800
rect 19300 24760 19306 24772
rect 19889 24769 19901 24772
rect 19935 24769 19947 24803
rect 22462 24800 22468 24812
rect 21298 24772 22468 24800
rect 19889 24763 19947 24769
rect 22462 24760 22468 24772
rect 22520 24760 22526 24812
rect 17405 24695 17463 24701
rect 17604 24704 18092 24732
rect 17497 24667 17555 24673
rect 17497 24664 17509 24667
rect 16356 24636 16712 24664
rect 16776 24636 17509 24664
rect 16356 24624 16362 24636
rect 15194 24596 15200 24608
rect 14476 24568 15200 24596
rect 15194 24556 15200 24568
rect 15252 24556 15258 24608
rect 15378 24556 15384 24608
rect 15436 24596 15442 24608
rect 16776 24596 16804 24636
rect 17497 24633 17509 24636
rect 17543 24633 17555 24667
rect 17497 24627 17555 24633
rect 15436 24568 16804 24596
rect 15436 24556 15442 24568
rect 16850 24556 16856 24608
rect 16908 24596 16914 24608
rect 17313 24599 17371 24605
rect 17313 24596 17325 24599
rect 16908 24568 17325 24596
rect 16908 24556 16914 24568
rect 17313 24565 17325 24568
rect 17359 24565 17371 24599
rect 17313 24559 17371 24565
rect 17402 24556 17408 24608
rect 17460 24596 17466 24608
rect 17604 24605 17632 24704
rect 19150 24692 19156 24744
rect 19208 24692 19214 24744
rect 20165 24735 20223 24741
rect 20165 24701 20177 24735
rect 20211 24732 20223 24735
rect 21358 24732 21364 24744
rect 20211 24704 21364 24732
rect 20211 24701 20223 24704
rect 20165 24695 20223 24701
rect 21358 24692 21364 24704
rect 21416 24692 21422 24744
rect 21637 24735 21695 24741
rect 21637 24701 21649 24735
rect 21683 24732 21695 24735
rect 22278 24732 22284 24744
rect 21683 24704 22284 24732
rect 21683 24701 21695 24704
rect 21637 24695 21695 24701
rect 22278 24692 22284 24704
rect 22336 24732 22342 24744
rect 22373 24735 22431 24741
rect 22373 24732 22385 24735
rect 22336 24704 22385 24732
rect 22336 24692 22342 24704
rect 22373 24701 22385 24704
rect 22419 24732 22431 24735
rect 22572 24732 22600 24831
rect 22419 24704 22600 24732
rect 22419 24701 22431 24704
rect 22373 24695 22431 24701
rect 17678 24624 17684 24676
rect 17736 24664 17742 24676
rect 17773 24667 17831 24673
rect 17773 24664 17785 24667
rect 17736 24636 17785 24664
rect 17736 24624 17742 24636
rect 17773 24633 17785 24636
rect 17819 24633 17831 24667
rect 17773 24627 17831 24633
rect 21542 24624 21548 24676
rect 21600 24664 21606 24676
rect 21600 24636 21956 24664
rect 21600 24624 21606 24636
rect 17589 24599 17647 24605
rect 17589 24596 17601 24599
rect 17460 24568 17601 24596
rect 17460 24556 17466 24568
rect 17589 24565 17601 24568
rect 17635 24565 17647 24599
rect 17589 24559 17647 24565
rect 17862 24556 17868 24608
rect 17920 24596 17926 24608
rect 18601 24599 18659 24605
rect 18601 24596 18613 24599
rect 17920 24568 18613 24596
rect 17920 24556 17926 24568
rect 18601 24565 18613 24568
rect 18647 24565 18659 24599
rect 18601 24559 18659 24565
rect 21726 24556 21732 24608
rect 21784 24596 21790 24608
rect 21821 24599 21879 24605
rect 21821 24596 21833 24599
rect 21784 24568 21833 24596
rect 21784 24556 21790 24568
rect 21821 24565 21833 24568
rect 21867 24565 21879 24599
rect 21928 24596 21956 24636
rect 22002 24624 22008 24676
rect 22060 24664 22066 24676
rect 22756 24664 22784 24831
rect 23014 24760 23020 24812
rect 23072 24760 23078 24812
rect 23201 24803 23259 24809
rect 23201 24769 23213 24803
rect 23247 24800 23259 24803
rect 23768 24800 23796 24896
rect 25682 24868 25688 24880
rect 25148 24840 25688 24868
rect 25148 24812 25176 24840
rect 25682 24828 25688 24840
rect 25740 24868 25746 24880
rect 25869 24871 25927 24877
rect 25869 24868 25881 24871
rect 25740 24840 25881 24868
rect 25740 24828 25746 24840
rect 25869 24837 25881 24840
rect 25915 24837 25927 24871
rect 25976 24868 26004 24908
rect 26237 24905 26249 24939
rect 26283 24936 26295 24939
rect 26418 24936 26424 24948
rect 26283 24908 26424 24936
rect 26283 24905 26295 24908
rect 26237 24899 26295 24905
rect 26418 24896 26424 24908
rect 26476 24936 26482 24948
rect 27154 24936 27160 24948
rect 26476 24908 27160 24936
rect 26476 24896 26482 24908
rect 27154 24896 27160 24908
rect 27212 24896 27218 24948
rect 26085 24871 26143 24877
rect 26085 24868 26097 24871
rect 25976 24840 26097 24868
rect 25869 24831 25927 24837
rect 26085 24837 26097 24840
rect 26131 24868 26143 24871
rect 26131 24840 26648 24868
rect 26131 24837 26143 24840
rect 26085 24831 26143 24837
rect 23247 24772 23796 24800
rect 23247 24769 23259 24772
rect 23201 24763 23259 24769
rect 24854 24760 24860 24812
rect 24912 24800 24918 24812
rect 24949 24803 25007 24809
rect 24949 24800 24961 24803
rect 24912 24772 24961 24800
rect 24912 24760 24918 24772
rect 24949 24769 24961 24772
rect 24995 24769 25007 24803
rect 24949 24763 25007 24769
rect 25041 24803 25099 24809
rect 25041 24769 25053 24803
rect 25087 24769 25099 24803
rect 25041 24763 25099 24769
rect 25056 24732 25084 24763
rect 25130 24760 25136 24812
rect 25188 24760 25194 24812
rect 26620 24809 26648 24840
rect 25777 24803 25835 24809
rect 25777 24769 25789 24803
rect 25823 24800 25835 24803
rect 26329 24803 26387 24809
rect 26329 24800 26341 24803
rect 25823 24772 26341 24800
rect 25823 24769 25835 24772
rect 25777 24763 25835 24769
rect 26329 24769 26341 24772
rect 26375 24769 26387 24803
rect 26329 24763 26387 24769
rect 26513 24803 26571 24809
rect 26513 24769 26525 24803
rect 26559 24769 26571 24803
rect 26513 24763 26571 24769
rect 26605 24803 26663 24809
rect 26605 24769 26617 24803
rect 26651 24769 26663 24803
rect 26605 24763 26663 24769
rect 26528 24732 26556 24763
rect 26970 24760 26976 24812
rect 27028 24760 27034 24812
rect 27154 24760 27160 24812
rect 27212 24760 27218 24812
rect 27801 24803 27859 24809
rect 27801 24769 27813 24803
rect 27847 24800 27859 24803
rect 27890 24800 27896 24812
rect 27847 24772 27896 24800
rect 27847 24769 27859 24772
rect 27801 24763 27859 24769
rect 27890 24760 27896 24772
rect 27948 24760 27954 24812
rect 25056 24704 25820 24732
rect 22060 24636 22784 24664
rect 22060 24624 22066 24636
rect 25792 24608 25820 24704
rect 26206 24704 26556 24732
rect 22741 24599 22799 24605
rect 22741 24596 22753 24599
rect 21928 24568 22753 24596
rect 21821 24559 21879 24565
rect 22741 24565 22753 24568
rect 22787 24565 22799 24599
rect 22741 24559 22799 24565
rect 25774 24556 25780 24608
rect 25832 24596 25838 24608
rect 26053 24599 26111 24605
rect 26053 24596 26065 24599
rect 25832 24568 26065 24596
rect 25832 24556 25838 24568
rect 26053 24565 26065 24568
rect 26099 24596 26111 24599
rect 26206 24596 26234 24704
rect 26326 24624 26332 24676
rect 26384 24624 26390 24676
rect 26099 24568 26234 24596
rect 26099 24565 26111 24568
rect 26053 24559 26111 24565
rect 26786 24556 26792 24608
rect 26844 24596 26850 24608
rect 26973 24599 27031 24605
rect 26973 24596 26985 24599
rect 26844 24568 26985 24596
rect 26844 24556 26850 24568
rect 26973 24565 26985 24568
rect 27019 24565 27031 24599
rect 26973 24559 27031 24565
rect 27709 24599 27767 24605
rect 27709 24565 27721 24599
rect 27755 24596 27767 24599
rect 27982 24596 27988 24608
rect 27755 24568 27988 24596
rect 27755 24565 27767 24568
rect 27709 24559 27767 24565
rect 27982 24556 27988 24568
rect 28040 24556 28046 24608
rect 1104 24506 28704 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 28704 24506
rect 1104 24432 28704 24454
rect 8665 24395 8723 24401
rect 8665 24361 8677 24395
rect 8711 24392 8723 24395
rect 8754 24392 8760 24404
rect 8711 24364 8760 24392
rect 8711 24361 8723 24364
rect 8665 24355 8723 24361
rect 8754 24352 8760 24364
rect 8812 24352 8818 24404
rect 10410 24352 10416 24404
rect 10468 24392 10474 24404
rect 10689 24395 10747 24401
rect 10689 24392 10701 24395
rect 10468 24364 10701 24392
rect 10468 24352 10474 24364
rect 10689 24361 10701 24364
rect 10735 24361 10747 24395
rect 10689 24355 10747 24361
rect 11054 24352 11060 24404
rect 11112 24392 11118 24404
rect 12989 24395 13047 24401
rect 12989 24392 13001 24395
rect 11112 24364 13001 24392
rect 11112 24352 11118 24364
rect 12989 24361 13001 24364
rect 13035 24392 13047 24395
rect 13814 24392 13820 24404
rect 13035 24364 13820 24392
rect 13035 24361 13047 24364
rect 12989 24355 13047 24361
rect 13814 24352 13820 24364
rect 13872 24352 13878 24404
rect 14090 24352 14096 24404
rect 14148 24392 14154 24404
rect 15286 24392 15292 24404
rect 14148 24364 15292 24392
rect 14148 24352 14154 24364
rect 15286 24352 15292 24364
rect 15344 24392 15350 24404
rect 16206 24392 16212 24404
rect 15344 24364 16212 24392
rect 15344 24352 15350 24364
rect 16206 24352 16212 24364
rect 16264 24352 16270 24404
rect 16301 24395 16359 24401
rect 16301 24361 16313 24395
rect 16347 24392 16359 24395
rect 16942 24392 16948 24404
rect 16347 24364 16948 24392
rect 16347 24361 16359 24364
rect 16301 24355 16359 24361
rect 16942 24352 16948 24364
rect 17000 24352 17006 24404
rect 17402 24392 17408 24404
rect 17236 24364 17408 24392
rect 12802 24284 12808 24336
rect 12860 24284 12866 24336
rect 15838 24284 15844 24336
rect 15896 24324 15902 24336
rect 16117 24327 16175 24333
rect 16117 24324 16129 24327
rect 15896 24296 16129 24324
rect 15896 24284 15902 24296
rect 16117 24293 16129 24296
rect 16163 24293 16175 24327
rect 16117 24287 16175 24293
rect 16669 24327 16727 24333
rect 16669 24293 16681 24327
rect 16715 24324 16727 24327
rect 17034 24324 17040 24336
rect 16715 24296 17040 24324
rect 16715 24293 16727 24296
rect 16669 24287 16727 24293
rect 5442 24216 5448 24268
rect 5500 24256 5506 24268
rect 6914 24256 6920 24268
rect 5500 24228 6920 24256
rect 5500 24216 5506 24228
rect 6914 24216 6920 24228
rect 6972 24256 6978 24268
rect 8941 24259 8999 24265
rect 8941 24256 8953 24259
rect 6972 24228 8953 24256
rect 6972 24216 6978 24228
rect 8941 24225 8953 24228
rect 8987 24256 8999 24259
rect 9582 24256 9588 24268
rect 8987 24228 9588 24256
rect 8987 24225 8999 24228
rect 8941 24219 8999 24225
rect 9582 24216 9588 24228
rect 9640 24216 9646 24268
rect 10686 24216 10692 24268
rect 10744 24256 10750 24268
rect 10965 24259 11023 24265
rect 10965 24256 10977 24259
rect 10744 24228 10977 24256
rect 10744 24216 10750 24228
rect 10965 24225 10977 24228
rect 11011 24256 11023 24259
rect 11790 24256 11796 24268
rect 11011 24228 11796 24256
rect 11011 24225 11023 24228
rect 10965 24219 11023 24225
rect 11790 24216 11796 24228
rect 11848 24256 11854 24268
rect 13078 24256 13084 24268
rect 11848 24228 13084 24256
rect 11848 24216 11854 24228
rect 13078 24216 13084 24228
rect 13136 24216 13142 24268
rect 13262 24216 13268 24268
rect 13320 24256 13326 24268
rect 14277 24259 14335 24265
rect 14277 24256 14289 24259
rect 13320 24228 14289 24256
rect 13320 24216 13326 24228
rect 14277 24225 14289 24228
rect 14323 24256 14335 24259
rect 15194 24256 15200 24268
rect 14323 24228 15200 24256
rect 14323 24225 14335 24228
rect 14277 24219 14335 24225
rect 15194 24216 15200 24228
rect 15252 24216 15258 24268
rect 16022 24216 16028 24268
rect 16080 24256 16086 24268
rect 16684 24256 16712 24287
rect 17034 24284 17040 24296
rect 17092 24284 17098 24336
rect 16080 24228 16712 24256
rect 16080 24216 16086 24228
rect 12912 24160 13216 24188
rect 7190 24080 7196 24132
rect 7248 24080 7254 24132
rect 7300 24092 7682 24120
rect 5902 24012 5908 24064
rect 5960 24052 5966 24064
rect 7300 24052 7328 24092
rect 9214 24080 9220 24132
rect 9272 24080 9278 24132
rect 10442 24092 11192 24120
rect 5960 24024 7328 24052
rect 11164 24052 11192 24092
rect 11238 24080 11244 24132
rect 11296 24080 11302 24132
rect 11698 24120 11704 24132
rect 11348 24092 11704 24120
rect 11348 24052 11376 24092
rect 11698 24080 11704 24092
rect 11756 24080 11762 24132
rect 11164 24024 11376 24052
rect 5960 24012 5966 24024
rect 11606 24012 11612 24064
rect 11664 24052 11670 24064
rect 12713 24055 12771 24061
rect 12713 24052 12725 24055
rect 11664 24024 12725 24052
rect 11664 24012 11670 24024
rect 12713 24021 12725 24024
rect 12759 24052 12771 24055
rect 12912 24052 12940 24160
rect 12986 24129 12992 24132
rect 12973 24123 12992 24129
rect 12973 24089 12985 24123
rect 12973 24083 12992 24089
rect 12986 24080 12992 24083
rect 13044 24080 13050 24132
rect 13188 24129 13216 24160
rect 15654 24148 15660 24200
rect 15712 24148 15718 24200
rect 16206 24148 16212 24200
rect 16264 24188 16270 24200
rect 17236 24188 17264 24364
rect 17402 24352 17408 24364
rect 17460 24352 17466 24404
rect 19150 24352 19156 24404
rect 19208 24392 19214 24404
rect 19245 24395 19303 24401
rect 19245 24392 19257 24395
rect 19208 24364 19257 24392
rect 19208 24352 19214 24364
rect 19245 24361 19257 24364
rect 19291 24361 19303 24395
rect 19245 24355 19303 24361
rect 21266 24352 21272 24404
rect 21324 24392 21330 24404
rect 21729 24395 21787 24401
rect 21729 24392 21741 24395
rect 21324 24364 21741 24392
rect 21324 24352 21330 24364
rect 21729 24361 21741 24364
rect 21775 24361 21787 24395
rect 21729 24355 21787 24361
rect 26421 24395 26479 24401
rect 26421 24361 26433 24395
rect 26467 24392 26479 24395
rect 26970 24392 26976 24404
rect 26467 24364 26976 24392
rect 26467 24361 26479 24364
rect 26421 24355 26479 24361
rect 26970 24352 26976 24364
rect 27028 24352 27034 24404
rect 21450 24284 21456 24336
rect 21508 24324 21514 24336
rect 22002 24324 22008 24336
rect 21508 24296 22008 24324
rect 21508 24284 21514 24296
rect 22002 24284 22008 24296
rect 22060 24324 22066 24336
rect 22419 24327 22477 24333
rect 22419 24324 22431 24327
rect 22060 24296 22431 24324
rect 22060 24284 22066 24296
rect 22419 24293 22431 24296
rect 22465 24293 22477 24327
rect 22419 24287 22477 24293
rect 26234 24284 26240 24336
rect 26292 24284 26298 24336
rect 17313 24259 17371 24265
rect 17313 24225 17325 24259
rect 17359 24256 17371 24259
rect 17586 24256 17592 24268
rect 17359 24228 17592 24256
rect 17359 24225 17371 24228
rect 17313 24219 17371 24225
rect 17586 24216 17592 24228
rect 17644 24216 17650 24268
rect 19518 24216 19524 24268
rect 19576 24256 19582 24268
rect 19797 24259 19855 24265
rect 19797 24256 19809 24259
rect 19576 24228 19809 24256
rect 19576 24216 19582 24228
rect 19797 24225 19809 24228
rect 19843 24225 19855 24259
rect 19797 24219 19855 24225
rect 21174 24216 21180 24268
rect 21232 24256 21238 24268
rect 21269 24259 21327 24265
rect 21269 24256 21281 24259
rect 21232 24228 21281 24256
rect 21232 24216 21238 24228
rect 21269 24225 21281 24228
rect 21315 24256 21327 24259
rect 21913 24259 21971 24265
rect 21913 24256 21925 24259
rect 21315 24228 21925 24256
rect 21315 24225 21327 24228
rect 21269 24219 21327 24225
rect 21913 24225 21925 24228
rect 21959 24225 21971 24259
rect 21913 24219 21971 24225
rect 24026 24216 24032 24268
rect 24084 24256 24090 24268
rect 24213 24259 24271 24265
rect 24213 24256 24225 24259
rect 24084 24228 24225 24256
rect 24084 24216 24090 24228
rect 24213 24225 24225 24228
rect 24259 24225 24271 24259
rect 24213 24219 24271 24225
rect 25501 24259 25559 24265
rect 25501 24225 25513 24259
rect 25547 24225 25559 24259
rect 25501 24219 25559 24225
rect 16264 24160 17264 24188
rect 16264 24148 16270 24160
rect 20162 24148 20168 24200
rect 20220 24188 20226 24200
rect 20625 24191 20683 24197
rect 20625 24188 20637 24191
rect 20220 24160 20637 24188
rect 20220 24148 20226 24160
rect 20625 24157 20637 24160
rect 20671 24157 20683 24191
rect 20625 24151 20683 24157
rect 20993 24191 21051 24197
rect 20993 24157 21005 24191
rect 21039 24157 21051 24191
rect 20993 24151 21051 24157
rect 13173 24123 13231 24129
rect 13173 24089 13185 24123
rect 13219 24089 13231 24123
rect 13173 24083 13231 24089
rect 14550 24080 14556 24132
rect 14608 24080 14614 24132
rect 12759 24024 12940 24052
rect 12759 24021 12771 24024
rect 12713 24015 12771 24021
rect 13354 24012 13360 24064
rect 13412 24052 13418 24064
rect 15672 24052 15700 24148
rect 16298 24080 16304 24132
rect 16356 24080 16362 24132
rect 17589 24123 17647 24129
rect 17589 24089 17601 24123
rect 17635 24089 17647 24123
rect 17589 24083 17647 24089
rect 13412 24024 15700 24052
rect 17604 24052 17632 24083
rect 18046 24080 18052 24132
rect 18104 24080 18110 24132
rect 20073 24123 20131 24129
rect 20073 24120 20085 24123
rect 18892 24092 20085 24120
rect 18892 24052 18920 24092
rect 20073 24089 20085 24092
rect 20119 24089 20131 24123
rect 21008 24120 21036 24151
rect 21082 24148 21088 24200
rect 21140 24148 21146 24200
rect 21361 24191 21419 24197
rect 21361 24157 21373 24191
rect 21407 24157 21419 24191
rect 21361 24151 21419 24157
rect 20073 24083 20131 24089
rect 20180 24092 21036 24120
rect 17604 24024 18920 24052
rect 19061 24055 19119 24061
rect 13412 24012 13418 24024
rect 19061 24021 19073 24055
rect 19107 24052 19119 24055
rect 19426 24052 19432 24064
rect 19107 24024 19432 24052
rect 19107 24021 19119 24024
rect 19061 24015 19119 24021
rect 19426 24012 19432 24024
rect 19484 24012 19490 24064
rect 19610 24012 19616 24064
rect 19668 24012 19674 24064
rect 19702 24012 19708 24064
rect 19760 24052 19766 24064
rect 20180 24052 20208 24092
rect 21266 24080 21272 24132
rect 21324 24120 21330 24132
rect 21376 24120 21404 24151
rect 21450 24148 21456 24200
rect 21508 24148 21514 24200
rect 21542 24148 21548 24200
rect 21600 24148 21606 24200
rect 21726 24148 21732 24200
rect 21784 24148 21790 24200
rect 22005 24191 22063 24197
rect 22005 24157 22017 24191
rect 22051 24157 22063 24191
rect 22005 24151 22063 24157
rect 21324 24092 21404 24120
rect 21560 24120 21588 24148
rect 22020 24120 22048 24151
rect 22278 24148 22284 24200
rect 22336 24148 22342 24200
rect 23845 24191 23903 24197
rect 23845 24157 23857 24191
rect 23891 24188 23903 24191
rect 25516 24188 25544 24219
rect 25590 24216 25596 24268
rect 25648 24256 25654 24268
rect 25961 24259 26019 24265
rect 25961 24256 25973 24259
rect 25648 24228 25973 24256
rect 25648 24216 25654 24228
rect 25961 24225 25973 24228
rect 26007 24225 26019 24259
rect 26252 24256 26280 24284
rect 26510 24256 26516 24268
rect 26252 24228 26516 24256
rect 25961 24219 26019 24225
rect 26510 24216 26516 24228
rect 26568 24216 26574 24268
rect 26786 24216 26792 24268
rect 26844 24216 26850 24268
rect 23891 24160 25544 24188
rect 25685 24191 25743 24197
rect 23891 24157 23903 24160
rect 23845 24151 23903 24157
rect 25685 24157 25697 24191
rect 25731 24157 25743 24191
rect 25685 24151 25743 24157
rect 25777 24191 25835 24197
rect 25777 24157 25789 24191
rect 25823 24157 25835 24191
rect 25777 24151 25835 24157
rect 21560 24092 22048 24120
rect 21324 24080 21330 24092
rect 22830 24080 22836 24132
rect 22888 24080 22894 24132
rect 19760 24024 20208 24052
rect 20809 24055 20867 24061
rect 19760 24012 19766 24024
rect 20809 24021 20821 24055
rect 20855 24052 20867 24055
rect 20990 24052 20996 24064
rect 20855 24024 20996 24052
rect 20855 24021 20867 24024
rect 20809 24015 20867 24021
rect 20990 24012 20996 24024
rect 21048 24012 21054 24064
rect 21634 24012 21640 24064
rect 21692 24052 21698 24064
rect 22189 24055 22247 24061
rect 22189 24052 22201 24055
rect 21692 24024 22201 24052
rect 21692 24012 21698 24024
rect 22189 24021 22201 24024
rect 22235 24021 22247 24055
rect 25700 24052 25728 24151
rect 25792 24120 25820 24151
rect 25866 24148 25872 24200
rect 25924 24148 25930 24200
rect 26237 24191 26295 24197
rect 26237 24157 26249 24191
rect 26283 24188 26295 24191
rect 26283 24160 26317 24188
rect 26283 24157 26295 24160
rect 26237 24151 26295 24157
rect 26252 24120 26280 24151
rect 26418 24148 26424 24200
rect 26476 24148 26482 24200
rect 25792 24092 26280 24120
rect 26142 24052 26148 24064
rect 25700 24024 26148 24052
rect 22189 24015 22247 24021
rect 26142 24012 26148 24024
rect 26200 24012 26206 24064
rect 26252 24052 26280 24092
rect 27798 24080 27804 24132
rect 27856 24080 27862 24132
rect 26418 24052 26424 24064
rect 26252 24024 26424 24052
rect 26418 24012 26424 24024
rect 26476 24052 26482 24064
rect 28261 24055 28319 24061
rect 28261 24052 28273 24055
rect 26476 24024 28273 24052
rect 26476 24012 26482 24024
rect 28261 24021 28273 24024
rect 28307 24021 28319 24055
rect 28261 24015 28319 24021
rect 1104 23962 28704 23984
rect 1104 23910 4874 23962
rect 4926 23910 4938 23962
rect 4990 23910 5002 23962
rect 5054 23910 5066 23962
rect 5118 23910 5130 23962
rect 5182 23910 28704 23962
rect 1104 23888 28704 23910
rect 9214 23808 9220 23860
rect 9272 23808 9278 23860
rect 10042 23808 10048 23860
rect 10100 23848 10106 23860
rect 12253 23851 12311 23857
rect 12253 23848 12265 23851
rect 10100 23820 12265 23848
rect 10100 23808 10106 23820
rect 12253 23817 12265 23820
rect 12299 23817 12311 23851
rect 12253 23811 12311 23817
rect 14182 23808 14188 23860
rect 14240 23848 14246 23860
rect 15197 23851 15255 23857
rect 15197 23848 15209 23851
rect 14240 23820 15209 23848
rect 14240 23808 14246 23820
rect 15197 23817 15209 23820
rect 15243 23817 15255 23851
rect 15197 23811 15255 23817
rect 15933 23851 15991 23857
rect 15933 23817 15945 23851
rect 15979 23848 15991 23851
rect 16206 23848 16212 23860
rect 15979 23820 16212 23848
rect 15979 23817 15991 23820
rect 15933 23811 15991 23817
rect 16206 23808 16212 23820
rect 16264 23808 16270 23860
rect 16758 23808 16764 23860
rect 16816 23808 16822 23860
rect 19337 23851 19395 23857
rect 19337 23817 19349 23851
rect 19383 23848 19395 23851
rect 19702 23848 19708 23860
rect 19383 23820 19708 23848
rect 19383 23817 19395 23820
rect 19337 23811 19395 23817
rect 19702 23808 19708 23820
rect 19760 23808 19766 23860
rect 20162 23808 20168 23860
rect 20220 23808 20226 23860
rect 21082 23808 21088 23860
rect 21140 23848 21146 23860
rect 22557 23851 22615 23857
rect 22557 23848 22569 23851
rect 21140 23820 22569 23848
rect 21140 23808 21146 23820
rect 22557 23817 22569 23820
rect 22603 23848 22615 23851
rect 25590 23848 25596 23860
rect 22603 23820 25596 23848
rect 22603 23817 22615 23820
rect 22557 23811 22615 23817
rect 25590 23808 25596 23820
rect 25648 23808 25654 23860
rect 25866 23808 25872 23860
rect 25924 23848 25930 23860
rect 27065 23851 27123 23857
rect 27065 23848 27077 23851
rect 25924 23820 27077 23848
rect 25924 23808 25930 23820
rect 27065 23817 27077 23820
rect 27111 23817 27123 23851
rect 27065 23811 27123 23817
rect 8941 23783 8999 23789
rect 8941 23749 8953 23783
rect 8987 23780 8999 23783
rect 9858 23780 9864 23792
rect 8987 23752 9864 23780
rect 8987 23749 8999 23752
rect 8941 23743 8999 23749
rect 9858 23740 9864 23752
rect 9916 23780 9922 23792
rect 13446 23780 13452 23792
rect 9916 23752 11928 23780
rect 9916 23740 9922 23752
rect 9122 23672 9128 23724
rect 9180 23672 9186 23724
rect 9217 23715 9275 23721
rect 9217 23681 9229 23715
rect 9263 23712 9275 23715
rect 9766 23712 9772 23724
rect 9263 23684 9772 23712
rect 9263 23681 9275 23684
rect 9217 23675 9275 23681
rect 9766 23672 9772 23684
rect 9824 23672 9830 23724
rect 10980 23721 11008 23752
rect 10965 23715 11023 23721
rect 10965 23681 10977 23715
rect 11011 23681 11023 23715
rect 10965 23675 11023 23681
rect 11054 23672 11060 23724
rect 11112 23672 11118 23724
rect 11241 23715 11299 23721
rect 11241 23681 11253 23715
rect 11287 23712 11299 23715
rect 11606 23712 11612 23724
rect 11287 23684 11612 23712
rect 11287 23681 11299 23684
rect 11241 23675 11299 23681
rect 11606 23672 11612 23684
rect 11664 23672 11670 23724
rect 11900 23721 11928 23752
rect 12176 23752 13452 23780
rect 12176 23724 12204 23752
rect 13446 23740 13452 23752
rect 13504 23740 13510 23792
rect 17862 23740 17868 23792
rect 17920 23740 17926 23792
rect 17954 23740 17960 23792
rect 18012 23780 18018 23792
rect 18012 23752 18354 23780
rect 18012 23740 18018 23752
rect 19610 23740 19616 23792
rect 19668 23780 19674 23792
rect 20257 23783 20315 23789
rect 20257 23780 20269 23783
rect 19668 23752 20269 23780
rect 19668 23740 19674 23752
rect 20257 23749 20269 23752
rect 20303 23749 20315 23783
rect 21266 23780 21272 23792
rect 20257 23743 20315 23749
rect 20364 23752 21272 23780
rect 11885 23715 11943 23721
rect 11885 23681 11897 23715
rect 11931 23681 11943 23715
rect 11885 23675 11943 23681
rect 12158 23672 12164 23724
rect 12216 23672 12222 23724
rect 12345 23715 12403 23721
rect 12345 23681 12357 23715
rect 12391 23712 12403 23715
rect 12986 23712 12992 23724
rect 12391 23684 12992 23712
rect 12391 23681 12403 23684
rect 12345 23675 12403 23681
rect 9140 23576 9168 23672
rect 11149 23647 11207 23653
rect 11149 23613 11161 23647
rect 11195 23644 11207 23647
rect 11701 23647 11759 23653
rect 11701 23644 11713 23647
rect 11195 23616 11713 23644
rect 11195 23613 11207 23616
rect 11149 23607 11207 23613
rect 11701 23613 11713 23616
rect 11747 23644 11759 23647
rect 11974 23644 11980 23656
rect 11747 23616 11980 23644
rect 11747 23613 11759 23616
rect 11701 23607 11759 23613
rect 11974 23604 11980 23616
rect 12032 23604 12038 23656
rect 12069 23647 12127 23653
rect 12069 23613 12081 23647
rect 12115 23644 12127 23647
rect 12360 23644 12388 23675
rect 12986 23672 12992 23684
rect 13044 23672 13050 23724
rect 15841 23715 15899 23721
rect 15841 23681 15853 23715
rect 15887 23712 15899 23715
rect 16022 23712 16028 23724
rect 15887 23684 16028 23712
rect 15887 23681 15899 23684
rect 15841 23675 15899 23681
rect 16022 23672 16028 23684
rect 16080 23672 16086 23724
rect 16114 23672 16120 23724
rect 16172 23672 16178 23724
rect 16298 23672 16304 23724
rect 16356 23672 16362 23724
rect 16669 23715 16727 23721
rect 16669 23681 16681 23715
rect 16715 23681 16727 23715
rect 16669 23675 16727 23681
rect 12115 23616 12388 23644
rect 16132 23644 16160 23672
rect 16684 23644 16712 23675
rect 16850 23672 16856 23724
rect 16908 23672 16914 23724
rect 19426 23672 19432 23724
rect 19484 23712 19490 23724
rect 19705 23715 19763 23721
rect 19705 23712 19717 23715
rect 19484 23684 19717 23712
rect 19484 23672 19490 23684
rect 19705 23681 19717 23684
rect 19751 23681 19763 23715
rect 19705 23675 19763 23681
rect 16132 23616 16712 23644
rect 12115 23613 12127 23616
rect 12069 23607 12127 23613
rect 17586 23604 17592 23656
rect 17644 23604 17650 23656
rect 19521 23647 19579 23653
rect 19521 23644 19533 23647
rect 17696 23616 19533 23644
rect 11514 23576 11520 23588
rect 9140 23548 11520 23576
rect 11514 23536 11520 23548
rect 11572 23576 11578 23588
rect 12158 23576 12164 23588
rect 11572 23548 12164 23576
rect 11572 23536 11578 23548
rect 12158 23536 12164 23548
rect 12216 23536 12222 23588
rect 17126 23536 17132 23588
rect 17184 23576 17190 23588
rect 17696 23576 17724 23616
rect 19521 23613 19533 23616
rect 19567 23644 19579 23647
rect 19610 23644 19616 23656
rect 19567 23616 19616 23644
rect 19567 23613 19579 23616
rect 19521 23607 19579 23613
rect 19610 23604 19616 23616
rect 19668 23604 19674 23656
rect 19720 23644 19748 23675
rect 19794 23672 19800 23724
rect 19852 23672 19858 23724
rect 20364 23644 20392 23752
rect 21266 23740 21272 23752
rect 21324 23740 21330 23792
rect 22922 23780 22928 23792
rect 22296 23752 22928 23780
rect 20990 23672 20996 23724
rect 21048 23672 21054 23724
rect 21174 23721 21180 23724
rect 21141 23715 21180 23721
rect 21141 23681 21153 23715
rect 21141 23675 21180 23681
rect 21174 23672 21180 23675
rect 21232 23672 21238 23724
rect 21358 23672 21364 23724
rect 21416 23672 21422 23724
rect 21499 23715 21557 23721
rect 21499 23681 21511 23715
rect 21545 23712 21557 23715
rect 21634 23712 21640 23724
rect 21545 23684 21640 23712
rect 21545 23681 21557 23684
rect 21499 23675 21557 23681
rect 21634 23672 21640 23684
rect 21692 23672 21698 23724
rect 22296 23721 22324 23752
rect 22922 23740 22928 23752
rect 22980 23740 22986 23792
rect 26326 23740 26332 23792
rect 26384 23780 26390 23792
rect 26384 23752 26648 23780
rect 26384 23740 26390 23752
rect 22281 23715 22339 23721
rect 22281 23681 22293 23715
rect 22327 23681 22339 23715
rect 22281 23675 22339 23681
rect 22649 23715 22707 23721
rect 22649 23681 22661 23715
rect 22695 23681 22707 23715
rect 22649 23675 22707 23681
rect 19720 23616 20392 23644
rect 20806 23604 20812 23656
rect 20864 23604 20870 23656
rect 22002 23604 22008 23656
rect 22060 23644 22066 23656
rect 22664 23644 22692 23675
rect 25682 23672 25688 23724
rect 25740 23672 25746 23724
rect 26418 23672 26424 23724
rect 26476 23672 26482 23724
rect 26620 23721 26648 23752
rect 27982 23740 27988 23792
rect 28040 23780 28046 23792
rect 28040 23752 28212 23780
rect 28040 23740 28046 23752
rect 26605 23715 26663 23721
rect 26605 23681 26617 23715
rect 26651 23681 26663 23715
rect 26605 23675 26663 23681
rect 26789 23715 26847 23721
rect 26789 23681 26801 23715
rect 26835 23712 26847 23715
rect 27154 23712 27160 23724
rect 26835 23684 27160 23712
rect 26835 23681 26847 23684
rect 26789 23675 26847 23681
rect 27154 23672 27160 23684
rect 27212 23712 27218 23724
rect 28184 23721 28212 23752
rect 28169 23715 28227 23721
rect 27212 23684 28120 23712
rect 27212 23672 27218 23684
rect 22060 23616 22692 23644
rect 27709 23647 27767 23653
rect 22060 23604 22066 23616
rect 27709 23613 27721 23647
rect 27755 23644 27767 23647
rect 27890 23644 27896 23656
rect 27755 23616 27896 23644
rect 27755 23613 27767 23616
rect 27709 23607 27767 23613
rect 27890 23604 27896 23616
rect 27948 23604 27954 23656
rect 28092 23653 28120 23684
rect 28169 23681 28181 23715
rect 28215 23681 28227 23715
rect 28169 23675 28227 23681
rect 28077 23647 28135 23653
rect 28077 23613 28089 23647
rect 28123 23613 28135 23647
rect 28077 23607 28135 23613
rect 17184 23548 17724 23576
rect 17184 23536 17190 23548
rect 26878 23536 26884 23588
rect 26936 23576 26942 23588
rect 27801 23579 27859 23585
rect 27801 23576 27813 23579
rect 26936 23548 27813 23576
rect 26936 23536 26942 23548
rect 27801 23545 27813 23548
rect 27847 23545 27859 23579
rect 27801 23539 27859 23545
rect 10781 23511 10839 23517
rect 10781 23477 10793 23511
rect 10827 23508 10839 23511
rect 11146 23508 11152 23520
rect 10827 23480 11152 23508
rect 10827 23477 10839 23480
rect 10781 23471 10839 23477
rect 11146 23468 11152 23480
rect 11204 23468 11210 23520
rect 21634 23468 21640 23520
rect 21692 23468 21698 23520
rect 22094 23468 22100 23520
rect 22152 23508 22158 23520
rect 22189 23511 22247 23517
rect 22189 23508 22201 23511
rect 22152 23480 22201 23508
rect 22152 23468 22158 23480
rect 22189 23477 22201 23480
rect 22235 23477 22247 23511
rect 22189 23471 22247 23477
rect 25038 23468 25044 23520
rect 25096 23508 25102 23520
rect 25593 23511 25651 23517
rect 25593 23508 25605 23511
rect 25096 23480 25605 23508
rect 25096 23468 25102 23480
rect 25593 23477 25605 23480
rect 25639 23477 25651 23511
rect 25593 23471 25651 23477
rect 1104 23418 28704 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 28704 23418
rect 1104 23344 28704 23366
rect 11238 23264 11244 23316
rect 11296 23304 11302 23316
rect 11333 23307 11391 23313
rect 11333 23304 11345 23307
rect 11296 23276 11345 23304
rect 11296 23264 11302 23276
rect 11333 23273 11345 23276
rect 11379 23273 11391 23307
rect 11333 23267 11391 23273
rect 19794 23264 19800 23316
rect 19852 23304 19858 23316
rect 20165 23307 20223 23313
rect 20165 23304 20177 23307
rect 19852 23276 20177 23304
rect 19852 23264 19858 23276
rect 20165 23273 20177 23276
rect 20211 23273 20223 23307
rect 20165 23267 20223 23273
rect 27890 23264 27896 23316
rect 27948 23304 27954 23316
rect 28261 23307 28319 23313
rect 28261 23304 28273 23307
rect 27948 23276 28273 23304
rect 27948 23264 27954 23276
rect 28261 23273 28273 23276
rect 28307 23273 28319 23307
rect 28261 23267 28319 23273
rect 15289 23239 15347 23245
rect 15289 23205 15301 23239
rect 15335 23236 15347 23239
rect 15378 23236 15384 23248
rect 15335 23208 15384 23236
rect 15335 23205 15347 23208
rect 15289 23199 15347 23205
rect 15378 23196 15384 23208
rect 15436 23196 15442 23248
rect 18969 23239 19027 23245
rect 18969 23205 18981 23239
rect 19015 23236 19027 23239
rect 20806 23236 20812 23248
rect 19015 23208 20812 23236
rect 19015 23205 19027 23208
rect 18969 23199 19027 23205
rect 20806 23196 20812 23208
rect 20864 23196 20870 23248
rect 10962 23128 10968 23180
rect 11020 23128 11026 23180
rect 15746 23128 15752 23180
rect 15804 23168 15810 23180
rect 16025 23171 16083 23177
rect 16025 23168 16037 23171
rect 15804 23140 16037 23168
rect 15804 23128 15810 23140
rect 16025 23137 16037 23140
rect 16071 23168 16083 23171
rect 17126 23168 17132 23180
rect 16071 23140 17132 23168
rect 16071 23137 16083 23140
rect 16025 23131 16083 23137
rect 17126 23128 17132 23140
rect 17184 23128 17190 23180
rect 17221 23171 17279 23177
rect 17221 23137 17233 23171
rect 17267 23168 17279 23171
rect 17586 23168 17592 23180
rect 17267 23140 17592 23168
rect 17267 23137 17279 23140
rect 17221 23131 17279 23137
rect 17586 23128 17592 23140
rect 17644 23128 17650 23180
rect 21726 23128 21732 23180
rect 21784 23168 21790 23180
rect 21913 23171 21971 23177
rect 21913 23168 21925 23171
rect 21784 23140 21925 23168
rect 21784 23128 21790 23140
rect 21913 23137 21925 23140
rect 21959 23137 21971 23171
rect 21913 23131 21971 23137
rect 26510 23128 26516 23180
rect 26568 23128 26574 23180
rect 26789 23171 26847 23177
rect 26789 23137 26801 23171
rect 26835 23168 26847 23171
rect 26878 23168 26884 23180
rect 26835 23140 26884 23168
rect 26835 23137 26847 23140
rect 26789 23131 26847 23137
rect 26878 23128 26884 23140
rect 26936 23128 26942 23180
rect 11146 23060 11152 23112
rect 11204 23060 11210 23112
rect 15013 23103 15071 23109
rect 15013 23069 15025 23103
rect 15059 23100 15071 23103
rect 15102 23100 15108 23112
rect 15059 23072 15108 23100
rect 15059 23069 15071 23072
rect 15013 23063 15071 23069
rect 15102 23060 15108 23072
rect 15160 23060 15166 23112
rect 15838 23060 15844 23112
rect 15896 23060 15902 23112
rect 16114 23060 16120 23112
rect 16172 23060 16178 23112
rect 19334 23060 19340 23112
rect 19392 23100 19398 23112
rect 19521 23103 19579 23109
rect 19521 23100 19533 23103
rect 19392 23072 19533 23100
rect 19392 23060 19398 23072
rect 19521 23069 19533 23072
rect 19567 23069 19579 23103
rect 19521 23063 19579 23069
rect 21634 23060 21640 23112
rect 21692 23060 21698 23112
rect 21821 23103 21879 23109
rect 21821 23069 21833 23103
rect 21867 23069 21879 23103
rect 21821 23063 21879 23069
rect 22005 23103 22063 23109
rect 22005 23069 22017 23103
rect 22051 23100 22063 23103
rect 22094 23100 22100 23112
rect 22051 23072 22100 23100
rect 22051 23069 22063 23072
rect 22005 23063 22063 23069
rect 15286 22992 15292 23044
rect 15344 22992 15350 23044
rect 17494 22992 17500 23044
rect 17552 22992 17558 23044
rect 17954 22992 17960 23044
rect 18012 22992 18018 23044
rect 20990 22992 20996 23044
rect 21048 23032 21054 23044
rect 21358 23032 21364 23044
rect 21048 23004 21364 23032
rect 21048 22992 21054 23004
rect 21358 22992 21364 23004
rect 21416 23032 21422 23044
rect 21836 23032 21864 23063
rect 22094 23060 22100 23072
rect 22152 23060 22158 23112
rect 22189 23103 22247 23109
rect 22189 23069 22201 23103
rect 22235 23100 22247 23103
rect 22830 23100 22836 23112
rect 22235 23072 22836 23100
rect 22235 23069 22247 23072
rect 22189 23063 22247 23069
rect 22830 23060 22836 23072
rect 22888 23060 22894 23112
rect 26237 23103 26295 23109
rect 26237 23069 26249 23103
rect 26283 23100 26295 23103
rect 26418 23100 26424 23112
rect 26283 23072 26424 23100
rect 26283 23069 26295 23072
rect 26237 23063 26295 23069
rect 26418 23060 26424 23072
rect 26476 23060 26482 23112
rect 21416 23004 21864 23032
rect 21416 22992 21422 23004
rect 27798 22992 27804 23044
rect 27856 22992 27862 23044
rect 15105 22967 15163 22973
rect 15105 22933 15117 22967
rect 15151 22964 15163 22967
rect 15562 22964 15568 22976
rect 15151 22936 15568 22964
rect 15151 22933 15163 22936
rect 15105 22927 15163 22933
rect 15562 22924 15568 22936
rect 15620 22924 15626 22976
rect 22373 22967 22431 22973
rect 22373 22933 22385 22967
rect 22419 22964 22431 22967
rect 23934 22964 23940 22976
rect 22419 22936 23940 22964
rect 22419 22933 22431 22936
rect 22373 22927 22431 22933
rect 23934 22924 23940 22936
rect 23992 22924 23998 22976
rect 26326 22924 26332 22976
rect 26384 22924 26390 22976
rect 1104 22874 28704 22896
rect 1104 22822 4874 22874
rect 4926 22822 4938 22874
rect 4990 22822 5002 22874
rect 5054 22822 5066 22874
rect 5118 22822 5130 22874
rect 5182 22822 28704 22874
rect 1104 22800 28704 22822
rect 15286 22720 15292 22772
rect 15344 22760 15350 22772
rect 15657 22763 15715 22769
rect 15657 22760 15669 22763
rect 15344 22732 15669 22760
rect 15344 22720 15350 22732
rect 15657 22729 15669 22732
rect 15703 22729 15715 22763
rect 15657 22723 15715 22729
rect 17954 22720 17960 22772
rect 18012 22760 18018 22772
rect 18874 22760 18880 22772
rect 18012 22732 18880 22760
rect 18012 22720 18018 22732
rect 18874 22720 18880 22732
rect 18932 22720 18938 22772
rect 7837 22695 7895 22701
rect 7837 22661 7849 22695
rect 7883 22692 7895 22695
rect 8110 22692 8116 22704
rect 7883 22664 8116 22692
rect 7883 22661 7895 22664
rect 7837 22655 7895 22661
rect 8110 22652 8116 22664
rect 8168 22652 8174 22704
rect 13262 22652 13268 22704
rect 13320 22652 13326 22704
rect 14921 22695 14979 22701
rect 14921 22661 14933 22695
rect 14967 22692 14979 22695
rect 15838 22692 15844 22704
rect 14967 22664 15844 22692
rect 14967 22661 14979 22664
rect 14921 22655 14979 22661
rect 15838 22652 15844 22664
rect 15896 22652 15902 22704
rect 22094 22652 22100 22704
rect 22152 22692 22158 22704
rect 24305 22695 24363 22701
rect 22152 22664 24072 22692
rect 22152 22652 22158 22664
rect 7469 22627 7527 22633
rect 7469 22593 7481 22627
rect 7515 22593 7527 22627
rect 7469 22587 7527 22593
rect 7484 22556 7512 22587
rect 7742 22584 7748 22636
rect 7800 22584 7806 22636
rect 8021 22627 8079 22633
rect 8021 22593 8033 22627
rect 8067 22624 8079 22627
rect 9674 22624 9680 22636
rect 8067 22596 9680 22624
rect 8067 22593 8079 22596
rect 8021 22587 8079 22593
rect 9674 22584 9680 22596
rect 9732 22584 9738 22636
rect 12161 22627 12219 22633
rect 12161 22593 12173 22627
rect 12207 22624 12219 22627
rect 13078 22624 13084 22636
rect 12207 22596 13084 22624
rect 12207 22593 12219 22596
rect 12161 22587 12219 22593
rect 13078 22584 13084 22596
rect 13136 22584 13142 22636
rect 14090 22584 14096 22636
rect 14148 22584 14154 22636
rect 15105 22627 15163 22633
rect 15105 22593 15117 22627
rect 15151 22593 15163 22627
rect 15105 22587 15163 22593
rect 15197 22627 15255 22633
rect 15197 22593 15209 22627
rect 15243 22593 15255 22627
rect 15197 22587 15255 22593
rect 14277 22559 14335 22565
rect 7484 22528 7880 22556
rect 7852 22500 7880 22528
rect 14277 22525 14289 22559
rect 14323 22556 14335 22559
rect 15010 22556 15016 22568
rect 14323 22528 15016 22556
rect 14323 22525 14335 22528
rect 14277 22519 14335 22525
rect 15010 22516 15016 22528
rect 15068 22516 15074 22568
rect 7834 22448 7840 22500
rect 7892 22448 7898 22500
rect 15120 22488 15148 22587
rect 15212 22556 15240 22587
rect 15286 22584 15292 22636
rect 15344 22584 15350 22636
rect 15378 22584 15384 22636
rect 15436 22624 15442 22636
rect 17221 22627 17279 22633
rect 17221 22624 17233 22627
rect 15436 22596 17233 22624
rect 15436 22584 15442 22596
rect 17221 22593 17233 22596
rect 17267 22593 17279 22627
rect 17221 22587 17279 22593
rect 23934 22584 23940 22636
rect 23992 22584 23998 22636
rect 24044 22633 24072 22664
rect 24305 22661 24317 22695
rect 24351 22692 24363 22695
rect 24578 22692 24584 22704
rect 24351 22664 24584 22692
rect 24351 22661 24363 22664
rect 24305 22655 24363 22661
rect 24578 22652 24584 22664
rect 24636 22692 24642 22704
rect 26237 22695 26295 22701
rect 24636 22664 24900 22692
rect 24636 22652 24642 22664
rect 24872 22633 24900 22664
rect 26237 22661 26249 22695
rect 26283 22692 26295 22695
rect 28350 22692 28356 22704
rect 26283 22664 28356 22692
rect 26283 22661 26295 22664
rect 26237 22655 26295 22661
rect 28350 22652 28356 22664
rect 28408 22652 28414 22704
rect 24030 22627 24088 22633
rect 24030 22593 24042 22627
rect 24076 22593 24088 22627
rect 24030 22587 24088 22593
rect 24213 22627 24271 22633
rect 24213 22593 24225 22627
rect 24259 22593 24271 22627
rect 24213 22587 24271 22593
rect 24402 22627 24460 22633
rect 24402 22593 24414 22627
rect 24448 22624 24460 22627
rect 24673 22627 24731 22633
rect 24673 22624 24685 22627
rect 24448 22596 24532 22624
rect 24448 22593 24460 22596
rect 24402 22587 24460 22593
rect 15930 22556 15936 22568
rect 15212 22528 15936 22556
rect 15930 22516 15936 22528
rect 15988 22556 15994 22568
rect 16209 22559 16267 22565
rect 16209 22556 16221 22559
rect 15988 22528 16221 22556
rect 15988 22516 15994 22528
rect 16209 22525 16221 22528
rect 16255 22525 16267 22559
rect 16209 22519 16267 22525
rect 20346 22516 20352 22568
rect 20404 22516 20410 22568
rect 22370 22516 22376 22568
rect 22428 22516 22434 22568
rect 23474 22516 23480 22568
rect 23532 22556 23538 22568
rect 23753 22559 23811 22565
rect 23753 22556 23765 22559
rect 23532 22528 23765 22556
rect 23532 22516 23538 22528
rect 23753 22525 23765 22528
rect 23799 22525 23811 22559
rect 23753 22519 23811 22525
rect 15562 22488 15568 22500
rect 15120 22460 15568 22488
rect 15562 22448 15568 22460
rect 15620 22488 15626 22500
rect 16482 22488 16488 22500
rect 15620 22460 16488 22488
rect 15620 22448 15626 22460
rect 16482 22448 16488 22460
rect 16540 22448 16546 22500
rect 22830 22448 22836 22500
rect 22888 22488 22894 22500
rect 24228 22488 24256 22587
rect 22888 22460 24256 22488
rect 22888 22448 22894 22460
rect 8021 22423 8079 22429
rect 8021 22389 8033 22423
rect 8067 22420 8079 22423
rect 9030 22420 9036 22432
rect 8067 22392 9036 22420
rect 8067 22389 8079 22392
rect 8021 22383 8079 22389
rect 9030 22380 9036 22392
rect 9088 22380 9094 22432
rect 11977 22423 12035 22429
rect 11977 22389 11989 22423
rect 12023 22420 12035 22423
rect 12066 22420 12072 22432
rect 12023 22392 12072 22420
rect 12023 22389 12035 22392
rect 11977 22383 12035 22389
rect 12066 22380 12072 22392
rect 12124 22380 12130 22432
rect 14366 22380 14372 22432
rect 14424 22420 14430 22432
rect 14829 22423 14887 22429
rect 14829 22420 14841 22423
rect 14424 22392 14841 22420
rect 14424 22380 14430 22392
rect 14829 22389 14841 22392
rect 14875 22389 14887 22423
rect 14829 22383 14887 22389
rect 15194 22380 15200 22432
rect 15252 22380 15258 22432
rect 15470 22380 15476 22432
rect 15528 22380 15534 22432
rect 16666 22380 16672 22432
rect 16724 22380 16730 22432
rect 19518 22380 19524 22432
rect 19576 22420 19582 22432
rect 19797 22423 19855 22429
rect 19797 22420 19809 22423
rect 19576 22392 19809 22420
rect 19576 22380 19582 22392
rect 19797 22389 19809 22392
rect 19843 22389 19855 22423
rect 19797 22383 19855 22389
rect 21818 22380 21824 22432
rect 21876 22380 21882 22432
rect 23014 22380 23020 22432
rect 23072 22420 23078 22432
rect 23201 22423 23259 22429
rect 23201 22420 23213 22423
rect 23072 22392 23213 22420
rect 23072 22380 23078 22392
rect 23201 22389 23213 22392
rect 23247 22389 23259 22423
rect 24504 22420 24532 22596
rect 24596 22596 24685 22624
rect 24596 22497 24624 22596
rect 24673 22593 24685 22596
rect 24719 22593 24731 22627
rect 24673 22587 24731 22593
rect 24857 22627 24915 22633
rect 24857 22593 24869 22627
rect 24903 22593 24915 22627
rect 24857 22587 24915 22593
rect 24946 22584 24952 22636
rect 25004 22584 25010 22636
rect 25222 22584 25228 22636
rect 25280 22584 25286 22636
rect 26418 22584 26424 22636
rect 26476 22584 26482 22636
rect 26513 22627 26571 22633
rect 26513 22593 26525 22627
rect 26559 22593 26571 22627
rect 26513 22587 26571 22593
rect 26789 22627 26847 22633
rect 26789 22593 26801 22627
rect 26835 22624 26847 22627
rect 27709 22627 27767 22633
rect 27709 22624 27721 22627
rect 26835 22596 27721 22624
rect 26835 22593 26847 22596
rect 26789 22587 26847 22593
rect 27709 22593 27721 22596
rect 27755 22624 27767 22627
rect 27890 22624 27896 22636
rect 27755 22596 27896 22624
rect 27755 22593 27767 22596
rect 27709 22587 27767 22593
rect 25038 22516 25044 22568
rect 25096 22516 25102 22568
rect 25590 22516 25596 22568
rect 25648 22516 25654 22568
rect 26326 22516 26332 22568
rect 26384 22556 26390 22568
rect 26528 22556 26556 22587
rect 27890 22584 27896 22596
rect 27948 22584 27954 22636
rect 27430 22556 27436 22568
rect 26384 22528 27436 22556
rect 26384 22516 26390 22528
rect 27430 22516 27436 22528
rect 27488 22516 27494 22568
rect 27614 22516 27620 22568
rect 27672 22516 27678 22568
rect 24581 22491 24639 22497
rect 24581 22457 24593 22491
rect 24627 22457 24639 22491
rect 24581 22451 24639 22457
rect 25409 22491 25467 22497
rect 25409 22457 25421 22491
rect 25455 22488 25467 22491
rect 26602 22488 26608 22500
rect 25455 22460 26608 22488
rect 25455 22457 25467 22460
rect 25409 22451 25467 22457
rect 26602 22448 26608 22460
rect 26660 22448 26666 22500
rect 26697 22491 26755 22497
rect 26697 22457 26709 22491
rect 26743 22488 26755 22491
rect 27982 22488 27988 22500
rect 26743 22460 27988 22488
rect 26743 22457 26755 22460
rect 26697 22451 26755 22457
rect 27982 22448 27988 22460
rect 28040 22448 28046 22500
rect 24854 22420 24860 22432
rect 24504 22392 24860 22420
rect 23201 22383 23259 22389
rect 24854 22380 24860 22392
rect 24912 22380 24918 22432
rect 26142 22380 26148 22432
rect 26200 22380 26206 22432
rect 26970 22380 26976 22432
rect 27028 22380 27034 22432
rect 28074 22380 28080 22432
rect 28132 22420 28138 22432
rect 28353 22423 28411 22429
rect 28353 22420 28365 22423
rect 28132 22392 28365 22420
rect 28132 22380 28138 22392
rect 28353 22389 28365 22392
rect 28399 22389 28411 22423
rect 28353 22383 28411 22389
rect 1104 22330 28704 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 28704 22330
rect 1104 22256 28704 22278
rect 15930 22176 15936 22228
rect 15988 22176 15994 22228
rect 16209 22219 16267 22225
rect 16209 22185 16221 22219
rect 16255 22216 16267 22219
rect 16482 22216 16488 22228
rect 16255 22188 16488 22216
rect 16255 22185 16267 22188
rect 16209 22179 16267 22185
rect 16482 22176 16488 22188
rect 16540 22176 16546 22228
rect 19518 22225 19524 22228
rect 19508 22219 19524 22225
rect 19508 22185 19520 22219
rect 19508 22179 19524 22185
rect 19518 22176 19524 22179
rect 19576 22176 19582 22228
rect 21348 22219 21406 22225
rect 21348 22185 21360 22219
rect 21394 22216 21406 22219
rect 21818 22216 21824 22228
rect 21394 22188 21824 22216
rect 21394 22185 21406 22188
rect 21348 22179 21406 22185
rect 21818 22176 21824 22188
rect 21876 22176 21882 22228
rect 22830 22176 22836 22228
rect 22888 22176 22894 22228
rect 25979 22219 26037 22225
rect 25979 22185 25991 22219
rect 26025 22216 26037 22219
rect 26142 22216 26148 22228
rect 26025 22188 26148 22216
rect 26025 22185 26037 22188
rect 25979 22179 26037 22185
rect 26142 22176 26148 22188
rect 26200 22176 26206 22228
rect 26592 22219 26650 22225
rect 26592 22185 26604 22219
rect 26638 22216 26650 22219
rect 26970 22216 26976 22228
rect 26638 22188 26976 22216
rect 26638 22185 26650 22188
rect 26592 22179 26650 22185
rect 26970 22176 26976 22188
rect 27028 22176 27034 22228
rect 16114 22108 16120 22160
rect 16172 22148 16178 22160
rect 16393 22151 16451 22157
rect 16393 22148 16405 22151
rect 16172 22120 16405 22148
rect 16172 22108 16178 22120
rect 16393 22117 16405 22120
rect 16439 22117 16451 22151
rect 16393 22111 16451 22117
rect 5813 22083 5871 22089
rect 5813 22049 5825 22083
rect 5859 22080 5871 22083
rect 5997 22083 6055 22089
rect 5997 22080 6009 22083
rect 5859 22052 6009 22080
rect 5859 22049 5871 22052
rect 5813 22043 5871 22049
rect 5997 22049 6009 22052
rect 6043 22080 6055 22083
rect 6914 22080 6920 22092
rect 6043 22052 6920 22080
rect 6043 22049 6055 22052
rect 5997 22043 6055 22049
rect 6914 22040 6920 22052
rect 6972 22080 6978 22092
rect 7926 22080 7932 22092
rect 6972 22052 7932 22080
rect 6972 22040 6978 22052
rect 7926 22040 7932 22052
rect 7984 22040 7990 22092
rect 8110 22040 8116 22092
rect 8168 22080 8174 22092
rect 9217 22083 9275 22089
rect 9217 22080 9229 22083
rect 8168 22052 9229 22080
rect 8168 22040 8174 22052
rect 9217 22049 9229 22052
rect 9263 22080 9275 22083
rect 11241 22083 11299 22089
rect 11241 22080 11253 22083
rect 9263 22052 11253 22080
rect 9263 22049 9275 22052
rect 9217 22043 9275 22049
rect 11241 22049 11253 22052
rect 11287 22049 11299 22083
rect 11241 22043 11299 22049
rect 12161 22083 12219 22089
rect 12161 22049 12173 22083
rect 12207 22080 12219 22083
rect 13170 22080 13176 22092
rect 12207 22052 13176 22080
rect 12207 22049 12219 22052
rect 12161 22043 12219 22049
rect 8570 22012 8576 22024
rect 7406 21984 8576 22012
rect 8570 21972 8576 21984
rect 8628 21972 8634 22024
rect 9309 22015 9367 22021
rect 9309 21981 9321 22015
rect 9355 22012 9367 22015
rect 10962 22012 10968 22024
rect 9355 21984 10968 22012
rect 9355 21981 9367 21984
rect 9309 21975 9367 21981
rect 10962 21972 10968 21984
rect 11020 22012 11026 22024
rect 11149 22015 11207 22021
rect 11149 22012 11161 22015
rect 11020 21984 11161 22012
rect 11020 21972 11026 21984
rect 11149 21981 11161 21984
rect 11195 21981 11207 22015
rect 11149 21975 11207 21981
rect 4798 21904 4804 21956
rect 4856 21904 4862 21956
rect 5534 21904 5540 21956
rect 5592 21904 5598 21956
rect 6270 21904 6276 21956
rect 6328 21904 6334 21956
rect 7834 21904 7840 21956
rect 7892 21904 7898 21956
rect 7926 21904 7932 21956
rect 7984 21944 7990 21956
rect 8665 21947 8723 21953
rect 8665 21944 8677 21947
rect 7984 21916 8677 21944
rect 7984 21904 7990 21916
rect 8665 21913 8677 21916
rect 8711 21944 8723 21947
rect 9582 21944 9588 21956
rect 8711 21916 9588 21944
rect 8711 21913 8723 21916
rect 8665 21907 8723 21913
rect 9582 21904 9588 21916
rect 9640 21904 9646 21956
rect 11256 21944 11284 22043
rect 13170 22040 13176 22052
rect 13228 22080 13234 22092
rect 14185 22083 14243 22089
rect 14185 22080 14197 22083
rect 13228 22052 14197 22080
rect 13228 22040 13234 22052
rect 14185 22049 14197 22052
rect 14231 22049 14243 22083
rect 14185 22043 14243 22049
rect 14461 22083 14519 22089
rect 14461 22049 14473 22083
rect 14507 22080 14519 22083
rect 16577 22083 16635 22089
rect 16577 22080 16589 22083
rect 14507 22052 16589 22080
rect 14507 22049 14519 22052
rect 14461 22043 14519 22049
rect 16577 22049 16589 22052
rect 16623 22049 16635 22083
rect 16577 22043 16635 22049
rect 17313 22083 17371 22089
rect 17313 22049 17325 22083
rect 17359 22080 17371 22083
rect 17586 22080 17592 22092
rect 17359 22052 17592 22080
rect 17359 22049 17371 22052
rect 17313 22043 17371 22049
rect 17586 22040 17592 22052
rect 17644 22080 17650 22092
rect 19242 22080 19248 22092
rect 17644 22052 19248 22080
rect 17644 22040 17650 22052
rect 19242 22040 19248 22052
rect 19300 22080 19306 22092
rect 21085 22083 21143 22089
rect 21085 22080 21097 22083
rect 19300 22052 21097 22080
rect 19300 22040 19306 22052
rect 21085 22049 21097 22052
rect 21131 22049 21143 22083
rect 21085 22043 21143 22049
rect 23937 22083 23995 22089
rect 23937 22049 23949 22083
rect 23983 22049 23995 22083
rect 23937 22043 23995 22049
rect 11422 21972 11428 22024
rect 11480 21972 11486 22024
rect 12066 21972 12072 22024
rect 12124 21972 12130 22024
rect 16114 21972 16120 22024
rect 16172 22012 16178 22024
rect 16485 22015 16543 22021
rect 16485 22012 16497 22015
rect 16172 21984 16497 22012
rect 16172 21972 16178 21984
rect 16485 21981 16497 21984
rect 16531 21981 16543 22015
rect 16485 21975 16543 21981
rect 16666 21972 16672 22024
rect 16724 21972 16730 22024
rect 23952 22012 23980 22043
rect 24026 22040 24032 22092
rect 24084 22080 24090 22092
rect 26237 22083 26295 22089
rect 26237 22080 26249 22083
rect 24084 22052 26249 22080
rect 24084 22040 24090 22052
rect 26237 22049 26249 22052
rect 26283 22080 26295 22083
rect 26329 22083 26387 22089
rect 26329 22080 26341 22083
rect 26283 22052 26341 22080
rect 26283 22049 26295 22052
rect 26237 22043 26295 22049
rect 26329 22049 26341 22052
rect 26375 22049 26387 22083
rect 26329 22043 26387 22049
rect 24210 22012 24216 22024
rect 23952 21984 24216 22012
rect 24210 21972 24216 21984
rect 24268 21972 24274 22024
rect 11256 21916 12020 21944
rect 4062 21836 4068 21888
rect 4120 21836 4126 21888
rect 7006 21836 7012 21888
rect 7064 21876 7070 21888
rect 7745 21879 7803 21885
rect 7745 21876 7757 21879
rect 7064 21848 7757 21876
rect 7064 21836 7070 21848
rect 7745 21845 7757 21848
rect 7791 21845 7803 21879
rect 7745 21839 7803 21845
rect 8941 21879 8999 21885
rect 8941 21845 8953 21879
rect 8987 21876 8999 21879
rect 9122 21876 9128 21888
rect 8987 21848 9128 21876
rect 8987 21845 8999 21848
rect 8941 21839 8999 21845
rect 9122 21836 9128 21848
rect 9180 21836 9186 21888
rect 11609 21879 11667 21885
rect 11609 21845 11621 21879
rect 11655 21876 11667 21879
rect 11790 21876 11796 21888
rect 11655 21848 11796 21876
rect 11655 21845 11667 21848
rect 11609 21839 11667 21845
rect 11790 21836 11796 21848
rect 11848 21836 11854 21888
rect 11882 21836 11888 21888
rect 11940 21836 11946 21888
rect 11992 21876 12020 21916
rect 12434 21904 12440 21956
rect 12492 21904 12498 21956
rect 12894 21904 12900 21956
rect 12952 21904 12958 21956
rect 15470 21904 15476 21956
rect 15528 21904 15534 21956
rect 15930 21904 15936 21956
rect 15988 21944 15994 21956
rect 16025 21947 16083 21953
rect 16025 21944 16037 21947
rect 15988 21916 16037 21944
rect 15988 21904 15994 21916
rect 16025 21913 16037 21916
rect 16071 21913 16083 21947
rect 16025 21907 16083 21913
rect 17586 21904 17592 21956
rect 17644 21904 17650 21956
rect 18874 21944 18880 21956
rect 18814 21916 18880 21944
rect 18874 21904 18880 21916
rect 18932 21944 18938 21956
rect 19794 21944 19800 21956
rect 18932 21916 19800 21944
rect 18932 21904 18938 21916
rect 19794 21904 19800 21916
rect 19852 21904 19858 21956
rect 20530 21904 20536 21956
rect 20588 21904 20594 21956
rect 23753 21947 23811 21953
rect 22586 21916 22784 21944
rect 22756 21888 22784 21916
rect 23753 21913 23765 21947
rect 23799 21944 23811 21947
rect 24578 21944 24584 21956
rect 23799 21916 24584 21944
rect 23799 21913 23811 21916
rect 23753 21907 23811 21913
rect 24578 21904 24584 21916
rect 24636 21904 24642 21956
rect 25498 21904 25504 21956
rect 25556 21904 25562 21956
rect 26344 21944 26372 22043
rect 26510 21944 26516 21956
rect 26344 21916 26516 21944
rect 26510 21904 26516 21916
rect 26568 21904 26574 21956
rect 28442 21944 28448 21956
rect 27830 21916 28448 21944
rect 28442 21904 28448 21916
rect 28500 21904 28506 21956
rect 12710 21876 12716 21888
rect 11992 21848 12716 21876
rect 12710 21836 12716 21848
rect 12768 21836 12774 21888
rect 13909 21879 13967 21885
rect 13909 21845 13921 21879
rect 13955 21876 13967 21879
rect 15102 21876 15108 21888
rect 13955 21848 15108 21876
rect 13955 21845 13967 21848
rect 13909 21839 13967 21845
rect 15102 21836 15108 21848
rect 15160 21876 15166 21888
rect 16225 21879 16283 21885
rect 16225 21876 16237 21879
rect 15160 21848 16237 21876
rect 15160 21836 15166 21848
rect 16225 21845 16237 21848
rect 16271 21845 16283 21879
rect 16225 21839 16283 21845
rect 19061 21879 19119 21885
rect 19061 21845 19073 21879
rect 19107 21876 19119 21879
rect 19334 21876 19340 21888
rect 19107 21848 19340 21876
rect 19107 21845 19119 21848
rect 19061 21839 19119 21845
rect 19334 21836 19340 21848
rect 19392 21836 19398 21888
rect 20990 21836 20996 21888
rect 21048 21836 21054 21888
rect 22738 21836 22744 21888
rect 22796 21876 22802 21888
rect 23106 21876 23112 21888
rect 22796 21848 23112 21876
rect 22796 21836 22802 21848
rect 23106 21836 23112 21848
rect 23164 21836 23170 21888
rect 23293 21879 23351 21885
rect 23293 21845 23305 21879
rect 23339 21876 23351 21879
rect 23474 21876 23480 21888
rect 23339 21848 23480 21876
rect 23339 21845 23351 21848
rect 23293 21839 23351 21845
rect 23474 21836 23480 21848
rect 23532 21836 23538 21888
rect 23658 21836 23664 21888
rect 23716 21836 23722 21888
rect 24489 21879 24547 21885
rect 24489 21845 24501 21879
rect 24535 21876 24547 21879
rect 25222 21876 25228 21888
rect 24535 21848 25228 21876
rect 24535 21845 24547 21848
rect 24489 21839 24547 21845
rect 25222 21836 25228 21848
rect 25280 21836 25286 21888
rect 27338 21836 27344 21888
rect 27396 21876 27402 21888
rect 28077 21879 28135 21885
rect 28077 21876 28089 21879
rect 27396 21848 28089 21876
rect 27396 21836 27402 21848
rect 28077 21845 28089 21848
rect 28123 21845 28135 21879
rect 28077 21839 28135 21845
rect 1104 21786 28704 21808
rect 1104 21734 4874 21786
rect 4926 21734 4938 21786
rect 4990 21734 5002 21786
rect 5054 21734 5066 21786
rect 5118 21734 5130 21786
rect 5182 21734 28704 21786
rect 1104 21712 28704 21734
rect 4893 21675 4951 21681
rect 4893 21641 4905 21675
rect 4939 21672 4951 21675
rect 5534 21672 5540 21684
rect 4939 21644 5540 21672
rect 4939 21641 4951 21644
rect 4893 21635 4951 21641
rect 5534 21632 5540 21644
rect 5592 21632 5598 21684
rect 6457 21675 6515 21681
rect 6457 21672 6469 21675
rect 5920 21644 6469 21672
rect 4982 21564 4988 21616
rect 5040 21604 5046 21616
rect 5920 21613 5948 21644
rect 6457 21641 6469 21644
rect 6503 21641 6515 21675
rect 6457 21635 6515 21641
rect 7834 21632 7840 21684
rect 7892 21672 7898 21684
rect 14090 21672 14096 21684
rect 7892 21644 14096 21672
rect 7892 21632 7898 21644
rect 14090 21632 14096 21644
rect 14148 21632 14154 21684
rect 16482 21672 16488 21684
rect 14752 21644 16488 21672
rect 5675 21607 5733 21613
rect 5675 21604 5687 21607
rect 5040 21576 5687 21604
rect 5040 21564 5046 21576
rect 5675 21573 5687 21576
rect 5721 21573 5733 21607
rect 5675 21567 5733 21573
rect 5905 21607 5963 21613
rect 5905 21573 5917 21607
rect 5951 21573 5963 21607
rect 9125 21607 9183 21613
rect 9125 21604 9137 21607
rect 5905 21567 5963 21573
rect 6012 21576 9137 21604
rect 4062 21496 4068 21548
rect 4120 21536 4126 21548
rect 4433 21539 4491 21545
rect 4433 21536 4445 21539
rect 4120 21508 4445 21536
rect 4120 21496 4126 21508
rect 4433 21505 4445 21508
rect 4479 21505 4491 21539
rect 4433 21499 4491 21505
rect 4341 21471 4399 21477
rect 4341 21437 4353 21471
rect 4387 21437 4399 21471
rect 4448 21468 4476 21499
rect 5074 21496 5080 21548
rect 5132 21496 5138 21548
rect 5169 21539 5227 21545
rect 5169 21505 5181 21539
rect 5215 21505 5227 21539
rect 5169 21499 5227 21505
rect 5261 21539 5319 21545
rect 5261 21505 5273 21539
rect 5307 21536 5319 21539
rect 5350 21536 5356 21548
rect 5307 21508 5356 21536
rect 5307 21505 5319 21508
rect 5261 21499 5319 21505
rect 5184 21468 5212 21499
rect 5350 21496 5356 21508
rect 5408 21496 5414 21548
rect 5445 21539 5503 21545
rect 5445 21505 5457 21539
rect 5491 21536 5503 21539
rect 5491 21508 5672 21536
rect 5491 21505 5503 21508
rect 5445 21499 5503 21505
rect 5537 21471 5595 21477
rect 5537 21468 5549 21471
rect 4448 21440 5549 21468
rect 4341 21431 4399 21437
rect 5537 21437 5549 21440
rect 5583 21437 5595 21471
rect 5644 21468 5672 21508
rect 5810 21496 5816 21548
rect 5868 21496 5874 21548
rect 6012 21545 6040 21576
rect 9125 21573 9137 21576
rect 9171 21573 9183 21607
rect 11698 21604 11704 21616
rect 11086 21576 11704 21604
rect 9125 21567 9183 21573
rect 11698 21564 11704 21576
rect 11756 21564 11762 21616
rect 11790 21564 11796 21616
rect 11848 21564 11854 21616
rect 5997 21539 6055 21545
rect 5997 21505 6009 21539
rect 6043 21505 6055 21539
rect 5997 21499 6055 21505
rect 6086 21496 6092 21548
rect 6144 21536 6150 21548
rect 6825 21539 6883 21545
rect 6825 21536 6837 21539
rect 6144 21508 6837 21536
rect 6144 21496 6150 21508
rect 6825 21505 6837 21508
rect 6871 21536 6883 21539
rect 6914 21536 6920 21548
rect 6871 21508 6920 21536
rect 6871 21505 6883 21508
rect 6825 21499 6883 21505
rect 6914 21496 6920 21508
rect 6972 21496 6978 21548
rect 7558 21496 7564 21548
rect 7616 21536 7622 21548
rect 8849 21539 8907 21545
rect 8849 21536 8861 21539
rect 7616 21508 8861 21536
rect 7616 21496 7622 21508
rect 8849 21505 8861 21508
rect 8895 21536 8907 21539
rect 9214 21536 9220 21548
rect 8895 21508 9220 21536
rect 8895 21505 8907 21508
rect 8849 21499 8907 21505
rect 9214 21496 9220 21508
rect 9272 21496 9278 21548
rect 9401 21539 9459 21545
rect 9401 21505 9413 21539
rect 9447 21505 9459 21539
rect 9401 21499 9459 21505
rect 5718 21468 5724 21480
rect 5644 21440 5724 21468
rect 5537 21431 5595 21437
rect 4356 21332 4384 21431
rect 4801 21403 4859 21409
rect 4801 21369 4813 21403
rect 4847 21400 4859 21403
rect 5350 21400 5356 21412
rect 4847 21372 5356 21400
rect 4847 21369 4859 21372
rect 4801 21363 4859 21369
rect 5350 21360 5356 21372
rect 5408 21360 5414 21412
rect 5552 21400 5580 21431
rect 5718 21428 5724 21440
rect 5776 21428 5782 21480
rect 6733 21471 6791 21477
rect 5828 21440 6224 21468
rect 5828 21400 5856 21440
rect 5552 21372 5856 21400
rect 6196 21400 6224 21440
rect 6733 21437 6745 21471
rect 6779 21468 6791 21471
rect 8662 21468 8668 21480
rect 6779 21440 8668 21468
rect 6779 21437 6791 21440
rect 6733 21431 6791 21437
rect 8662 21428 8668 21440
rect 8720 21468 8726 21480
rect 9125 21471 9183 21477
rect 9125 21468 9137 21471
rect 8720 21440 9137 21468
rect 8720 21428 8726 21440
rect 9125 21437 9137 21440
rect 9171 21437 9183 21471
rect 9125 21431 9183 21437
rect 7190 21400 7196 21412
rect 6196 21372 7196 21400
rect 6086 21332 6092 21344
rect 4356 21304 6092 21332
rect 6086 21292 6092 21304
rect 6144 21292 6150 21344
rect 6178 21292 6184 21344
rect 6236 21292 6242 21344
rect 6840 21341 6868 21372
rect 7190 21360 7196 21372
rect 7248 21400 7254 21412
rect 9416 21400 9444 21499
rect 9582 21496 9588 21548
rect 9640 21496 9646 21548
rect 12894 21496 12900 21548
rect 12952 21496 12958 21548
rect 13262 21496 13268 21548
rect 13320 21536 13326 21548
rect 13449 21539 13507 21545
rect 13449 21536 13461 21539
rect 13320 21508 13461 21536
rect 13320 21496 13326 21508
rect 13449 21505 13461 21508
rect 13495 21536 13507 21539
rect 14277 21539 14335 21545
rect 13495 21508 13584 21536
rect 13495 21505 13507 21508
rect 13449 21499 13507 21505
rect 9858 21428 9864 21480
rect 9916 21428 9922 21480
rect 11517 21471 11575 21477
rect 11517 21437 11529 21471
rect 11563 21468 11575 21471
rect 13556 21468 13584 21508
rect 14277 21505 14289 21539
rect 14323 21536 14335 21539
rect 14752 21536 14780 21644
rect 16482 21632 16488 21644
rect 16540 21632 16546 21684
rect 20073 21675 20131 21681
rect 20073 21641 20085 21675
rect 20119 21672 20131 21675
rect 20346 21672 20352 21684
rect 20119 21644 20352 21672
rect 20119 21641 20131 21644
rect 20073 21635 20131 21641
rect 20346 21632 20352 21644
rect 20404 21632 20410 21684
rect 20533 21675 20591 21681
rect 20533 21641 20545 21675
rect 20579 21672 20591 21675
rect 20990 21672 20996 21684
rect 20579 21644 20996 21672
rect 20579 21641 20591 21644
rect 20533 21635 20591 21641
rect 20990 21632 20996 21644
rect 21048 21632 21054 21684
rect 21821 21675 21879 21681
rect 21821 21641 21833 21675
rect 21867 21672 21879 21675
rect 22370 21672 22376 21684
rect 21867 21644 22376 21672
rect 21867 21641 21879 21644
rect 21821 21635 21879 21641
rect 22370 21632 22376 21644
rect 22428 21632 22434 21684
rect 24026 21672 24032 21684
rect 22756 21644 24032 21672
rect 16298 21604 16304 21616
rect 16238 21576 16304 21604
rect 16298 21564 16304 21576
rect 16356 21604 16362 21616
rect 18874 21604 18880 21616
rect 16356 21576 18880 21604
rect 16356 21564 16362 21576
rect 18874 21564 18880 21576
rect 18932 21564 18938 21616
rect 19242 21564 19248 21616
rect 19300 21604 19306 21616
rect 19797 21607 19855 21613
rect 19797 21604 19809 21607
rect 19300 21576 19809 21604
rect 19300 21564 19306 21576
rect 19797 21573 19809 21576
rect 19843 21573 19855 21607
rect 19797 21567 19855 21573
rect 22281 21607 22339 21613
rect 22281 21573 22293 21607
rect 22327 21604 22339 21607
rect 22646 21604 22652 21616
rect 22327 21576 22652 21604
rect 22327 21573 22339 21576
rect 22281 21567 22339 21573
rect 22646 21564 22652 21576
rect 22704 21564 22710 21616
rect 14323 21508 14780 21536
rect 19061 21539 19119 21545
rect 14323 21505 14335 21508
rect 14277 21499 14335 21505
rect 19061 21505 19073 21539
rect 19107 21536 19119 21539
rect 19334 21536 19340 21548
rect 19107 21508 19340 21536
rect 19107 21505 19119 21508
rect 19061 21499 19119 21505
rect 19334 21496 19340 21508
rect 19392 21496 19398 21548
rect 20441 21539 20499 21545
rect 20441 21505 20453 21539
rect 20487 21536 20499 21539
rect 20901 21539 20959 21545
rect 20901 21536 20913 21539
rect 20487 21508 20913 21536
rect 20487 21505 20499 21508
rect 20441 21499 20499 21505
rect 20901 21505 20913 21508
rect 20947 21505 20959 21539
rect 20901 21499 20959 21505
rect 22186 21496 22192 21548
rect 22244 21496 22250 21548
rect 22756 21480 22784 21644
rect 24026 21632 24032 21644
rect 24084 21632 24090 21684
rect 24489 21675 24547 21681
rect 24489 21641 24501 21675
rect 24535 21672 24547 21675
rect 24578 21672 24584 21684
rect 24535 21644 24584 21672
rect 24535 21641 24547 21644
rect 24489 21635 24547 21641
rect 24578 21632 24584 21644
rect 24636 21632 24642 21684
rect 25498 21672 25504 21684
rect 24688 21644 25504 21672
rect 23014 21564 23020 21616
rect 23072 21564 23078 21616
rect 24688 21604 24716 21644
rect 25498 21632 25504 21644
rect 25556 21632 25562 21684
rect 25590 21632 25596 21684
rect 25648 21672 25654 21684
rect 25685 21675 25743 21681
rect 25685 21672 25697 21675
rect 25648 21644 25697 21672
rect 25648 21632 25654 21644
rect 25685 21641 25697 21644
rect 25731 21641 25743 21675
rect 25685 21635 25743 21641
rect 26418 21632 26424 21684
rect 26476 21672 26482 21684
rect 26476 21644 27292 21672
rect 26476 21632 26482 21644
rect 24242 21576 24716 21604
rect 25038 21564 25044 21616
rect 25096 21604 25102 21616
rect 27264 21604 27292 21644
rect 27338 21604 27344 21616
rect 25096 21576 27108 21604
rect 27264 21576 27344 21604
rect 25096 21564 25102 21576
rect 25317 21539 25375 21545
rect 25317 21505 25329 21539
rect 25363 21536 25375 21539
rect 25777 21539 25835 21545
rect 25777 21536 25789 21539
rect 25363 21508 25789 21536
rect 25363 21505 25375 21508
rect 25317 21499 25375 21505
rect 25777 21505 25789 21508
rect 25823 21505 25835 21539
rect 25777 21499 25835 21505
rect 26602 21496 26608 21548
rect 26660 21536 26666 21548
rect 27080 21545 27108 21576
rect 27338 21564 27344 21576
rect 27396 21564 27402 21616
rect 26973 21539 27031 21545
rect 26973 21536 26985 21539
rect 26660 21508 26985 21536
rect 26660 21496 26666 21508
rect 26973 21505 26985 21508
rect 27019 21505 27031 21539
rect 26973 21499 27031 21505
rect 27066 21539 27124 21545
rect 27066 21505 27078 21539
rect 27112 21505 27124 21539
rect 27066 21499 27124 21505
rect 27249 21539 27307 21545
rect 27249 21505 27261 21539
rect 27295 21505 27307 21539
rect 27249 21499 27307 21505
rect 11563 21440 13584 21468
rect 11563 21437 11575 21440
rect 11517 21431 11575 21437
rect 7248 21372 9444 21400
rect 7248 21360 7254 21372
rect 10962 21360 10968 21412
rect 11020 21400 11026 21412
rect 11333 21403 11391 21409
rect 11333 21400 11345 21403
rect 11020 21372 11345 21400
rect 11020 21360 11026 21372
rect 11333 21369 11345 21372
rect 11379 21369 11391 21403
rect 11333 21363 11391 21369
rect 6825 21335 6883 21341
rect 6825 21301 6837 21335
rect 6871 21301 6883 21335
rect 6825 21295 6883 21301
rect 6914 21292 6920 21344
rect 6972 21332 6978 21344
rect 9309 21335 9367 21341
rect 9309 21332 9321 21335
rect 6972 21304 9321 21332
rect 6972 21292 6978 21304
rect 9309 21301 9321 21304
rect 9355 21301 9367 21335
rect 11348 21332 11376 21363
rect 13078 21360 13084 21412
rect 13136 21400 13142 21412
rect 13265 21403 13323 21409
rect 13265 21400 13277 21403
rect 13136 21372 13277 21400
rect 13136 21360 13142 21372
rect 13265 21369 13277 21372
rect 13311 21369 13323 21403
rect 13556 21400 13584 21440
rect 14366 21428 14372 21480
rect 14424 21428 14430 21480
rect 14737 21471 14795 21477
rect 14737 21437 14749 21471
rect 14783 21437 14795 21471
rect 14737 21431 14795 21437
rect 15013 21471 15071 21477
rect 15013 21437 15025 21471
rect 15059 21468 15071 21471
rect 15470 21468 15476 21480
rect 15059 21440 15476 21468
rect 15059 21437 15071 21440
rect 15013 21431 15071 21437
rect 14752 21400 14780 21431
rect 15470 21428 15476 21440
rect 15528 21428 15534 21480
rect 19610 21428 19616 21480
rect 19668 21468 19674 21480
rect 20625 21471 20683 21477
rect 20625 21468 20637 21471
rect 19668 21440 20637 21468
rect 19668 21428 19674 21440
rect 20625 21437 20637 21440
rect 20671 21437 20683 21471
rect 20625 21431 20683 21437
rect 13556 21372 14780 21400
rect 20640 21400 20668 21431
rect 21450 21428 21456 21480
rect 21508 21428 21514 21480
rect 22465 21471 22523 21477
rect 22465 21437 22477 21471
rect 22511 21437 22523 21471
rect 22465 21431 22523 21437
rect 22480 21400 22508 21431
rect 22738 21428 22744 21480
rect 22796 21428 22802 21480
rect 24210 21468 24216 21480
rect 22848 21440 24216 21468
rect 22848 21400 22876 21440
rect 24210 21428 24216 21440
rect 24268 21468 24274 21480
rect 25133 21471 25191 21477
rect 25133 21468 25145 21471
rect 24268 21440 25145 21468
rect 24268 21428 24274 21440
rect 25133 21437 25145 21440
rect 25179 21437 25191 21471
rect 25133 21431 25191 21437
rect 20640 21372 22876 21400
rect 13265 21363 13323 21369
rect 12894 21332 12900 21344
rect 11348 21304 12900 21332
rect 9309 21295 9367 21301
rect 12894 21292 12900 21304
rect 12952 21292 12958 21344
rect 14645 21335 14703 21341
rect 14645 21301 14657 21335
rect 14691 21332 14703 21335
rect 14826 21332 14832 21344
rect 14691 21304 14832 21332
rect 14691 21301 14703 21304
rect 14645 21295 14703 21301
rect 14826 21292 14832 21304
rect 14884 21292 14890 21344
rect 25148 21332 25176 21431
rect 25222 21428 25228 21480
rect 25280 21428 25286 21480
rect 26326 21428 26332 21480
rect 26384 21428 26390 21480
rect 27264 21468 27292 21499
rect 27430 21496 27436 21548
rect 27488 21545 27494 21548
rect 27488 21536 27496 21545
rect 27488 21508 27533 21536
rect 27488 21499 27496 21508
rect 27488 21496 27494 21499
rect 26436 21440 27292 21468
rect 25240 21400 25268 21428
rect 26436 21400 26464 21440
rect 28258 21428 28264 21480
rect 28316 21428 28322 21480
rect 25240 21372 26464 21400
rect 26786 21360 26792 21412
rect 26844 21400 26850 21412
rect 27709 21403 27767 21409
rect 27709 21400 27721 21403
rect 26844 21372 27721 21400
rect 26844 21360 26850 21372
rect 27709 21369 27721 21372
rect 27755 21369 27767 21403
rect 27709 21363 27767 21369
rect 27154 21332 27160 21344
rect 25148 21304 27160 21332
rect 27154 21292 27160 21304
rect 27212 21292 27218 21344
rect 27617 21335 27675 21341
rect 27617 21301 27629 21335
rect 27663 21332 27675 21335
rect 28166 21332 28172 21344
rect 27663 21304 28172 21332
rect 27663 21301 27675 21304
rect 27617 21295 27675 21301
rect 28166 21292 28172 21304
rect 28224 21292 28230 21344
rect 1104 21242 28704 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 28704 21242
rect 1104 21168 28704 21190
rect 4985 21131 5043 21137
rect 4985 21097 4997 21131
rect 5031 21128 5043 21131
rect 5718 21128 5724 21140
rect 5031 21100 5724 21128
rect 5031 21097 5043 21100
rect 4985 21091 5043 21097
rect 5718 21088 5724 21100
rect 5776 21088 5782 21140
rect 6270 21088 6276 21140
rect 6328 21128 6334 21140
rect 6733 21131 6791 21137
rect 6733 21128 6745 21131
rect 6328 21100 6745 21128
rect 6328 21088 6334 21100
rect 6733 21097 6745 21100
rect 6779 21097 6791 21131
rect 6733 21091 6791 21097
rect 11422 21088 11428 21140
rect 11480 21128 11486 21140
rect 12069 21131 12127 21137
rect 12069 21128 12081 21131
rect 11480 21100 12081 21128
rect 11480 21088 11486 21100
rect 12069 21097 12081 21100
rect 12115 21097 12127 21131
rect 12069 21091 12127 21097
rect 12161 21131 12219 21137
rect 12161 21097 12173 21131
rect 12207 21128 12219 21131
rect 12434 21128 12440 21140
rect 12207 21100 12440 21128
rect 12207 21097 12219 21100
rect 12161 21091 12219 21097
rect 8956 21032 9720 21060
rect 5074 20952 5080 21004
rect 5132 20992 5138 21004
rect 5132 20964 5948 20992
rect 5132 20952 5138 20964
rect 5166 20884 5172 20936
rect 5224 20884 5230 20936
rect 5350 20884 5356 20936
rect 5408 20884 5414 20936
rect 5534 20884 5540 20936
rect 5592 20924 5598 20936
rect 5810 20924 5816 20936
rect 5592 20896 5816 20924
rect 5592 20884 5598 20896
rect 5810 20884 5816 20896
rect 5868 20884 5874 20936
rect 5920 20868 5948 20964
rect 6178 20884 6184 20936
rect 6236 20884 6242 20936
rect 6549 20927 6607 20933
rect 6549 20924 6561 20927
rect 6288 20896 6561 20924
rect 4706 20816 4712 20868
rect 4764 20856 4770 20868
rect 4982 20856 4988 20868
rect 4764 20828 4988 20856
rect 4764 20816 4770 20828
rect 4982 20816 4988 20828
rect 5040 20856 5046 20868
rect 5261 20859 5319 20865
rect 5261 20856 5273 20859
rect 5040 20828 5273 20856
rect 5040 20816 5046 20828
rect 5261 20825 5273 20828
rect 5307 20825 5319 20859
rect 5261 20819 5319 20825
rect 5902 20816 5908 20868
rect 5960 20856 5966 20868
rect 6288 20856 6316 20896
rect 6549 20893 6561 20896
rect 6595 20893 6607 20927
rect 6549 20887 6607 20893
rect 6917 20927 6975 20933
rect 6917 20893 6929 20927
rect 6963 20924 6975 20927
rect 7834 20924 7840 20936
rect 6963 20896 7840 20924
rect 6963 20893 6975 20896
rect 6917 20887 6975 20893
rect 7834 20884 7840 20896
rect 7892 20884 7898 20936
rect 8386 20884 8392 20936
rect 8444 20924 8450 20936
rect 8956 20933 8984 21032
rect 9214 20952 9220 21004
rect 9272 20992 9278 21004
rect 9585 20995 9643 21001
rect 9585 20992 9597 20995
rect 9272 20964 9597 20992
rect 9272 20952 9278 20964
rect 9585 20961 9597 20964
rect 9631 20961 9643 20995
rect 9692 20992 9720 21032
rect 11333 20995 11391 21001
rect 9692 20964 11192 20992
rect 9585 20955 9643 20961
rect 11164 20936 11192 20964
rect 11333 20961 11345 20995
rect 11379 20992 11391 20995
rect 11425 20995 11483 21001
rect 11425 20992 11437 20995
rect 11379 20964 11437 20992
rect 11379 20961 11391 20964
rect 11333 20955 11391 20961
rect 11425 20961 11437 20964
rect 11471 20961 11483 20995
rect 12084 20992 12112 21091
rect 12434 21088 12440 21100
rect 12492 21088 12498 21140
rect 15470 21088 15476 21140
rect 15528 21088 15534 21140
rect 17494 21088 17500 21140
rect 17552 21088 17558 21140
rect 23658 21088 23664 21140
rect 23716 21128 23722 21140
rect 24213 21131 24271 21137
rect 24213 21128 24225 21131
rect 23716 21100 24225 21128
rect 23716 21088 23722 21100
rect 24213 21097 24225 21100
rect 24259 21097 24271 21131
rect 24213 21091 24271 21097
rect 12084 20964 12572 20992
rect 11425 20955 11483 20961
rect 8665 20927 8723 20933
rect 8665 20924 8677 20927
rect 8444 20896 8677 20924
rect 8444 20884 8450 20896
rect 8665 20893 8677 20896
rect 8711 20893 8723 20927
rect 8665 20887 8723 20893
rect 8941 20927 8999 20933
rect 8941 20893 8953 20927
rect 8987 20893 8999 20927
rect 8941 20887 8999 20893
rect 5960 20828 6316 20856
rect 5960 20816 5966 20828
rect 6362 20816 6368 20868
rect 6420 20816 6426 20868
rect 6457 20859 6515 20865
rect 6457 20825 6469 20859
rect 6503 20856 6515 20859
rect 7006 20856 7012 20868
rect 6503 20828 7012 20856
rect 6503 20825 6515 20828
rect 6457 20819 6515 20825
rect 7006 20816 7012 20828
rect 7064 20816 7070 20868
rect 7558 20816 7564 20868
rect 7616 20856 7622 20868
rect 7653 20859 7711 20865
rect 7653 20856 7665 20859
rect 7616 20828 7665 20856
rect 7616 20816 7622 20828
rect 7653 20825 7665 20828
rect 7699 20825 7711 20859
rect 7653 20819 7711 20825
rect 8113 20791 8171 20797
rect 8113 20757 8125 20791
rect 8159 20788 8171 20791
rect 8202 20788 8208 20800
rect 8159 20760 8208 20788
rect 8159 20757 8171 20760
rect 8113 20751 8171 20757
rect 8202 20748 8208 20760
rect 8260 20748 8266 20800
rect 8680 20788 8708 20887
rect 9122 20884 9128 20936
rect 9180 20884 9186 20936
rect 9306 20884 9312 20936
rect 9364 20884 9370 20936
rect 11146 20884 11152 20936
rect 11204 20924 11210 20936
rect 11882 20924 11888 20936
rect 11204 20896 11888 20924
rect 11204 20884 11210 20896
rect 11882 20884 11888 20896
rect 11940 20924 11946 20936
rect 12544 20933 12572 20964
rect 14826 20952 14832 21004
rect 14884 20952 14890 21004
rect 19242 20952 19248 21004
rect 19300 20992 19306 21004
rect 19889 20995 19947 21001
rect 19889 20992 19901 20995
rect 19300 20964 19901 20992
rect 19300 20952 19306 20964
rect 12345 20927 12403 20933
rect 12345 20924 12357 20927
rect 11940 20896 12357 20924
rect 11940 20884 11946 20896
rect 12345 20893 12357 20896
rect 12391 20893 12403 20927
rect 12345 20887 12403 20893
rect 12529 20927 12587 20933
rect 12529 20893 12541 20927
rect 12575 20893 12587 20927
rect 12529 20887 12587 20893
rect 12621 20927 12679 20933
rect 12621 20893 12633 20927
rect 12667 20893 12679 20927
rect 12621 20887 12679 20893
rect 9217 20859 9275 20865
rect 9217 20825 9229 20859
rect 9263 20856 9275 20859
rect 9861 20859 9919 20865
rect 9861 20856 9873 20859
rect 9263 20828 9873 20856
rect 9263 20825 9275 20828
rect 9217 20819 9275 20825
rect 9861 20825 9873 20828
rect 9907 20856 9919 20859
rect 9950 20856 9956 20868
rect 9907 20828 9956 20856
rect 9907 20825 9919 20828
rect 9861 20819 9919 20825
rect 9950 20816 9956 20828
rect 10008 20816 10014 20868
rect 12636 20856 12664 20887
rect 12710 20884 12716 20936
rect 12768 20884 12774 20936
rect 12894 20884 12900 20936
rect 12952 20884 12958 20936
rect 15194 20884 15200 20936
rect 15252 20924 15258 20936
rect 15565 20927 15623 20933
rect 15565 20924 15577 20927
rect 15252 20896 15577 20924
rect 15252 20884 15258 20896
rect 15565 20893 15577 20896
rect 15611 20893 15623 20927
rect 15565 20887 15623 20893
rect 15838 20884 15844 20936
rect 15896 20884 15902 20936
rect 17681 20927 17739 20933
rect 17681 20893 17693 20927
rect 17727 20893 17739 20927
rect 17681 20887 17739 20893
rect 12805 20859 12863 20865
rect 12805 20856 12817 20859
rect 11086 20828 12434 20856
rect 12636 20828 12817 20856
rect 9306 20788 9312 20800
rect 8680 20760 9312 20788
rect 9306 20748 9312 20760
rect 9364 20748 9370 20800
rect 9493 20791 9551 20797
rect 9493 20757 9505 20791
rect 9539 20788 9551 20791
rect 9766 20788 9772 20800
rect 9539 20760 9772 20788
rect 9539 20757 9551 20760
rect 9493 20751 9551 20757
rect 9766 20748 9772 20760
rect 9824 20748 9830 20800
rect 12406 20788 12434 20828
rect 12805 20825 12817 20828
rect 12851 20825 12863 20859
rect 12805 20819 12863 20825
rect 14366 20816 14372 20868
rect 14424 20856 14430 20868
rect 15657 20859 15715 20865
rect 15657 20856 15669 20859
rect 14424 20828 15669 20856
rect 14424 20816 14430 20828
rect 15657 20825 15669 20828
rect 15703 20825 15715 20859
rect 17696 20856 17724 20887
rect 17954 20884 17960 20936
rect 18012 20884 18018 20936
rect 19352 20933 19380 20964
rect 19889 20961 19901 20964
rect 19935 20961 19947 20995
rect 19889 20955 19947 20961
rect 21729 20995 21787 21001
rect 21729 20961 21741 20995
rect 21775 20992 21787 20995
rect 22738 20992 22744 21004
rect 21775 20964 22744 20992
rect 21775 20961 21787 20964
rect 21729 20955 21787 20961
rect 22738 20952 22744 20964
rect 22796 20952 22802 21004
rect 23477 20995 23535 21001
rect 23477 20961 23489 20995
rect 23523 20992 23535 20995
rect 23569 20995 23627 21001
rect 23569 20992 23581 20995
rect 23523 20964 23581 20992
rect 23523 20961 23535 20964
rect 23477 20955 23535 20961
rect 23569 20961 23581 20964
rect 23615 20961 23627 20995
rect 23569 20955 23627 20961
rect 24026 20952 24032 21004
rect 24084 20992 24090 21004
rect 24762 20992 24768 21004
rect 24084 20964 24768 20992
rect 24084 20952 24090 20964
rect 24762 20952 24768 20964
rect 24820 20992 24826 21004
rect 25133 20995 25191 21001
rect 25133 20992 25145 20995
rect 24820 20964 25145 20992
rect 24820 20952 24826 20964
rect 25133 20961 25145 20964
rect 25179 20992 25191 20995
rect 26513 20995 26571 21001
rect 26513 20992 26525 20995
rect 25179 20964 26525 20992
rect 25179 20961 25191 20964
rect 25133 20955 25191 20961
rect 26513 20961 26525 20964
rect 26559 20961 26571 20995
rect 26513 20955 26571 20961
rect 26786 20952 26792 21004
rect 26844 20952 26850 21004
rect 19337 20927 19395 20933
rect 19337 20893 19349 20927
rect 19383 20924 19395 20927
rect 19383 20896 19417 20924
rect 19383 20893 19395 20896
rect 19337 20887 19395 20893
rect 23106 20884 23112 20936
rect 23164 20924 23170 20936
rect 25498 20924 25504 20936
rect 23164 20896 25504 20924
rect 23164 20884 23170 20896
rect 25498 20884 25504 20896
rect 25556 20884 25562 20936
rect 18414 20856 18420 20868
rect 17696 20828 18420 20856
rect 15657 20819 15715 20825
rect 18414 20816 18420 20828
rect 18472 20816 18478 20868
rect 20162 20816 20168 20868
rect 20220 20816 20226 20868
rect 20622 20816 20628 20868
rect 20680 20816 20686 20868
rect 22005 20859 22063 20865
rect 22005 20825 22017 20859
rect 22051 20856 22063 20859
rect 22278 20856 22284 20868
rect 22051 20828 22284 20856
rect 22051 20825 22063 20828
rect 22005 20819 22063 20825
rect 22278 20816 22284 20828
rect 22336 20816 22342 20868
rect 24394 20816 24400 20868
rect 24452 20816 24458 20868
rect 26786 20816 26792 20868
rect 26844 20856 26850 20868
rect 26844 20828 27278 20856
rect 26844 20816 26850 20828
rect 12710 20788 12716 20800
rect 12406 20760 12716 20788
rect 12710 20748 12716 20760
rect 12768 20788 12774 20800
rect 12986 20788 12992 20800
rect 12768 20760 12992 20788
rect 12768 20748 12774 20760
rect 12986 20748 12992 20760
rect 13044 20748 13050 20800
rect 15930 20748 15936 20800
rect 15988 20788 15994 20800
rect 16025 20791 16083 20797
rect 16025 20788 16037 20791
rect 15988 20760 16037 20788
rect 15988 20748 15994 20760
rect 16025 20757 16037 20760
rect 16071 20757 16083 20791
rect 16025 20751 16083 20757
rect 17402 20748 17408 20800
rect 17460 20788 17466 20800
rect 17865 20791 17923 20797
rect 17865 20788 17877 20791
rect 17460 20760 17877 20788
rect 17460 20748 17466 20760
rect 17865 20757 17877 20760
rect 17911 20757 17923 20791
rect 17865 20751 17923 20757
rect 21634 20748 21640 20800
rect 21692 20748 21698 20800
rect 27798 20748 27804 20800
rect 27856 20788 27862 20800
rect 28261 20791 28319 20797
rect 28261 20788 28273 20791
rect 27856 20760 28273 20788
rect 27856 20748 27862 20760
rect 28261 20757 28273 20760
rect 28307 20757 28319 20791
rect 28261 20751 28319 20757
rect 1104 20698 28704 20720
rect 1104 20646 4874 20698
rect 4926 20646 4938 20698
rect 4990 20646 5002 20698
rect 5054 20646 5066 20698
rect 5118 20646 5130 20698
rect 5182 20646 28704 20698
rect 1104 20624 28704 20646
rect 4798 20544 4804 20596
rect 4856 20584 4862 20596
rect 5902 20584 5908 20596
rect 4856 20556 5212 20584
rect 4856 20544 4862 20556
rect 5184 20516 5212 20556
rect 5736 20556 5908 20584
rect 5442 20516 5448 20528
rect 5106 20488 5448 20516
rect 5442 20476 5448 20488
rect 5500 20476 5506 20528
rect 5736 20516 5764 20556
rect 5902 20544 5908 20556
rect 5960 20544 5966 20596
rect 7469 20587 7527 20593
rect 7469 20553 7481 20587
rect 7515 20584 7527 20587
rect 8110 20584 8116 20596
rect 7515 20556 8116 20584
rect 7515 20553 7527 20556
rect 7469 20547 7527 20553
rect 8110 20544 8116 20556
rect 8168 20544 8174 20596
rect 9398 20544 9404 20596
rect 9456 20584 9462 20596
rect 9585 20587 9643 20593
rect 9585 20584 9597 20587
rect 9456 20556 9597 20584
rect 9456 20544 9462 20556
rect 9585 20553 9597 20556
rect 9631 20553 9643 20587
rect 9585 20547 9643 20553
rect 9858 20544 9864 20596
rect 9916 20584 9922 20596
rect 10321 20587 10379 20593
rect 10321 20584 10333 20587
rect 9916 20556 10333 20584
rect 9916 20544 9922 20556
rect 10321 20553 10333 20556
rect 10367 20553 10379 20587
rect 14090 20584 14096 20596
rect 10321 20547 10379 20553
rect 13464 20556 14096 20584
rect 5644 20488 5764 20516
rect 5644 20457 5672 20488
rect 5810 20476 5816 20528
rect 5868 20516 5874 20528
rect 6362 20516 6368 20528
rect 5868 20488 6368 20516
rect 5868 20476 5874 20488
rect 6362 20476 6368 20488
rect 6420 20516 6426 20528
rect 6420 20488 6868 20516
rect 6420 20476 6426 20488
rect 5629 20451 5687 20457
rect 5629 20417 5641 20451
rect 5675 20417 5687 20451
rect 5629 20411 5687 20417
rect 5718 20408 5724 20460
rect 5776 20408 5782 20460
rect 5997 20451 6055 20457
rect 5997 20417 6009 20451
rect 6043 20417 6055 20451
rect 6840 20448 6868 20488
rect 6914 20476 6920 20528
rect 6972 20516 6978 20528
rect 7009 20519 7067 20525
rect 7009 20516 7021 20519
rect 6972 20488 7021 20516
rect 6972 20476 6978 20488
rect 7009 20485 7021 20488
rect 7055 20485 7067 20519
rect 8386 20516 8392 20528
rect 7009 20479 7067 20485
rect 7300 20488 8392 20516
rect 7300 20460 7328 20488
rect 8386 20476 8392 20488
rect 8444 20476 8450 20528
rect 8570 20476 8576 20528
rect 8628 20476 8634 20528
rect 10045 20519 10103 20525
rect 10045 20485 10057 20519
rect 10091 20516 10103 20519
rect 10962 20516 10968 20528
rect 10091 20488 10968 20516
rect 10091 20485 10103 20488
rect 10045 20479 10103 20485
rect 10962 20476 10968 20488
rect 11020 20476 11026 20528
rect 13464 20525 13492 20556
rect 14090 20544 14096 20556
rect 14148 20584 14154 20596
rect 16390 20584 16396 20596
rect 14148 20556 16396 20584
rect 14148 20544 14154 20556
rect 16390 20544 16396 20556
rect 16448 20544 16454 20596
rect 19242 20584 19248 20596
rect 18156 20556 19248 20584
rect 13449 20519 13507 20525
rect 13449 20485 13461 20519
rect 13495 20485 13507 20519
rect 16298 20516 16304 20528
rect 16146 20488 16304 20516
rect 13449 20479 13507 20485
rect 16298 20476 16304 20488
rect 16356 20476 16362 20528
rect 6840 20420 7144 20448
rect 5997 20411 6055 20417
rect 3602 20340 3608 20392
rect 3660 20340 3666 20392
rect 3881 20383 3939 20389
rect 3881 20349 3893 20383
rect 3927 20380 3939 20383
rect 3927 20352 5488 20380
rect 3927 20349 3939 20352
rect 3881 20343 3939 20349
rect 5460 20321 5488 20352
rect 5534 20340 5540 20392
rect 5592 20380 5598 20392
rect 6012 20380 6040 20411
rect 5592 20352 6040 20380
rect 5592 20340 5598 20352
rect 5445 20315 5503 20321
rect 5445 20281 5457 20315
rect 5491 20281 5503 20315
rect 5445 20275 5503 20281
rect 5258 20204 5264 20256
rect 5316 20244 5322 20256
rect 5353 20247 5411 20253
rect 5353 20244 5365 20247
rect 5316 20216 5365 20244
rect 5316 20204 5322 20216
rect 5353 20213 5365 20216
rect 5399 20244 5411 20247
rect 5626 20244 5632 20256
rect 5399 20216 5632 20244
rect 5399 20213 5411 20216
rect 5353 20207 5411 20213
rect 5626 20204 5632 20216
rect 5684 20204 5690 20256
rect 7006 20204 7012 20256
rect 7064 20204 7070 20256
rect 7116 20244 7144 20420
rect 7190 20408 7196 20460
rect 7248 20408 7254 20460
rect 7282 20408 7288 20460
rect 7340 20408 7346 20460
rect 9766 20408 9772 20460
rect 9824 20408 9830 20460
rect 9953 20451 10011 20457
rect 9953 20417 9965 20451
rect 9999 20417 10011 20451
rect 9953 20411 10011 20417
rect 10137 20451 10195 20457
rect 10137 20417 10149 20451
rect 10183 20448 10195 20451
rect 10686 20448 10692 20460
rect 10183 20420 10692 20448
rect 10183 20417 10195 20420
rect 10137 20411 10195 20417
rect 7558 20340 7564 20392
rect 7616 20380 7622 20392
rect 7837 20383 7895 20389
rect 7837 20380 7849 20383
rect 7616 20352 7849 20380
rect 7616 20340 7622 20352
rect 7837 20349 7849 20352
rect 7883 20349 7895 20383
rect 7837 20343 7895 20349
rect 8110 20340 8116 20392
rect 8168 20340 8174 20392
rect 8570 20340 8576 20392
rect 8628 20380 8634 20392
rect 9582 20380 9588 20392
rect 8628 20352 9588 20380
rect 8628 20340 8634 20352
rect 9582 20340 9588 20352
rect 9640 20340 9646 20392
rect 8294 20244 8300 20256
rect 7116 20216 8300 20244
rect 8294 20204 8300 20216
rect 8352 20244 8358 20256
rect 9582 20244 9588 20256
rect 8352 20216 9588 20244
rect 8352 20204 8358 20216
rect 9582 20204 9588 20216
rect 9640 20244 9646 20256
rect 9968 20244 9996 20411
rect 10686 20408 10692 20420
rect 10744 20408 10750 20460
rect 12345 20451 12403 20457
rect 12345 20417 12357 20451
rect 12391 20417 12403 20451
rect 12345 20411 12403 20417
rect 13357 20451 13415 20457
rect 13357 20417 13369 20451
rect 13403 20417 13415 20451
rect 13357 20411 13415 20417
rect 11606 20272 11612 20324
rect 11664 20312 11670 20324
rect 12161 20315 12219 20321
rect 12161 20312 12173 20315
rect 11664 20284 12173 20312
rect 11664 20272 11670 20284
rect 12161 20281 12173 20284
rect 12207 20281 12219 20315
rect 12161 20275 12219 20281
rect 9640 20216 9996 20244
rect 12360 20244 12388 20411
rect 13372 20380 13400 20411
rect 16482 20408 16488 20460
rect 16540 20448 16546 20460
rect 18156 20457 18184 20556
rect 19242 20544 19248 20556
rect 19300 20544 19306 20596
rect 19889 20587 19947 20593
rect 19889 20553 19901 20587
rect 19935 20584 19947 20587
rect 21450 20584 21456 20596
rect 19935 20556 21456 20584
rect 19935 20553 19947 20556
rect 19889 20547 19947 20553
rect 21450 20544 21456 20556
rect 21508 20544 21514 20596
rect 22186 20544 22192 20596
rect 22244 20584 22250 20596
rect 22649 20587 22707 20593
rect 22649 20584 22661 20587
rect 22244 20556 22661 20584
rect 22244 20544 22250 20556
rect 22649 20553 22661 20556
rect 22695 20553 22707 20587
rect 22649 20547 22707 20553
rect 25225 20587 25283 20593
rect 25225 20553 25237 20587
rect 25271 20584 25283 20587
rect 26326 20584 26332 20596
rect 25271 20556 26332 20584
rect 25271 20553 25283 20556
rect 25225 20547 25283 20553
rect 26326 20544 26332 20556
rect 26384 20544 26390 20596
rect 26973 20587 27031 20593
rect 26973 20553 26985 20587
rect 27019 20584 27031 20587
rect 27614 20584 27620 20596
rect 27019 20556 27620 20584
rect 27019 20553 27031 20556
rect 26973 20547 27031 20553
rect 27614 20544 27620 20556
rect 27672 20544 27678 20596
rect 19794 20516 19800 20528
rect 19642 20488 19800 20516
rect 19794 20476 19800 20488
rect 19852 20516 19858 20528
rect 20622 20516 20628 20528
rect 19852 20488 20628 20516
rect 19852 20476 19858 20488
rect 20622 20476 20628 20488
rect 20680 20516 20686 20528
rect 21085 20519 21143 20525
rect 21085 20516 21097 20519
rect 20680 20488 21097 20516
rect 20680 20476 20686 20488
rect 21085 20485 21097 20488
rect 21131 20485 21143 20519
rect 25498 20516 25504 20528
rect 24978 20488 25504 20516
rect 21085 20479 21143 20485
rect 25498 20476 25504 20488
rect 25556 20476 25562 20528
rect 27430 20476 27436 20528
rect 27488 20476 27494 20528
rect 28074 20476 28080 20528
rect 28132 20476 28138 20528
rect 28166 20476 28172 20528
rect 28224 20476 28230 20528
rect 17313 20451 17371 20457
rect 17313 20448 17325 20451
rect 16540 20420 17325 20448
rect 16540 20408 16546 20420
rect 17313 20417 17325 20420
rect 17359 20417 17371 20451
rect 17313 20411 17371 20417
rect 18141 20451 18199 20457
rect 18141 20417 18153 20451
rect 18187 20417 18199 20451
rect 18141 20411 18199 20417
rect 20530 20408 20536 20460
rect 20588 20448 20594 20460
rect 21450 20448 21456 20460
rect 20588 20420 21456 20448
rect 20588 20408 20594 20420
rect 21450 20408 21456 20420
rect 21508 20408 21514 20460
rect 21634 20408 21640 20460
rect 21692 20448 21698 20460
rect 22005 20451 22063 20457
rect 22005 20448 22017 20451
rect 21692 20420 22017 20448
rect 21692 20408 21698 20420
rect 22005 20417 22017 20420
rect 22051 20417 22063 20451
rect 22005 20411 22063 20417
rect 26789 20451 26847 20457
rect 26789 20417 26801 20451
rect 26835 20448 26847 20451
rect 27341 20451 27399 20457
rect 27341 20448 27353 20451
rect 26835 20420 27353 20448
rect 26835 20417 26847 20420
rect 26789 20411 26847 20417
rect 27341 20417 27353 20420
rect 27387 20417 27399 20451
rect 27341 20411 27399 20417
rect 27982 20408 27988 20460
rect 28040 20408 28046 20460
rect 28350 20408 28356 20460
rect 28408 20408 28414 20460
rect 14182 20380 14188 20392
rect 13372 20352 14188 20380
rect 14182 20340 14188 20352
rect 14240 20380 14246 20392
rect 14645 20383 14703 20389
rect 14645 20380 14657 20383
rect 14240 20352 14657 20380
rect 14240 20340 14246 20352
rect 14645 20349 14657 20352
rect 14691 20349 14703 20383
rect 14645 20343 14703 20349
rect 14921 20383 14979 20389
rect 14921 20349 14933 20383
rect 14967 20380 14979 20383
rect 15930 20380 15936 20392
rect 14967 20352 15936 20380
rect 14967 20349 14979 20352
rect 14921 20343 14979 20349
rect 15930 20340 15936 20352
rect 15988 20340 15994 20392
rect 17034 20340 17040 20392
rect 17092 20380 17098 20392
rect 17221 20383 17279 20389
rect 17221 20380 17233 20383
rect 17092 20352 17233 20380
rect 17092 20340 17098 20352
rect 17221 20349 17233 20352
rect 17267 20349 17279 20383
rect 17221 20343 17279 20349
rect 18417 20383 18475 20389
rect 18417 20349 18429 20383
rect 18463 20380 18475 20383
rect 18874 20380 18880 20392
rect 18463 20352 18880 20380
rect 18463 20349 18475 20352
rect 18417 20343 18475 20349
rect 18874 20340 18880 20352
rect 18932 20340 18938 20392
rect 23474 20340 23480 20392
rect 23532 20340 23538 20392
rect 23750 20340 23756 20392
rect 23808 20340 23814 20392
rect 26237 20383 26295 20389
rect 26237 20349 26249 20383
rect 26283 20380 26295 20383
rect 26694 20380 26700 20392
rect 26283 20352 26700 20380
rect 26283 20349 26295 20352
rect 26237 20343 26295 20349
rect 26694 20340 26700 20352
rect 26752 20340 26758 20392
rect 27246 20340 27252 20392
rect 27304 20380 27310 20392
rect 27525 20383 27583 20389
rect 27525 20380 27537 20383
rect 27304 20352 27537 20380
rect 27304 20340 27310 20352
rect 27525 20349 27537 20352
rect 27571 20349 27583 20383
rect 27525 20343 27583 20349
rect 19426 20272 19432 20324
rect 19484 20312 19490 20324
rect 19484 20284 23612 20312
rect 19484 20272 19490 20284
rect 16206 20244 16212 20256
rect 12360 20216 16212 20244
rect 9640 20204 9646 20216
rect 16206 20204 16212 20216
rect 16264 20244 16270 20256
rect 16393 20247 16451 20253
rect 16393 20244 16405 20247
rect 16264 20216 16405 20244
rect 16264 20204 16270 20216
rect 16393 20213 16405 20216
rect 16439 20213 16451 20247
rect 16393 20207 16451 20213
rect 17681 20247 17739 20253
rect 17681 20213 17693 20247
rect 17727 20244 17739 20247
rect 18230 20244 18236 20256
rect 17727 20216 18236 20244
rect 17727 20213 17739 20216
rect 17681 20207 17739 20213
rect 18230 20204 18236 20216
rect 18288 20204 18294 20256
rect 23584 20244 23612 20284
rect 25498 20272 25504 20324
rect 25556 20312 25562 20324
rect 28442 20312 28448 20324
rect 25556 20284 28448 20312
rect 25556 20272 25562 20284
rect 28442 20272 28448 20284
rect 28500 20272 28506 20324
rect 24394 20244 24400 20256
rect 23584 20216 24400 20244
rect 24394 20204 24400 20216
rect 24452 20204 24458 20256
rect 27801 20247 27859 20253
rect 27801 20213 27813 20247
rect 27847 20244 27859 20247
rect 27982 20244 27988 20256
rect 27847 20216 27988 20244
rect 27847 20213 27859 20216
rect 27801 20207 27859 20213
rect 27982 20204 27988 20216
rect 28040 20204 28046 20256
rect 1104 20154 28704 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 28704 20154
rect 1104 20080 28704 20102
rect 7190 20049 7196 20052
rect 7147 20043 7196 20049
rect 7147 20009 7159 20043
rect 7193 20009 7196 20043
rect 7147 20003 7196 20009
rect 7190 20000 7196 20003
rect 7248 20000 7254 20052
rect 7377 20043 7435 20049
rect 7377 20009 7389 20043
rect 7423 20040 7435 20043
rect 7742 20040 7748 20052
rect 7423 20012 7748 20040
rect 7423 20009 7435 20012
rect 7377 20003 7435 20009
rect 7742 20000 7748 20012
rect 7800 20000 7806 20052
rect 7929 20043 7987 20049
rect 7929 20009 7941 20043
rect 7975 20040 7987 20043
rect 8110 20040 8116 20052
rect 7975 20012 8116 20040
rect 7975 20009 7987 20012
rect 7929 20003 7987 20009
rect 8110 20000 8116 20012
rect 8168 20000 8174 20052
rect 8662 20000 8668 20052
rect 8720 20000 8726 20052
rect 12618 20000 12624 20052
rect 12676 20040 12682 20052
rect 13633 20043 13691 20049
rect 13633 20040 13645 20043
rect 12676 20012 13645 20040
rect 12676 20000 12682 20012
rect 13633 20009 13645 20012
rect 13679 20009 13691 20043
rect 13633 20003 13691 20009
rect 17402 20000 17408 20052
rect 17460 20000 17466 20052
rect 17586 20000 17592 20052
rect 17644 20040 17650 20052
rect 17773 20043 17831 20049
rect 17773 20040 17785 20043
rect 17644 20012 17785 20040
rect 17644 20000 17650 20012
rect 17773 20009 17785 20012
rect 17819 20009 17831 20043
rect 17773 20003 17831 20009
rect 19889 20043 19947 20049
rect 19889 20009 19901 20043
rect 19935 20040 19947 20043
rect 20162 20040 20168 20052
rect 19935 20012 20168 20040
rect 19935 20009 19947 20012
rect 19889 20003 19947 20009
rect 20162 20000 20168 20012
rect 20220 20000 20226 20052
rect 26694 20000 26700 20052
rect 26752 20040 26758 20052
rect 26789 20043 26847 20049
rect 26789 20040 26801 20043
rect 26752 20012 26801 20040
rect 26752 20000 26758 20012
rect 26789 20009 26801 20012
rect 26835 20009 26847 20043
rect 26789 20003 26847 20009
rect 27801 20043 27859 20049
rect 27801 20009 27813 20043
rect 27847 20040 27859 20043
rect 28258 20040 28264 20052
rect 27847 20012 28264 20040
rect 27847 20009 27859 20012
rect 27801 20003 27859 20009
rect 28258 20000 28264 20012
rect 28316 20000 28322 20052
rect 6914 19932 6920 19984
rect 6972 19972 6978 19984
rect 7285 19975 7343 19981
rect 7285 19972 7297 19975
rect 6972 19944 7297 19972
rect 6972 19932 6978 19944
rect 7285 19941 7297 19944
rect 7331 19941 7343 19975
rect 12636 19972 12664 20000
rect 15746 19972 15752 19984
rect 7285 19935 7343 19941
rect 11900 19944 12664 19972
rect 13832 19944 15752 19972
rect 5902 19864 5908 19916
rect 5960 19904 5966 19916
rect 8941 19907 8999 19913
rect 8941 19904 8953 19907
rect 5960 19876 7788 19904
rect 5960 19864 5966 19876
rect 7760 19848 7788 19876
rect 8496 19876 8953 19904
rect 7006 19796 7012 19848
rect 7064 19796 7070 19848
rect 7282 19796 7288 19848
rect 7340 19836 7346 19848
rect 7469 19839 7527 19845
rect 7469 19836 7481 19839
rect 7340 19808 7481 19836
rect 7340 19796 7346 19808
rect 7469 19805 7481 19808
rect 7515 19805 7527 19839
rect 7469 19799 7527 19805
rect 7742 19796 7748 19848
rect 7800 19836 7806 19848
rect 8113 19839 8171 19845
rect 8113 19836 8125 19839
rect 7800 19808 8125 19836
rect 7800 19796 7806 19808
rect 8113 19805 8125 19808
rect 8159 19805 8171 19839
rect 8113 19799 8171 19805
rect 8202 19796 8208 19848
rect 8260 19796 8266 19848
rect 8496 19845 8524 19876
rect 8941 19873 8953 19876
rect 8987 19873 8999 19907
rect 8941 19867 8999 19873
rect 11238 19864 11244 19916
rect 11296 19904 11302 19916
rect 11900 19904 11928 19944
rect 13832 19913 13860 19944
rect 15746 19932 15752 19944
rect 15804 19932 15810 19984
rect 17034 19932 17040 19984
rect 17092 19972 17098 19984
rect 24118 19972 24124 19984
rect 17092 19944 20668 19972
rect 17092 19932 17098 19944
rect 11296 19876 11928 19904
rect 11296 19864 11302 19876
rect 8481 19839 8539 19845
rect 8481 19805 8493 19839
rect 8527 19805 8539 19839
rect 8481 19799 8539 19805
rect 8757 19839 8815 19845
rect 8757 19805 8769 19839
rect 8803 19805 8815 19839
rect 8757 19799 8815 19805
rect 3602 19660 3608 19712
rect 3660 19700 3666 19712
rect 6822 19700 6828 19712
rect 3660 19672 6828 19700
rect 3660 19660 3666 19672
rect 6822 19660 6828 19672
rect 6880 19660 6886 19712
rect 7024 19700 7052 19796
rect 8294 19728 8300 19780
rect 8352 19728 8358 19780
rect 8772 19768 8800 19799
rect 9030 19796 9036 19848
rect 9088 19836 9094 19848
rect 9125 19839 9183 19845
rect 9125 19836 9137 19839
rect 9088 19808 9137 19836
rect 9088 19796 9094 19808
rect 9125 19805 9137 19808
rect 9171 19805 9183 19839
rect 9125 19799 9183 19805
rect 9401 19839 9459 19845
rect 9401 19805 9413 19839
rect 9447 19805 9459 19839
rect 9401 19799 9459 19805
rect 11517 19839 11575 19845
rect 11517 19805 11529 19839
rect 11563 19836 11575 19839
rect 11698 19836 11704 19848
rect 11563 19808 11704 19836
rect 11563 19805 11575 19808
rect 11517 19799 11575 19805
rect 9416 19768 9444 19799
rect 11698 19796 11704 19808
rect 11756 19796 11762 19848
rect 11900 19845 11928 19876
rect 12069 19907 12127 19913
rect 12069 19873 12081 19907
rect 12115 19904 12127 19907
rect 12452 19904 12756 19912
rect 13817 19907 13875 19913
rect 12115 19884 13584 19904
rect 12115 19876 12480 19884
rect 12728 19876 13584 19884
rect 12115 19873 12127 19876
rect 12069 19867 12127 19873
rect 12529 19849 12587 19855
rect 11885 19839 11943 19845
rect 11885 19805 11897 19839
rect 11931 19805 11943 19839
rect 11885 19799 11943 19805
rect 12437 19839 12495 19845
rect 12437 19805 12449 19839
rect 12483 19805 12495 19839
rect 12529 19815 12541 19849
rect 12575 19836 12587 19849
rect 12618 19836 12624 19848
rect 12575 19815 12624 19836
rect 12529 19809 12624 19815
rect 12544 19808 12624 19809
rect 12437 19799 12495 19805
rect 8772 19740 9444 19768
rect 12452 19768 12480 19799
rect 12618 19796 12624 19808
rect 12676 19796 12682 19848
rect 12897 19839 12955 19845
rect 12897 19805 12909 19839
rect 12943 19836 12955 19839
rect 13262 19836 13268 19848
rect 12943 19808 13268 19836
rect 12943 19805 12955 19808
rect 12897 19799 12955 19805
rect 12526 19768 12532 19780
rect 12452 19740 12532 19768
rect 8772 19700 8800 19740
rect 12526 19728 12532 19740
rect 12584 19768 12590 19780
rect 12912 19768 12940 19799
rect 13262 19796 13268 19808
rect 13320 19796 13326 19848
rect 13556 19845 13584 19876
rect 13817 19873 13829 19907
rect 13863 19873 13875 19907
rect 14185 19907 14243 19913
rect 14185 19904 14197 19907
rect 13817 19867 13875 19873
rect 13924 19876 14197 19904
rect 13541 19839 13599 19845
rect 13541 19805 13553 19839
rect 13587 19836 13599 19839
rect 13924 19836 13952 19876
rect 14185 19873 14197 19876
rect 14231 19873 14243 19907
rect 14185 19867 14243 19873
rect 16482 19864 16488 19916
rect 16540 19904 16546 19916
rect 16761 19907 16819 19913
rect 16761 19904 16773 19907
rect 16540 19876 16773 19904
rect 16540 19864 16546 19876
rect 16761 19873 16773 19876
rect 16807 19873 16819 19907
rect 18506 19904 18512 19916
rect 16761 19867 16819 19873
rect 17880 19876 18512 19904
rect 13587 19808 13952 19836
rect 14093 19839 14151 19845
rect 13587 19805 13599 19808
rect 13541 19799 13599 19805
rect 14093 19805 14105 19839
rect 14139 19805 14151 19839
rect 14093 19799 14151 19805
rect 15841 19839 15899 19845
rect 15841 19805 15853 19839
rect 15887 19836 15899 19839
rect 16022 19836 16028 19848
rect 15887 19808 16028 19836
rect 15887 19805 15899 19808
rect 15841 19799 15899 19805
rect 12584 19740 12940 19768
rect 13449 19771 13507 19777
rect 12584 19728 12590 19740
rect 13449 19737 13461 19771
rect 13495 19768 13507 19771
rect 14108 19768 14136 19799
rect 16022 19796 16028 19808
rect 16080 19836 16086 19848
rect 17880 19836 17908 19876
rect 18506 19864 18512 19876
rect 18564 19864 18570 19916
rect 20349 19907 20407 19913
rect 20349 19904 20361 19907
rect 19628 19876 20361 19904
rect 17954 19845 17960 19848
rect 16080 19808 17908 19836
rect 16080 19796 16086 19808
rect 17952 19799 17960 19845
rect 17954 19796 17960 19799
rect 18012 19796 18018 19848
rect 18230 19796 18236 19848
rect 18288 19845 18294 19848
rect 18288 19839 18327 19845
rect 18315 19805 18327 19839
rect 18288 19799 18327 19805
rect 18288 19796 18294 19799
rect 18414 19796 18420 19848
rect 18472 19836 18478 19848
rect 19242 19836 19248 19848
rect 18472 19808 19248 19836
rect 18472 19796 18478 19808
rect 19242 19796 19248 19808
rect 19300 19796 19306 19848
rect 19426 19845 19432 19848
rect 19393 19839 19432 19845
rect 19393 19805 19405 19839
rect 19393 19799 19432 19805
rect 19426 19796 19432 19799
rect 19484 19796 19490 19848
rect 19628 19845 19656 19876
rect 20349 19873 20361 19876
rect 20395 19904 20407 19907
rect 20530 19904 20536 19916
rect 20395 19876 20536 19904
rect 20395 19873 20407 19876
rect 20349 19867 20407 19873
rect 20530 19864 20536 19876
rect 20588 19864 20594 19916
rect 19613 19839 19671 19845
rect 19613 19805 19625 19839
rect 19659 19805 19671 19839
rect 19613 19799 19671 19805
rect 19702 19796 19708 19848
rect 19760 19845 19766 19848
rect 19760 19836 19768 19845
rect 20441 19839 20499 19845
rect 19760 19808 19805 19836
rect 19760 19799 19768 19808
rect 20441 19805 20453 19839
rect 20487 19836 20499 19839
rect 20640 19836 20668 19944
rect 23308 19944 24124 19972
rect 20809 19907 20867 19913
rect 20809 19873 20821 19907
rect 20855 19904 20867 19907
rect 21910 19904 21916 19916
rect 20855 19876 21916 19904
rect 20855 19873 20867 19876
rect 20809 19867 20867 19873
rect 21910 19864 21916 19876
rect 21968 19864 21974 19916
rect 22094 19864 22100 19916
rect 22152 19864 22158 19916
rect 22373 19907 22431 19913
rect 22373 19873 22385 19907
rect 22419 19904 22431 19907
rect 23198 19904 23204 19916
rect 22419 19876 23204 19904
rect 22419 19873 22431 19876
rect 22373 19867 22431 19873
rect 23198 19864 23204 19876
rect 23256 19864 23262 19916
rect 22005 19839 22063 19845
rect 22005 19836 22017 19839
rect 20487 19808 22017 19836
rect 20487 19805 20499 19808
rect 20441 19799 20499 19805
rect 22005 19805 22017 19808
rect 22051 19836 22063 19839
rect 23308 19836 23336 19944
rect 24118 19932 24124 19944
rect 24176 19932 24182 19984
rect 23474 19904 23480 19916
rect 23400 19876 23480 19904
rect 23400 19845 23428 19876
rect 23474 19864 23480 19876
rect 23532 19904 23538 19916
rect 23532 19876 25084 19904
rect 23532 19864 23538 19876
rect 25056 19848 25084 19876
rect 27246 19864 27252 19916
rect 27304 19864 27310 19916
rect 27341 19907 27399 19913
rect 27341 19873 27353 19907
rect 27387 19904 27399 19907
rect 27798 19904 27804 19916
rect 27387 19876 27804 19904
rect 27387 19873 27399 19876
rect 27341 19867 27399 19873
rect 27798 19864 27804 19876
rect 27856 19864 27862 19916
rect 22051 19808 23336 19836
rect 23385 19839 23443 19845
rect 22051 19805 22063 19808
rect 22005 19799 22063 19805
rect 23385 19805 23397 19839
rect 23431 19805 23443 19839
rect 23569 19839 23627 19845
rect 23569 19836 23581 19839
rect 23385 19799 23443 19805
rect 23492 19808 23581 19836
rect 19760 19796 19766 19799
rect 13495 19740 14136 19768
rect 13495 19737 13507 19740
rect 13449 19731 13507 19737
rect 7024 19672 8800 19700
rect 8846 19660 8852 19712
rect 8904 19700 8910 19712
rect 9309 19703 9367 19709
rect 9309 19700 9321 19703
rect 8904 19672 9321 19700
rect 8904 19660 8910 19672
rect 9309 19669 9321 19672
rect 9355 19669 9367 19703
rect 9309 19663 9367 19669
rect 9582 19660 9588 19712
rect 9640 19700 9646 19712
rect 11609 19703 11667 19709
rect 11609 19700 11621 19703
rect 9640 19672 11621 19700
rect 9640 19660 9646 19672
rect 11609 19669 11621 19672
rect 11655 19669 11667 19703
rect 11609 19663 11667 19669
rect 12713 19703 12771 19709
rect 12713 19669 12725 19703
rect 12759 19700 12771 19703
rect 12894 19700 12900 19712
rect 12759 19672 12900 19700
rect 12759 19669 12771 19672
rect 12713 19663 12771 19669
rect 12894 19660 12900 19672
rect 12952 19660 12958 19712
rect 13538 19660 13544 19712
rect 13596 19700 13602 19712
rect 13817 19703 13875 19709
rect 13817 19700 13829 19703
rect 13596 19672 13829 19700
rect 13596 19660 13602 19672
rect 13817 19669 13829 19672
rect 13863 19669 13875 19703
rect 13817 19663 13875 19669
rect 15657 19703 15715 19709
rect 15657 19669 15669 19703
rect 15703 19700 15715 19703
rect 15746 19700 15752 19712
rect 15703 19672 15752 19700
rect 15703 19669 15715 19672
rect 15657 19663 15715 19669
rect 15746 19660 15752 19672
rect 15804 19660 15810 19712
rect 17972 19700 18000 19796
rect 23492 19780 23520 19808
rect 23569 19805 23581 19808
rect 23615 19805 23627 19839
rect 23569 19799 23627 19805
rect 23662 19839 23720 19845
rect 23662 19805 23674 19839
rect 23708 19805 23720 19839
rect 23662 19799 23720 19805
rect 24075 19839 24133 19845
rect 24075 19805 24087 19839
rect 24121 19836 24133 19839
rect 24210 19836 24216 19848
rect 24121 19808 24216 19836
rect 24121 19805 24133 19808
rect 24075 19799 24133 19805
rect 18046 19728 18052 19780
rect 18104 19728 18110 19780
rect 18141 19771 18199 19777
rect 18141 19737 18153 19771
rect 18187 19768 18199 19771
rect 18598 19768 18604 19780
rect 18187 19740 18604 19768
rect 18187 19737 18199 19740
rect 18141 19731 18199 19737
rect 18598 19728 18604 19740
rect 18656 19768 18662 19780
rect 19521 19771 19579 19777
rect 19521 19768 19533 19771
rect 18656 19740 19533 19768
rect 18656 19728 18662 19740
rect 19521 19737 19533 19740
rect 19567 19768 19579 19771
rect 19567 19740 19748 19768
rect 19567 19737 19579 19740
rect 19521 19731 19579 19737
rect 18690 19700 18696 19712
rect 17972 19672 18696 19700
rect 18690 19660 18696 19672
rect 18748 19660 18754 19712
rect 19720 19700 19748 19740
rect 23474 19728 23480 19780
rect 23532 19728 23538 19780
rect 23676 19768 23704 19799
rect 24210 19796 24216 19808
rect 24268 19796 24274 19848
rect 24762 19796 24768 19848
rect 24820 19796 24826 19848
rect 25038 19796 25044 19848
rect 25096 19796 25102 19848
rect 27706 19796 27712 19848
rect 27764 19836 27770 19848
rect 27985 19839 28043 19845
rect 27985 19836 27997 19839
rect 27764 19808 27997 19836
rect 27764 19796 27770 19808
rect 27985 19805 27997 19808
rect 28031 19836 28043 19839
rect 28074 19836 28080 19848
rect 28031 19808 28080 19836
rect 28031 19805 28043 19808
rect 27985 19799 28043 19805
rect 28074 19796 28080 19808
rect 28132 19796 28138 19848
rect 28353 19839 28411 19845
rect 28353 19805 28365 19839
rect 28399 19836 28411 19839
rect 28442 19836 28448 19848
rect 28399 19808 28448 19836
rect 28399 19805 28411 19808
rect 28353 19799 28411 19805
rect 28442 19796 28448 19808
rect 28500 19796 28506 19848
rect 23676 19740 23796 19768
rect 22002 19700 22008 19712
rect 19720 19672 22008 19700
rect 22002 19660 22008 19672
rect 22060 19660 22066 19712
rect 23768 19700 23796 19740
rect 23842 19728 23848 19780
rect 23900 19728 23906 19780
rect 23934 19728 23940 19780
rect 23992 19728 23998 19780
rect 25317 19771 25375 19777
rect 25317 19768 25329 19771
rect 24228 19740 25329 19768
rect 24026 19700 24032 19712
rect 23768 19672 24032 19700
rect 24026 19660 24032 19672
rect 24084 19660 24090 19712
rect 24228 19709 24256 19740
rect 25317 19737 25329 19740
rect 25363 19737 25375 19771
rect 26786 19768 26792 19780
rect 26542 19740 26792 19768
rect 25317 19731 25375 19737
rect 26786 19728 26792 19740
rect 26844 19728 26850 19780
rect 24213 19703 24271 19709
rect 24213 19669 24225 19703
rect 24259 19669 24271 19703
rect 24213 19663 24271 19669
rect 27433 19703 27491 19709
rect 27433 19669 27445 19703
rect 27479 19700 27491 19703
rect 27706 19700 27712 19712
rect 27479 19672 27712 19700
rect 27479 19669 27491 19672
rect 27433 19663 27491 19669
rect 27706 19660 27712 19672
rect 27764 19660 27770 19712
rect 1104 19610 28704 19632
rect 1104 19558 4874 19610
rect 4926 19558 4938 19610
rect 4990 19558 5002 19610
rect 5054 19558 5066 19610
rect 5118 19558 5130 19610
rect 5182 19558 28704 19610
rect 1104 19536 28704 19558
rect 5905 19499 5963 19505
rect 5905 19496 5917 19499
rect 5092 19468 5917 19496
rect 4706 19388 4712 19440
rect 4764 19428 4770 19440
rect 4867 19431 4925 19437
rect 4867 19428 4879 19431
rect 4764 19400 4879 19428
rect 4764 19388 4770 19400
rect 4867 19397 4879 19400
rect 4913 19428 4925 19431
rect 4913 19397 4936 19428
rect 4867 19391 4936 19397
rect 4709 19295 4767 19301
rect 4709 19261 4721 19295
rect 4755 19292 4767 19295
rect 4908 19292 4936 19391
rect 4982 19320 4988 19372
rect 5040 19320 5046 19372
rect 5092 19369 5120 19468
rect 5905 19465 5917 19468
rect 5951 19465 5963 19499
rect 5905 19459 5963 19465
rect 11238 19456 11244 19508
rect 11296 19456 11302 19508
rect 11698 19456 11704 19508
rect 11756 19456 11762 19508
rect 12023 19499 12081 19505
rect 12023 19465 12035 19499
rect 12069 19496 12081 19499
rect 12526 19496 12532 19508
rect 12069 19468 12532 19496
rect 12069 19465 12081 19468
rect 12023 19459 12081 19465
rect 12526 19456 12532 19468
rect 12584 19456 12590 19508
rect 16022 19456 16028 19508
rect 16080 19456 16086 19508
rect 18046 19456 18052 19508
rect 18104 19496 18110 19508
rect 18141 19499 18199 19505
rect 18141 19496 18153 19499
rect 18104 19468 18153 19496
rect 18104 19456 18110 19468
rect 18141 19465 18153 19468
rect 18187 19465 18199 19499
rect 18141 19459 18199 19465
rect 18598 19456 18604 19508
rect 18656 19456 18662 19508
rect 18874 19456 18880 19508
rect 18932 19456 18938 19508
rect 19242 19456 19248 19508
rect 19300 19496 19306 19508
rect 19300 19468 21496 19496
rect 19300 19456 19306 19468
rect 8110 19428 8116 19440
rect 5184 19400 5488 19428
rect 5184 19369 5212 19400
rect 5077 19363 5135 19369
rect 5077 19329 5089 19363
rect 5123 19329 5135 19363
rect 5077 19323 5135 19329
rect 5169 19363 5227 19369
rect 5169 19329 5181 19363
rect 5215 19329 5227 19363
rect 5169 19323 5227 19329
rect 5258 19320 5264 19372
rect 5316 19320 5322 19372
rect 5460 19369 5488 19400
rect 7576 19400 8116 19428
rect 7576 19372 7604 19400
rect 8110 19388 8116 19400
rect 8168 19388 8174 19440
rect 11514 19428 11520 19440
rect 11164 19400 11520 19428
rect 5445 19363 5503 19369
rect 5445 19329 5457 19363
rect 5491 19329 5503 19363
rect 5445 19323 5503 19329
rect 5534 19320 5540 19372
rect 5592 19320 5598 19372
rect 5626 19320 5632 19372
rect 5684 19320 5690 19372
rect 5813 19363 5871 19369
rect 5813 19329 5825 19363
rect 5859 19329 5871 19363
rect 5813 19323 5871 19329
rect 5276 19292 5304 19320
rect 4755 19264 4844 19292
rect 4908 19264 5304 19292
rect 5353 19295 5411 19301
rect 4755 19261 4767 19264
rect 4709 19255 4767 19261
rect 4816 19236 4844 19264
rect 5353 19261 5365 19295
rect 5399 19292 5411 19295
rect 5552 19292 5580 19320
rect 5399 19264 5580 19292
rect 5828 19292 5856 19323
rect 5902 19320 5908 19372
rect 5960 19320 5966 19372
rect 6086 19320 6092 19372
rect 6144 19320 6150 19372
rect 6822 19320 6828 19372
rect 6880 19360 6886 19372
rect 7558 19360 7564 19372
rect 6880 19332 7564 19360
rect 6880 19320 6886 19332
rect 7558 19320 7564 19332
rect 7616 19320 7622 19372
rect 8938 19320 8944 19372
rect 8996 19320 9002 19372
rect 11164 19369 11192 19400
rect 11514 19388 11520 19400
rect 11572 19388 11578 19440
rect 11716 19428 11744 19456
rect 11716 19400 12388 19428
rect 11149 19363 11207 19369
rect 11149 19329 11161 19363
rect 11195 19329 11207 19363
rect 11149 19323 11207 19329
rect 11330 19320 11336 19372
rect 11388 19320 11394 19372
rect 11422 19320 11428 19372
rect 11480 19360 11486 19372
rect 11885 19363 11943 19369
rect 11885 19360 11897 19363
rect 11480 19332 11897 19360
rect 11480 19320 11486 19332
rect 11885 19329 11897 19332
rect 11931 19329 11943 19363
rect 12360 19360 12388 19400
rect 12710 19388 12716 19440
rect 12768 19388 12774 19440
rect 18414 19428 18420 19440
rect 18248 19400 18420 19428
rect 13449 19363 13507 19369
rect 12360 19332 12434 19360
rect 11885 19323 11943 19329
rect 6104 19292 6132 19320
rect 7837 19295 7895 19301
rect 7837 19292 7849 19295
rect 5828 19264 6132 19292
rect 7668 19264 7849 19292
rect 5399 19261 5411 19264
rect 5353 19255 5411 19261
rect 4798 19184 4804 19236
rect 4856 19184 4862 19236
rect 7558 19184 7564 19236
rect 7616 19224 7622 19236
rect 7668 19224 7696 19264
rect 7837 19261 7849 19264
rect 7883 19261 7895 19295
rect 7837 19255 7895 19261
rect 7616 19196 7696 19224
rect 7616 19184 7622 19196
rect 4062 19116 4068 19168
rect 4120 19156 4126 19168
rect 5442 19156 5448 19168
rect 4120 19128 5448 19156
rect 4120 19116 4126 19128
rect 5442 19116 5448 19128
rect 5500 19156 5506 19168
rect 8938 19156 8944 19168
rect 5500 19128 8944 19156
rect 5500 19116 5506 19128
rect 8938 19116 8944 19128
rect 8996 19116 9002 19168
rect 9306 19116 9312 19168
rect 9364 19116 9370 19168
rect 11900 19156 11928 19323
rect 12406 19292 12434 19332
rect 13449 19329 13461 19363
rect 13495 19360 13507 19363
rect 13538 19360 13544 19372
rect 13495 19332 13544 19360
rect 13495 19329 13507 19332
rect 13449 19323 13507 19329
rect 13538 19320 13544 19332
rect 13596 19320 13602 19372
rect 16206 19320 16212 19372
rect 16264 19320 16270 19372
rect 17034 19320 17040 19372
rect 17092 19360 17098 19372
rect 17954 19360 17960 19372
rect 17092 19332 17960 19360
rect 17092 19320 17098 19332
rect 17954 19320 17960 19332
rect 18012 19320 18018 19372
rect 18248 19369 18276 19400
rect 18414 19388 18420 19400
rect 18472 19388 18478 19440
rect 18509 19431 18567 19437
rect 18509 19397 18521 19431
rect 18555 19428 18567 19431
rect 18616 19428 18644 19456
rect 18555 19400 18644 19428
rect 18555 19397 18567 19400
rect 18509 19391 18567 19397
rect 18233 19363 18291 19369
rect 18233 19329 18245 19363
rect 18279 19329 18291 19363
rect 18233 19323 18291 19329
rect 18326 19363 18384 19369
rect 18326 19329 18338 19363
rect 18372 19329 18384 19363
rect 18326 19323 18384 19329
rect 12986 19292 12992 19304
rect 12406 19264 12992 19292
rect 12986 19252 12992 19264
rect 13044 19252 13050 19304
rect 13817 19295 13875 19301
rect 13817 19261 13829 19295
rect 13863 19292 13875 19295
rect 14182 19292 14188 19304
rect 13863 19264 14188 19292
rect 13863 19261 13875 19264
rect 13817 19255 13875 19261
rect 14182 19252 14188 19264
rect 14240 19252 14246 19304
rect 15562 19252 15568 19304
rect 15620 19292 15626 19304
rect 15749 19295 15807 19301
rect 15749 19292 15761 19295
rect 15620 19264 15761 19292
rect 15620 19252 15626 19264
rect 15749 19261 15761 19264
rect 15795 19292 15807 19295
rect 16482 19292 16488 19304
rect 15795 19264 16488 19292
rect 15795 19261 15807 19264
rect 15749 19255 15807 19261
rect 16482 19252 16488 19264
rect 16540 19252 16546 19304
rect 17129 19295 17187 19301
rect 17129 19261 17141 19295
rect 17175 19292 17187 19295
rect 17494 19292 17500 19304
rect 17175 19264 17500 19292
rect 17175 19261 17187 19264
rect 17129 19255 17187 19261
rect 17494 19252 17500 19264
rect 17552 19252 17558 19304
rect 17405 19227 17463 19233
rect 14476 19196 16160 19224
rect 14476 19156 14504 19196
rect 11900 19128 14504 19156
rect 14550 19116 14556 19168
rect 14608 19156 14614 19168
rect 15105 19159 15163 19165
rect 15105 19156 15117 19159
rect 14608 19128 15117 19156
rect 14608 19116 14614 19128
rect 15105 19125 15117 19128
rect 15151 19125 15163 19159
rect 16132 19156 16160 19196
rect 17405 19193 17417 19227
rect 17451 19224 17463 19227
rect 18340 19224 18368 19323
rect 18598 19320 18604 19372
rect 18656 19320 18662 19372
rect 18690 19320 18696 19372
rect 18748 19369 18754 19372
rect 18748 19363 18797 19369
rect 18748 19329 18751 19363
rect 18785 19360 18797 19363
rect 19702 19360 19708 19372
rect 18785 19332 19708 19360
rect 18785 19329 18797 19332
rect 18748 19323 18797 19329
rect 18748 19320 18754 19323
rect 19702 19320 19708 19332
rect 19760 19320 19766 19372
rect 20438 19320 20444 19372
rect 20496 19360 20502 19372
rect 21269 19363 21327 19369
rect 21269 19360 21281 19363
rect 20496 19332 21281 19360
rect 20496 19320 20502 19332
rect 21269 19329 21281 19332
rect 21315 19329 21327 19363
rect 21468 19360 21496 19468
rect 22278 19456 22284 19508
rect 22336 19496 22342 19508
rect 22465 19499 22523 19505
rect 22465 19496 22477 19499
rect 22336 19468 22477 19496
rect 22336 19456 22342 19468
rect 22465 19465 22477 19468
rect 22511 19465 22523 19499
rect 22465 19459 22523 19465
rect 23124 19468 23612 19496
rect 22002 19388 22008 19440
rect 22060 19428 22066 19440
rect 22189 19431 22247 19437
rect 22060 19400 22140 19428
rect 22060 19388 22066 19400
rect 21821 19363 21879 19369
rect 21821 19360 21833 19363
rect 21468 19332 21833 19360
rect 21269 19323 21327 19329
rect 21821 19329 21833 19332
rect 21867 19329 21879 19363
rect 21821 19323 21879 19329
rect 21837 19292 21865 19323
rect 21910 19320 21916 19372
rect 21968 19360 21974 19372
rect 22112 19369 22140 19400
rect 22189 19397 22201 19431
rect 22235 19428 22247 19431
rect 22557 19431 22615 19437
rect 22557 19428 22569 19431
rect 22235 19400 22569 19428
rect 22235 19397 22247 19400
rect 22189 19391 22247 19397
rect 22557 19397 22569 19400
rect 22603 19397 22615 19431
rect 22557 19391 22615 19397
rect 22097 19363 22155 19369
rect 21968 19332 22013 19360
rect 21968 19320 21974 19332
rect 22097 19329 22109 19363
rect 22143 19360 22155 19363
rect 22143 19332 22237 19360
rect 22143 19329 22155 19332
rect 22097 19323 22155 19329
rect 22209 19292 22237 19332
rect 22278 19320 22284 19372
rect 22336 19369 22342 19372
rect 22336 19360 22344 19369
rect 23124 19360 23152 19468
rect 23198 19388 23204 19440
rect 23256 19428 23262 19440
rect 23256 19400 23428 19428
rect 23256 19388 23262 19400
rect 23400 19369 23428 19400
rect 23584 19372 23612 19468
rect 23750 19456 23756 19508
rect 23808 19496 23814 19508
rect 23937 19499 23995 19505
rect 23937 19496 23949 19499
rect 23808 19468 23949 19496
rect 23808 19456 23814 19468
rect 23937 19465 23949 19468
rect 23983 19465 23995 19499
rect 23937 19459 23995 19465
rect 27706 19456 27712 19508
rect 27764 19456 27770 19508
rect 24210 19428 24216 19440
rect 23812 19400 24216 19428
rect 23812 19372 23840 19400
rect 24210 19388 24216 19400
rect 24268 19388 24274 19440
rect 24305 19431 24363 19437
rect 24305 19397 24317 19431
rect 24351 19428 24363 19431
rect 24394 19428 24400 19440
rect 24351 19400 24400 19428
rect 24351 19397 24363 19400
rect 24305 19391 24363 19397
rect 24394 19388 24400 19400
rect 24452 19388 24458 19440
rect 22336 19332 22381 19360
rect 22480 19332 23152 19360
rect 23293 19363 23351 19369
rect 22336 19323 22344 19332
rect 22336 19320 22342 19323
rect 22480 19292 22508 19332
rect 23293 19329 23305 19363
rect 23339 19329 23351 19363
rect 23293 19323 23351 19329
rect 23386 19363 23444 19369
rect 23386 19329 23398 19363
rect 23432 19329 23444 19363
rect 23386 19323 23444 19329
rect 21837 19264 22094 19292
rect 22209 19264 22508 19292
rect 17451 19196 18368 19224
rect 17451 19193 17463 19196
rect 17405 19187 17463 19193
rect 18046 19156 18052 19168
rect 16132 19128 18052 19156
rect 15105 19119 15163 19125
rect 18046 19116 18052 19128
rect 18104 19116 18110 19168
rect 22066 19156 22094 19264
rect 23198 19252 23204 19304
rect 23256 19252 23262 19304
rect 23308 19292 23336 19323
rect 23566 19320 23572 19372
rect 23624 19320 23630 19372
rect 23658 19320 23664 19372
rect 23716 19320 23722 19372
rect 23750 19320 23756 19372
rect 23808 19360 23840 19372
rect 24228 19360 24256 19388
rect 24946 19360 24952 19372
rect 23808 19332 23853 19360
rect 24228 19332 24952 19360
rect 23808 19323 23816 19332
rect 23808 19320 23814 19323
rect 24946 19320 24952 19332
rect 25004 19320 25010 19372
rect 23474 19292 23480 19304
rect 23308 19264 23480 19292
rect 23474 19252 23480 19264
rect 23532 19292 23538 19304
rect 24486 19292 24492 19304
rect 23532 19264 24492 19292
rect 23532 19252 23538 19264
rect 24486 19252 24492 19264
rect 24544 19252 24550 19304
rect 25038 19252 25044 19304
rect 25096 19292 25102 19304
rect 25133 19295 25191 19301
rect 25133 19292 25145 19295
rect 25096 19264 25145 19292
rect 25096 19252 25102 19264
rect 25133 19261 25145 19264
rect 25179 19292 25191 19295
rect 26142 19292 26148 19304
rect 25179 19264 26148 19292
rect 25179 19261 25191 19264
rect 25133 19255 25191 19261
rect 26142 19252 26148 19264
rect 26200 19252 26206 19304
rect 27890 19252 27896 19304
rect 27948 19292 27954 19304
rect 28261 19295 28319 19301
rect 28261 19292 28273 19295
rect 27948 19264 28273 19292
rect 27948 19252 27954 19264
rect 28261 19261 28273 19264
rect 28307 19261 28319 19295
rect 28261 19255 28319 19261
rect 23492 19156 23520 19252
rect 22066 19128 23520 19156
rect 1104 19066 28704 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 28704 19066
rect 1104 18992 28704 19014
rect 5442 18912 5448 18964
rect 5500 18952 5506 18964
rect 5537 18955 5595 18961
rect 5537 18952 5549 18955
rect 5500 18924 5549 18952
rect 5500 18912 5506 18924
rect 5537 18921 5549 18924
rect 5583 18921 5595 18955
rect 5537 18915 5595 18921
rect 6086 18912 6092 18964
rect 6144 18952 6150 18964
rect 6273 18955 6331 18961
rect 6273 18952 6285 18955
rect 6144 18924 6285 18952
rect 6144 18912 6150 18924
rect 6273 18921 6285 18924
rect 6319 18921 6331 18955
rect 6273 18915 6331 18921
rect 8938 18912 8944 18964
rect 8996 18952 9002 18964
rect 9033 18955 9091 18961
rect 9033 18952 9045 18955
rect 8996 18924 9045 18952
rect 8996 18912 9002 18924
rect 9033 18921 9045 18924
rect 9079 18921 9091 18955
rect 9033 18915 9091 18921
rect 11330 18912 11336 18964
rect 11388 18952 11394 18964
rect 11885 18955 11943 18961
rect 11885 18952 11897 18955
rect 11388 18924 11897 18952
rect 11388 18912 11394 18924
rect 11885 18921 11897 18924
rect 11931 18921 11943 18955
rect 14461 18955 14519 18961
rect 14461 18952 14473 18955
rect 11885 18915 11943 18921
rect 12406 18924 14473 18952
rect 5258 18844 5264 18896
rect 5316 18884 5322 18896
rect 5721 18887 5779 18893
rect 5721 18884 5733 18887
rect 5316 18856 5733 18884
rect 5316 18844 5322 18856
rect 5721 18853 5733 18856
rect 5767 18884 5779 18887
rect 5767 18856 6500 18884
rect 5767 18853 5779 18856
rect 5721 18847 5779 18853
rect 5902 18816 5908 18828
rect 5644 18788 5908 18816
rect 4798 18708 4804 18760
rect 4856 18748 4862 18760
rect 5353 18751 5411 18757
rect 5353 18748 5365 18751
rect 4856 18720 5365 18748
rect 4856 18708 4862 18720
rect 5353 18717 5365 18720
rect 5399 18717 5411 18751
rect 5353 18711 5411 18717
rect 5445 18751 5503 18757
rect 5445 18717 5457 18751
rect 5491 18748 5503 18751
rect 5534 18748 5540 18760
rect 5491 18720 5540 18748
rect 5491 18717 5503 18720
rect 5445 18711 5503 18717
rect 4430 18640 4436 18692
rect 4488 18680 4494 18692
rect 5368 18680 5396 18711
rect 5534 18708 5540 18720
rect 5592 18708 5598 18760
rect 5644 18680 5672 18788
rect 5902 18776 5908 18788
rect 5960 18816 5966 18828
rect 5960 18788 6132 18816
rect 5960 18776 5966 18788
rect 5718 18708 5724 18760
rect 5776 18708 5782 18760
rect 5994 18708 6000 18760
rect 6052 18708 6058 18760
rect 6104 18757 6132 18788
rect 6472 18757 6500 18856
rect 11422 18844 11428 18896
rect 11480 18844 11486 18896
rect 12406 18884 12434 18924
rect 14461 18921 14473 18924
rect 14507 18952 14519 18955
rect 14829 18955 14887 18961
rect 14829 18952 14841 18955
rect 14507 18924 14841 18952
rect 14507 18921 14519 18924
rect 14461 18915 14519 18921
rect 14829 18921 14841 18924
rect 14875 18921 14887 18955
rect 15838 18952 15844 18964
rect 14829 18915 14887 18921
rect 14936 18924 15844 18952
rect 12802 18884 12808 18896
rect 11532 18856 12434 18884
rect 12544 18856 12808 18884
rect 10962 18816 10968 18828
rect 6564 18788 10968 18816
rect 6089 18751 6147 18757
rect 6089 18717 6101 18751
rect 6135 18717 6147 18751
rect 6089 18711 6147 18717
rect 6457 18751 6515 18757
rect 6457 18717 6469 18751
rect 6503 18717 6515 18751
rect 6457 18711 6515 18717
rect 6564 18680 6592 18788
rect 10962 18776 10968 18788
rect 11020 18816 11026 18828
rect 11532 18816 11560 18856
rect 11020 18788 11560 18816
rect 11020 18776 11026 18788
rect 11974 18776 11980 18828
rect 12032 18816 12038 18828
rect 12544 18825 12572 18856
rect 12802 18844 12808 18856
rect 12860 18844 12866 18896
rect 13817 18887 13875 18893
rect 13817 18853 13829 18887
rect 13863 18884 13875 18887
rect 14936 18884 14964 18924
rect 15838 18912 15844 18924
rect 15896 18952 15902 18964
rect 18230 18952 18236 18964
rect 15896 18924 18236 18952
rect 15896 18912 15902 18924
rect 18230 18912 18236 18924
rect 18288 18912 18294 18964
rect 18417 18955 18475 18961
rect 18417 18921 18429 18955
rect 18463 18952 18475 18955
rect 18598 18952 18604 18964
rect 18463 18924 18604 18952
rect 18463 18921 18475 18924
rect 18417 18915 18475 18921
rect 18598 18912 18604 18924
rect 18656 18912 18662 18964
rect 23658 18912 23664 18964
rect 23716 18952 23722 18964
rect 23937 18955 23995 18961
rect 23937 18952 23949 18955
rect 23716 18924 23949 18952
rect 23716 18912 23722 18924
rect 23937 18921 23949 18924
rect 23983 18921 23995 18955
rect 23937 18915 23995 18921
rect 27890 18912 27896 18964
rect 27948 18912 27954 18964
rect 13863 18856 14964 18884
rect 18325 18887 18383 18893
rect 13863 18853 13875 18856
rect 13817 18847 13875 18853
rect 18325 18853 18337 18887
rect 18371 18884 18383 18887
rect 19426 18884 19432 18896
rect 18371 18856 19432 18884
rect 18371 18853 18383 18856
rect 18325 18847 18383 18853
rect 12161 18819 12219 18825
rect 12161 18816 12173 18819
rect 12032 18788 12173 18816
rect 12032 18776 12038 18788
rect 12161 18785 12173 18788
rect 12207 18785 12219 18819
rect 12161 18779 12219 18785
rect 12529 18819 12587 18825
rect 12529 18785 12541 18819
rect 12575 18785 12587 18819
rect 12894 18816 12900 18828
rect 12529 18779 12587 18785
rect 12820 18788 12900 18816
rect 8570 18708 8576 18760
rect 8628 18748 8634 18760
rect 9309 18751 9367 18757
rect 9309 18748 9321 18751
rect 8628 18720 9321 18748
rect 8628 18708 8634 18720
rect 9309 18717 9321 18720
rect 9355 18717 9367 18751
rect 9309 18711 9367 18717
rect 9769 18751 9827 18757
rect 9769 18717 9781 18751
rect 9815 18748 9827 18751
rect 9858 18748 9864 18760
rect 9815 18720 9864 18748
rect 9815 18717 9827 18720
rect 9769 18711 9827 18717
rect 9858 18708 9864 18720
rect 9916 18708 9922 18760
rect 11146 18708 11152 18760
rect 11204 18748 11210 18760
rect 11241 18751 11299 18757
rect 11241 18748 11253 18751
rect 11204 18720 11253 18748
rect 11204 18708 11210 18720
rect 11241 18717 11253 18720
rect 11287 18717 11299 18751
rect 11241 18711 11299 18717
rect 11425 18751 11483 18757
rect 11425 18717 11437 18751
rect 11471 18717 11483 18751
rect 11425 18711 11483 18717
rect 4488 18652 4660 18680
rect 5368 18652 5672 18680
rect 5736 18652 6592 18680
rect 4488 18640 4494 18652
rect 4249 18615 4307 18621
rect 4249 18581 4261 18615
rect 4295 18612 4307 18615
rect 4522 18612 4528 18624
rect 4295 18584 4528 18612
rect 4295 18581 4307 18584
rect 4249 18575 4307 18581
rect 4522 18572 4528 18584
rect 4580 18572 4586 18624
rect 4632 18612 4660 18652
rect 5736 18612 5764 18652
rect 7742 18640 7748 18692
rect 7800 18680 7806 18692
rect 9876 18680 9904 18708
rect 11440 18680 11468 18711
rect 11606 18708 11612 18760
rect 11664 18708 11670 18760
rect 11698 18708 11704 18760
rect 11756 18748 11762 18760
rect 12820 18757 12848 18788
rect 12894 18776 12900 18788
rect 12952 18816 12958 18828
rect 13832 18816 13860 18847
rect 19426 18844 19432 18856
rect 19484 18844 19490 18896
rect 23198 18844 23204 18896
rect 23256 18844 23262 18896
rect 12952 18788 13860 18816
rect 12952 18776 12958 18788
rect 14182 18776 14188 18828
rect 14240 18816 14246 18828
rect 15105 18819 15163 18825
rect 15105 18816 15117 18819
rect 14240 18788 15117 18816
rect 14240 18776 14246 18788
rect 15105 18785 15117 18788
rect 15151 18785 15163 18819
rect 15105 18779 15163 18785
rect 16853 18819 16911 18825
rect 16853 18785 16865 18819
rect 16899 18816 16911 18819
rect 17494 18816 17500 18828
rect 16899 18788 17500 18816
rect 16899 18785 16911 18788
rect 16853 18779 16911 18785
rect 17494 18776 17500 18788
rect 17552 18776 17558 18828
rect 18049 18819 18107 18825
rect 18049 18785 18061 18819
rect 18095 18816 18107 18819
rect 18598 18816 18604 18828
rect 18095 18788 18604 18816
rect 18095 18785 18107 18788
rect 18049 18779 18107 18785
rect 18598 18776 18604 18788
rect 18656 18816 18662 18828
rect 18969 18819 19027 18825
rect 18969 18816 18981 18819
rect 18656 18788 18981 18816
rect 18656 18776 18662 18788
rect 18969 18785 18981 18788
rect 19015 18785 19027 18819
rect 18969 18779 19027 18785
rect 20165 18819 20223 18825
rect 20165 18785 20177 18819
rect 20211 18816 20223 18819
rect 20438 18816 20444 18828
rect 20211 18788 20444 18816
rect 20211 18785 20223 18788
rect 20165 18779 20223 18785
rect 20438 18776 20444 18788
rect 20496 18776 20502 18828
rect 22094 18776 22100 18828
rect 22152 18816 22158 18828
rect 22189 18819 22247 18825
rect 22189 18816 22201 18819
rect 22152 18788 22201 18816
rect 22152 18776 22158 18788
rect 22189 18785 22201 18788
rect 22235 18816 22247 18819
rect 22925 18819 22983 18825
rect 22925 18816 22937 18819
rect 22235 18788 22937 18816
rect 22235 18785 22247 18788
rect 22189 18779 22247 18785
rect 22925 18785 22937 18788
rect 22971 18816 22983 18819
rect 23216 18816 23244 18844
rect 23382 18816 23388 18828
rect 22971 18788 23388 18816
rect 22971 18785 22983 18788
rect 22925 18779 22983 18785
rect 23382 18776 23388 18788
rect 23440 18776 23446 18828
rect 23566 18776 23572 18828
rect 23624 18816 23630 18828
rect 23842 18816 23848 18828
rect 23624 18788 23848 18816
rect 23624 18776 23630 18788
rect 23842 18776 23848 18788
rect 23900 18816 23906 18828
rect 24489 18819 24547 18825
rect 24489 18816 24501 18819
rect 23900 18788 24501 18816
rect 23900 18776 23906 18788
rect 24489 18785 24501 18788
rect 24535 18785 24547 18819
rect 24489 18779 24547 18785
rect 12069 18751 12127 18757
rect 12069 18748 12081 18751
rect 11756 18720 12081 18748
rect 11756 18708 11762 18720
rect 12069 18717 12081 18720
rect 12115 18717 12127 18751
rect 12069 18711 12127 18717
rect 12805 18751 12863 18757
rect 12805 18717 12817 18751
rect 12851 18717 12863 18751
rect 12805 18711 12863 18717
rect 12986 18708 12992 18760
rect 13044 18748 13050 18760
rect 13081 18751 13139 18757
rect 13081 18748 13093 18751
rect 13044 18720 13093 18748
rect 13044 18708 13050 18720
rect 13081 18717 13093 18720
rect 13127 18717 13139 18751
rect 13081 18711 13139 18717
rect 11793 18683 11851 18689
rect 11793 18680 11805 18683
rect 7800 18652 9812 18680
rect 9876 18652 11805 18680
rect 7800 18640 7806 18652
rect 4632 18584 5764 18612
rect 5810 18572 5816 18624
rect 5868 18572 5874 18624
rect 8846 18572 8852 18624
rect 8904 18612 8910 18624
rect 9585 18615 9643 18621
rect 9585 18612 9597 18615
rect 8904 18584 9597 18612
rect 8904 18572 8910 18584
rect 9585 18581 9597 18584
rect 9631 18581 9643 18615
rect 9784 18612 9812 18652
rect 11793 18649 11805 18652
rect 11839 18680 11851 18683
rect 13096 18680 13124 18711
rect 13262 18708 13268 18760
rect 13320 18748 13326 18760
rect 13357 18751 13415 18757
rect 13357 18748 13369 18751
rect 13320 18720 13369 18748
rect 13320 18708 13326 18720
rect 13357 18717 13369 18720
rect 13403 18717 13415 18751
rect 13357 18711 13415 18717
rect 13541 18751 13599 18757
rect 13541 18717 13553 18751
rect 13587 18717 13599 18751
rect 13541 18711 13599 18717
rect 14277 18751 14335 18757
rect 14277 18717 14289 18751
rect 14323 18748 14335 18751
rect 14458 18748 14464 18760
rect 14323 18720 14464 18748
rect 14323 18717 14335 18720
rect 14277 18711 14335 18717
rect 13556 18680 13584 18711
rect 14458 18708 14464 18720
rect 14516 18708 14522 18760
rect 14550 18708 14556 18760
rect 14608 18708 14614 18760
rect 14645 18751 14703 18757
rect 14645 18717 14657 18751
rect 14691 18717 14703 18751
rect 14645 18711 14703 18717
rect 14660 18680 14688 18711
rect 16482 18708 16488 18760
rect 16540 18708 16546 18760
rect 17954 18708 17960 18760
rect 18012 18708 18018 18760
rect 23198 18708 23204 18760
rect 23256 18748 23262 18760
rect 23293 18751 23351 18757
rect 23293 18748 23305 18751
rect 23256 18720 23305 18748
rect 23256 18708 23262 18720
rect 23293 18717 23305 18720
rect 23339 18717 23351 18751
rect 23293 18711 23351 18717
rect 24673 18751 24731 18757
rect 24673 18717 24685 18751
rect 24719 18717 24731 18751
rect 24673 18711 24731 18717
rect 11839 18652 12756 18680
rect 13096 18652 13584 18680
rect 13648 18652 14228 18680
rect 11839 18649 11851 18652
rect 11793 18643 11851 18649
rect 12728 18624 12756 18652
rect 11422 18612 11428 18624
rect 9784 18584 11428 18612
rect 9585 18575 9643 18581
rect 11422 18572 11428 18584
rect 11480 18572 11486 18624
rect 12618 18572 12624 18624
rect 12676 18572 12682 18624
rect 12710 18572 12716 18624
rect 12768 18572 12774 18624
rect 13262 18572 13268 18624
rect 13320 18612 13326 18624
rect 13648 18621 13676 18652
rect 13633 18615 13691 18621
rect 13633 18612 13645 18615
rect 13320 18584 13645 18612
rect 13320 18572 13326 18584
rect 13633 18581 13645 18584
rect 13679 18581 13691 18615
rect 13633 18575 13691 18581
rect 14090 18572 14096 18624
rect 14148 18572 14154 18624
rect 14200 18612 14228 18652
rect 14384 18652 14688 18680
rect 14384 18612 14412 18652
rect 15378 18640 15384 18692
rect 15436 18640 15442 18692
rect 19334 18680 19340 18692
rect 16684 18652 19340 18680
rect 14200 18584 14412 18612
rect 14458 18572 14464 18624
rect 14516 18612 14522 18624
rect 15194 18612 15200 18624
rect 14516 18584 15200 18612
rect 14516 18572 14522 18584
rect 15194 18572 15200 18584
rect 15252 18612 15258 18624
rect 16206 18612 16212 18624
rect 15252 18584 16212 18612
rect 15252 18572 15258 18584
rect 16206 18572 16212 18584
rect 16264 18572 16270 18624
rect 16390 18572 16396 18624
rect 16448 18612 16454 18624
rect 16684 18612 16712 18652
rect 19334 18640 19340 18652
rect 19392 18640 19398 18692
rect 20717 18683 20775 18689
rect 20717 18649 20729 18683
rect 20763 18680 20775 18683
rect 20806 18680 20812 18692
rect 20763 18652 20812 18680
rect 20763 18649 20775 18652
rect 20717 18643 20775 18649
rect 20806 18640 20812 18652
rect 20864 18640 20870 18692
rect 21174 18640 21180 18692
rect 21232 18640 21238 18692
rect 22002 18640 22008 18692
rect 22060 18680 22066 18692
rect 22281 18683 22339 18689
rect 22281 18680 22293 18683
rect 22060 18652 22293 18680
rect 22060 18640 22066 18652
rect 22281 18649 22293 18652
rect 22327 18649 22339 18683
rect 24688 18680 24716 18711
rect 24854 18708 24860 18760
rect 24912 18708 24918 18760
rect 26142 18708 26148 18760
rect 26200 18708 26206 18760
rect 25038 18680 25044 18692
rect 24688 18652 25044 18680
rect 22281 18643 22339 18649
rect 25038 18640 25044 18652
rect 25096 18640 25102 18692
rect 25774 18640 25780 18692
rect 25832 18680 25838 18692
rect 26421 18683 26479 18689
rect 26421 18680 26433 18683
rect 25832 18652 26433 18680
rect 25832 18640 25838 18652
rect 26421 18649 26433 18652
rect 26467 18649 26479 18683
rect 26421 18643 26479 18649
rect 26878 18640 26884 18692
rect 26936 18640 26942 18692
rect 16448 18584 16712 18612
rect 16448 18572 16454 18584
rect 16942 18572 16948 18624
rect 17000 18572 17006 18624
rect 18138 18572 18144 18624
rect 18196 18612 18202 18624
rect 22370 18612 22376 18624
rect 18196 18584 22376 18612
rect 18196 18572 18202 18584
rect 22370 18572 22376 18584
rect 22428 18572 22434 18624
rect 1104 18522 28704 18544
rect 1104 18470 4874 18522
rect 4926 18470 4938 18522
rect 4990 18470 5002 18522
rect 5054 18470 5066 18522
rect 5118 18470 5130 18522
rect 5182 18470 28704 18522
rect 1104 18448 28704 18470
rect 3881 18411 3939 18417
rect 3881 18377 3893 18411
rect 3927 18408 3939 18411
rect 4798 18408 4804 18420
rect 3927 18380 4804 18408
rect 3927 18377 3939 18380
rect 3881 18371 3939 18377
rect 4798 18368 4804 18380
rect 4856 18368 4862 18420
rect 5074 18368 5080 18420
rect 5132 18408 5138 18420
rect 5442 18408 5448 18420
rect 5132 18380 5448 18408
rect 5132 18368 5138 18380
rect 5442 18368 5448 18380
rect 5500 18368 5506 18420
rect 5810 18408 5816 18420
rect 5552 18380 5816 18408
rect 3694 18340 3700 18352
rect 3634 18312 3700 18340
rect 3694 18300 3700 18312
rect 3752 18340 3758 18352
rect 4062 18340 4068 18352
rect 3752 18312 4068 18340
rect 3752 18300 3758 18312
rect 4062 18300 4068 18312
rect 4120 18300 4126 18352
rect 4617 18343 4675 18349
rect 4617 18340 4629 18343
rect 4172 18312 4629 18340
rect 4172 18281 4200 18312
rect 4617 18309 4629 18312
rect 4663 18309 4675 18343
rect 5552 18340 5580 18380
rect 5810 18368 5816 18380
rect 5868 18368 5874 18420
rect 7558 18368 7564 18420
rect 7616 18368 7622 18420
rect 8205 18411 8263 18417
rect 8205 18408 8217 18411
rect 8128 18380 8217 18408
rect 4617 18303 4675 18309
rect 5000 18312 5580 18340
rect 4157 18275 4215 18281
rect 4157 18241 4169 18275
rect 4203 18241 4215 18275
rect 4157 18235 4215 18241
rect 4249 18275 4307 18281
rect 4249 18241 4261 18275
rect 4295 18272 4307 18275
rect 4295 18244 4476 18272
rect 4295 18241 4307 18244
rect 4249 18235 4307 18241
rect 2133 18207 2191 18213
rect 2133 18173 2145 18207
rect 2179 18173 2191 18207
rect 2133 18167 2191 18173
rect 2409 18207 2467 18213
rect 2409 18173 2421 18207
rect 2455 18204 2467 18207
rect 3973 18207 4031 18213
rect 3973 18204 3985 18207
rect 2455 18176 3985 18204
rect 2455 18173 2467 18176
rect 2409 18167 2467 18173
rect 3973 18173 3985 18176
rect 4019 18173 4031 18207
rect 4448 18204 4476 18244
rect 4522 18232 4528 18284
rect 4580 18232 4586 18284
rect 4798 18232 4804 18284
rect 4856 18232 4862 18284
rect 5000 18281 5028 18312
rect 4985 18275 5043 18281
rect 4985 18241 4997 18275
rect 5031 18241 5043 18275
rect 4985 18235 5043 18241
rect 5077 18275 5135 18281
rect 5077 18241 5089 18275
rect 5123 18272 5135 18275
rect 5258 18272 5264 18284
rect 5123 18244 5264 18272
rect 5123 18241 5135 18244
rect 5077 18235 5135 18241
rect 5258 18232 5264 18244
rect 5316 18232 5322 18284
rect 5442 18232 5448 18284
rect 5500 18272 5506 18284
rect 5537 18275 5595 18281
rect 5537 18272 5549 18275
rect 5500 18244 5549 18272
rect 5500 18232 5506 18244
rect 5537 18241 5549 18244
rect 5583 18241 5595 18275
rect 5537 18235 5595 18241
rect 5813 18275 5871 18281
rect 5813 18241 5825 18275
rect 5859 18272 5871 18275
rect 5902 18272 5908 18284
rect 5859 18244 5908 18272
rect 5859 18241 5871 18244
rect 5813 18235 5871 18241
rect 5902 18232 5908 18244
rect 5960 18232 5966 18284
rect 7742 18232 7748 18284
rect 7800 18232 7806 18284
rect 8128 18281 8156 18380
rect 8205 18377 8217 18380
rect 8251 18377 8263 18411
rect 8205 18371 8263 18377
rect 10873 18411 10931 18417
rect 10873 18377 10885 18411
rect 10919 18408 10931 18411
rect 14274 18408 14280 18420
rect 10919 18380 14280 18408
rect 10919 18377 10931 18380
rect 10873 18371 10931 18377
rect 14274 18368 14280 18380
rect 14332 18368 14338 18420
rect 15378 18368 15384 18420
rect 15436 18408 15442 18420
rect 15749 18411 15807 18417
rect 15749 18408 15761 18411
rect 15436 18380 15761 18408
rect 15436 18368 15442 18380
rect 15749 18377 15761 18380
rect 15795 18377 15807 18411
rect 15749 18371 15807 18377
rect 16117 18411 16175 18417
rect 16117 18377 16129 18411
rect 16163 18408 16175 18411
rect 16942 18408 16948 18420
rect 16163 18380 16948 18408
rect 16163 18377 16175 18380
rect 16117 18371 16175 18377
rect 16942 18368 16948 18380
rect 17000 18368 17006 18420
rect 17144 18380 18184 18408
rect 11330 18340 11336 18352
rect 8220 18312 8984 18340
rect 10442 18312 11336 18340
rect 8220 18284 8248 18312
rect 7837 18275 7895 18281
rect 7837 18241 7849 18275
rect 7883 18241 7895 18275
rect 7837 18235 7895 18241
rect 7929 18275 7987 18281
rect 7929 18241 7941 18275
rect 7975 18272 7987 18275
rect 8113 18275 8171 18281
rect 7975 18244 8064 18272
rect 7975 18241 7987 18244
rect 7929 18235 7987 18241
rect 4614 18204 4620 18216
rect 4448 18176 4620 18204
rect 3973 18167 4031 18173
rect 1854 18028 1860 18080
rect 1912 18068 1918 18080
rect 2148 18068 2176 18167
rect 4614 18164 4620 18176
rect 4672 18164 4678 18216
rect 4890 18164 4896 18216
rect 4948 18204 4954 18216
rect 5169 18207 5227 18213
rect 5169 18204 5181 18207
rect 4948 18176 5181 18204
rect 4948 18164 4954 18176
rect 5169 18173 5181 18176
rect 5215 18204 5227 18207
rect 5629 18207 5687 18213
rect 5629 18204 5641 18207
rect 5215 18176 5641 18204
rect 5215 18173 5227 18176
rect 5169 18167 5227 18173
rect 4154 18096 4160 18148
rect 4212 18136 4218 18148
rect 4430 18136 4436 18148
rect 4212 18108 4436 18136
rect 4212 18096 4218 18108
rect 4430 18096 4436 18108
rect 4488 18136 4494 18148
rect 4798 18136 4804 18148
rect 4488 18108 4804 18136
rect 4488 18096 4494 18108
rect 4798 18096 4804 18108
rect 4856 18096 4862 18148
rect 3602 18068 3608 18080
rect 1912 18040 3608 18068
rect 1912 18028 1918 18040
rect 3602 18028 3608 18040
rect 3660 18028 3666 18080
rect 5258 18028 5264 18080
rect 5316 18028 5322 18080
rect 5350 18028 5356 18080
rect 5408 18028 5414 18080
rect 5460 18068 5488 18176
rect 5629 18173 5641 18176
rect 5675 18173 5687 18207
rect 7852 18204 7880 18235
rect 7852 18176 7972 18204
rect 5629 18167 5687 18173
rect 5644 18136 5672 18167
rect 5810 18136 5816 18148
rect 5644 18108 5816 18136
rect 5810 18096 5816 18108
rect 5868 18096 5874 18148
rect 5534 18068 5540 18080
rect 5460 18040 5540 18068
rect 5534 18028 5540 18040
rect 5592 18028 5598 18080
rect 5626 18028 5632 18080
rect 5684 18028 5690 18080
rect 5997 18071 6055 18077
rect 5997 18037 6009 18071
rect 6043 18068 6055 18071
rect 6638 18068 6644 18080
rect 6043 18040 6644 18068
rect 6043 18037 6055 18040
rect 5997 18031 6055 18037
rect 6638 18028 6644 18040
rect 6696 18028 6702 18080
rect 7944 18068 7972 18176
rect 8036 18136 8064 18244
rect 8113 18241 8125 18275
rect 8159 18241 8171 18275
rect 8113 18235 8171 18241
rect 8202 18232 8208 18284
rect 8260 18232 8266 18284
rect 8481 18275 8539 18281
rect 8481 18241 8493 18275
rect 8527 18272 8539 18275
rect 8662 18272 8668 18284
rect 8527 18244 8668 18272
rect 8527 18241 8539 18244
rect 8481 18235 8539 18241
rect 8662 18232 8668 18244
rect 8720 18232 8726 18284
rect 8956 18281 8984 18312
rect 11330 18300 11336 18312
rect 11388 18300 11394 18352
rect 12802 18300 12808 18352
rect 12860 18340 12866 18352
rect 12860 18312 14582 18340
rect 12860 18300 12866 18312
rect 15838 18300 15844 18352
rect 15896 18340 15902 18352
rect 17144 18349 17172 18380
rect 17129 18343 17187 18349
rect 17129 18340 17141 18343
rect 15896 18312 17141 18340
rect 15896 18300 15902 18312
rect 17129 18309 17141 18312
rect 17175 18309 17187 18343
rect 17129 18303 17187 18309
rect 17310 18300 17316 18352
rect 17368 18349 17374 18352
rect 17368 18343 17387 18349
rect 17375 18309 17387 18343
rect 18156 18340 18184 18380
rect 19150 18368 19156 18420
rect 19208 18408 19214 18420
rect 20549 18411 20607 18417
rect 20549 18408 20561 18411
rect 19208 18380 20561 18408
rect 19208 18368 19214 18380
rect 20549 18377 20561 18380
rect 20595 18377 20607 18411
rect 20549 18371 20607 18377
rect 20717 18411 20775 18417
rect 20717 18377 20729 18411
rect 20763 18377 20775 18411
rect 20717 18371 20775 18377
rect 20346 18340 20352 18352
rect 18156 18312 20352 18340
rect 17368 18303 17387 18309
rect 17368 18300 17374 18303
rect 20346 18300 20352 18312
rect 20404 18300 20410 18352
rect 8941 18275 8999 18281
rect 8941 18241 8953 18275
rect 8987 18241 8999 18275
rect 8941 18235 8999 18241
rect 10781 18275 10839 18281
rect 10781 18241 10793 18275
rect 10827 18272 10839 18275
rect 10870 18272 10876 18284
rect 10827 18244 10876 18272
rect 10827 18241 10839 18244
rect 10781 18235 10839 18241
rect 10870 18232 10876 18244
rect 10928 18232 10934 18284
rect 10962 18232 10968 18284
rect 11020 18232 11026 18284
rect 11422 18232 11428 18284
rect 11480 18272 11486 18284
rect 11517 18275 11575 18281
rect 11517 18272 11529 18275
rect 11480 18244 11529 18272
rect 11480 18232 11486 18244
rect 11517 18241 11529 18244
rect 11563 18241 11575 18275
rect 11517 18235 11575 18241
rect 11885 18275 11943 18281
rect 11885 18241 11897 18275
rect 11931 18241 11943 18275
rect 11885 18235 11943 18241
rect 12345 18275 12403 18281
rect 12345 18241 12357 18275
rect 12391 18272 12403 18275
rect 12618 18272 12624 18284
rect 12391 18244 12624 18272
rect 12391 18241 12403 18244
rect 12345 18235 12403 18241
rect 8294 18164 8300 18216
rect 8352 18164 8358 18216
rect 8386 18164 8392 18216
rect 8444 18164 8450 18216
rect 8757 18207 8815 18213
rect 8757 18173 8769 18207
rect 8803 18173 8815 18207
rect 8757 18167 8815 18173
rect 8312 18136 8340 18164
rect 8570 18136 8576 18148
rect 8036 18108 8576 18136
rect 8570 18096 8576 18108
rect 8628 18096 8634 18148
rect 8294 18068 8300 18080
rect 7944 18040 8300 18068
rect 8294 18028 8300 18040
rect 8352 18028 8358 18080
rect 8772 18068 8800 18167
rect 8846 18164 8852 18216
rect 8904 18164 8910 18216
rect 9214 18164 9220 18216
rect 9272 18164 9278 18216
rect 10686 18164 10692 18216
rect 10744 18204 10750 18216
rect 11900 18204 11928 18235
rect 12618 18232 12624 18244
rect 12676 18232 12682 18284
rect 15930 18232 15936 18284
rect 15988 18232 15994 18284
rect 16206 18232 16212 18284
rect 16264 18272 16270 18284
rect 17865 18275 17923 18281
rect 17865 18272 17877 18275
rect 16264 18244 17877 18272
rect 16264 18232 16270 18244
rect 17865 18241 17877 18244
rect 17911 18241 17923 18275
rect 17865 18235 17923 18241
rect 18138 18232 18144 18284
rect 18196 18232 18202 18284
rect 19058 18232 19064 18284
rect 19116 18232 19122 18284
rect 19337 18275 19395 18281
rect 19337 18241 19349 18275
rect 19383 18241 19395 18275
rect 20732 18272 20760 18371
rect 20806 18368 20812 18420
rect 20864 18368 20870 18420
rect 21177 18411 21235 18417
rect 21177 18377 21189 18411
rect 21223 18408 21235 18411
rect 22002 18408 22008 18420
rect 21223 18380 22008 18408
rect 21223 18377 21235 18380
rect 21177 18371 21235 18377
rect 22002 18368 22008 18380
rect 22060 18368 22066 18420
rect 24486 18368 24492 18420
rect 24544 18368 24550 18420
rect 24670 18408 24676 18420
rect 24596 18380 24676 18408
rect 22281 18343 22339 18349
rect 22281 18309 22293 18343
rect 22327 18340 22339 18343
rect 22741 18343 22799 18349
rect 22741 18340 22753 18343
rect 22327 18312 22753 18340
rect 22327 18309 22339 18312
rect 22281 18303 22339 18309
rect 22741 18309 22753 18312
rect 22787 18309 22799 18343
rect 24596 18340 24624 18380
rect 24670 18368 24676 18380
rect 24728 18368 24734 18420
rect 25774 18368 25780 18420
rect 25832 18368 25838 18420
rect 22741 18303 22799 18309
rect 24136 18312 24624 18340
rect 24136 18284 24164 18312
rect 24854 18300 24860 18352
rect 24912 18340 24918 18352
rect 24912 18312 25544 18340
rect 24912 18300 24918 18312
rect 20993 18275 21051 18281
rect 20993 18272 21005 18275
rect 20732 18244 21005 18272
rect 19337 18235 19395 18241
rect 20993 18241 21005 18244
rect 21039 18241 21051 18275
rect 20993 18235 21051 18241
rect 21269 18275 21327 18281
rect 21269 18241 21281 18275
rect 21315 18241 21327 18275
rect 21269 18235 21327 18241
rect 10744 18176 11928 18204
rect 10744 18164 10750 18176
rect 11900 18136 11928 18176
rect 13817 18207 13875 18213
rect 13817 18173 13829 18207
rect 13863 18173 13875 18207
rect 13817 18167 13875 18173
rect 12161 18139 12219 18145
rect 12161 18136 12173 18139
rect 11900 18108 12173 18136
rect 12161 18105 12173 18108
rect 12207 18105 12219 18139
rect 12161 18099 12219 18105
rect 9766 18068 9772 18080
rect 8772 18040 9772 18068
rect 9766 18028 9772 18040
rect 9824 18068 9830 18080
rect 10594 18068 10600 18080
rect 9824 18040 10600 18068
rect 9824 18028 9830 18040
rect 10594 18028 10600 18040
rect 10652 18068 10658 18080
rect 10689 18071 10747 18077
rect 10689 18068 10701 18071
rect 10652 18040 10701 18068
rect 10652 18028 10658 18040
rect 10689 18037 10701 18040
rect 10735 18037 10747 18071
rect 13832 18068 13860 18167
rect 14090 18164 14096 18216
rect 14148 18164 14154 18216
rect 15562 18164 15568 18216
rect 15620 18164 15626 18216
rect 15672 18176 17632 18204
rect 14182 18068 14188 18080
rect 13832 18040 14188 18068
rect 10689 18031 10747 18037
rect 14182 18028 14188 18040
rect 14240 18028 14246 18080
rect 14274 18028 14280 18080
rect 14332 18068 14338 18080
rect 15672 18068 15700 18176
rect 17604 18136 17632 18176
rect 19352 18136 19380 18235
rect 21284 18204 21312 18235
rect 22094 18232 22100 18284
rect 22152 18232 22158 18284
rect 22370 18232 22376 18284
rect 22428 18272 22434 18284
rect 23661 18275 23719 18281
rect 22428 18244 22784 18272
rect 22428 18232 22434 18244
rect 22756 18216 22784 18244
rect 23661 18241 23673 18275
rect 23707 18272 23719 18275
rect 24118 18272 24124 18284
rect 23707 18244 24124 18272
rect 23707 18241 23719 18244
rect 23661 18235 23719 18241
rect 24118 18232 24124 18244
rect 24176 18232 24182 18284
rect 25130 18232 25136 18284
rect 25188 18232 25194 18284
rect 25314 18232 25320 18284
rect 25372 18232 25378 18284
rect 25516 18281 25544 18312
rect 25409 18275 25467 18281
rect 25409 18241 25421 18275
rect 25455 18241 25467 18275
rect 25409 18235 25467 18241
rect 25501 18275 25559 18281
rect 25501 18241 25513 18275
rect 25547 18272 25559 18275
rect 25590 18272 25596 18284
rect 25547 18244 25596 18272
rect 25547 18241 25559 18244
rect 25501 18235 25559 18241
rect 17604 18108 19380 18136
rect 19536 18176 21312 18204
rect 19536 18080 19564 18176
rect 22738 18164 22744 18216
rect 22796 18164 22802 18216
rect 23198 18164 23204 18216
rect 23256 18204 23262 18216
rect 23293 18207 23351 18213
rect 23293 18204 23305 18207
rect 23256 18176 23305 18204
rect 23256 18164 23262 18176
rect 23293 18173 23305 18176
rect 23339 18204 23351 18207
rect 23569 18207 23627 18213
rect 23569 18204 23581 18207
rect 23339 18176 23581 18204
rect 23339 18173 23351 18176
rect 23293 18167 23351 18173
rect 23569 18173 23581 18176
rect 23615 18173 23627 18207
rect 23569 18167 23627 18173
rect 24026 18164 24032 18216
rect 24084 18164 24090 18216
rect 25424 18204 25452 18235
rect 25590 18232 25596 18244
rect 25648 18232 25654 18284
rect 25866 18204 25872 18216
rect 25424 18176 25872 18204
rect 25866 18164 25872 18176
rect 25924 18164 25930 18216
rect 14332 18040 15700 18068
rect 17313 18071 17371 18077
rect 14332 18028 14338 18040
rect 17313 18037 17325 18071
rect 17359 18068 17371 18071
rect 17402 18068 17408 18080
rect 17359 18040 17408 18068
rect 17359 18037 17371 18040
rect 17313 18031 17371 18037
rect 17402 18028 17408 18040
rect 17460 18028 17466 18080
rect 17494 18028 17500 18080
rect 17552 18028 17558 18080
rect 18877 18071 18935 18077
rect 18877 18037 18889 18071
rect 18923 18068 18935 18071
rect 19150 18068 19156 18080
rect 18923 18040 19156 18068
rect 18923 18037 18935 18040
rect 18877 18031 18935 18037
rect 19150 18028 19156 18040
rect 19208 18028 19214 18080
rect 19518 18028 19524 18080
rect 19576 18028 19582 18080
rect 20530 18028 20536 18080
rect 20588 18028 20594 18080
rect 21726 18028 21732 18080
rect 21784 18068 21790 18080
rect 21913 18071 21971 18077
rect 21913 18068 21925 18071
rect 21784 18040 21925 18068
rect 21784 18028 21790 18040
rect 21913 18037 21925 18040
rect 21959 18037 21971 18071
rect 21913 18031 21971 18037
rect 24673 18071 24731 18077
rect 24673 18037 24685 18071
rect 24719 18068 24731 18071
rect 25038 18068 25044 18080
rect 24719 18040 25044 18068
rect 24719 18037 24731 18040
rect 24673 18031 24731 18037
rect 25038 18028 25044 18040
rect 25096 18028 25102 18080
rect 1104 17978 28704 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 28704 17978
rect 1104 17904 28704 17926
rect 4062 17824 4068 17876
rect 4120 17864 4126 17876
rect 4157 17867 4215 17873
rect 4157 17864 4169 17867
rect 4120 17836 4169 17864
rect 4120 17824 4126 17836
rect 4157 17833 4169 17836
rect 4203 17833 4215 17867
rect 4157 17827 4215 17833
rect 4341 17867 4399 17873
rect 4341 17833 4353 17867
rect 4387 17864 4399 17867
rect 4614 17864 4620 17876
rect 4387 17836 4620 17864
rect 4387 17833 4399 17836
rect 4341 17827 4399 17833
rect 4614 17824 4620 17836
rect 4672 17824 4678 17876
rect 5350 17824 5356 17876
rect 5408 17824 5414 17876
rect 5442 17824 5448 17876
rect 5500 17864 5506 17876
rect 5629 17867 5687 17873
rect 5629 17864 5641 17867
rect 5500 17836 5641 17864
rect 5500 17824 5506 17836
rect 5629 17833 5641 17836
rect 5675 17833 5687 17867
rect 5629 17827 5687 17833
rect 5994 17824 6000 17876
rect 6052 17824 6058 17876
rect 6914 17824 6920 17876
rect 6972 17864 6978 17876
rect 7101 17867 7159 17873
rect 7101 17864 7113 17867
rect 6972 17836 7113 17864
rect 6972 17824 6978 17836
rect 7101 17833 7113 17836
rect 7147 17833 7159 17867
rect 7101 17827 7159 17833
rect 8386 17824 8392 17876
rect 8444 17864 8450 17876
rect 8481 17867 8539 17873
rect 8481 17864 8493 17867
rect 8444 17836 8493 17864
rect 8444 17824 8450 17836
rect 8481 17833 8493 17836
rect 8527 17833 8539 17867
rect 8481 17827 8539 17833
rect 8662 17824 8668 17876
rect 8720 17864 8726 17876
rect 9401 17867 9459 17873
rect 9401 17864 9413 17867
rect 8720 17836 9413 17864
rect 8720 17824 8726 17836
rect 9401 17833 9413 17836
rect 9447 17833 9459 17867
rect 9858 17864 9864 17876
rect 9401 17827 9459 17833
rect 9600 17836 9864 17864
rect 4893 17799 4951 17805
rect 4893 17796 4905 17799
rect 3988 17768 4905 17796
rect 1854 17688 1860 17740
rect 1912 17688 1918 17740
rect 2133 17731 2191 17737
rect 2133 17697 2145 17731
rect 2179 17728 2191 17731
rect 3789 17731 3847 17737
rect 3789 17728 3801 17731
rect 2179 17700 3801 17728
rect 2179 17697 2191 17700
rect 2133 17691 2191 17697
rect 3789 17697 3801 17700
rect 3835 17697 3847 17731
rect 3789 17691 3847 17697
rect 3694 17660 3700 17672
rect 3266 17632 3700 17660
rect 3694 17620 3700 17632
rect 3752 17620 3758 17672
rect 3988 17669 4016 17768
rect 4893 17765 4905 17768
rect 4939 17765 4951 17799
rect 5368 17796 5396 17824
rect 9600 17796 9628 17836
rect 9858 17824 9864 17836
rect 9916 17824 9922 17876
rect 15562 17824 15568 17876
rect 15620 17864 15626 17876
rect 15657 17867 15715 17873
rect 15657 17864 15669 17867
rect 15620 17836 15669 17864
rect 15620 17824 15626 17836
rect 15657 17833 15669 17836
rect 15703 17833 15715 17867
rect 15657 17827 15715 17833
rect 15841 17867 15899 17873
rect 15841 17833 15853 17867
rect 15887 17864 15899 17867
rect 15930 17864 15936 17876
rect 15887 17836 15936 17864
rect 15887 17833 15899 17836
rect 15841 17827 15899 17833
rect 15930 17824 15936 17836
rect 15988 17824 15994 17876
rect 18598 17824 18604 17876
rect 18656 17864 18662 17876
rect 18877 17867 18935 17873
rect 18877 17864 18889 17867
rect 18656 17836 18889 17864
rect 18656 17824 18662 17836
rect 18877 17833 18889 17836
rect 18923 17833 18935 17867
rect 18877 17827 18935 17833
rect 20530 17824 20536 17876
rect 20588 17864 20594 17876
rect 20993 17867 21051 17873
rect 20993 17864 21005 17867
rect 20588 17836 21005 17864
rect 20588 17824 20594 17836
rect 20993 17833 21005 17836
rect 21039 17833 21051 17867
rect 20993 17827 21051 17833
rect 22094 17824 22100 17876
rect 22152 17864 22158 17876
rect 23293 17867 23351 17873
rect 23293 17864 23305 17867
rect 22152 17836 23305 17864
rect 22152 17824 22158 17836
rect 23293 17833 23305 17836
rect 23339 17833 23351 17867
rect 23293 17827 23351 17833
rect 23382 17824 23388 17876
rect 23440 17864 23446 17876
rect 23477 17867 23535 17873
rect 23477 17864 23489 17867
rect 23440 17836 23489 17864
rect 23440 17824 23446 17836
rect 23477 17833 23489 17836
rect 23523 17833 23535 17867
rect 23477 17827 23535 17833
rect 24857 17867 24915 17873
rect 24857 17833 24869 17867
rect 24903 17864 24915 17867
rect 25130 17864 25136 17876
rect 24903 17836 25136 17864
rect 24903 17833 24915 17836
rect 24857 17827 24915 17833
rect 25130 17824 25136 17836
rect 25188 17824 25194 17876
rect 25314 17824 25320 17876
rect 25372 17824 25378 17876
rect 5368 17768 5672 17796
rect 4893 17759 4951 17765
rect 4982 17688 4988 17740
rect 5040 17728 5046 17740
rect 5040 17700 5304 17728
rect 5040 17688 5046 17700
rect 3973 17663 4031 17669
rect 3973 17629 3985 17663
rect 4019 17629 4031 17663
rect 3973 17623 4031 17629
rect 4249 17663 4307 17669
rect 4249 17629 4261 17663
rect 4295 17629 4307 17663
rect 4249 17623 4307 17629
rect 4525 17663 4583 17669
rect 4525 17629 4537 17663
rect 4571 17660 4583 17663
rect 4614 17660 4620 17672
rect 4571 17632 4620 17660
rect 4571 17629 4583 17632
rect 4525 17623 4583 17629
rect 4264 17592 4292 17623
rect 4614 17620 4620 17632
rect 4672 17620 4678 17672
rect 4706 17620 4712 17672
rect 4764 17620 4770 17672
rect 4801 17663 4859 17669
rect 4801 17629 4813 17663
rect 4847 17660 4859 17663
rect 4890 17660 4896 17672
rect 4847 17632 4896 17660
rect 4847 17629 4859 17632
rect 4801 17623 4859 17629
rect 4816 17592 4844 17623
rect 4890 17620 4896 17632
rect 4948 17620 4954 17672
rect 5074 17669 5080 17672
rect 5072 17623 5080 17669
rect 5132 17660 5138 17672
rect 5276 17660 5304 17700
rect 5444 17663 5502 17669
rect 5444 17660 5456 17663
rect 5132 17632 5172 17660
rect 5276 17632 5456 17660
rect 5074 17620 5080 17623
rect 5132 17620 5138 17632
rect 5444 17629 5456 17632
rect 5490 17629 5502 17663
rect 5444 17623 5502 17629
rect 3620 17564 4844 17592
rect 5169 17595 5227 17601
rect 3620 17533 3648 17564
rect 5169 17561 5181 17595
rect 5215 17561 5227 17595
rect 5169 17555 5227 17561
rect 3605 17527 3663 17533
rect 3605 17493 3617 17527
rect 3651 17493 3663 17527
rect 3605 17487 3663 17493
rect 4706 17484 4712 17536
rect 4764 17524 4770 17536
rect 5074 17524 5080 17536
rect 4764 17496 5080 17524
rect 4764 17484 4770 17496
rect 5074 17484 5080 17496
rect 5132 17484 5138 17536
rect 5184 17524 5212 17555
rect 5258 17552 5264 17604
rect 5316 17552 5322 17604
rect 5460 17592 5488 17623
rect 5534 17620 5540 17672
rect 5592 17620 5598 17672
rect 5644 17669 5672 17768
rect 6380 17768 9628 17796
rect 5629 17663 5687 17669
rect 5629 17629 5641 17663
rect 5675 17660 5687 17663
rect 5718 17660 5724 17672
rect 5675 17632 5724 17660
rect 5675 17629 5687 17632
rect 5629 17623 5687 17629
rect 5718 17620 5724 17632
rect 5776 17620 5782 17672
rect 5810 17620 5816 17672
rect 5868 17620 5874 17672
rect 6178 17592 6184 17604
rect 5460 17564 6184 17592
rect 6178 17552 6184 17564
rect 6236 17552 6242 17604
rect 6380 17524 6408 17768
rect 9674 17756 9680 17808
rect 9732 17796 9738 17808
rect 24213 17799 24271 17805
rect 9732 17768 9904 17796
rect 9732 17756 9738 17768
rect 9306 17728 9312 17740
rect 8496 17700 9312 17728
rect 6546 17620 6552 17672
rect 6604 17620 6610 17672
rect 6638 17620 6644 17672
rect 6696 17620 6702 17672
rect 6822 17620 6828 17672
rect 6880 17620 6886 17672
rect 6917 17663 6975 17669
rect 6917 17629 6929 17663
rect 6963 17660 6975 17663
rect 7006 17660 7012 17672
rect 6963 17632 7012 17660
rect 6963 17629 6975 17632
rect 6917 17623 6975 17629
rect 7006 17620 7012 17632
rect 7064 17620 7070 17672
rect 8386 17552 8392 17604
rect 8444 17592 8450 17604
rect 8496 17601 8524 17700
rect 9306 17688 9312 17700
rect 9364 17728 9370 17740
rect 9769 17731 9827 17737
rect 9769 17728 9781 17731
rect 9364 17700 9781 17728
rect 9364 17688 9370 17700
rect 9769 17697 9781 17700
rect 9815 17697 9827 17731
rect 9769 17691 9827 17697
rect 8757 17663 8815 17669
rect 8757 17629 8769 17663
rect 8803 17660 8815 17663
rect 9122 17660 9128 17672
rect 8803 17632 9128 17660
rect 8803 17629 8815 17632
rect 8757 17623 8815 17629
rect 9122 17620 9128 17632
rect 9180 17660 9186 17672
rect 9876 17669 9904 17768
rect 24213 17765 24225 17799
rect 24259 17796 24271 17799
rect 25332 17796 25360 17824
rect 24259 17768 25360 17796
rect 24259 17765 24271 17768
rect 24213 17759 24271 17765
rect 10594 17688 10600 17740
rect 10652 17728 10658 17740
rect 11149 17731 11207 17737
rect 11149 17728 11161 17731
rect 10652 17700 11161 17728
rect 10652 17688 10658 17700
rect 11149 17697 11161 17700
rect 11195 17697 11207 17731
rect 11149 17691 11207 17697
rect 16853 17731 16911 17737
rect 16853 17697 16865 17731
rect 16899 17728 16911 17731
rect 17862 17728 17868 17740
rect 16899 17700 17868 17728
rect 16899 17697 16911 17700
rect 16853 17691 16911 17697
rect 17862 17688 17868 17700
rect 17920 17728 17926 17740
rect 19245 17731 19303 17737
rect 19245 17728 19257 17731
rect 17920 17700 19257 17728
rect 17920 17688 17926 17700
rect 19245 17697 19257 17700
rect 19291 17728 19303 17731
rect 20530 17728 20536 17740
rect 19291 17700 20536 17728
rect 19291 17697 19303 17700
rect 19245 17691 19303 17697
rect 20530 17688 20536 17700
rect 20588 17728 20594 17740
rect 21453 17731 21511 17737
rect 21453 17728 21465 17731
rect 20588 17700 21465 17728
rect 20588 17688 20594 17700
rect 21453 17697 21465 17700
rect 21499 17697 21511 17731
rect 21453 17691 21511 17697
rect 21726 17688 21732 17740
rect 21784 17688 21790 17740
rect 22094 17688 22100 17740
rect 22152 17728 22158 17740
rect 22152 17700 23704 17728
rect 22152 17688 22158 17700
rect 9585 17663 9643 17669
rect 9585 17660 9597 17663
rect 9180 17632 9597 17660
rect 9180 17620 9186 17632
rect 9585 17629 9597 17632
rect 9631 17629 9643 17663
rect 9585 17623 9643 17629
rect 9677 17663 9735 17669
rect 9677 17629 9689 17663
rect 9723 17629 9735 17663
rect 9677 17623 9735 17629
rect 9861 17663 9919 17669
rect 9861 17629 9873 17663
rect 9907 17660 9919 17663
rect 10870 17660 10876 17672
rect 9907 17632 10876 17660
rect 9907 17629 9919 17632
rect 9861 17623 9919 17629
rect 8481 17595 8539 17601
rect 8481 17592 8493 17595
rect 8444 17564 8493 17592
rect 8444 17552 8450 17564
rect 8481 17561 8493 17564
rect 8527 17561 8539 17595
rect 8481 17555 8539 17561
rect 8665 17595 8723 17601
rect 8665 17561 8677 17595
rect 8711 17592 8723 17595
rect 9692 17592 9720 17623
rect 10870 17620 10876 17632
rect 10928 17620 10934 17672
rect 10965 17663 11023 17669
rect 10965 17629 10977 17663
rect 11011 17629 11023 17663
rect 10965 17623 11023 17629
rect 10134 17592 10140 17604
rect 8711 17564 10140 17592
rect 8711 17561 8723 17564
rect 8665 17555 8723 17561
rect 10134 17552 10140 17564
rect 10192 17552 10198 17604
rect 10980 17592 11008 17623
rect 11238 17620 11244 17672
rect 11296 17620 11302 17672
rect 11422 17620 11428 17672
rect 11480 17620 11486 17672
rect 23382 17660 23388 17672
rect 22862 17632 23388 17660
rect 23382 17620 23388 17632
rect 23440 17620 23446 17672
rect 11054 17592 11060 17604
rect 10980 17564 11060 17592
rect 11054 17552 11060 17564
rect 11112 17592 11118 17604
rect 11974 17592 11980 17604
rect 11112 17564 11980 17592
rect 11112 17552 11118 17564
rect 11974 17552 11980 17564
rect 12032 17552 12038 17604
rect 15473 17595 15531 17601
rect 15473 17561 15485 17595
rect 15519 17592 15531 17595
rect 15838 17592 15844 17604
rect 15519 17564 15844 17592
rect 15519 17561 15531 17564
rect 15473 17555 15531 17561
rect 15838 17552 15844 17564
rect 15896 17552 15902 17604
rect 17129 17595 17187 17601
rect 17129 17561 17141 17595
rect 17175 17592 17187 17595
rect 17402 17592 17408 17604
rect 17175 17564 17408 17592
rect 17175 17561 17187 17564
rect 17129 17555 17187 17561
rect 17402 17552 17408 17564
rect 17460 17552 17466 17604
rect 18354 17564 18460 17592
rect 5184 17496 6408 17524
rect 10042 17484 10048 17536
rect 10100 17484 10106 17536
rect 10226 17484 10232 17536
rect 10284 17524 10290 17536
rect 10781 17527 10839 17533
rect 10781 17524 10793 17527
rect 10284 17496 10793 17524
rect 10284 17484 10290 17496
rect 10781 17493 10793 17496
rect 10827 17493 10839 17527
rect 10781 17487 10839 17493
rect 11333 17527 11391 17533
rect 11333 17493 11345 17527
rect 11379 17524 11391 17527
rect 12342 17524 12348 17536
rect 11379 17496 12348 17524
rect 11379 17493 11391 17496
rect 11333 17487 11391 17493
rect 12342 17484 12348 17496
rect 12400 17484 12406 17536
rect 15562 17484 15568 17536
rect 15620 17524 15626 17536
rect 15673 17527 15731 17533
rect 15673 17524 15685 17527
rect 15620 17496 15685 17524
rect 15620 17484 15626 17496
rect 15673 17493 15685 17496
rect 15719 17493 15731 17527
rect 15673 17487 15731 17493
rect 16482 17484 16488 17536
rect 16540 17524 16546 17536
rect 18432 17524 18460 17564
rect 18506 17552 18512 17604
rect 18564 17592 18570 17604
rect 18693 17595 18751 17601
rect 18693 17592 18705 17595
rect 18564 17564 18705 17592
rect 18564 17552 18570 17564
rect 18693 17561 18705 17564
rect 18739 17561 18751 17595
rect 18693 17555 18751 17561
rect 18909 17595 18967 17601
rect 18909 17561 18921 17595
rect 18955 17592 18967 17595
rect 19150 17592 19156 17604
rect 18955 17564 19156 17592
rect 18955 17561 18967 17564
rect 18909 17555 18967 17561
rect 19150 17552 19156 17564
rect 19208 17552 19214 17604
rect 19426 17552 19432 17604
rect 19484 17592 19490 17604
rect 19521 17595 19579 17601
rect 19521 17592 19533 17595
rect 19484 17564 19533 17592
rect 19484 17552 19490 17564
rect 19521 17561 19533 17564
rect 19567 17561 19579 17595
rect 21174 17592 21180 17604
rect 20746 17564 21180 17592
rect 19521 17555 19579 17561
rect 21174 17552 21180 17564
rect 21232 17552 21238 17604
rect 23676 17601 23704 17700
rect 23952 17700 24440 17728
rect 23952 17672 23980 17700
rect 23934 17620 23940 17672
rect 23992 17620 23998 17672
rect 24118 17620 24124 17672
rect 24176 17620 24182 17672
rect 24412 17669 24440 17700
rect 25314 17688 25320 17740
rect 25372 17728 25378 17740
rect 26142 17728 26148 17740
rect 25372 17700 26148 17728
rect 25372 17688 25378 17700
rect 26142 17688 26148 17700
rect 26200 17728 26206 17740
rect 26513 17731 26571 17737
rect 26513 17728 26525 17731
rect 26200 17700 26525 17728
rect 26200 17688 26206 17700
rect 26513 17697 26525 17700
rect 26559 17697 26571 17731
rect 26513 17691 26571 17697
rect 24213 17663 24271 17669
rect 24213 17629 24225 17663
rect 24259 17629 24271 17663
rect 24213 17623 24271 17629
rect 24397 17663 24455 17669
rect 24397 17629 24409 17663
rect 24443 17629 24455 17663
rect 24397 17623 24455 17629
rect 23661 17595 23719 17601
rect 23661 17561 23673 17595
rect 23707 17561 23719 17595
rect 24228 17592 24256 17623
rect 24670 17620 24676 17672
rect 24728 17620 24734 17672
rect 25130 17620 25136 17672
rect 25188 17620 25194 17672
rect 25225 17663 25283 17669
rect 25225 17629 25237 17663
rect 25271 17660 25283 17663
rect 25501 17663 25559 17669
rect 25501 17660 25513 17663
rect 25271 17632 25513 17660
rect 25271 17629 25283 17632
rect 25225 17623 25283 17629
rect 25501 17629 25513 17632
rect 25547 17629 25559 17663
rect 25501 17623 25559 17629
rect 24489 17595 24547 17601
rect 24489 17592 24501 17595
rect 24228 17564 24501 17592
rect 23661 17555 23719 17561
rect 24489 17561 24501 17564
rect 24535 17592 24547 17595
rect 25240 17592 25268 17623
rect 25590 17620 25596 17672
rect 25648 17620 25654 17672
rect 25869 17663 25927 17669
rect 25869 17629 25881 17663
rect 25915 17629 25927 17663
rect 25869 17623 25927 17629
rect 24535 17564 25268 17592
rect 24535 17561 24547 17564
rect 24489 17555 24547 17561
rect 25884 17536 25912 17623
rect 26786 17552 26792 17604
rect 26844 17552 26850 17604
rect 26878 17552 26884 17604
rect 26936 17592 26942 17604
rect 26936 17564 27278 17592
rect 26936 17552 26942 17564
rect 18782 17524 18788 17536
rect 16540 17496 18788 17524
rect 16540 17484 16546 17496
rect 18782 17484 18788 17496
rect 18840 17484 18846 17536
rect 19061 17527 19119 17533
rect 19061 17493 19073 17527
rect 19107 17524 19119 17527
rect 19242 17524 19248 17536
rect 19107 17496 19248 17524
rect 19107 17493 19119 17496
rect 19061 17487 19119 17493
rect 19242 17484 19248 17496
rect 19300 17484 19306 17536
rect 22370 17484 22376 17536
rect 22428 17524 22434 17536
rect 23198 17524 23204 17536
rect 22428 17496 23204 17524
rect 22428 17484 22434 17496
rect 23198 17484 23204 17496
rect 23256 17484 23262 17536
rect 23290 17484 23296 17536
rect 23348 17524 23354 17536
rect 23451 17527 23509 17533
rect 23451 17524 23463 17527
rect 23348 17496 23463 17524
rect 23348 17484 23354 17496
rect 23451 17493 23463 17496
rect 23497 17493 23509 17527
rect 23451 17487 23509 17493
rect 25038 17484 25044 17536
rect 25096 17484 25102 17536
rect 25130 17484 25136 17536
rect 25188 17524 25194 17536
rect 25774 17524 25780 17536
rect 25188 17496 25780 17524
rect 25188 17484 25194 17496
rect 25774 17484 25780 17496
rect 25832 17484 25838 17536
rect 25866 17484 25872 17536
rect 25924 17524 25930 17536
rect 28258 17524 28264 17536
rect 25924 17496 28264 17524
rect 25924 17484 25930 17496
rect 28258 17484 28264 17496
rect 28316 17484 28322 17536
rect 1104 17434 28704 17456
rect 1104 17382 4874 17434
rect 4926 17382 4938 17434
rect 4990 17382 5002 17434
rect 5054 17382 5066 17434
rect 5118 17382 5130 17434
rect 5182 17382 28704 17434
rect 1104 17360 28704 17382
rect 5258 17280 5264 17332
rect 5316 17280 5322 17332
rect 5534 17280 5540 17332
rect 5592 17320 5598 17332
rect 8754 17320 8760 17332
rect 5592 17292 8760 17320
rect 5592 17280 5598 17292
rect 8754 17280 8760 17292
rect 8812 17320 8818 17332
rect 8941 17323 8999 17329
rect 8812 17292 8892 17320
rect 8812 17280 8818 17292
rect 5994 17252 6000 17264
rect 5368 17224 6000 17252
rect 5169 17187 5227 17193
rect 5169 17153 5181 17187
rect 5215 17184 5227 17187
rect 5258 17184 5264 17196
rect 5215 17156 5264 17184
rect 5215 17153 5227 17156
rect 5169 17147 5227 17153
rect 5258 17144 5264 17156
rect 5316 17144 5322 17196
rect 5368 17193 5396 17224
rect 5994 17212 6000 17224
rect 6052 17212 6058 17264
rect 6546 17212 6552 17264
rect 6604 17252 6610 17264
rect 8297 17255 8355 17261
rect 8297 17252 8309 17255
rect 6604 17224 8309 17252
rect 6604 17212 6610 17224
rect 5353 17187 5411 17193
rect 5353 17153 5365 17187
rect 5399 17153 5411 17187
rect 5353 17147 5411 17153
rect 5442 17144 5448 17196
rect 5500 17184 5506 17196
rect 6748 17193 6776 17224
rect 8297 17221 8309 17224
rect 8343 17221 8355 17255
rect 8297 17215 8355 17221
rect 8386 17212 8392 17264
rect 8444 17252 8450 17264
rect 8864 17252 8892 17292
rect 8941 17289 8953 17323
rect 8987 17320 8999 17323
rect 9214 17320 9220 17332
rect 8987 17292 9220 17320
rect 8987 17289 8999 17292
rect 8941 17283 8999 17289
rect 9214 17280 9220 17292
rect 9272 17280 9278 17332
rect 10134 17280 10140 17332
rect 10192 17280 10198 17332
rect 17402 17280 17408 17332
rect 17460 17280 17466 17332
rect 18506 17280 18512 17332
rect 18564 17320 18570 17332
rect 18564 17292 22094 17320
rect 18564 17280 18570 17292
rect 10042 17252 10048 17264
rect 8444 17224 8800 17252
rect 8864 17224 9168 17252
rect 8444 17212 8450 17224
rect 5629 17187 5687 17193
rect 5629 17184 5641 17187
rect 5500 17156 5641 17184
rect 5500 17144 5506 17156
rect 5629 17153 5641 17156
rect 5675 17153 5687 17187
rect 5629 17147 5687 17153
rect 6733 17187 6791 17193
rect 6733 17153 6745 17187
rect 6779 17153 6791 17187
rect 6733 17147 6791 17153
rect 6914 17144 6920 17196
rect 6972 17144 6978 17196
rect 7006 17144 7012 17196
rect 7064 17144 7070 17196
rect 8478 17144 8484 17196
rect 8536 17144 8542 17196
rect 8772 17193 8800 17224
rect 9140 17193 9168 17224
rect 9232 17224 10048 17252
rect 9232 17193 9260 17224
rect 10042 17212 10048 17224
rect 10100 17212 10106 17264
rect 11054 17252 11060 17264
rect 10152 17224 11060 17252
rect 8573 17187 8631 17193
rect 8573 17153 8585 17187
rect 8619 17153 8631 17187
rect 8573 17147 8631 17153
rect 8757 17187 8815 17193
rect 8757 17153 8769 17187
rect 8803 17153 8815 17187
rect 8757 17147 8815 17153
rect 8849 17187 8907 17193
rect 8849 17153 8861 17187
rect 8895 17153 8907 17187
rect 8849 17147 8907 17153
rect 9101 17187 9168 17193
rect 9101 17153 9113 17187
rect 9147 17156 9168 17187
rect 9217 17187 9275 17193
rect 9147 17153 9159 17156
rect 9101 17147 9159 17153
rect 9217 17153 9229 17187
rect 9263 17153 9275 17187
rect 9217 17147 9275 17153
rect 5718 17076 5724 17128
rect 5776 17116 5782 17128
rect 6549 17119 6607 17125
rect 6549 17116 6561 17119
rect 5776 17088 6561 17116
rect 5776 17076 5782 17088
rect 6549 17085 6561 17088
rect 6595 17085 6607 17119
rect 6549 17079 6607 17085
rect 5997 17051 6055 17057
rect 5997 17017 6009 17051
rect 6043 17048 6055 17051
rect 6454 17048 6460 17060
rect 6043 17020 6460 17048
rect 6043 17017 6055 17020
rect 5997 17011 6055 17017
rect 6454 17008 6460 17020
rect 6512 17008 6518 17060
rect 8588 16980 8616 17147
rect 8864 17116 8892 17147
rect 9306 17144 9312 17196
rect 9364 17144 9370 17196
rect 9490 17144 9496 17196
rect 9548 17144 9554 17196
rect 9766 17144 9772 17196
rect 9824 17144 9830 17196
rect 9953 17187 10011 17193
rect 9953 17153 9965 17187
rect 9999 17184 10011 17187
rect 10152 17184 10180 17224
rect 11054 17212 11060 17224
rect 11112 17212 11118 17264
rect 17773 17255 17831 17261
rect 17773 17221 17785 17255
rect 17819 17252 17831 17255
rect 18233 17255 18291 17261
rect 18233 17252 18245 17255
rect 17819 17224 18245 17252
rect 17819 17221 17831 17224
rect 17773 17215 17831 17221
rect 18233 17221 18245 17224
rect 18279 17221 18291 17255
rect 18233 17215 18291 17221
rect 19061 17255 19119 17261
rect 19061 17221 19073 17255
rect 19107 17252 19119 17255
rect 20073 17255 20131 17261
rect 20073 17252 20085 17255
rect 19107 17224 20085 17252
rect 19107 17221 19119 17224
rect 19061 17215 19119 17221
rect 20073 17221 20085 17224
rect 20119 17221 20131 17255
rect 22066 17252 22094 17292
rect 22278 17280 22284 17332
rect 22336 17320 22342 17332
rect 22399 17323 22457 17329
rect 22399 17320 22411 17323
rect 22336 17292 22411 17320
rect 22336 17280 22342 17292
rect 22399 17289 22411 17292
rect 22445 17320 22457 17323
rect 23290 17320 23296 17332
rect 22445 17292 23296 17320
rect 22445 17289 22457 17292
rect 22399 17283 22457 17289
rect 23290 17280 23296 17292
rect 23348 17280 23354 17332
rect 22189 17255 22247 17261
rect 22189 17252 22201 17255
rect 22066 17224 22201 17252
rect 20073 17215 20131 17221
rect 22189 17221 22201 17224
rect 22235 17221 22247 17255
rect 22189 17215 22247 17221
rect 9999 17156 10180 17184
rect 9999 17153 10011 17156
rect 9953 17147 10011 17153
rect 10226 17144 10232 17196
rect 10284 17144 10290 17196
rect 12342 17144 12348 17196
rect 12400 17144 12406 17196
rect 12434 17144 12440 17196
rect 12492 17184 12498 17196
rect 12802 17184 12808 17196
rect 12492 17156 12808 17184
rect 12492 17144 12498 17156
rect 12802 17144 12808 17156
rect 12860 17144 12866 17196
rect 15289 17187 15347 17193
rect 15289 17153 15301 17187
rect 15335 17184 15347 17187
rect 15838 17184 15844 17196
rect 15335 17156 15844 17184
rect 15335 17153 15347 17156
rect 15289 17147 15347 17153
rect 15838 17144 15844 17156
rect 15896 17144 15902 17196
rect 16022 17144 16028 17196
rect 16080 17184 16086 17196
rect 17221 17187 17279 17193
rect 17221 17184 17233 17187
rect 16080 17156 17233 17184
rect 16080 17144 16086 17156
rect 17221 17153 17233 17156
rect 17267 17153 17279 17187
rect 17221 17147 17279 17153
rect 17494 17144 17500 17196
rect 17552 17184 17558 17196
rect 17589 17187 17647 17193
rect 17589 17184 17601 17187
rect 17552 17156 17601 17184
rect 17552 17144 17558 17156
rect 17589 17153 17601 17156
rect 17635 17153 17647 17187
rect 17589 17147 17647 17153
rect 17865 17187 17923 17193
rect 17865 17153 17877 17187
rect 17911 17184 17923 17187
rect 18138 17184 18144 17196
rect 17911 17156 18144 17184
rect 17911 17153 17923 17156
rect 17865 17147 17923 17153
rect 18138 17144 18144 17156
rect 18196 17184 18202 17196
rect 18506 17184 18512 17196
rect 18196 17156 18512 17184
rect 18196 17144 18202 17156
rect 18506 17144 18512 17156
rect 18564 17144 18570 17196
rect 18598 17144 18604 17196
rect 18656 17184 18662 17196
rect 18785 17187 18843 17193
rect 18785 17184 18797 17187
rect 18656 17156 18797 17184
rect 18656 17144 18662 17156
rect 18785 17153 18797 17156
rect 18831 17153 18843 17187
rect 18785 17147 18843 17153
rect 18969 17187 19027 17193
rect 18969 17153 18981 17187
rect 19015 17153 19027 17187
rect 18969 17147 19027 17153
rect 10244 17116 10272 17144
rect 8864 17088 10272 17116
rect 12360 17116 12388 17144
rect 12360 17088 12940 17116
rect 8754 17008 8760 17060
rect 8812 17048 8818 17060
rect 10594 17048 10600 17060
rect 8812 17020 10600 17048
rect 8812 17008 8818 17020
rect 10594 17008 10600 17020
rect 10652 17008 10658 17060
rect 9582 16980 9588 16992
rect 8588 16952 9588 16980
rect 9582 16940 9588 16952
rect 9640 16940 9646 16992
rect 12158 16940 12164 16992
rect 12216 16940 12222 16992
rect 12437 16983 12495 16989
rect 12437 16949 12449 16983
rect 12483 16980 12495 16983
rect 12802 16980 12808 16992
rect 12483 16952 12808 16980
rect 12483 16949 12495 16952
rect 12437 16943 12495 16949
rect 12802 16940 12808 16952
rect 12860 16940 12866 16992
rect 12912 16980 12940 17088
rect 13906 17076 13912 17128
rect 13964 17076 13970 17128
rect 14182 17076 14188 17128
rect 14240 17076 14246 17128
rect 15565 17119 15623 17125
rect 15565 17085 15577 17119
rect 15611 17116 15623 17119
rect 16669 17119 16727 17125
rect 16669 17116 16681 17119
rect 15611 17088 16681 17116
rect 15611 17085 15623 17088
rect 15565 17079 15623 17085
rect 16669 17085 16681 17088
rect 16715 17085 16727 17119
rect 18984 17116 19012 17147
rect 19242 17144 19248 17196
rect 19300 17144 19306 17196
rect 19426 17144 19432 17196
rect 19484 17144 19490 17196
rect 20622 17144 20628 17196
rect 20680 17184 20686 17196
rect 20717 17187 20775 17193
rect 20717 17184 20729 17187
rect 20680 17156 20729 17184
rect 20680 17144 20686 17156
rect 20717 17153 20729 17156
rect 20763 17153 20775 17187
rect 22204 17184 22232 17215
rect 22646 17212 22652 17264
rect 22704 17252 22710 17264
rect 22893 17255 22951 17261
rect 22893 17252 22905 17255
rect 22704 17224 22905 17252
rect 22704 17212 22710 17224
rect 22893 17221 22905 17224
rect 22939 17221 22951 17255
rect 22893 17215 22951 17221
rect 23109 17255 23167 17261
rect 23109 17221 23121 17255
rect 23155 17221 23167 17255
rect 23109 17215 23167 17221
rect 23124 17184 23152 17215
rect 26878 17212 26884 17264
rect 26936 17252 26942 17264
rect 27709 17255 27767 17261
rect 27709 17252 27721 17255
rect 26936 17224 27721 17252
rect 26936 17212 26942 17224
rect 27709 17221 27721 17224
rect 27755 17221 27767 17255
rect 27709 17215 27767 17221
rect 28074 17212 28080 17264
rect 28132 17212 28138 17264
rect 22204 17156 23152 17184
rect 20717 17147 20775 17153
rect 25590 17144 25596 17196
rect 25648 17144 25654 17196
rect 19518 17116 19524 17128
rect 18984 17088 19524 17116
rect 16669 17079 16727 17085
rect 19518 17076 19524 17088
rect 19576 17116 19582 17128
rect 19978 17116 19984 17128
rect 19576 17088 19984 17116
rect 19576 17076 19582 17088
rect 19978 17076 19984 17088
rect 20036 17076 20042 17128
rect 25317 17119 25375 17125
rect 25317 17085 25329 17119
rect 25363 17116 25375 17119
rect 25406 17116 25412 17128
rect 25363 17088 25412 17116
rect 25363 17085 25375 17088
rect 25317 17079 25375 17085
rect 25406 17076 25412 17088
rect 25464 17076 25470 17128
rect 25501 17119 25559 17125
rect 25501 17085 25513 17119
rect 25547 17116 25559 17119
rect 25866 17116 25872 17128
rect 25547 17088 25872 17116
rect 25547 17085 25559 17088
rect 25501 17079 25559 17085
rect 25866 17076 25872 17088
rect 25924 17076 25930 17128
rect 14108 17020 17356 17048
rect 14108 16980 14136 17020
rect 17328 16992 17356 17020
rect 22462 17008 22468 17060
rect 22520 17048 22526 17060
rect 22741 17051 22799 17057
rect 22741 17048 22753 17051
rect 22520 17020 22753 17048
rect 22520 17008 22526 17020
rect 22741 17017 22753 17020
rect 22787 17017 22799 17051
rect 22741 17011 22799 17017
rect 12912 16952 14136 16980
rect 14734 16940 14740 16992
rect 14792 16980 14798 16992
rect 15105 16983 15163 16989
rect 15105 16980 15117 16983
rect 14792 16952 15117 16980
rect 14792 16940 14798 16952
rect 15105 16949 15117 16952
rect 15151 16949 15163 16983
rect 15105 16943 15163 16949
rect 15470 16940 15476 16992
rect 15528 16940 15534 16992
rect 17310 16940 17316 16992
rect 17368 16980 17374 16992
rect 22278 16980 22284 16992
rect 17368 16952 22284 16980
rect 17368 16940 17374 16952
rect 22278 16940 22284 16952
rect 22336 16940 22342 16992
rect 22370 16940 22376 16992
rect 22428 16940 22434 16992
rect 22554 16940 22560 16992
rect 22612 16940 22618 16992
rect 22925 16983 22983 16989
rect 22925 16949 22937 16983
rect 22971 16980 22983 16983
rect 23934 16980 23940 16992
rect 22971 16952 23940 16980
rect 22971 16949 22983 16952
rect 22925 16943 22983 16949
rect 23934 16940 23940 16952
rect 23992 16940 23998 16992
rect 25038 16940 25044 16992
rect 25096 16980 25102 16992
rect 25409 16983 25467 16989
rect 25409 16980 25421 16983
rect 25096 16952 25421 16980
rect 25096 16940 25102 16952
rect 25409 16949 25421 16952
rect 25455 16949 25467 16983
rect 25409 16943 25467 16949
rect 1104 16890 28704 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 28704 16890
rect 1104 16816 28704 16838
rect 4798 16736 4804 16788
rect 4856 16776 4862 16788
rect 5626 16776 5632 16788
rect 4856 16748 5632 16776
rect 4856 16736 4862 16748
rect 5626 16736 5632 16748
rect 5684 16736 5690 16788
rect 8662 16736 8668 16788
rect 8720 16776 8726 16788
rect 9306 16776 9312 16788
rect 8720 16748 9312 16776
rect 8720 16736 8726 16748
rect 9306 16736 9312 16748
rect 9364 16736 9370 16788
rect 15470 16736 15476 16788
rect 15528 16776 15534 16788
rect 16206 16776 16212 16788
rect 15528 16748 16212 16776
rect 15528 16736 15534 16748
rect 16206 16736 16212 16748
rect 16264 16776 16270 16788
rect 19058 16776 19064 16788
rect 16264 16748 19064 16776
rect 16264 16736 16270 16748
rect 19058 16736 19064 16748
rect 19116 16776 19122 16788
rect 22646 16776 22652 16788
rect 19116 16748 22652 16776
rect 19116 16736 19122 16748
rect 22646 16736 22652 16748
rect 22704 16736 22710 16788
rect 25038 16736 25044 16788
rect 25096 16736 25102 16788
rect 26786 16736 26792 16788
rect 26844 16776 26850 16788
rect 27157 16779 27215 16785
rect 27157 16776 27169 16779
rect 26844 16748 27169 16776
rect 26844 16736 26850 16748
rect 27157 16745 27169 16748
rect 27203 16745 27215 16779
rect 27157 16739 27215 16745
rect 6089 16711 6147 16717
rect 6089 16677 6101 16711
rect 6135 16677 6147 16711
rect 26878 16708 26884 16720
rect 6089 16671 6147 16677
rect 26712 16680 26884 16708
rect 4430 16600 4436 16652
rect 4488 16640 4494 16652
rect 5442 16640 5448 16652
rect 4488 16612 5448 16640
rect 4488 16600 4494 16612
rect 5442 16600 5448 16612
rect 5500 16640 5506 16652
rect 5537 16643 5595 16649
rect 5537 16640 5549 16643
rect 5500 16612 5549 16640
rect 5500 16600 5506 16612
rect 5537 16609 5549 16612
rect 5583 16609 5595 16643
rect 5537 16603 5595 16609
rect 5813 16575 5871 16581
rect 5813 16541 5825 16575
rect 5859 16572 5871 16575
rect 6104 16572 6132 16671
rect 6178 16600 6184 16652
rect 6236 16640 6242 16652
rect 7742 16640 7748 16652
rect 6236 16612 6592 16640
rect 6236 16600 6242 16612
rect 6564 16584 6592 16612
rect 6748 16612 7748 16640
rect 6748 16584 6776 16612
rect 7742 16600 7748 16612
rect 7800 16600 7806 16652
rect 9401 16643 9459 16649
rect 9401 16609 9413 16643
rect 9447 16640 9459 16643
rect 10134 16640 10140 16652
rect 9447 16612 10140 16640
rect 9447 16609 9459 16612
rect 9401 16603 9459 16609
rect 10134 16600 10140 16612
rect 10192 16600 10198 16652
rect 12434 16640 12440 16652
rect 11440 16612 12440 16640
rect 5859 16544 6132 16572
rect 6268 16575 6326 16581
rect 5859 16541 5871 16544
rect 5813 16535 5871 16541
rect 6268 16541 6280 16575
rect 6314 16541 6326 16575
rect 6268 16535 6326 16541
rect 5994 16396 6000 16448
rect 6052 16396 6058 16448
rect 6288 16436 6316 16535
rect 6454 16532 6460 16584
rect 6512 16532 6518 16584
rect 6546 16532 6552 16584
rect 6604 16581 6610 16584
rect 6604 16575 6643 16581
rect 6631 16541 6643 16575
rect 6604 16535 6643 16541
rect 6604 16532 6610 16535
rect 6730 16532 6736 16584
rect 6788 16532 6794 16584
rect 9030 16532 9036 16584
rect 9088 16532 9094 16584
rect 9231 16575 9289 16581
rect 9231 16541 9243 16575
rect 9277 16572 9289 16575
rect 9582 16572 9588 16584
rect 9277 16544 9588 16572
rect 9277 16541 9289 16544
rect 9231 16535 9289 16541
rect 9582 16532 9588 16544
rect 9640 16532 9646 16584
rect 11330 16532 11336 16584
rect 11388 16572 11394 16584
rect 11440 16572 11468 16612
rect 12434 16600 12440 16612
rect 12492 16600 12498 16652
rect 12713 16643 12771 16649
rect 12713 16609 12725 16643
rect 12759 16640 12771 16643
rect 14182 16640 14188 16652
rect 12759 16612 14188 16640
rect 12759 16609 12771 16612
rect 12713 16603 12771 16609
rect 14182 16600 14188 16612
rect 14240 16640 14246 16652
rect 14461 16643 14519 16649
rect 14461 16640 14473 16643
rect 14240 16612 14473 16640
rect 14240 16600 14246 16612
rect 14461 16609 14473 16612
rect 14507 16609 14519 16643
rect 14461 16603 14519 16609
rect 14734 16600 14740 16652
rect 14792 16600 14798 16652
rect 23753 16643 23811 16649
rect 23753 16609 23765 16643
rect 23799 16640 23811 16643
rect 23934 16640 23940 16652
rect 23799 16612 23940 16640
rect 23799 16609 23811 16612
rect 23753 16603 23811 16609
rect 23934 16600 23940 16612
rect 23992 16600 23998 16652
rect 25130 16600 25136 16652
rect 25188 16600 25194 16652
rect 25222 16600 25228 16652
rect 25280 16600 25286 16652
rect 11388 16544 11468 16572
rect 11388 16532 11394 16544
rect 12802 16532 12808 16584
rect 12860 16532 12866 16584
rect 13817 16575 13875 16581
rect 13817 16541 13829 16575
rect 13863 16572 13875 16575
rect 14274 16572 14280 16584
rect 13863 16544 14280 16572
rect 13863 16541 13875 16544
rect 13817 16535 13875 16541
rect 14274 16532 14280 16544
rect 14332 16532 14338 16584
rect 18046 16532 18052 16584
rect 18104 16572 18110 16584
rect 18509 16575 18567 16581
rect 18509 16572 18521 16575
rect 18104 16544 18521 16572
rect 18104 16532 18110 16544
rect 18509 16541 18521 16544
rect 18555 16541 18567 16575
rect 18509 16535 18567 16541
rect 22373 16575 22431 16581
rect 22373 16541 22385 16575
rect 22419 16572 22431 16575
rect 22554 16572 22560 16584
rect 22419 16544 22560 16572
rect 22419 16541 22431 16544
rect 22373 16535 22431 16541
rect 22554 16532 22560 16544
rect 22612 16532 22618 16584
rect 22646 16532 22652 16584
rect 22704 16532 22710 16584
rect 24857 16575 24915 16581
rect 24857 16541 24869 16575
rect 24903 16572 24915 16575
rect 24903 16544 25084 16572
rect 24903 16541 24915 16544
rect 24857 16535 24915 16541
rect 6365 16507 6423 16513
rect 6365 16473 6377 16507
rect 6411 16504 6423 16507
rect 8846 16504 8852 16516
rect 6411 16476 8852 16504
rect 6411 16473 6423 16476
rect 6365 16467 6423 16473
rect 8846 16464 8852 16476
rect 8904 16464 8910 16516
rect 9048 16504 9076 16532
rect 11146 16504 11152 16516
rect 9048 16476 11152 16504
rect 11146 16464 11152 16476
rect 11204 16464 11210 16516
rect 12434 16464 12440 16516
rect 12492 16464 12498 16516
rect 16482 16504 16488 16516
rect 15962 16476 16488 16504
rect 16482 16464 16488 16476
rect 16540 16464 16546 16516
rect 8386 16436 8392 16448
rect 6288 16408 8392 16436
rect 8386 16396 8392 16408
rect 8444 16396 8450 16448
rect 8938 16396 8944 16448
rect 8996 16436 9002 16448
rect 9033 16439 9091 16445
rect 9033 16436 9045 16439
rect 8996 16408 9045 16436
rect 8996 16396 9002 16408
rect 9033 16405 9045 16408
rect 9079 16405 9091 16439
rect 9033 16399 9091 16405
rect 10965 16439 11023 16445
rect 10965 16405 10977 16439
rect 11011 16436 11023 16439
rect 11422 16436 11428 16448
rect 11011 16408 11428 16436
rect 11011 16405 11023 16408
rect 10965 16399 11023 16405
rect 11422 16396 11428 16408
rect 11480 16396 11486 16448
rect 13170 16396 13176 16448
rect 13228 16436 13234 16448
rect 13449 16439 13507 16445
rect 13449 16436 13461 16439
rect 13228 16408 13461 16436
rect 13228 16396 13234 16408
rect 13449 16405 13461 16408
rect 13495 16405 13507 16439
rect 13449 16399 13507 16405
rect 13538 16396 13544 16448
rect 13596 16436 13602 16448
rect 13633 16439 13691 16445
rect 13633 16436 13645 16439
rect 13596 16408 13645 16436
rect 13596 16396 13602 16408
rect 13633 16405 13645 16408
rect 13679 16436 13691 16439
rect 15102 16436 15108 16448
rect 13679 16408 15108 16436
rect 13679 16405 13691 16408
rect 13633 16399 13691 16405
rect 15102 16396 15108 16408
rect 15160 16396 15166 16448
rect 16022 16396 16028 16448
rect 16080 16436 16086 16448
rect 16209 16439 16267 16445
rect 16209 16436 16221 16439
rect 16080 16408 16221 16436
rect 16080 16396 16086 16408
rect 16209 16405 16221 16408
rect 16255 16405 16267 16439
rect 16209 16399 16267 16405
rect 18690 16396 18696 16448
rect 18748 16396 18754 16448
rect 22186 16396 22192 16448
rect 22244 16396 22250 16448
rect 22557 16439 22615 16445
rect 22557 16405 22569 16439
rect 22603 16436 22615 16439
rect 23109 16439 23167 16445
rect 23109 16436 23121 16439
rect 22603 16408 23121 16436
rect 22603 16405 22615 16408
rect 22557 16399 22615 16405
rect 23109 16405 23121 16408
rect 23155 16405 23167 16439
rect 23109 16399 23167 16405
rect 24670 16396 24676 16448
rect 24728 16396 24734 16448
rect 24854 16396 24860 16448
rect 24912 16436 24918 16448
rect 25056 16436 25084 16544
rect 26602 16532 26608 16584
rect 26660 16572 26666 16584
rect 26712 16572 26740 16680
rect 26878 16668 26884 16680
rect 26936 16668 26942 16720
rect 27709 16643 27767 16649
rect 27709 16640 27721 16643
rect 26660 16544 26740 16572
rect 26804 16612 27721 16640
rect 26660 16532 26666 16544
rect 25498 16464 25504 16516
rect 25556 16464 25562 16516
rect 26804 16436 26832 16612
rect 27709 16609 27721 16612
rect 27755 16609 27767 16643
rect 28258 16640 28264 16652
rect 27709 16603 27767 16609
rect 27816 16612 28264 16640
rect 27617 16575 27675 16581
rect 27617 16541 27629 16575
rect 27663 16572 27675 16575
rect 27816 16572 27844 16612
rect 28258 16600 28264 16612
rect 28316 16600 28322 16652
rect 27663 16544 27844 16572
rect 27663 16541 27675 16544
rect 27617 16535 27675 16541
rect 24912 16408 26832 16436
rect 24912 16396 24918 16408
rect 26970 16396 26976 16448
rect 27028 16436 27034 16448
rect 27525 16439 27583 16445
rect 27525 16436 27537 16439
rect 27028 16408 27537 16436
rect 27028 16396 27034 16408
rect 27525 16405 27537 16408
rect 27571 16405 27583 16439
rect 27525 16399 27583 16405
rect 1104 16346 28704 16368
rect 1104 16294 4874 16346
rect 4926 16294 4938 16346
rect 4990 16294 5002 16346
rect 5054 16294 5066 16346
rect 5118 16294 5130 16346
rect 5182 16294 28704 16346
rect 1104 16272 28704 16294
rect 4430 16192 4436 16244
rect 4488 16192 4494 16244
rect 4614 16192 4620 16244
rect 4672 16232 4678 16244
rect 5534 16232 5540 16244
rect 4672 16204 5540 16232
rect 4672 16192 4678 16204
rect 5534 16192 5540 16204
rect 5592 16232 5598 16244
rect 6730 16232 6736 16244
rect 5592 16204 6736 16232
rect 5592 16192 5598 16204
rect 6730 16192 6736 16204
rect 6788 16192 6794 16244
rect 6914 16192 6920 16244
rect 6972 16232 6978 16244
rect 7745 16235 7803 16241
rect 7745 16232 7757 16235
rect 6972 16204 7757 16232
rect 6972 16192 6978 16204
rect 7745 16201 7757 16204
rect 7791 16201 7803 16235
rect 7745 16195 7803 16201
rect 8113 16235 8171 16241
rect 8113 16201 8125 16235
rect 8159 16232 8171 16235
rect 8938 16232 8944 16244
rect 8159 16204 8944 16232
rect 8159 16201 8171 16204
rect 8113 16195 8171 16201
rect 8938 16192 8944 16204
rect 8996 16232 9002 16244
rect 9214 16232 9220 16244
rect 8996 16204 9220 16232
rect 8996 16192 9002 16204
rect 9214 16192 9220 16204
rect 9272 16192 9278 16244
rect 9309 16235 9367 16241
rect 9309 16201 9321 16235
rect 9355 16232 9367 16235
rect 9490 16232 9496 16244
rect 9355 16204 9496 16232
rect 9355 16201 9367 16204
rect 9309 16195 9367 16201
rect 9490 16192 9496 16204
rect 9548 16192 9554 16244
rect 12802 16192 12808 16244
rect 12860 16192 12866 16244
rect 12986 16192 12992 16244
rect 13044 16192 13050 16244
rect 16022 16232 16028 16244
rect 14108 16204 16028 16232
rect 3694 16124 3700 16176
rect 3752 16164 3758 16176
rect 5905 16167 5963 16173
rect 3752 16136 4738 16164
rect 3752 16124 3758 16136
rect 5905 16133 5917 16167
rect 5951 16164 5963 16167
rect 5994 16164 6000 16176
rect 5951 16136 6000 16164
rect 5951 16133 5963 16136
rect 5905 16127 5963 16133
rect 5994 16124 6000 16136
rect 6052 16124 6058 16176
rect 9033 16167 9091 16173
rect 9033 16133 9045 16167
rect 9079 16164 9091 16167
rect 9953 16167 10011 16173
rect 9953 16164 9965 16167
rect 9079 16136 9965 16164
rect 9079 16133 9091 16136
rect 9033 16127 9091 16133
rect 9953 16133 9965 16136
rect 9999 16133 10011 16167
rect 12820 16164 12848 16192
rect 13004 16164 13032 16192
rect 13722 16164 13728 16176
rect 9953 16127 10011 16133
rect 12636 16136 12848 16164
rect 12912 16136 13728 16164
rect 8386 16056 8392 16108
rect 8444 16056 8450 16108
rect 8846 16105 8852 16108
rect 8823 16099 8852 16105
rect 8823 16065 8835 16099
rect 8823 16059 8852 16065
rect 8846 16056 8852 16059
rect 8904 16056 8910 16108
rect 8938 16056 8944 16108
rect 8996 16056 9002 16108
rect 9122 16056 9128 16108
rect 9180 16056 9186 16108
rect 9214 16056 9220 16108
rect 9272 16096 9278 16108
rect 9401 16099 9459 16105
rect 9401 16096 9413 16099
rect 9272 16068 9413 16096
rect 9272 16056 9278 16068
rect 9401 16065 9413 16068
rect 9447 16065 9459 16099
rect 9401 16059 9459 16065
rect 9493 16099 9551 16105
rect 9493 16065 9505 16099
rect 9539 16065 9551 16099
rect 9493 16059 9551 16065
rect 9677 16099 9735 16105
rect 9677 16065 9689 16099
rect 9723 16065 9735 16099
rect 9677 16059 9735 16065
rect 7926 16037 7932 16040
rect 6181 16031 6239 16037
rect 6181 15997 6193 16031
rect 6227 15997 6239 16031
rect 6181 15991 6239 15997
rect 7904 16031 7932 16037
rect 7904 15997 7916 16031
rect 7904 15991 7932 15997
rect 5350 15852 5356 15904
rect 5408 15892 5414 15904
rect 6196 15892 6224 15991
rect 7926 15988 7932 15991
rect 7984 15988 7990 16040
rect 8018 15988 8024 16040
rect 8076 15988 8082 16040
rect 8570 15988 8576 16040
rect 8628 16028 8634 16040
rect 8665 16031 8723 16037
rect 8665 16028 8677 16031
rect 8628 16000 8677 16028
rect 8628 15988 8634 16000
rect 8665 15997 8677 16000
rect 8711 15997 8723 16031
rect 9508 16028 9536 16059
rect 9582 16028 9588 16040
rect 8665 15991 8723 15997
rect 9416 16000 9588 16028
rect 8478 15920 8484 15972
rect 8536 15960 8542 15972
rect 9416 15960 9444 16000
rect 9582 15988 9588 16000
rect 9640 15988 9646 16040
rect 9692 16028 9720 16059
rect 9766 16056 9772 16108
rect 9824 16056 9830 16108
rect 12636 16105 12664 16136
rect 12616 16099 12674 16105
rect 12616 16065 12628 16099
rect 12662 16065 12674 16099
rect 12616 16059 12674 16065
rect 12710 16056 12716 16108
rect 12768 16056 12774 16108
rect 12805 16099 12863 16105
rect 12805 16065 12817 16099
rect 12851 16096 12863 16099
rect 12912 16096 12940 16136
rect 13722 16124 13728 16136
rect 13780 16124 13786 16176
rect 12851 16068 12940 16096
rect 12851 16065 12863 16068
rect 12805 16059 12863 16065
rect 12986 16056 12992 16108
rect 13044 16056 13050 16108
rect 13081 16099 13139 16105
rect 13081 16065 13093 16099
rect 13127 16096 13139 16099
rect 13446 16096 13452 16108
rect 13127 16068 13452 16096
rect 13127 16065 13139 16068
rect 13081 16059 13139 16065
rect 13446 16056 13452 16068
rect 13504 16056 13510 16108
rect 13538 16056 13544 16108
rect 13596 16056 13602 16108
rect 13817 16099 13875 16105
rect 13817 16065 13829 16099
rect 13863 16065 13875 16099
rect 13817 16059 13875 16065
rect 13955 16099 14013 16105
rect 13955 16065 13967 16099
rect 14001 16096 14013 16099
rect 14108 16096 14136 16204
rect 16022 16192 16028 16204
rect 16080 16192 16086 16244
rect 23569 16235 23627 16241
rect 23569 16201 23581 16235
rect 23615 16232 23627 16235
rect 23934 16232 23940 16244
rect 23615 16204 23940 16232
rect 23615 16201 23627 16204
rect 23569 16195 23627 16201
rect 23934 16192 23940 16204
rect 23992 16192 23998 16244
rect 24854 16192 24860 16244
rect 24912 16192 24918 16244
rect 25317 16235 25375 16241
rect 25317 16201 25329 16235
rect 25363 16232 25375 16235
rect 25498 16232 25504 16244
rect 25363 16204 25504 16232
rect 25363 16201 25375 16204
rect 25317 16195 25375 16201
rect 25498 16192 25504 16204
rect 25556 16192 25562 16244
rect 25774 16192 25780 16244
rect 25832 16192 25838 16244
rect 16298 16164 16304 16176
rect 16238 16136 16304 16164
rect 16298 16124 16304 16136
rect 16356 16164 16362 16176
rect 16482 16164 16488 16176
rect 16356 16136 16488 16164
rect 16356 16124 16362 16136
rect 16482 16124 16488 16136
rect 16540 16124 16546 16176
rect 18782 16124 18788 16176
rect 18840 16124 18846 16176
rect 22097 16167 22155 16173
rect 22097 16133 22109 16167
rect 22143 16164 22155 16167
rect 22186 16164 22192 16176
rect 22143 16136 22192 16164
rect 22143 16133 22155 16136
rect 22097 16127 22155 16133
rect 22186 16124 22192 16136
rect 22244 16124 22250 16176
rect 23382 16164 23388 16176
rect 23322 16136 23388 16164
rect 23382 16124 23388 16136
rect 23440 16124 23446 16176
rect 26605 16167 26663 16173
rect 26605 16164 26617 16167
rect 25424 16136 26617 16164
rect 25424 16108 25452 16136
rect 26605 16133 26617 16136
rect 26651 16133 26663 16167
rect 26605 16127 26663 16133
rect 14001 16068 14136 16096
rect 14001 16065 14013 16068
rect 13955 16059 14013 16065
rect 9858 16028 9864 16040
rect 9692 16000 9864 16028
rect 9858 15988 9864 16000
rect 9916 15988 9922 16040
rect 11422 15988 11428 16040
rect 11480 16028 11486 16040
rect 11517 16031 11575 16037
rect 11517 16028 11529 16031
rect 11480 16000 11529 16028
rect 11480 15988 11486 16000
rect 11517 15997 11529 16000
rect 11563 15997 11575 16031
rect 13832 16028 13860 16059
rect 14182 16056 14188 16108
rect 14240 16096 14246 16108
rect 14737 16099 14795 16105
rect 14737 16096 14749 16099
rect 14240 16068 14749 16096
rect 14240 16056 14246 16068
rect 14737 16065 14749 16068
rect 14783 16065 14795 16099
rect 14737 16059 14795 16065
rect 17862 16056 17868 16108
rect 17920 16056 17926 16108
rect 20622 16056 20628 16108
rect 20680 16096 20686 16108
rect 21085 16099 21143 16105
rect 21085 16096 21097 16099
rect 20680 16068 21097 16096
rect 20680 16056 20686 16068
rect 21085 16065 21097 16068
rect 21131 16065 21143 16099
rect 21085 16059 21143 16065
rect 25041 16099 25099 16105
rect 25041 16065 25053 16099
rect 25087 16065 25099 16099
rect 25041 16059 25099 16065
rect 25225 16099 25283 16105
rect 25225 16065 25237 16099
rect 25271 16096 25283 16099
rect 25406 16096 25412 16108
rect 25271 16068 25412 16096
rect 25271 16065 25283 16068
rect 25225 16059 25283 16065
rect 13832 16000 14228 16028
rect 11517 15991 11575 15997
rect 8536 15932 9444 15960
rect 8536 15920 8542 15932
rect 5408 15864 6224 15892
rect 5408 15852 5414 15864
rect 8294 15852 8300 15904
rect 8352 15892 8358 15904
rect 8846 15892 8852 15904
rect 8352 15864 8852 15892
rect 8352 15852 8358 15864
rect 8846 15852 8852 15864
rect 8904 15892 8910 15904
rect 9398 15892 9404 15904
rect 8904 15864 9404 15892
rect 8904 15852 8910 15864
rect 9398 15852 9404 15864
rect 9456 15852 9462 15904
rect 11790 15852 11796 15904
rect 11848 15892 11854 15904
rect 12161 15895 12219 15901
rect 12161 15892 12173 15895
rect 11848 15864 12173 15892
rect 11848 15852 11854 15864
rect 12161 15861 12173 15864
rect 12207 15861 12219 15895
rect 12161 15855 12219 15861
rect 12437 15895 12495 15901
rect 12437 15861 12449 15895
rect 12483 15892 12495 15895
rect 12526 15892 12532 15904
rect 12483 15864 12532 15892
rect 12483 15861 12495 15864
rect 12437 15855 12495 15861
rect 12526 15852 12532 15864
rect 12584 15852 12590 15904
rect 13446 15852 13452 15904
rect 13504 15892 13510 15904
rect 14093 15895 14151 15901
rect 14093 15892 14105 15895
rect 13504 15864 14105 15892
rect 13504 15852 13510 15864
rect 14093 15861 14105 15864
rect 14139 15861 14151 15895
rect 14200 15892 14228 16000
rect 15010 15988 15016 16040
rect 15068 15988 15074 16040
rect 15654 15988 15660 16040
rect 15712 16028 15718 16040
rect 16485 16031 16543 16037
rect 16485 16028 16497 16031
rect 15712 16000 16497 16028
rect 15712 15988 15718 16000
rect 16485 15997 16497 16000
rect 16531 16028 16543 16031
rect 17221 16031 17279 16037
rect 17221 16028 17233 16031
rect 16531 16000 17233 16028
rect 16531 15997 16543 16000
rect 16485 15991 16543 15997
rect 17221 15997 17233 16000
rect 17267 15997 17279 16031
rect 17221 15991 17279 15997
rect 18141 16031 18199 16037
rect 18141 15997 18153 16031
rect 18187 16028 18199 16031
rect 18230 16028 18236 16040
rect 18187 16000 18236 16028
rect 18187 15997 18199 16000
rect 18141 15991 18199 15997
rect 18230 15988 18236 16000
rect 18288 15988 18294 16040
rect 19613 16031 19671 16037
rect 19613 15997 19625 16031
rect 19659 16028 19671 16031
rect 20257 16031 20315 16037
rect 20257 16028 20269 16031
rect 19659 16000 20269 16028
rect 19659 15997 19671 16000
rect 19613 15991 19671 15997
rect 20257 15997 20269 16000
rect 20303 16028 20315 16031
rect 20438 16028 20444 16040
rect 20303 16000 20444 16028
rect 20303 15997 20315 16000
rect 20257 15991 20315 15997
rect 20438 15988 20444 16000
rect 20496 15988 20502 16040
rect 21358 15988 21364 16040
rect 21416 15988 21422 16040
rect 21818 15988 21824 16040
rect 21876 15988 21882 16040
rect 19150 15920 19156 15972
rect 19208 15960 19214 15972
rect 21269 15963 21327 15969
rect 21269 15960 21281 15963
rect 19208 15932 21281 15960
rect 19208 15920 19214 15932
rect 21269 15929 21281 15932
rect 21315 15929 21327 15963
rect 25056 15960 25084 16059
rect 25406 16056 25412 16068
rect 25464 16056 25470 16108
rect 25590 16056 25596 16108
rect 25648 16096 25654 16108
rect 25685 16099 25743 16105
rect 25685 16096 25697 16099
rect 25648 16068 25697 16096
rect 25648 16056 25654 16068
rect 25685 16065 25697 16068
rect 25731 16096 25743 16099
rect 26970 16096 26976 16108
rect 25731 16068 26976 16096
rect 25731 16065 25743 16068
rect 25685 16059 25743 16065
rect 26970 16056 26976 16068
rect 27028 16056 27034 16108
rect 28350 16056 28356 16108
rect 28408 16056 28414 16108
rect 25961 16031 26019 16037
rect 25961 15997 25973 16031
rect 26007 16028 26019 16031
rect 26145 16031 26203 16037
rect 26145 16028 26157 16031
rect 26007 16000 26157 16028
rect 26007 15997 26019 16000
rect 25961 15991 26019 15997
rect 26145 15997 26157 16000
rect 26191 15997 26203 16031
rect 26145 15991 26203 15997
rect 26237 15963 26295 15969
rect 26237 15960 26249 15963
rect 25056 15932 26249 15960
rect 21269 15923 21327 15929
rect 26160 15904 26188 15932
rect 26237 15929 26249 15932
rect 26283 15929 26295 15963
rect 26237 15923 26295 15929
rect 15746 15892 15752 15904
rect 14200 15864 15752 15892
rect 14093 15855 14151 15861
rect 15746 15852 15752 15864
rect 15804 15852 15810 15904
rect 16666 15852 16672 15904
rect 16724 15852 16730 15904
rect 19702 15852 19708 15904
rect 19760 15852 19766 15904
rect 20898 15852 20904 15904
rect 20956 15852 20962 15904
rect 26142 15852 26148 15904
rect 26200 15852 26206 15904
rect 27614 15852 27620 15904
rect 27672 15892 27678 15904
rect 28169 15895 28227 15901
rect 28169 15892 28181 15895
rect 27672 15864 28181 15892
rect 27672 15852 27678 15864
rect 28169 15861 28181 15864
rect 28215 15861 28227 15895
rect 28169 15855 28227 15861
rect 1104 15802 28704 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 28704 15802
rect 1104 15728 28704 15750
rect 9033 15691 9091 15697
rect 9033 15657 9045 15691
rect 9079 15688 9091 15691
rect 9122 15688 9128 15700
rect 9079 15660 9128 15688
rect 9079 15657 9091 15660
rect 9033 15651 9091 15657
rect 9122 15648 9128 15660
rect 9180 15648 9186 15700
rect 12253 15691 12311 15697
rect 12253 15657 12265 15691
rect 12299 15688 12311 15691
rect 12434 15688 12440 15700
rect 12299 15660 12440 15688
rect 12299 15657 12311 15660
rect 12253 15651 12311 15657
rect 12434 15648 12440 15660
rect 12492 15648 12498 15700
rect 12897 15691 12955 15697
rect 12897 15657 12909 15691
rect 12943 15688 12955 15691
rect 13078 15688 13084 15700
rect 12943 15660 13084 15688
rect 12943 15657 12955 15660
rect 12897 15651 12955 15657
rect 13078 15648 13084 15660
rect 13136 15648 13142 15700
rect 13633 15691 13691 15697
rect 13633 15657 13645 15691
rect 13679 15688 13691 15691
rect 13906 15688 13912 15700
rect 13679 15660 13912 15688
rect 13679 15657 13691 15660
rect 13633 15651 13691 15657
rect 13906 15648 13912 15660
rect 13964 15648 13970 15700
rect 15010 15648 15016 15700
rect 15068 15688 15074 15700
rect 15933 15691 15991 15697
rect 15933 15688 15945 15691
rect 15068 15660 15945 15688
rect 15068 15648 15074 15660
rect 15933 15657 15945 15660
rect 15979 15657 15991 15691
rect 15933 15651 15991 15657
rect 16206 15648 16212 15700
rect 16264 15688 16270 15700
rect 16301 15691 16359 15697
rect 16301 15688 16313 15691
rect 16264 15660 16313 15688
rect 16264 15648 16270 15660
rect 16301 15657 16313 15660
rect 16347 15657 16359 15691
rect 16301 15651 16359 15657
rect 18230 15648 18236 15700
rect 18288 15648 18294 15700
rect 20622 15648 20628 15700
rect 20680 15648 20686 15700
rect 20714 15648 20720 15700
rect 20772 15688 20778 15700
rect 21085 15691 21143 15697
rect 21085 15688 21097 15691
rect 20772 15660 21097 15688
rect 20772 15648 20778 15660
rect 21085 15657 21097 15660
rect 21131 15688 21143 15691
rect 21174 15688 21180 15700
rect 21131 15660 21180 15688
rect 21131 15657 21143 15660
rect 21085 15651 21143 15657
rect 21174 15648 21180 15660
rect 21232 15648 21238 15700
rect 21358 15648 21364 15700
rect 21416 15648 21422 15700
rect 22186 15688 22192 15700
rect 22066 15660 22192 15688
rect 13096 15620 13124 15648
rect 14090 15620 14096 15632
rect 13096 15592 14096 15620
rect 14090 15580 14096 15592
rect 14148 15580 14154 15632
rect 15838 15580 15844 15632
rect 15896 15580 15902 15632
rect 18690 15580 18696 15632
rect 18748 15620 18754 15632
rect 22066 15620 22094 15660
rect 22186 15648 22192 15660
rect 22244 15648 22250 15700
rect 23382 15648 23388 15700
rect 23440 15688 23446 15700
rect 23440 15660 25820 15688
rect 23440 15648 23446 15660
rect 18748 15592 22094 15620
rect 18748 15580 18754 15592
rect 8478 15512 8484 15564
rect 8536 15552 8542 15564
rect 10042 15552 10048 15564
rect 8536 15524 10048 15552
rect 8536 15512 8542 15524
rect 10042 15512 10048 15524
rect 10100 15552 10106 15564
rect 10137 15555 10195 15561
rect 10137 15552 10149 15555
rect 10100 15524 10149 15552
rect 10100 15512 10106 15524
rect 10137 15521 10149 15524
rect 10183 15521 10195 15555
rect 11698 15552 11704 15564
rect 10137 15515 10195 15521
rect 10428 15524 11704 15552
rect 10428 15496 10456 15524
rect 11698 15512 11704 15524
rect 11756 15512 11762 15564
rect 11790 15512 11796 15564
rect 11848 15512 11854 15564
rect 12158 15552 12164 15564
rect 11900 15524 12164 15552
rect 9214 15444 9220 15496
rect 9272 15444 9278 15496
rect 9766 15444 9772 15496
rect 9824 15444 9830 15496
rect 9861 15487 9919 15493
rect 9861 15453 9873 15487
rect 9907 15453 9919 15487
rect 9861 15447 9919 15453
rect 9674 15376 9680 15428
rect 9732 15416 9738 15428
rect 9876 15416 9904 15447
rect 10410 15444 10416 15496
rect 10468 15444 10474 15496
rect 11238 15444 11244 15496
rect 11296 15484 11302 15496
rect 11900 15493 11928 15524
rect 12158 15512 12164 15524
rect 12216 15552 12222 15564
rect 12216 15524 13124 15552
rect 12216 15512 12222 15524
rect 11885 15487 11943 15493
rect 11885 15484 11897 15487
rect 11296 15456 11897 15484
rect 11296 15444 11302 15456
rect 11885 15453 11897 15456
rect 11931 15453 11943 15487
rect 11885 15447 11943 15453
rect 12069 15487 12127 15493
rect 12069 15453 12081 15487
rect 12115 15484 12127 15487
rect 12526 15484 12532 15496
rect 12115 15456 12532 15484
rect 12115 15453 12127 15456
rect 12069 15447 12127 15453
rect 12526 15444 12532 15456
rect 12584 15444 12590 15496
rect 13096 15484 13124 15524
rect 13170 15512 13176 15564
rect 13228 15512 13234 15564
rect 13265 15555 13323 15561
rect 13265 15521 13277 15555
rect 13311 15552 13323 15555
rect 16206 15552 16212 15564
rect 13311 15524 16212 15552
rect 13311 15521 13323 15524
rect 13265 15515 13323 15521
rect 13280 15484 13308 15515
rect 16206 15512 16212 15524
rect 16264 15512 16270 15564
rect 16393 15555 16451 15561
rect 16393 15521 16405 15555
rect 16439 15552 16451 15555
rect 16666 15552 16672 15564
rect 16439 15524 16672 15552
rect 16439 15521 16451 15524
rect 16393 15515 16451 15521
rect 16666 15512 16672 15524
rect 16724 15512 16730 15564
rect 13096 15456 13308 15484
rect 13446 15444 13452 15496
rect 13504 15444 13510 15496
rect 15194 15444 15200 15496
rect 15252 15444 15258 15496
rect 15378 15493 15384 15496
rect 15345 15487 15384 15493
rect 15345 15453 15357 15487
rect 15345 15447 15384 15453
rect 15378 15444 15384 15447
rect 15436 15444 15442 15496
rect 15654 15444 15660 15496
rect 15712 15493 15718 15496
rect 15712 15484 15720 15493
rect 15712 15456 15757 15484
rect 15712 15447 15720 15456
rect 15712 15444 15718 15447
rect 15930 15444 15936 15496
rect 15988 15484 15994 15496
rect 16117 15487 16175 15493
rect 16117 15484 16129 15487
rect 15988 15456 16129 15484
rect 15988 15444 15994 15456
rect 16117 15453 16129 15456
rect 16163 15453 16175 15487
rect 16117 15447 16175 15453
rect 18417 15487 18475 15493
rect 18417 15453 18429 15487
rect 18463 15484 18475 15487
rect 18800 15484 18828 15592
rect 18877 15555 18935 15561
rect 18877 15521 18889 15555
rect 18923 15552 18935 15555
rect 19702 15552 19708 15564
rect 18923 15524 19708 15552
rect 18923 15521 18935 15524
rect 18877 15515 18935 15521
rect 19702 15512 19708 15524
rect 19760 15512 19766 15564
rect 18463 15456 18828 15484
rect 18463 15453 18475 15456
rect 18417 15447 18475 15453
rect 19426 15444 19432 15496
rect 19484 15484 19490 15496
rect 19797 15487 19855 15493
rect 19797 15484 19809 15487
rect 19484 15456 19809 15484
rect 19484 15444 19490 15456
rect 19797 15453 19809 15456
rect 19843 15453 19855 15487
rect 19797 15447 19855 15453
rect 19978 15444 19984 15496
rect 20036 15444 20042 15496
rect 20272 15493 20300 15592
rect 21818 15512 21824 15564
rect 21876 15552 21882 15564
rect 22097 15555 22155 15561
rect 22097 15552 22109 15555
rect 21876 15524 22109 15552
rect 21876 15512 21882 15524
rect 22097 15521 22109 15524
rect 22143 15552 22155 15555
rect 24397 15555 24455 15561
rect 24397 15552 24409 15555
rect 22143 15524 24409 15552
rect 22143 15521 22155 15524
rect 22097 15515 22155 15521
rect 24397 15521 24409 15524
rect 24443 15552 24455 15555
rect 25222 15552 25228 15564
rect 24443 15524 25228 15552
rect 24443 15521 24455 15524
rect 24397 15515 24455 15521
rect 25222 15512 25228 15524
rect 25280 15512 25286 15564
rect 20074 15487 20132 15493
rect 20074 15453 20086 15487
rect 20120 15453 20132 15487
rect 20074 15447 20132 15453
rect 20257 15487 20315 15493
rect 20257 15453 20269 15487
rect 20303 15453 20315 15487
rect 20257 15447 20315 15453
rect 12989 15419 13047 15425
rect 12989 15416 13001 15419
rect 9732 15388 9904 15416
rect 12544 15388 13001 15416
rect 9732 15376 9738 15388
rect 12544 15360 12572 15388
rect 12989 15385 13001 15388
rect 13035 15385 13047 15419
rect 12989 15379 13047 15385
rect 13722 15376 13728 15428
rect 13780 15416 13786 15428
rect 15470 15416 15476 15428
rect 13780 15388 15476 15416
rect 13780 15376 13786 15388
rect 15470 15376 15476 15388
rect 15528 15376 15534 15428
rect 15565 15419 15623 15425
rect 15565 15385 15577 15419
rect 15611 15416 15623 15419
rect 15746 15416 15752 15428
rect 15611 15388 15752 15416
rect 15611 15385 15623 15388
rect 15565 15379 15623 15385
rect 15746 15376 15752 15388
rect 15804 15376 15810 15428
rect 18322 15376 18328 15428
rect 18380 15416 18386 15428
rect 18509 15419 18567 15425
rect 18509 15416 18521 15419
rect 18380 15388 18521 15416
rect 18380 15376 18386 15388
rect 18509 15385 18521 15388
rect 18555 15385 18567 15419
rect 18509 15379 18567 15385
rect 18601 15419 18659 15425
rect 18601 15385 18613 15419
rect 18647 15385 18659 15419
rect 18601 15379 18659 15385
rect 6546 15308 6552 15360
rect 6604 15348 6610 15360
rect 7466 15348 7472 15360
rect 6604 15320 7472 15348
rect 6604 15308 6610 15320
rect 7466 15308 7472 15320
rect 7524 15308 7530 15360
rect 12526 15308 12532 15360
rect 12584 15308 12590 15360
rect 18616 15348 18644 15379
rect 18690 15376 18696 15428
rect 18748 15425 18754 15428
rect 18748 15419 18777 15425
rect 18765 15385 18777 15419
rect 19444 15416 19472 15444
rect 18748 15379 18777 15385
rect 18892 15388 19472 15416
rect 18748 15376 18754 15379
rect 18892 15348 18920 15388
rect 18616 15320 18920 15348
rect 18966 15308 18972 15360
rect 19024 15348 19030 15360
rect 19245 15351 19303 15357
rect 19245 15348 19257 15351
rect 19024 15320 19257 15348
rect 19024 15308 19030 15320
rect 19245 15317 19257 15320
rect 19291 15317 19303 15351
rect 19245 15311 19303 15317
rect 19334 15308 19340 15360
rect 19392 15348 19398 15360
rect 20088 15348 20116 15447
rect 20438 15444 20444 15496
rect 20496 15493 20502 15496
rect 20496 15484 20504 15493
rect 20496 15456 20541 15484
rect 20640 15456 20944 15484
rect 20496 15447 20504 15456
rect 20496 15444 20502 15447
rect 20346 15376 20352 15428
rect 20404 15416 20410 15428
rect 20640 15416 20668 15456
rect 20404 15388 20668 15416
rect 20809 15419 20867 15425
rect 20404 15376 20410 15388
rect 20809 15385 20821 15419
rect 20855 15385 20867 15419
rect 20916 15416 20944 15456
rect 21910 15444 21916 15496
rect 21968 15444 21974 15496
rect 24118 15444 24124 15496
rect 24176 15444 24182 15496
rect 25792 15484 25820 15660
rect 26142 15648 26148 15700
rect 26200 15648 26206 15700
rect 26602 15484 26608 15496
rect 25792 15470 26608 15484
rect 25806 15456 26608 15470
rect 26602 15444 26608 15456
rect 26660 15444 26666 15496
rect 27798 15444 27804 15496
rect 27856 15444 27862 15496
rect 22094 15416 22100 15428
rect 20916 15388 22100 15416
rect 20809 15379 20867 15385
rect 19392 15320 20116 15348
rect 20824 15348 20852 15379
rect 22094 15376 22100 15388
rect 22152 15376 22158 15428
rect 22370 15376 22376 15428
rect 22428 15376 22434 15428
rect 23382 15376 23388 15428
rect 23440 15376 23446 15428
rect 24670 15376 24676 15428
rect 24728 15376 24734 15428
rect 27890 15416 27896 15428
rect 25994 15388 27896 15416
rect 21450 15348 21456 15360
rect 20824 15320 21456 15348
rect 19392 15308 19398 15320
rect 21450 15308 21456 15320
rect 21508 15348 21514 15360
rect 25994 15348 26022 15388
rect 27890 15376 27896 15388
rect 27948 15376 27954 15428
rect 28077 15419 28135 15425
rect 28077 15385 28089 15419
rect 28123 15416 28135 15419
rect 28166 15416 28172 15428
rect 28123 15388 28172 15416
rect 28123 15385 28135 15388
rect 28077 15379 28135 15385
rect 28166 15376 28172 15388
rect 28224 15376 28230 15428
rect 21508 15320 26022 15348
rect 21508 15308 21514 15320
rect 27154 15308 27160 15360
rect 27212 15348 27218 15360
rect 27617 15351 27675 15357
rect 27617 15348 27629 15351
rect 27212 15320 27629 15348
rect 27212 15308 27218 15320
rect 27617 15317 27629 15320
rect 27663 15317 27675 15351
rect 27617 15311 27675 15317
rect 1104 15258 28704 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 28704 15258
rect 1104 15184 28704 15206
rect 7466 15104 7472 15156
rect 7524 15144 7530 15156
rect 9030 15144 9036 15156
rect 7524 15116 9036 15144
rect 7524 15104 7530 15116
rect 9030 15104 9036 15116
rect 9088 15104 9094 15156
rect 9582 15104 9588 15156
rect 9640 15104 9646 15156
rect 11885 15147 11943 15153
rect 11885 15113 11897 15147
rect 11931 15144 11943 15147
rect 12618 15144 12624 15156
rect 11931 15116 12624 15144
rect 11931 15113 11943 15116
rect 11885 15107 11943 15113
rect 12618 15104 12624 15116
rect 12676 15144 12682 15156
rect 12986 15144 12992 15156
rect 12676 15116 12992 15144
rect 12676 15104 12682 15116
rect 12986 15104 12992 15116
rect 13044 15104 13050 15156
rect 17862 15104 17868 15156
rect 17920 15144 17926 15156
rect 21637 15147 21695 15153
rect 17920 15116 19932 15144
rect 17920 15104 17926 15116
rect 6270 15036 6276 15088
rect 6328 15076 6334 15088
rect 8481 15079 8539 15085
rect 8481 15076 8493 15079
rect 6328 15048 8493 15076
rect 6328 15036 6334 15048
rect 8481 15045 8493 15048
rect 8527 15076 8539 15079
rect 9490 15076 9496 15088
rect 8527 15048 9496 15076
rect 8527 15045 8539 15048
rect 8481 15039 8539 15045
rect 9490 15036 9496 15048
rect 9548 15036 9554 15088
rect 12894 15036 12900 15088
rect 12952 15076 12958 15088
rect 13725 15079 13783 15085
rect 13725 15076 13737 15079
rect 12952 15048 13737 15076
rect 12952 15036 12958 15048
rect 13725 15045 13737 15048
rect 13771 15045 13783 15079
rect 13725 15039 13783 15045
rect 14090 15036 14096 15088
rect 14148 15036 14154 15088
rect 7006 14968 7012 15020
rect 7064 14968 7070 15020
rect 7193 15011 7251 15017
rect 7193 14977 7205 15011
rect 7239 15008 7251 15011
rect 7742 15008 7748 15020
rect 7239 14980 7748 15008
rect 7239 14977 7251 14980
rect 7193 14971 7251 14977
rect 7742 14968 7748 14980
rect 7800 15008 7806 15020
rect 8018 15008 8024 15020
rect 7800 14980 8024 15008
rect 7800 14968 7806 14980
rect 8018 14968 8024 14980
rect 8076 14968 8082 15020
rect 8386 14968 8392 15020
rect 8444 14968 8450 15020
rect 8665 15011 8723 15017
rect 8665 14977 8677 15011
rect 8711 15008 8723 15011
rect 9122 15008 9128 15020
rect 8711 14980 9128 15008
rect 8711 14977 8723 14980
rect 8665 14971 8723 14977
rect 7024 14940 7052 14968
rect 7650 14940 7656 14952
rect 7024 14912 7656 14940
rect 7650 14900 7656 14912
rect 7708 14900 7714 14952
rect 8680 14940 8708 14971
rect 9122 14968 9128 14980
rect 9180 14968 9186 15020
rect 9309 15011 9367 15017
rect 9309 14977 9321 15011
rect 9355 14977 9367 15011
rect 9309 14971 9367 14977
rect 8036 14912 8708 14940
rect 8036 14872 8064 14912
rect 9214 14900 9220 14952
rect 9272 14900 9278 14952
rect 9324 14940 9352 14971
rect 9582 14968 9588 15020
rect 9640 15008 9646 15020
rect 9674 15008 9680 15020
rect 9640 14980 9680 15008
rect 9640 14968 9646 14980
rect 9674 14968 9680 14980
rect 9732 14968 9738 15020
rect 9766 14968 9772 15020
rect 9824 14968 9830 15020
rect 10042 14968 10048 15020
rect 10100 14968 10106 15020
rect 15838 14968 15844 15020
rect 15896 14968 15902 15020
rect 16025 15011 16083 15017
rect 16025 14977 16037 15011
rect 16071 15008 16083 15011
rect 16206 15008 16212 15020
rect 16071 14980 16212 15008
rect 16071 14977 16083 14980
rect 16025 14971 16083 14977
rect 16206 14968 16212 14980
rect 16264 14968 16270 15020
rect 16482 14968 16488 15020
rect 16540 15008 16546 15020
rect 17221 15011 17279 15017
rect 17221 15008 17233 15011
rect 16540 14980 17233 15008
rect 16540 14968 16546 14980
rect 17221 14977 17233 14980
rect 17267 14977 17279 15011
rect 17221 14971 17279 14977
rect 17862 14968 17868 15020
rect 17920 14968 17926 15020
rect 19904 15017 19932 15116
rect 21637 15113 21649 15147
rect 21683 15144 21695 15147
rect 21910 15144 21916 15156
rect 21683 15116 21916 15144
rect 21683 15113 21695 15116
rect 21637 15107 21695 15113
rect 21910 15104 21916 15116
rect 21968 15104 21974 15156
rect 22189 15147 22247 15153
rect 22189 15113 22201 15147
rect 22235 15144 22247 15147
rect 22370 15144 22376 15156
rect 22235 15116 22376 15144
rect 22235 15113 22247 15116
rect 22189 15107 22247 15113
rect 22370 15104 22376 15116
rect 22428 15104 22434 15156
rect 22557 15147 22615 15153
rect 22557 15113 22569 15147
rect 22603 15144 22615 15147
rect 24118 15144 24124 15156
rect 22603 15116 24124 15144
rect 22603 15113 22615 15116
rect 22557 15107 22615 15113
rect 24118 15104 24124 15116
rect 24176 15104 24182 15156
rect 27801 15147 27859 15153
rect 27801 15113 27813 15147
rect 27847 15144 27859 15147
rect 28074 15144 28080 15156
rect 27847 15116 28080 15144
rect 27847 15113 27859 15116
rect 27801 15107 27859 15113
rect 28074 15104 28080 15116
rect 28132 15104 28138 15156
rect 23382 15076 23388 15088
rect 21390 15048 23388 15076
rect 23382 15036 23388 15048
rect 23440 15036 23446 15088
rect 27890 15036 27896 15088
rect 27948 15036 27954 15088
rect 19889 15011 19947 15017
rect 19274 14994 19748 15008
rect 19260 14980 19748 14994
rect 10060 14940 10088 14968
rect 9324 14912 10088 14940
rect 13354 14900 13360 14952
rect 13412 14900 13418 14952
rect 13633 14943 13691 14949
rect 13633 14909 13645 14943
rect 13679 14940 13691 14943
rect 13814 14940 13820 14952
rect 13679 14912 13820 14940
rect 13679 14909 13691 14912
rect 13633 14903 13691 14909
rect 13814 14900 13820 14912
rect 13872 14900 13878 14952
rect 16117 14943 16175 14949
rect 16117 14909 16129 14943
rect 16163 14940 16175 14943
rect 16669 14943 16727 14949
rect 16669 14940 16681 14943
rect 16163 14912 16681 14940
rect 16163 14909 16175 14912
rect 16117 14903 16175 14909
rect 16669 14909 16681 14912
rect 16715 14909 16727 14943
rect 16669 14903 16727 14909
rect 18141 14943 18199 14949
rect 18141 14909 18153 14943
rect 18187 14940 18199 14943
rect 18230 14940 18236 14952
rect 18187 14912 18236 14940
rect 18187 14909 18199 14912
rect 18141 14903 18199 14909
rect 18230 14900 18236 14912
rect 18288 14900 18294 14952
rect 18782 14900 18788 14952
rect 18840 14940 18846 14952
rect 19260 14940 19288 14980
rect 18840 14912 19288 14940
rect 18840 14900 18846 14912
rect 6840 14844 8064 14872
rect 6546 14764 6552 14816
rect 6604 14804 6610 14816
rect 6840 14813 6868 14844
rect 8110 14832 8116 14884
rect 8168 14872 8174 14884
rect 8849 14875 8907 14881
rect 8849 14872 8861 14875
rect 8168 14844 8861 14872
rect 8168 14832 8174 14844
rect 8849 14841 8861 14844
rect 8895 14872 8907 14875
rect 10318 14872 10324 14884
rect 8895 14844 10324 14872
rect 8895 14841 8907 14844
rect 8849 14835 8907 14841
rect 10318 14832 10324 14844
rect 10376 14832 10382 14884
rect 6825 14807 6883 14813
rect 6825 14804 6837 14807
rect 6604 14776 6837 14804
rect 6604 14764 6610 14776
rect 6825 14773 6837 14776
rect 6871 14773 6883 14807
rect 6825 14767 6883 14773
rect 7926 14764 7932 14816
rect 7984 14804 7990 14816
rect 8941 14807 8999 14813
rect 8941 14804 8953 14807
rect 7984 14776 8953 14804
rect 7984 14764 7990 14776
rect 8941 14773 8953 14776
rect 8987 14804 8999 14807
rect 9858 14804 9864 14816
rect 8987 14776 9864 14804
rect 8987 14773 8999 14776
rect 8941 14767 8999 14773
rect 9858 14764 9864 14776
rect 9916 14764 9922 14816
rect 9953 14807 10011 14813
rect 9953 14773 9965 14807
rect 9999 14804 10011 14807
rect 10042 14804 10048 14816
rect 9999 14776 10048 14804
rect 9999 14773 10011 14776
rect 9953 14767 10011 14773
rect 10042 14764 10048 14776
rect 10100 14804 10106 14816
rect 10410 14804 10416 14816
rect 10100 14776 10416 14804
rect 10100 14764 10106 14776
rect 10410 14764 10416 14776
rect 10468 14764 10474 14816
rect 15654 14764 15660 14816
rect 15712 14764 15718 14816
rect 19426 14764 19432 14816
rect 19484 14804 19490 14816
rect 19613 14807 19671 14813
rect 19613 14804 19625 14807
rect 19484 14776 19625 14804
rect 19484 14764 19490 14776
rect 19613 14773 19625 14776
rect 19659 14773 19671 14807
rect 19720 14804 19748 14980
rect 19889 14977 19901 15011
rect 19935 14977 19947 15011
rect 19889 14971 19947 14977
rect 22373 15011 22431 15017
rect 22373 14977 22385 15011
rect 22419 15008 22431 15011
rect 22462 15008 22468 15020
rect 22419 14980 22468 15008
rect 22419 14977 22431 14980
rect 22373 14971 22431 14977
rect 22462 14968 22468 14980
rect 22520 14968 22526 15020
rect 22646 14968 22652 15020
rect 22704 14968 22710 15020
rect 20165 14943 20223 14949
rect 20165 14909 20177 14943
rect 20211 14940 20223 14943
rect 20898 14940 20904 14952
rect 20211 14912 20904 14940
rect 20211 14909 20223 14912
rect 20165 14903 20223 14909
rect 20898 14900 20904 14912
rect 20956 14900 20962 14952
rect 20622 14804 20628 14816
rect 19720 14776 20628 14804
rect 19613 14767 19671 14773
rect 20622 14764 20628 14776
rect 20680 14764 20686 14816
rect 1104 14714 28704 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 28704 14714
rect 1104 14640 28704 14662
rect 6733 14603 6791 14609
rect 6733 14600 6745 14603
rect 5552 14572 6745 14600
rect 5442 14356 5448 14408
rect 5500 14356 5506 14408
rect 5552 14405 5580 14572
rect 6733 14569 6745 14572
rect 6779 14569 6791 14603
rect 6733 14563 6791 14569
rect 7006 14560 7012 14612
rect 7064 14600 7070 14612
rect 8294 14600 8300 14612
rect 7064 14572 8300 14600
rect 7064 14560 7070 14572
rect 8294 14560 8300 14572
rect 8352 14560 8358 14612
rect 8386 14560 8392 14612
rect 8444 14600 8450 14612
rect 8444 14572 9076 14600
rect 8444 14560 8450 14572
rect 8202 14492 8208 14544
rect 8260 14532 8266 14544
rect 8941 14535 8999 14541
rect 8941 14532 8953 14535
rect 8260 14504 8953 14532
rect 8260 14492 8266 14504
rect 8941 14501 8953 14504
rect 8987 14501 8999 14535
rect 9048 14532 9076 14572
rect 9766 14560 9772 14612
rect 9824 14600 9830 14612
rect 10229 14603 10287 14609
rect 10229 14600 10241 14603
rect 9824 14572 10241 14600
rect 9824 14560 9830 14572
rect 10229 14569 10241 14572
rect 10275 14569 10287 14603
rect 10229 14563 10287 14569
rect 11882 14560 11888 14612
rect 11940 14600 11946 14612
rect 13633 14603 13691 14609
rect 13633 14600 13645 14603
rect 11940 14572 13645 14600
rect 11940 14560 11946 14572
rect 13633 14569 13645 14572
rect 13679 14569 13691 14603
rect 13633 14563 13691 14569
rect 18230 14560 18236 14612
rect 18288 14560 18294 14612
rect 9048 14504 9812 14532
rect 8941 14495 8999 14501
rect 5626 14424 5632 14476
rect 5684 14464 5690 14476
rect 6457 14467 6515 14473
rect 6457 14464 6469 14467
rect 5684 14436 6469 14464
rect 5684 14424 5690 14436
rect 6457 14433 6469 14436
rect 6503 14464 6515 14467
rect 6638 14464 6644 14476
rect 6503 14436 6644 14464
rect 6503 14433 6515 14436
rect 6457 14427 6515 14433
rect 6638 14424 6644 14436
rect 6696 14424 6702 14476
rect 7466 14424 7472 14476
rect 7524 14424 7530 14476
rect 8294 14424 8300 14476
rect 8352 14464 8358 14476
rect 8352 14436 9260 14464
rect 8352 14424 8358 14436
rect 5537 14399 5595 14405
rect 5537 14365 5549 14399
rect 5583 14365 5595 14399
rect 5537 14359 5595 14365
rect 5813 14399 5871 14405
rect 5813 14365 5825 14399
rect 5859 14396 5871 14399
rect 5902 14396 5908 14408
rect 5859 14368 5908 14396
rect 5859 14365 5871 14368
rect 5813 14359 5871 14365
rect 5902 14356 5908 14368
rect 5960 14356 5966 14408
rect 6914 14356 6920 14408
rect 6972 14396 6978 14408
rect 7285 14399 7343 14405
rect 7285 14396 7297 14399
rect 6972 14368 7297 14396
rect 6972 14356 6978 14368
rect 7285 14365 7297 14368
rect 7331 14365 7343 14399
rect 7285 14359 7343 14365
rect 7650 14356 7656 14408
rect 7708 14356 7714 14408
rect 7742 14356 7748 14408
rect 7800 14356 7806 14408
rect 7926 14356 7932 14408
rect 7984 14356 7990 14408
rect 8110 14356 8116 14408
rect 8168 14356 8174 14408
rect 8202 14356 8208 14408
rect 8260 14356 8266 14408
rect 8478 14356 8484 14408
rect 8536 14356 8542 14408
rect 8570 14356 8576 14408
rect 8628 14356 8634 14408
rect 9232 14405 9260 14436
rect 9490 14424 9496 14476
rect 9548 14464 9554 14476
rect 9585 14467 9643 14473
rect 9585 14464 9597 14467
rect 9548 14436 9597 14464
rect 9548 14424 9554 14436
rect 9585 14433 9597 14436
rect 9631 14464 9643 14467
rect 9631 14436 9720 14464
rect 9631 14433 9643 14436
rect 9585 14427 9643 14433
rect 9125 14399 9183 14405
rect 9125 14365 9137 14399
rect 9171 14365 9183 14399
rect 9125 14359 9183 14365
rect 9217 14399 9275 14405
rect 9217 14365 9229 14399
rect 9263 14365 9275 14399
rect 9217 14359 9275 14365
rect 5629 14331 5687 14337
rect 5629 14297 5641 14331
rect 5675 14328 5687 14331
rect 8389 14331 8447 14337
rect 8389 14328 8401 14331
rect 5675 14300 8401 14328
rect 5675 14297 5687 14300
rect 5629 14291 5687 14297
rect 8389 14297 8401 14300
rect 8435 14328 8447 14331
rect 8662 14328 8668 14340
rect 8435 14300 8668 14328
rect 8435 14297 8447 14300
rect 8389 14291 8447 14297
rect 8662 14288 8668 14300
rect 8720 14288 8726 14340
rect 4706 14220 4712 14272
rect 4764 14260 4770 14272
rect 5261 14263 5319 14269
rect 5261 14260 5273 14263
rect 4764 14232 5273 14260
rect 4764 14220 4770 14232
rect 5261 14229 5273 14232
rect 5307 14229 5319 14263
rect 5261 14223 5319 14229
rect 5718 14220 5724 14272
rect 5776 14260 5782 14272
rect 5905 14263 5963 14269
rect 5905 14260 5917 14263
rect 5776 14232 5917 14260
rect 5776 14220 5782 14232
rect 5905 14229 5917 14232
rect 5951 14229 5963 14263
rect 5905 14223 5963 14229
rect 6270 14220 6276 14272
rect 6328 14220 6334 14272
rect 6362 14220 6368 14272
rect 6420 14220 6426 14272
rect 6822 14220 6828 14272
rect 6880 14260 6886 14272
rect 7469 14263 7527 14269
rect 7469 14260 7481 14263
rect 6880 14232 7481 14260
rect 6880 14220 6886 14232
rect 7469 14229 7481 14232
rect 7515 14229 7527 14263
rect 7469 14223 7527 14229
rect 8021 14263 8079 14269
rect 8021 14229 8033 14263
rect 8067 14260 8079 14263
rect 8294 14260 8300 14272
rect 8067 14232 8300 14260
rect 8067 14229 8079 14232
rect 8021 14223 8079 14229
rect 8294 14220 8300 14232
rect 8352 14220 8358 14272
rect 8754 14220 8760 14272
rect 8812 14220 8818 14272
rect 9140 14260 9168 14359
rect 9306 14356 9312 14408
rect 9364 14356 9370 14408
rect 9692 14405 9720 14436
rect 9677 14399 9735 14405
rect 9677 14365 9689 14399
rect 9723 14365 9735 14399
rect 9784 14396 9812 14504
rect 13354 14492 13360 14544
rect 13412 14532 13418 14544
rect 13449 14535 13507 14541
rect 13449 14532 13461 14535
rect 13412 14504 13461 14532
rect 13412 14492 13418 14504
rect 13449 14501 13461 14504
rect 13495 14501 13507 14535
rect 13449 14495 13507 14501
rect 18969 14535 19027 14541
rect 18969 14501 18981 14535
rect 19015 14501 19027 14535
rect 18969 14495 19027 14501
rect 9858 14424 9864 14476
rect 9916 14464 9922 14476
rect 11609 14467 11667 14473
rect 9916 14436 10548 14464
rect 9916 14424 9922 14436
rect 9784 14368 9904 14396
rect 9677 14359 9735 14365
rect 9398 14288 9404 14340
rect 9456 14337 9462 14340
rect 9876 14337 9904 14368
rect 9950 14356 9956 14408
rect 10008 14356 10014 14408
rect 10042 14356 10048 14408
rect 10100 14356 10106 14408
rect 10318 14356 10324 14408
rect 10376 14356 10382 14408
rect 10520 14405 10548 14436
rect 11609 14433 11621 14467
rect 11655 14464 11667 14467
rect 13814 14464 13820 14476
rect 11655 14436 13820 14464
rect 11655 14433 11667 14436
rect 11609 14427 11667 14433
rect 13814 14424 13820 14436
rect 13872 14424 13878 14476
rect 18984 14464 19012 14495
rect 19521 14467 19579 14473
rect 19521 14464 19533 14467
rect 18984 14436 19533 14464
rect 19521 14433 19533 14436
rect 19567 14433 19579 14467
rect 19521 14427 19579 14433
rect 26789 14467 26847 14473
rect 26789 14433 26801 14467
rect 26835 14464 26847 14467
rect 27982 14464 27988 14476
rect 26835 14436 27988 14464
rect 26835 14433 26847 14436
rect 26789 14427 26847 14433
rect 27982 14424 27988 14436
rect 28040 14424 28046 14476
rect 10505 14399 10563 14405
rect 10505 14365 10517 14399
rect 10551 14365 10563 14399
rect 10505 14359 10563 14365
rect 11330 14356 11336 14408
rect 11388 14356 11394 14408
rect 11514 14356 11520 14408
rect 11572 14356 11578 14408
rect 18138 14396 18144 14408
rect 13832 14368 18144 14396
rect 9456 14331 9485 14337
rect 9473 14297 9485 14331
rect 9456 14291 9485 14297
rect 9861 14331 9919 14337
rect 9861 14297 9873 14331
rect 9907 14328 9919 14331
rect 11425 14331 11483 14337
rect 9907 14300 10824 14328
rect 9907 14297 9919 14300
rect 9861 14291 9919 14297
rect 9456 14288 9462 14291
rect 10689 14263 10747 14269
rect 10689 14260 10701 14263
rect 9140 14232 10701 14260
rect 10689 14229 10701 14232
rect 10735 14229 10747 14263
rect 10796 14260 10824 14300
rect 11425 14297 11437 14331
rect 11471 14328 11483 14331
rect 11885 14331 11943 14337
rect 11885 14328 11897 14331
rect 11471 14300 11897 14328
rect 11471 14297 11483 14300
rect 11425 14291 11483 14297
rect 11885 14297 11897 14300
rect 11931 14297 11943 14331
rect 11885 14291 11943 14297
rect 12894 14288 12900 14340
rect 12952 14288 12958 14340
rect 13601 14331 13659 14337
rect 13601 14328 13613 14331
rect 13188 14300 13613 14328
rect 12158 14260 12164 14272
rect 10796 14232 12164 14260
rect 10689 14223 10747 14229
rect 12158 14220 12164 14232
rect 12216 14220 12222 14272
rect 12802 14220 12808 14272
rect 12860 14260 12866 14272
rect 13188 14260 13216 14300
rect 13601 14297 13613 14300
rect 13647 14297 13659 14331
rect 13601 14291 13659 14297
rect 13722 14288 13728 14340
rect 13780 14328 13786 14340
rect 13832 14337 13860 14368
rect 18138 14356 18144 14368
rect 18196 14356 18202 14408
rect 18325 14399 18383 14405
rect 18325 14365 18337 14399
rect 18371 14365 18383 14399
rect 18325 14359 18383 14365
rect 13817 14331 13875 14337
rect 13817 14328 13829 14331
rect 13780 14300 13829 14328
rect 13780 14288 13786 14300
rect 13817 14297 13829 14300
rect 13863 14297 13875 14331
rect 13817 14291 13875 14297
rect 15286 14288 15292 14340
rect 15344 14288 15350 14340
rect 18340 14328 18368 14359
rect 18690 14356 18696 14408
rect 18748 14356 18754 14408
rect 18785 14399 18843 14405
rect 18785 14365 18797 14399
rect 18831 14396 18843 14399
rect 18874 14396 18880 14408
rect 18831 14368 18880 14396
rect 18831 14365 18843 14368
rect 18785 14359 18843 14365
rect 18800 14328 18828 14359
rect 18874 14356 18880 14368
rect 18932 14356 18938 14408
rect 19242 14356 19248 14408
rect 19300 14356 19306 14408
rect 20622 14356 20628 14408
rect 20680 14356 20686 14408
rect 26510 14356 26516 14408
rect 26568 14356 26574 14408
rect 18340 14300 18828 14328
rect 18966 14288 18972 14340
rect 19024 14288 19030 14340
rect 28074 14328 28080 14340
rect 28014 14300 28080 14328
rect 28074 14288 28080 14300
rect 28132 14288 28138 14340
rect 12860 14232 13216 14260
rect 13357 14263 13415 14269
rect 12860 14220 12866 14232
rect 13357 14229 13369 14263
rect 13403 14260 13415 14263
rect 13446 14260 13452 14272
rect 13403 14232 13452 14260
rect 13403 14229 13415 14232
rect 13357 14223 13415 14229
rect 13446 14220 13452 14232
rect 13504 14220 13510 14272
rect 16390 14220 16396 14272
rect 16448 14260 16454 14272
rect 16577 14263 16635 14269
rect 16577 14260 16589 14263
rect 16448 14232 16589 14260
rect 16448 14220 16454 14232
rect 16577 14229 16589 14232
rect 16623 14229 16635 14263
rect 16577 14223 16635 14229
rect 20990 14220 20996 14272
rect 21048 14220 21054 14272
rect 27430 14220 27436 14272
rect 27488 14260 27494 14272
rect 28261 14263 28319 14269
rect 28261 14260 28273 14263
rect 27488 14232 28273 14260
rect 27488 14220 27494 14232
rect 28261 14229 28273 14232
rect 28307 14229 28319 14263
rect 28261 14223 28319 14229
rect 1104 14170 28704 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 28704 14170
rect 1104 14096 28704 14118
rect 5350 14056 5356 14068
rect 4448 14028 5356 14056
rect 4448 13929 4476 14028
rect 5350 14016 5356 14028
rect 5408 14016 5414 14068
rect 6181 14059 6239 14065
rect 6181 14025 6193 14059
rect 6227 14025 6239 14059
rect 6181 14019 6239 14025
rect 4706 13948 4712 14000
rect 4764 13948 4770 14000
rect 6196 13988 6224 14019
rect 6362 14016 6368 14068
rect 6420 14016 6426 14068
rect 11882 14016 11888 14068
rect 11940 14056 11946 14068
rect 12253 14059 12311 14065
rect 12253 14056 12265 14059
rect 11940 14028 12265 14056
rect 11940 14016 11946 14028
rect 12253 14025 12265 14028
rect 12299 14025 12311 14059
rect 12897 14059 12955 14065
rect 12897 14056 12909 14059
rect 12253 14019 12311 14025
rect 12452 14028 12909 14056
rect 6196 13960 6960 13988
rect 4433 13923 4491 13929
rect 4433 13889 4445 13923
rect 4479 13889 4491 13923
rect 4433 13883 4491 13889
rect 5810 13880 5816 13932
rect 5868 13880 5874 13932
rect 6546 13880 6552 13932
rect 6604 13880 6610 13932
rect 6641 13923 6699 13929
rect 6641 13889 6653 13923
rect 6687 13920 6699 13923
rect 6822 13920 6828 13932
rect 6687 13892 6828 13920
rect 6687 13889 6699 13892
rect 6641 13883 6699 13889
rect 6822 13880 6828 13892
rect 6880 13880 6886 13932
rect 6932 13864 6960 13960
rect 7006 13948 7012 14000
rect 7064 13948 7070 14000
rect 7742 13988 7748 14000
rect 7208 13960 7748 13988
rect 6914 13812 6920 13864
rect 6972 13812 6978 13864
rect 7208 13861 7236 13960
rect 7742 13948 7748 13960
rect 7800 13948 7806 14000
rect 8754 13948 8760 14000
rect 8812 13988 8818 14000
rect 8849 13991 8907 13997
rect 8849 13988 8861 13991
rect 8812 13960 8861 13988
rect 8812 13948 8818 13960
rect 8849 13957 8861 13960
rect 8895 13957 8907 13991
rect 8849 13951 8907 13957
rect 8938 13948 8944 14000
rect 8996 13988 9002 14000
rect 8996 13960 9338 13988
rect 8996 13948 9002 13960
rect 10134 13948 10140 14000
rect 10192 13988 10198 14000
rect 12452 13997 12480 14028
rect 12897 14025 12909 14028
rect 12943 14025 12955 14059
rect 12897 14019 12955 14025
rect 16482 14016 16488 14068
rect 16540 14016 16546 14068
rect 18966 14016 18972 14068
rect 19024 14016 19030 14068
rect 19978 14016 19984 14068
rect 20036 14056 20042 14068
rect 20622 14056 20628 14068
rect 20036 14028 20628 14056
rect 20036 14016 20042 14028
rect 20622 14016 20628 14028
rect 20680 14056 20686 14068
rect 26510 14056 26516 14068
rect 20680 14028 22508 14056
rect 20680 14016 20686 14028
rect 10597 13991 10655 13997
rect 10597 13988 10609 13991
rect 10192 13960 10609 13988
rect 10192 13948 10198 13960
rect 10597 13957 10609 13960
rect 10643 13957 10655 13991
rect 12437 13991 12495 13997
rect 12437 13988 12449 13991
rect 10597 13951 10655 13957
rect 12176 13960 12449 13988
rect 7561 13923 7619 13929
rect 7561 13920 7573 13923
rect 7300 13892 7573 13920
rect 7193 13855 7251 13861
rect 7193 13821 7205 13855
rect 7239 13821 7251 13855
rect 7193 13815 7251 13821
rect 6270 13744 6276 13796
rect 6328 13784 6334 13796
rect 6822 13784 6828 13796
rect 6328 13756 6828 13784
rect 6328 13744 6334 13756
rect 6822 13744 6828 13756
rect 6880 13784 6886 13796
rect 7300 13784 7328 13892
rect 7561 13889 7573 13892
rect 7607 13889 7619 13923
rect 8386 13920 8392 13932
rect 7561 13883 7619 13889
rect 7668 13892 8392 13920
rect 7668 13861 7696 13892
rect 8386 13880 8392 13892
rect 8444 13880 8450 13932
rect 11330 13880 11336 13932
rect 11388 13920 11394 13932
rect 12176 13929 12204 13960
rect 12437 13957 12449 13960
rect 12483 13957 12495 13991
rect 12437 13951 12495 13957
rect 12618 13948 12624 14000
rect 12676 13948 12682 14000
rect 12802 13948 12808 14000
rect 12860 13948 12866 14000
rect 13357 13991 13415 13997
rect 13357 13988 13369 13991
rect 12912 13960 13369 13988
rect 12161 13923 12219 13929
rect 12161 13920 12173 13923
rect 11388 13892 12173 13920
rect 11388 13880 11394 13892
rect 12161 13889 12173 13892
rect 12207 13889 12219 13923
rect 12161 13883 12219 13889
rect 12250 13880 12256 13932
rect 12308 13920 12314 13932
rect 12345 13923 12403 13929
rect 12345 13920 12357 13923
rect 12308 13892 12357 13920
rect 12308 13880 12314 13892
rect 12345 13889 12357 13892
rect 12391 13920 12403 13923
rect 12636 13920 12664 13948
rect 12391 13892 12664 13920
rect 12391 13889 12403 13892
rect 12345 13883 12403 13889
rect 7653 13855 7711 13861
rect 7653 13821 7665 13855
rect 7699 13821 7711 13855
rect 7653 13815 7711 13821
rect 8294 13812 8300 13864
rect 8352 13852 8358 13864
rect 8573 13855 8631 13861
rect 8573 13852 8585 13855
rect 8352 13824 8585 13852
rect 8352 13812 8358 13824
rect 8573 13821 8585 13824
rect 8619 13821 8631 13855
rect 8573 13815 8631 13821
rect 11514 13812 11520 13864
rect 11572 13852 11578 13864
rect 12912 13852 12940 13960
rect 13357 13957 13369 13960
rect 13403 13957 13415 13991
rect 16298 13988 16304 14000
rect 16238 13960 16304 13988
rect 13357 13951 13415 13957
rect 16298 13948 16304 13960
rect 16356 13948 16362 14000
rect 18690 13948 18696 14000
rect 18748 13988 18754 14000
rect 19889 13991 19947 13997
rect 19889 13988 19901 13991
rect 18748 13960 19901 13988
rect 18748 13948 18754 13960
rect 19889 13957 19901 13960
rect 19935 13957 19947 13991
rect 19889 13951 19947 13957
rect 22094 13948 22100 14000
rect 22152 13948 22158 14000
rect 13081 13923 13139 13929
rect 13081 13889 13093 13923
rect 13127 13889 13139 13923
rect 13081 13883 13139 13889
rect 13265 13923 13323 13929
rect 13265 13889 13277 13923
rect 13311 13920 13323 13923
rect 13538 13920 13544 13932
rect 13311 13892 13544 13920
rect 13311 13889 13323 13892
rect 13265 13883 13323 13889
rect 11572 13824 12940 13852
rect 11572 13812 11578 13824
rect 6880 13756 7328 13784
rect 6880 13744 6886 13756
rect 12158 13744 12164 13796
rect 12216 13784 12222 13796
rect 12894 13784 12900 13796
rect 12216 13756 12900 13784
rect 12216 13744 12222 13756
rect 12894 13744 12900 13756
rect 12952 13744 12958 13796
rect 13096 13784 13124 13883
rect 13538 13880 13544 13892
rect 13596 13920 13602 13932
rect 13633 13923 13691 13929
rect 13633 13920 13645 13923
rect 13596 13892 13645 13920
rect 13596 13880 13602 13892
rect 13633 13889 13645 13892
rect 13679 13889 13691 13923
rect 13633 13883 13691 13889
rect 13814 13880 13820 13932
rect 13872 13920 13878 13932
rect 14737 13923 14795 13929
rect 14737 13920 14749 13923
rect 13872 13892 14749 13920
rect 13872 13880 13878 13892
rect 14737 13889 14749 13892
rect 14783 13889 14795 13923
rect 14737 13883 14795 13889
rect 17678 13880 17684 13932
rect 17736 13880 17742 13932
rect 19245 13923 19303 13929
rect 19245 13889 19257 13923
rect 19291 13920 19303 13923
rect 19426 13920 19432 13932
rect 19291 13892 19432 13920
rect 19291 13889 19303 13892
rect 19245 13883 19303 13889
rect 19426 13880 19432 13892
rect 19484 13880 19490 13932
rect 21910 13880 21916 13932
rect 21968 13929 21974 13932
rect 21968 13923 22017 13929
rect 21968 13889 21971 13923
rect 22005 13889 22017 13923
rect 21968 13883 22017 13889
rect 21968 13880 21974 13883
rect 22186 13880 22192 13932
rect 22244 13880 22250 13932
rect 22480 13929 22508 14028
rect 24136 14028 26516 14056
rect 24136 13929 24164 14028
rect 26510 14016 26516 14028
rect 26568 14016 26574 14068
rect 27522 14016 27528 14068
rect 27580 14056 27586 14068
rect 27801 14059 27859 14065
rect 27801 14056 27813 14059
rect 27580 14028 27813 14056
rect 27580 14016 27586 14028
rect 27801 14025 27813 14028
rect 27847 14025 27859 14059
rect 27801 14019 27859 14025
rect 28258 14016 28264 14068
rect 28316 14016 28322 14068
rect 27062 13948 27068 14000
rect 27120 13988 27126 14000
rect 27120 13960 27568 13988
rect 27120 13948 27126 13960
rect 22317 13923 22375 13929
rect 22317 13920 22329 13923
rect 22296 13889 22329 13920
rect 22363 13889 22375 13923
rect 22296 13883 22375 13889
rect 22465 13923 22523 13929
rect 22465 13889 22477 13923
rect 22511 13889 22523 13923
rect 22465 13883 22523 13889
rect 24121 13923 24179 13929
rect 24121 13889 24133 13923
rect 24167 13889 24179 13923
rect 24121 13883 24179 13889
rect 13357 13855 13415 13861
rect 13357 13821 13369 13855
rect 13403 13852 13415 13855
rect 13722 13852 13728 13864
rect 13403 13824 13728 13852
rect 13403 13821 13415 13824
rect 13357 13815 13415 13821
rect 13722 13812 13728 13824
rect 13780 13812 13786 13864
rect 15013 13855 15071 13861
rect 15013 13821 15025 13855
rect 15059 13852 15071 13855
rect 15654 13852 15660 13864
rect 15059 13824 15660 13852
rect 15059 13821 15071 13824
rect 15013 13815 15071 13821
rect 15654 13812 15660 13824
rect 15712 13812 15718 13864
rect 16574 13812 16580 13864
rect 16632 13852 16638 13864
rect 16669 13855 16727 13861
rect 16669 13852 16681 13855
rect 16632 13824 16681 13852
rect 16632 13812 16638 13824
rect 16669 13821 16681 13824
rect 16715 13821 16727 13855
rect 16669 13815 16727 13821
rect 17313 13855 17371 13861
rect 17313 13821 17325 13855
rect 17359 13852 17371 13855
rect 17405 13855 17463 13861
rect 17405 13852 17417 13855
rect 17359 13824 17417 13852
rect 17359 13821 17371 13824
rect 17313 13815 17371 13821
rect 17405 13821 17417 13824
rect 17451 13821 17463 13855
rect 17405 13815 17463 13821
rect 17497 13855 17555 13861
rect 17497 13821 17509 13855
rect 17543 13852 17555 13855
rect 17543 13824 18092 13852
rect 17543 13821 17555 13824
rect 17497 13815 17555 13821
rect 18064 13784 18092 13824
rect 18138 13812 18144 13864
rect 18196 13852 18202 13864
rect 18969 13855 19027 13861
rect 18969 13852 18981 13855
rect 18196 13824 18981 13852
rect 18196 13812 18202 13824
rect 18969 13821 18981 13824
rect 19015 13821 19027 13855
rect 18969 13815 19027 13821
rect 19150 13812 19156 13864
rect 19208 13852 19214 13864
rect 20441 13855 20499 13861
rect 20441 13852 20453 13855
rect 19208 13824 20453 13852
rect 19208 13812 19214 13824
rect 20441 13821 20453 13824
rect 20487 13852 20499 13855
rect 20990 13852 20996 13864
rect 20487 13824 20996 13852
rect 20487 13821 20499 13824
rect 20441 13815 20499 13821
rect 20990 13812 20996 13824
rect 21048 13812 21054 13864
rect 22296 13852 22324 13883
rect 25498 13880 25504 13932
rect 25556 13880 25562 13932
rect 27249 13923 27307 13929
rect 27249 13889 27261 13923
rect 27295 13920 27307 13923
rect 27430 13920 27436 13932
rect 27295 13892 27436 13920
rect 27295 13889 27307 13892
rect 27249 13883 27307 13889
rect 27430 13880 27436 13892
rect 27488 13880 27494 13932
rect 27540 13929 27568 13960
rect 27525 13923 27583 13929
rect 27525 13889 27537 13923
rect 27571 13889 27583 13923
rect 27525 13883 27583 13889
rect 27982 13880 27988 13932
rect 28040 13880 28046 13932
rect 28077 13923 28135 13929
rect 28077 13889 28089 13923
rect 28123 13889 28135 13923
rect 28077 13883 28135 13889
rect 22112 13824 22324 13852
rect 18874 13784 18880 13796
rect 13096 13756 13400 13784
rect 18064 13756 18880 13784
rect 13372 13728 13400 13756
rect 18874 13744 18880 13756
rect 18932 13744 18938 13796
rect 13354 13676 13360 13728
rect 13412 13716 13418 13728
rect 13541 13719 13599 13725
rect 13541 13716 13553 13719
rect 13412 13688 13553 13716
rect 13412 13676 13418 13688
rect 13541 13685 13553 13688
rect 13587 13685 13599 13719
rect 13541 13679 13599 13685
rect 17586 13676 17592 13728
rect 17644 13716 17650 13728
rect 17865 13719 17923 13725
rect 17865 13716 17877 13719
rect 17644 13688 17877 13716
rect 17644 13676 17650 13688
rect 17865 13685 17877 13688
rect 17911 13685 17923 13719
rect 17865 13679 17923 13685
rect 19058 13676 19064 13728
rect 19116 13716 19122 13728
rect 19168 13725 19196 13812
rect 22112 13796 22140 13824
rect 25406 13812 25412 13864
rect 25464 13852 25470 13864
rect 25869 13855 25927 13861
rect 25869 13852 25881 13855
rect 25464 13824 25881 13852
rect 25464 13812 25470 13824
rect 25869 13821 25881 13824
rect 25915 13821 25927 13855
rect 25869 13815 25927 13821
rect 27338 13812 27344 13864
rect 27396 13812 27402 13864
rect 27709 13855 27767 13861
rect 27709 13821 27721 13855
rect 27755 13852 27767 13855
rect 28092 13852 28120 13883
rect 27755 13824 28120 13852
rect 27755 13821 27767 13824
rect 27709 13815 27767 13821
rect 22094 13744 22100 13796
rect 22152 13744 22158 13796
rect 27433 13787 27491 13793
rect 27433 13753 27445 13787
rect 27479 13784 27491 13787
rect 27614 13784 27620 13796
rect 27479 13756 27620 13784
rect 27479 13753 27491 13756
rect 27433 13747 27491 13753
rect 27614 13744 27620 13756
rect 27672 13744 27678 13796
rect 19153 13719 19211 13725
rect 19153 13716 19165 13719
rect 19116 13688 19165 13716
rect 19116 13676 19122 13688
rect 19153 13685 19165 13688
rect 19199 13685 19211 13719
rect 19153 13679 19211 13685
rect 21821 13719 21879 13725
rect 21821 13685 21833 13719
rect 21867 13716 21879 13719
rect 22002 13716 22008 13728
rect 21867 13688 22008 13716
rect 21867 13685 21879 13688
rect 21821 13679 21879 13685
rect 22002 13676 22008 13688
rect 22060 13676 22066 13728
rect 24384 13719 24442 13725
rect 24384 13685 24396 13719
rect 24430 13716 24442 13719
rect 24854 13716 24860 13728
rect 24430 13688 24860 13716
rect 24430 13685 24442 13688
rect 24384 13679 24442 13685
rect 24854 13676 24860 13688
rect 24912 13676 24918 13728
rect 1104 13626 28704 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 28704 13626
rect 1104 13552 28704 13574
rect 6822 13472 6828 13524
rect 6880 13472 6886 13524
rect 15930 13472 15936 13524
rect 15988 13472 15994 13524
rect 16117 13515 16175 13521
rect 16117 13481 16129 13515
rect 16163 13512 16175 13515
rect 16574 13512 16580 13524
rect 16163 13484 16580 13512
rect 16163 13481 16175 13484
rect 16117 13475 16175 13481
rect 16574 13472 16580 13484
rect 16632 13472 16638 13524
rect 16482 13404 16488 13456
rect 16540 13404 16546 13456
rect 5077 13379 5135 13385
rect 5077 13345 5089 13379
rect 5123 13376 5135 13379
rect 5350 13376 5356 13388
rect 5123 13348 5356 13376
rect 5123 13345 5135 13348
rect 5077 13339 5135 13345
rect 5350 13336 5356 13348
rect 5408 13336 5414 13388
rect 15654 13376 15660 13388
rect 15304 13348 15660 13376
rect 15194 13268 15200 13320
rect 15252 13308 15258 13320
rect 15304 13317 15332 13348
rect 15654 13336 15660 13348
rect 15712 13336 15718 13388
rect 16500 13376 16528 13404
rect 16408 13348 16528 13376
rect 15289 13311 15347 13317
rect 15289 13308 15301 13311
rect 15252 13280 15301 13308
rect 15252 13268 15258 13280
rect 15289 13277 15301 13280
rect 15335 13277 15347 13311
rect 15289 13271 15347 13277
rect 15382 13311 15440 13317
rect 15382 13277 15394 13311
rect 15428 13277 15440 13311
rect 15382 13271 15440 13277
rect 5353 13243 5411 13249
rect 5353 13209 5365 13243
rect 5399 13240 5411 13243
rect 5626 13240 5632 13252
rect 5399 13212 5632 13240
rect 5399 13209 5411 13212
rect 5353 13203 5411 13209
rect 5626 13200 5632 13212
rect 5684 13200 5690 13252
rect 5810 13240 5816 13252
rect 5736 13212 5816 13240
rect 4614 13132 4620 13184
rect 4672 13172 4678 13184
rect 5736 13172 5764 13212
rect 5810 13200 5816 13212
rect 5868 13200 5874 13252
rect 14458 13200 14464 13252
rect 14516 13240 14522 13252
rect 15396 13240 15424 13271
rect 15470 13268 15476 13320
rect 15528 13308 15534 13320
rect 15565 13311 15623 13317
rect 15565 13308 15577 13311
rect 15528 13280 15577 13308
rect 15528 13268 15534 13280
rect 15565 13277 15577 13280
rect 15611 13277 15623 13311
rect 15565 13271 15623 13277
rect 15795 13311 15853 13317
rect 15795 13277 15807 13311
rect 15841 13308 15853 13311
rect 16408 13308 16436 13348
rect 17586 13336 17592 13388
rect 17644 13336 17650 13388
rect 17865 13379 17923 13385
rect 17865 13345 17877 13379
rect 17911 13376 17923 13379
rect 19242 13376 19248 13388
rect 17911 13348 19248 13376
rect 17911 13345 17923 13348
rect 17865 13339 17923 13345
rect 19242 13336 19248 13348
rect 19300 13336 19306 13388
rect 26510 13336 26516 13388
rect 26568 13336 26574 13388
rect 26789 13379 26847 13385
rect 26789 13345 26801 13379
rect 26835 13376 26847 13379
rect 27798 13376 27804 13388
rect 26835 13348 27804 13376
rect 26835 13345 26847 13348
rect 26789 13339 26847 13345
rect 27798 13336 27804 13348
rect 27856 13336 27862 13388
rect 15841 13280 16436 13308
rect 15841 13277 15853 13280
rect 15795 13271 15853 13277
rect 21542 13268 21548 13320
rect 21600 13268 21606 13320
rect 23937 13311 23995 13317
rect 23937 13308 23949 13311
rect 23308 13280 23949 13308
rect 14516 13212 15424 13240
rect 15657 13243 15715 13249
rect 14516 13200 14522 13212
rect 15657 13209 15669 13243
rect 15703 13240 15715 13243
rect 15703 13212 15792 13240
rect 15703 13209 15715 13212
rect 15657 13203 15715 13209
rect 15764 13184 15792 13212
rect 17126 13200 17132 13252
rect 17184 13200 17190 13252
rect 21818 13200 21824 13252
rect 21876 13200 21882 13252
rect 23198 13240 23204 13252
rect 23046 13212 23204 13240
rect 23198 13200 23204 13212
rect 23256 13200 23262 13252
rect 4672 13144 5764 13172
rect 4672 13132 4678 13144
rect 15746 13132 15752 13184
rect 15804 13132 15810 13184
rect 22186 13132 22192 13184
rect 22244 13172 22250 13184
rect 23308 13181 23336 13280
rect 23937 13277 23949 13280
rect 23983 13277 23995 13311
rect 23937 13271 23995 13277
rect 27798 13200 27804 13252
rect 27856 13200 27862 13252
rect 23293 13175 23351 13181
rect 23293 13172 23305 13175
rect 22244 13144 23305 13172
rect 22244 13132 22250 13144
rect 23293 13141 23305 13144
rect 23339 13141 23351 13175
rect 23293 13135 23351 13141
rect 23382 13132 23388 13184
rect 23440 13132 23446 13184
rect 26970 13132 26976 13184
rect 27028 13172 27034 13184
rect 28261 13175 28319 13181
rect 28261 13172 28273 13175
rect 27028 13144 28273 13172
rect 27028 13132 27034 13144
rect 28261 13141 28273 13144
rect 28307 13141 28319 13175
rect 28261 13135 28319 13141
rect 1104 13082 28704 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 28704 13082
rect 1104 13008 28704 13030
rect 12894 12968 12900 12980
rect 12728 12940 12900 12968
rect 12250 12860 12256 12912
rect 12308 12900 12314 12912
rect 12728 12909 12756 12940
rect 12894 12928 12900 12940
rect 12952 12928 12958 12980
rect 13541 12971 13599 12977
rect 13541 12937 13553 12971
rect 13587 12968 13599 12971
rect 13722 12968 13728 12980
rect 13587 12940 13728 12968
rect 13587 12937 13599 12940
rect 13541 12931 13599 12937
rect 13722 12928 13728 12940
rect 13780 12928 13786 12980
rect 15378 12928 15384 12980
rect 15436 12968 15442 12980
rect 15565 12971 15623 12977
rect 15565 12968 15577 12971
rect 15436 12940 15577 12968
rect 15436 12928 15442 12940
rect 15565 12937 15577 12940
rect 15611 12937 15623 12971
rect 15565 12931 15623 12937
rect 15838 12928 15844 12980
rect 15896 12968 15902 12980
rect 16301 12971 16359 12977
rect 16301 12968 16313 12971
rect 15896 12940 16313 12968
rect 15896 12928 15902 12940
rect 16301 12937 16313 12940
rect 16347 12937 16359 12971
rect 16301 12931 16359 12937
rect 17678 12928 17684 12980
rect 17736 12968 17742 12980
rect 17773 12971 17831 12977
rect 17773 12968 17785 12971
rect 17736 12940 17785 12968
rect 17736 12928 17742 12940
rect 17773 12937 17785 12940
rect 17819 12937 17831 12971
rect 17773 12931 17831 12937
rect 21818 12928 21824 12980
rect 21876 12928 21882 12980
rect 27893 12971 27951 12977
rect 27893 12968 27905 12971
rect 27448 12940 27905 12968
rect 27448 12912 27476 12940
rect 27893 12937 27905 12940
rect 27939 12937 27951 12971
rect 27893 12931 27951 12937
rect 12621 12903 12679 12909
rect 12621 12900 12633 12903
rect 12308 12872 12633 12900
rect 12308 12860 12314 12872
rect 12621 12869 12633 12872
rect 12667 12869 12679 12903
rect 12621 12863 12679 12869
rect 12713 12903 12771 12909
rect 12713 12869 12725 12903
rect 12759 12869 12771 12903
rect 12713 12863 12771 12869
rect 12820 12872 14582 12900
rect 11606 12792 11612 12844
rect 11664 12832 11670 12844
rect 11885 12835 11943 12841
rect 11885 12832 11897 12835
rect 11664 12804 11897 12832
rect 11664 12792 11670 12804
rect 11885 12801 11897 12804
rect 11931 12801 11943 12835
rect 11885 12795 11943 12801
rect 12529 12835 12587 12841
rect 12529 12801 12541 12835
rect 12575 12801 12587 12835
rect 12529 12795 12587 12801
rect 11698 12724 11704 12776
rect 11756 12764 11762 12776
rect 12342 12764 12348 12776
rect 11756 12736 12348 12764
rect 11756 12724 11762 12736
rect 12342 12724 12348 12736
rect 12400 12764 12406 12776
rect 12544 12764 12572 12795
rect 12400 12736 12572 12764
rect 12400 12724 12406 12736
rect 10962 12656 10968 12708
rect 11020 12696 11026 12708
rect 12820 12696 12848 12872
rect 15470 12860 15476 12912
rect 15528 12900 15534 12912
rect 15933 12903 15991 12909
rect 15933 12900 15945 12903
rect 15528 12872 15945 12900
rect 15528 12860 15534 12872
rect 15933 12869 15945 12872
rect 15979 12869 15991 12903
rect 17405 12903 17463 12909
rect 15933 12863 15991 12869
rect 17144 12872 17356 12900
rect 12897 12835 12955 12841
rect 12897 12801 12909 12835
rect 12943 12801 12955 12835
rect 12897 12795 12955 12801
rect 12912 12764 12940 12795
rect 13078 12792 13084 12844
rect 13136 12832 13142 12844
rect 13725 12835 13783 12841
rect 13725 12832 13737 12835
rect 13136 12804 13737 12832
rect 13136 12792 13142 12804
rect 13725 12801 13737 12804
rect 13771 12801 13783 12835
rect 13725 12795 13783 12801
rect 13814 12792 13820 12844
rect 13872 12792 13878 12844
rect 15654 12792 15660 12844
rect 15712 12792 15718 12844
rect 15750 12835 15808 12841
rect 15750 12801 15762 12835
rect 15796 12801 15808 12835
rect 15750 12795 15808 12801
rect 13262 12764 13268 12776
rect 12912 12736 13268 12764
rect 13262 12724 13268 12736
rect 13320 12764 13326 12776
rect 13538 12764 13544 12776
rect 13320 12736 13544 12764
rect 13320 12724 13326 12736
rect 13538 12724 13544 12736
rect 13596 12724 13602 12776
rect 14090 12724 14096 12776
rect 14148 12724 14154 12776
rect 14550 12724 14556 12776
rect 14608 12764 14614 12776
rect 15764 12764 15792 12795
rect 15838 12792 15844 12844
rect 15896 12832 15902 12844
rect 16025 12835 16083 12841
rect 16025 12832 16037 12835
rect 15896 12804 16037 12832
rect 15896 12792 15902 12804
rect 16025 12801 16037 12804
rect 16071 12801 16083 12835
rect 16025 12795 16083 12801
rect 16163 12835 16221 12841
rect 16163 12801 16175 12835
rect 16209 12832 16221 12835
rect 16574 12832 16580 12844
rect 16209 12804 16580 12832
rect 16209 12801 16221 12804
rect 16163 12795 16221 12801
rect 16574 12792 16580 12804
rect 16632 12792 16638 12844
rect 17144 12841 17172 12872
rect 17129 12835 17187 12841
rect 17129 12801 17141 12835
rect 17175 12801 17187 12835
rect 17129 12795 17187 12801
rect 17222 12835 17280 12841
rect 17222 12801 17234 12835
rect 17268 12801 17280 12835
rect 17222 12795 17280 12801
rect 14608 12736 15792 12764
rect 14608 12724 14614 12736
rect 16482 12724 16488 12776
rect 16540 12764 16546 12776
rect 17236 12764 17264 12795
rect 16540 12736 17264 12764
rect 16540 12724 16546 12736
rect 11020 12668 12848 12696
rect 11020 12656 11026 12668
rect 5902 12588 5908 12640
rect 5960 12628 5966 12640
rect 11054 12628 11060 12640
rect 5960 12600 11060 12628
rect 5960 12588 5966 12600
rect 11054 12588 11060 12600
rect 11112 12588 11118 12640
rect 11422 12588 11428 12640
rect 11480 12628 11486 12640
rect 11701 12631 11759 12637
rect 11701 12628 11713 12631
rect 11480 12600 11713 12628
rect 11480 12588 11486 12600
rect 11701 12597 11713 12600
rect 11747 12597 11759 12631
rect 11701 12591 11759 12597
rect 12345 12631 12403 12637
rect 12345 12597 12357 12631
rect 12391 12628 12403 12631
rect 12434 12628 12440 12640
rect 12391 12600 12440 12628
rect 12391 12597 12403 12600
rect 12345 12591 12403 12597
rect 12434 12588 12440 12600
rect 12492 12628 12498 12640
rect 12802 12628 12808 12640
rect 12492 12600 12808 12628
rect 12492 12588 12498 12600
rect 12802 12588 12808 12600
rect 12860 12588 12866 12640
rect 17328 12628 17356 12872
rect 17405 12869 17417 12903
rect 17451 12900 17463 12903
rect 18690 12900 18696 12912
rect 17451 12872 18696 12900
rect 17451 12869 17463 12872
rect 17405 12863 17463 12869
rect 18690 12860 18696 12872
rect 18748 12860 18754 12912
rect 23382 12900 23388 12912
rect 22296 12872 23388 12900
rect 17497 12835 17555 12841
rect 17497 12801 17509 12835
rect 17543 12801 17555 12835
rect 17497 12795 17555 12801
rect 17635 12835 17693 12841
rect 17635 12801 17647 12835
rect 17681 12832 17693 12835
rect 19150 12832 19156 12844
rect 17681 12804 19156 12832
rect 17681 12801 17693 12804
rect 17635 12795 17693 12801
rect 17512 12764 17540 12795
rect 19150 12792 19156 12804
rect 19208 12832 19214 12844
rect 19521 12835 19579 12841
rect 19521 12832 19533 12835
rect 19208 12804 19533 12832
rect 19208 12792 19214 12804
rect 19521 12801 19533 12804
rect 19567 12801 19579 12835
rect 19521 12795 19579 12801
rect 20717 12835 20775 12841
rect 20717 12801 20729 12835
rect 20763 12832 20775 12835
rect 21174 12832 21180 12844
rect 20763 12804 21180 12832
rect 20763 12801 20775 12804
rect 20717 12795 20775 12801
rect 21174 12792 21180 12804
rect 21232 12792 21238 12844
rect 22002 12792 22008 12844
rect 22060 12792 22066 12844
rect 22296 12841 22324 12872
rect 23382 12860 23388 12872
rect 23440 12860 23446 12912
rect 26786 12900 26792 12912
rect 25714 12872 26792 12900
rect 26786 12860 26792 12872
rect 26844 12860 26850 12912
rect 27430 12860 27436 12912
rect 27488 12860 27494 12912
rect 22281 12835 22339 12841
rect 22281 12801 22293 12835
rect 22327 12801 22339 12835
rect 22554 12832 22560 12844
rect 22281 12795 22339 12801
rect 22388 12804 22560 12832
rect 18414 12764 18420 12776
rect 17512 12736 18420 12764
rect 18414 12724 18420 12736
rect 18472 12724 18478 12776
rect 19702 12724 19708 12776
rect 19760 12724 19766 12776
rect 20349 12767 20407 12773
rect 20349 12733 20361 12767
rect 20395 12764 20407 12767
rect 20441 12767 20499 12773
rect 20441 12764 20453 12767
rect 20395 12736 20453 12764
rect 20395 12733 20407 12736
rect 20349 12727 20407 12733
rect 20441 12733 20453 12736
rect 20487 12733 20499 12767
rect 22189 12767 22247 12773
rect 22189 12764 22201 12767
rect 20441 12727 20499 12733
rect 22066 12736 22201 12764
rect 18874 12656 18880 12708
rect 18932 12696 18938 12708
rect 20533 12699 20591 12705
rect 20533 12696 20545 12699
rect 18932 12668 20545 12696
rect 18932 12656 18938 12668
rect 20533 12665 20545 12668
rect 20579 12696 20591 12699
rect 22066 12696 22094 12736
rect 22189 12733 22201 12736
rect 22235 12764 22247 12767
rect 22388 12764 22416 12804
rect 22554 12792 22560 12804
rect 22612 12832 22618 12844
rect 22612 12804 22784 12832
rect 22612 12792 22618 12804
rect 22235 12736 22416 12764
rect 22465 12767 22523 12773
rect 22235 12733 22247 12736
rect 22189 12727 22247 12733
rect 22465 12733 22477 12767
rect 22511 12764 22523 12767
rect 22646 12764 22652 12776
rect 22511 12736 22652 12764
rect 22511 12733 22523 12736
rect 22465 12727 22523 12733
rect 22646 12724 22652 12736
rect 22704 12724 22710 12776
rect 22756 12764 22784 12804
rect 23290 12792 23296 12844
rect 23348 12792 23354 12844
rect 26421 12835 26479 12841
rect 26421 12801 26433 12835
rect 26467 12832 26479 12835
rect 26510 12832 26516 12844
rect 26467 12804 26516 12832
rect 26467 12801 26479 12804
rect 26421 12795 26479 12801
rect 26510 12792 26516 12804
rect 26568 12792 26574 12844
rect 26602 12792 26608 12844
rect 26660 12832 26666 12844
rect 27157 12835 27215 12841
rect 27157 12832 27169 12835
rect 26660 12804 27169 12832
rect 26660 12792 26666 12804
rect 27157 12801 27169 12804
rect 27203 12832 27215 12835
rect 27203 12804 27660 12832
rect 27203 12801 27215 12804
rect 27157 12795 27215 12801
rect 23569 12767 23627 12773
rect 22756 12736 23520 12764
rect 20579 12668 22094 12696
rect 20579 12665 20591 12668
rect 20533 12659 20591 12665
rect 22738 12656 22744 12708
rect 22796 12696 22802 12708
rect 23109 12699 23167 12705
rect 23109 12696 23121 12699
rect 22796 12668 23121 12696
rect 22796 12656 22802 12668
rect 23109 12665 23121 12668
rect 23155 12665 23167 12699
rect 23109 12659 23167 12665
rect 23492 12640 23520 12736
rect 23569 12733 23581 12767
rect 23615 12764 23627 12767
rect 23753 12767 23811 12773
rect 23753 12764 23765 12767
rect 23615 12736 23765 12764
rect 23615 12733 23627 12736
rect 23569 12727 23627 12733
rect 23753 12733 23765 12736
rect 23799 12733 23811 12767
rect 23753 12727 23811 12733
rect 24210 12724 24216 12776
rect 24268 12764 24274 12776
rect 24305 12767 24363 12773
rect 24305 12764 24317 12767
rect 24268 12736 24317 12764
rect 24268 12724 24274 12736
rect 24305 12733 24317 12736
rect 24351 12733 24363 12767
rect 24305 12727 24363 12733
rect 26145 12767 26203 12773
rect 26145 12733 26157 12767
rect 26191 12764 26203 12767
rect 27341 12767 27399 12773
rect 27341 12764 27353 12767
rect 26191 12736 27353 12764
rect 26191 12733 26203 12736
rect 26145 12727 26203 12733
rect 27341 12733 27353 12736
rect 27387 12764 27399 12767
rect 27522 12764 27528 12776
rect 27387 12736 27528 12764
rect 27387 12733 27399 12736
rect 27341 12727 27399 12733
rect 27522 12724 27528 12736
rect 27580 12724 27586 12776
rect 27632 12696 27660 12804
rect 28074 12792 28080 12844
rect 28132 12792 28138 12844
rect 28350 12792 28356 12844
rect 28408 12792 28414 12844
rect 28169 12699 28227 12705
rect 28169 12696 28181 12699
rect 27632 12668 28181 12696
rect 28169 12665 28181 12668
rect 28215 12665 28227 12699
rect 28169 12659 28227 12665
rect 18414 12628 18420 12640
rect 17328 12600 18420 12628
rect 18414 12588 18420 12600
rect 18472 12588 18478 12640
rect 18966 12588 18972 12640
rect 19024 12588 19030 12640
rect 20714 12588 20720 12640
rect 20772 12628 20778 12640
rect 20901 12631 20959 12637
rect 20901 12628 20913 12631
rect 20772 12600 20913 12628
rect 20772 12588 20778 12600
rect 20901 12597 20913 12600
rect 20947 12597 20959 12631
rect 20901 12591 20959 12597
rect 22278 12588 22284 12640
rect 22336 12628 22342 12640
rect 23017 12631 23075 12637
rect 23017 12628 23029 12631
rect 22336 12600 23029 12628
rect 22336 12588 22342 12600
rect 23017 12597 23029 12600
rect 23063 12597 23075 12631
rect 23017 12591 23075 12597
rect 23474 12588 23480 12640
rect 23532 12588 23538 12640
rect 24670 12588 24676 12640
rect 24728 12588 24734 12640
rect 26878 12588 26884 12640
rect 26936 12628 26942 12640
rect 26973 12631 27031 12637
rect 26973 12628 26985 12631
rect 26936 12600 26985 12628
rect 26936 12588 26942 12600
rect 26973 12597 26985 12600
rect 27019 12597 27031 12631
rect 26973 12591 27031 12597
rect 27154 12588 27160 12640
rect 27212 12588 27218 12640
rect 1104 12538 28704 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 28704 12538
rect 1104 12464 28704 12486
rect 5718 12384 5724 12436
rect 5776 12424 5782 12436
rect 5813 12427 5871 12433
rect 5813 12424 5825 12427
rect 5776 12396 5825 12424
rect 5776 12384 5782 12396
rect 5813 12393 5825 12396
rect 5859 12393 5871 12427
rect 12526 12424 12532 12436
rect 5813 12387 5871 12393
rect 10888 12396 12532 12424
rect 10888 12368 10916 12396
rect 12526 12384 12532 12396
rect 12584 12384 12590 12436
rect 12894 12384 12900 12436
rect 12952 12424 12958 12436
rect 13170 12424 13176 12436
rect 12952 12396 13176 12424
rect 12952 12384 12958 12396
rect 13170 12384 13176 12396
rect 13228 12384 13234 12436
rect 13725 12427 13783 12433
rect 13725 12393 13737 12427
rect 13771 12424 13783 12427
rect 13909 12427 13967 12433
rect 13771 12396 13860 12424
rect 13771 12393 13783 12396
rect 13725 12387 13783 12393
rect 10870 12316 10876 12368
rect 10928 12316 10934 12368
rect 11149 12359 11207 12365
rect 11149 12325 11161 12359
rect 11195 12325 11207 12359
rect 11149 12319 11207 12325
rect 11900 12328 12204 12356
rect 11164 12288 11192 12319
rect 10244 12260 11192 12288
rect 4798 12180 4804 12232
rect 4856 12220 4862 12232
rect 5261 12223 5319 12229
rect 5261 12220 5273 12223
rect 4856 12192 5273 12220
rect 4856 12180 4862 12192
rect 5261 12189 5273 12192
rect 5307 12189 5319 12223
rect 5261 12183 5319 12189
rect 5629 12223 5687 12229
rect 5629 12189 5641 12223
rect 5675 12220 5687 12223
rect 5810 12220 5816 12232
rect 5675 12192 5816 12220
rect 5675 12189 5687 12192
rect 5629 12183 5687 12189
rect 5276 12084 5304 12183
rect 5810 12180 5816 12192
rect 5868 12220 5874 12232
rect 5905 12223 5963 12229
rect 5905 12220 5917 12223
rect 5868 12192 5917 12220
rect 5868 12180 5874 12192
rect 5905 12189 5917 12192
rect 5951 12189 5963 12223
rect 5905 12183 5963 12189
rect 6089 12223 6147 12229
rect 6089 12189 6101 12223
rect 6135 12220 6147 12223
rect 6178 12220 6184 12232
rect 6135 12192 6184 12220
rect 6135 12189 6147 12192
rect 6089 12183 6147 12189
rect 6178 12180 6184 12192
rect 6236 12220 6242 12232
rect 10244 12229 10272 12260
rect 10229 12223 10287 12229
rect 6236 12192 10180 12220
rect 6236 12180 6242 12192
rect 5442 12112 5448 12164
rect 5500 12112 5506 12164
rect 5534 12112 5540 12164
rect 5592 12112 5598 12164
rect 5902 12084 5908 12096
rect 5276 12056 5908 12084
rect 5902 12044 5908 12056
rect 5960 12044 5966 12096
rect 5994 12044 6000 12096
rect 6052 12044 6058 12096
rect 9214 12044 9220 12096
rect 9272 12084 9278 12096
rect 10045 12087 10103 12093
rect 10045 12084 10057 12087
rect 9272 12056 10057 12084
rect 9272 12044 9278 12056
rect 10045 12053 10057 12056
rect 10091 12053 10103 12087
rect 10152 12084 10180 12192
rect 10229 12189 10241 12223
rect 10275 12189 10287 12223
rect 10229 12183 10287 12189
rect 10318 12180 10324 12232
rect 10376 12220 10382 12232
rect 10413 12223 10471 12229
rect 10413 12220 10425 12223
rect 10376 12192 10425 12220
rect 10376 12180 10382 12192
rect 10413 12189 10425 12192
rect 10459 12189 10471 12223
rect 10413 12183 10471 12189
rect 10505 12223 10563 12229
rect 10505 12189 10517 12223
rect 10551 12220 10563 12223
rect 10778 12220 10784 12232
rect 10551 12192 10784 12220
rect 10551 12189 10563 12192
rect 10505 12183 10563 12189
rect 10428 12152 10456 12183
rect 10778 12180 10784 12192
rect 10836 12180 10842 12232
rect 11330 12229 11336 12232
rect 11328 12220 11336 12229
rect 11291 12192 11336 12220
rect 11328 12183 11336 12192
rect 11330 12180 11336 12183
rect 11388 12180 11394 12232
rect 11422 12180 11428 12232
rect 11480 12180 11486 12232
rect 11698 12220 11704 12232
rect 11659 12192 11704 12220
rect 11698 12180 11704 12192
rect 11756 12180 11762 12232
rect 11793 12223 11851 12229
rect 11793 12189 11805 12223
rect 11839 12220 11851 12223
rect 11900 12220 11928 12328
rect 12176 12300 12204 12328
rect 12710 12316 12716 12368
rect 12768 12356 12774 12368
rect 13630 12356 13636 12368
rect 12768 12328 13636 12356
rect 12768 12316 12774 12328
rect 13630 12316 13636 12328
rect 13688 12316 13694 12368
rect 13832 12356 13860 12396
rect 13909 12393 13921 12427
rect 13955 12424 13967 12427
rect 14090 12424 14096 12436
rect 13955 12396 14096 12424
rect 13955 12393 13967 12396
rect 13909 12387 13967 12393
rect 14090 12384 14096 12396
rect 14148 12384 14154 12436
rect 18693 12427 18751 12433
rect 18693 12393 18705 12427
rect 18739 12424 18751 12427
rect 18874 12424 18880 12436
rect 18739 12396 18880 12424
rect 18739 12393 18751 12396
rect 18693 12387 18751 12393
rect 18874 12384 18880 12396
rect 18932 12384 18938 12436
rect 19150 12384 19156 12436
rect 19208 12424 19214 12436
rect 19245 12427 19303 12433
rect 19245 12424 19257 12427
rect 19208 12396 19257 12424
rect 19208 12384 19214 12396
rect 19245 12393 19257 12396
rect 19291 12393 19303 12427
rect 20622 12424 20628 12436
rect 19245 12387 19303 12393
rect 19720 12396 20628 12424
rect 14185 12359 14243 12365
rect 14185 12356 14197 12359
rect 13832 12328 14197 12356
rect 14185 12325 14197 12328
rect 14231 12325 14243 12359
rect 14185 12319 14243 12325
rect 18414 12316 18420 12368
rect 18472 12356 18478 12368
rect 19720 12356 19748 12396
rect 20622 12384 20628 12396
rect 20680 12384 20686 12436
rect 22373 12427 22431 12433
rect 22373 12393 22385 12427
rect 22419 12424 22431 12427
rect 23290 12424 23296 12436
rect 22419 12396 23296 12424
rect 22419 12393 22431 12396
rect 22373 12387 22431 12393
rect 23290 12384 23296 12396
rect 23348 12384 23354 12436
rect 18472 12328 19748 12356
rect 18472 12316 18478 12328
rect 12066 12248 12072 12300
rect 12124 12248 12130 12300
rect 12158 12248 12164 12300
rect 12216 12288 12222 12300
rect 15654 12288 15660 12300
rect 12216 12260 15660 12288
rect 12216 12248 12222 12260
rect 15654 12248 15660 12260
rect 15712 12248 15718 12300
rect 18601 12291 18659 12297
rect 18601 12257 18613 12291
rect 18647 12288 18659 12291
rect 18966 12288 18972 12300
rect 18647 12260 18972 12288
rect 18647 12257 18659 12260
rect 18601 12251 18659 12257
rect 18966 12248 18972 12260
rect 19024 12248 19030 12300
rect 19061 12291 19119 12297
rect 19061 12257 19073 12291
rect 19107 12288 19119 12291
rect 20717 12291 20775 12297
rect 20717 12288 20729 12291
rect 19107 12260 20729 12288
rect 19107 12257 19119 12260
rect 19061 12251 19119 12257
rect 20717 12257 20729 12260
rect 20763 12257 20775 12291
rect 22370 12288 22376 12300
rect 20717 12251 20775 12257
rect 22020 12260 22376 12288
rect 11839 12192 11928 12220
rect 11839 12189 11851 12192
rect 11793 12183 11851 12189
rect 11974 12180 11980 12232
rect 12032 12180 12038 12232
rect 12250 12180 12256 12232
rect 12308 12180 12314 12232
rect 12342 12180 12348 12232
rect 12400 12180 12406 12232
rect 12710 12220 12716 12232
rect 12452 12192 12716 12220
rect 11238 12152 11244 12164
rect 10428 12124 11244 12152
rect 11238 12112 11244 12124
rect 11296 12112 11302 12164
rect 11514 12112 11520 12164
rect 11572 12152 11578 12164
rect 11572 12124 12388 12152
rect 11572 12112 11578 12124
rect 12250 12084 12256 12096
rect 10152 12056 12256 12084
rect 10045 12047 10103 12053
rect 12250 12044 12256 12056
rect 12308 12044 12314 12096
rect 12360 12084 12388 12124
rect 12452 12084 12480 12192
rect 12710 12180 12716 12192
rect 12768 12180 12774 12232
rect 12802 12180 12808 12232
rect 12860 12180 12866 12232
rect 13078 12180 13084 12232
rect 13136 12180 13142 12232
rect 13262 12180 13268 12232
rect 13320 12180 13326 12232
rect 13354 12180 13360 12232
rect 13412 12180 13418 12232
rect 14274 12180 14280 12232
rect 14332 12220 14338 12232
rect 14369 12223 14427 12229
rect 14369 12220 14381 12223
rect 14332 12192 14381 12220
rect 14332 12180 14338 12192
rect 14369 12189 14381 12192
rect 14415 12189 14427 12223
rect 14369 12183 14427 12189
rect 14458 12180 14464 12232
rect 14516 12180 14522 12232
rect 14550 12180 14556 12232
rect 14608 12180 14614 12232
rect 14645 12223 14703 12229
rect 14645 12189 14657 12223
rect 14691 12220 14703 12223
rect 15378 12220 15384 12232
rect 14691 12192 15384 12220
rect 14691 12189 14703 12192
rect 14645 12183 14703 12189
rect 15378 12180 15384 12192
rect 15436 12180 15442 12232
rect 18874 12180 18880 12232
rect 18932 12180 18938 12232
rect 20990 12180 20996 12232
rect 21048 12220 21054 12232
rect 21542 12220 21548 12232
rect 21048 12192 21548 12220
rect 21048 12180 21054 12192
rect 21542 12180 21548 12192
rect 21600 12180 21606 12232
rect 21729 12223 21787 12229
rect 21729 12189 21741 12223
rect 21775 12189 21787 12223
rect 21729 12183 21787 12189
rect 12529 12155 12587 12161
rect 12529 12121 12541 12155
rect 12575 12152 12587 12155
rect 13170 12152 13176 12164
rect 12575 12124 13176 12152
rect 12575 12121 12587 12124
rect 12529 12115 12587 12121
rect 13170 12112 13176 12124
rect 13228 12112 13234 12164
rect 14476 12152 14504 12180
rect 14734 12152 14740 12164
rect 14476 12124 14740 12152
rect 14734 12112 14740 12124
rect 14792 12112 14798 12164
rect 20254 12112 20260 12164
rect 20312 12112 20318 12164
rect 20622 12112 20628 12164
rect 20680 12152 20686 12164
rect 21744 12152 21772 12183
rect 21818 12180 21824 12232
rect 21876 12180 21882 12232
rect 22020 12161 22048 12260
rect 22370 12248 22376 12260
rect 22428 12248 22434 12300
rect 22465 12291 22523 12297
rect 22465 12257 22477 12291
rect 22511 12288 22523 12291
rect 24394 12288 24400 12300
rect 22511 12260 24400 12288
rect 22511 12257 22523 12260
rect 22465 12251 22523 12257
rect 24394 12248 24400 12260
rect 24452 12288 24458 12300
rect 26234 12288 26240 12300
rect 24452 12260 26240 12288
rect 24452 12248 24458 12260
rect 26234 12248 26240 12260
rect 26292 12288 26298 12300
rect 26510 12288 26516 12300
rect 26292 12260 26516 12288
rect 26292 12248 26298 12260
rect 26510 12248 26516 12260
rect 26568 12248 26574 12300
rect 22186 12180 22192 12232
rect 22244 12229 22250 12232
rect 22244 12220 22252 12229
rect 22244 12192 22289 12220
rect 22244 12183 22252 12192
rect 22244 12180 22250 12183
rect 20680 12124 21772 12152
rect 22005 12155 22063 12161
rect 20680 12112 20686 12124
rect 22005 12121 22017 12155
rect 22051 12121 22063 12155
rect 22005 12115 22063 12121
rect 22097 12155 22155 12161
rect 22097 12121 22109 12155
rect 22143 12152 22155 12155
rect 22462 12152 22468 12164
rect 22143 12124 22468 12152
rect 22143 12121 22155 12124
rect 22097 12115 22155 12121
rect 12360 12056 12480 12084
rect 12621 12087 12679 12093
rect 12621 12053 12633 12087
rect 12667 12084 12679 12087
rect 12986 12084 12992 12096
rect 12667 12056 12992 12084
rect 12667 12053 12679 12056
rect 12621 12047 12679 12053
rect 12986 12044 12992 12056
rect 13044 12044 13050 12096
rect 13538 12044 13544 12096
rect 13596 12084 13602 12096
rect 13725 12087 13783 12093
rect 13725 12084 13737 12087
rect 13596 12056 13737 12084
rect 13596 12044 13602 12056
rect 13725 12053 13737 12056
rect 13771 12084 13783 12087
rect 15470 12084 15476 12096
rect 13771 12056 15476 12084
rect 13771 12053 13783 12056
rect 13725 12047 13783 12053
rect 15470 12044 15476 12056
rect 15528 12044 15534 12096
rect 18690 12044 18696 12096
rect 18748 12084 18754 12096
rect 22020 12084 22048 12115
rect 22462 12112 22468 12124
rect 22520 12112 22526 12164
rect 22738 12112 22744 12164
rect 22796 12112 22802 12164
rect 25498 12152 25504 12164
rect 23966 12124 25504 12152
rect 22186 12084 22192 12096
rect 18748 12056 22192 12084
rect 18748 12044 18754 12056
rect 22186 12044 22192 12056
rect 22244 12044 22250 12096
rect 23382 12044 23388 12096
rect 23440 12084 23446 12096
rect 24044 12084 24072 12124
rect 25498 12112 25504 12124
rect 25556 12112 25562 12164
rect 26513 12155 26571 12161
rect 26513 12121 26525 12155
rect 26559 12121 26571 12155
rect 27890 12152 27896 12164
rect 27738 12124 27896 12152
rect 26513 12115 26571 12121
rect 23440 12056 24072 12084
rect 23440 12044 23446 12056
rect 24210 12044 24216 12096
rect 24268 12044 24274 12096
rect 26528 12084 26556 12115
rect 27890 12112 27896 12124
rect 27948 12112 27954 12164
rect 27154 12084 27160 12096
rect 26528 12056 27160 12084
rect 27154 12044 27160 12056
rect 27212 12044 27218 12096
rect 27985 12087 28043 12093
rect 27985 12053 27997 12087
rect 28031 12084 28043 12087
rect 28166 12084 28172 12096
rect 28031 12056 28172 12084
rect 28031 12053 28043 12056
rect 27985 12047 28043 12053
rect 28166 12044 28172 12056
rect 28224 12044 28230 12096
rect 1104 11994 28704 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 28704 11994
rect 1104 11920 28704 11942
rect 5350 11880 5356 11892
rect 3344 11852 5356 11880
rect 3344 11753 3372 11852
rect 5350 11840 5356 11852
rect 5408 11840 5414 11892
rect 7742 11840 7748 11892
rect 7800 11880 7806 11892
rect 13630 11880 13636 11892
rect 7800 11852 13636 11880
rect 7800 11840 7806 11852
rect 4614 11772 4620 11824
rect 4672 11772 4678 11824
rect 5368 11812 5396 11840
rect 6825 11815 6883 11821
rect 6825 11812 6837 11815
rect 5368 11784 6837 11812
rect 6825 11781 6837 11784
rect 6871 11812 6883 11815
rect 6914 11812 6920 11824
rect 6871 11784 6920 11812
rect 6871 11781 6883 11784
rect 6825 11775 6883 11781
rect 6914 11772 6920 11784
rect 6972 11812 6978 11824
rect 8202 11812 8208 11824
rect 6972 11784 8208 11812
rect 6972 11772 6978 11784
rect 8202 11772 8208 11784
rect 8260 11772 8266 11824
rect 11992 11821 12020 11852
rect 13630 11840 13636 11852
rect 13688 11840 13694 11892
rect 18506 11840 18512 11892
rect 18564 11880 18570 11892
rect 18564 11852 18828 11880
rect 18564 11840 18570 11852
rect 11977 11815 12035 11821
rect 11977 11781 11989 11815
rect 12023 11781 12035 11815
rect 11977 11775 12035 11781
rect 12805 11815 12863 11821
rect 12805 11781 12817 11815
rect 12851 11812 12863 11815
rect 13725 11815 13783 11821
rect 13725 11812 13737 11815
rect 12851 11784 13737 11812
rect 12851 11781 12863 11784
rect 12805 11775 12863 11781
rect 13725 11781 13737 11784
rect 13771 11812 13783 11815
rect 13814 11812 13820 11824
rect 13771 11784 13820 11812
rect 13771 11781 13783 11784
rect 13725 11775 13783 11781
rect 3329 11747 3387 11753
rect 3329 11713 3341 11747
rect 3375 11713 3387 11747
rect 3329 11707 3387 11713
rect 5905 11747 5963 11753
rect 5905 11713 5917 11747
rect 5951 11713 5963 11747
rect 5905 11707 5963 11713
rect 3602 11636 3608 11688
rect 3660 11636 3666 11688
rect 5077 11679 5135 11685
rect 5077 11645 5089 11679
rect 5123 11676 5135 11679
rect 5810 11676 5816 11688
rect 5123 11648 5816 11676
rect 5123 11645 5135 11648
rect 5077 11639 5135 11645
rect 5810 11636 5816 11648
rect 5868 11636 5874 11688
rect 5920 11676 5948 11707
rect 6086 11704 6092 11756
rect 6144 11704 6150 11756
rect 6181 11747 6239 11753
rect 6181 11713 6193 11747
rect 6227 11744 6239 11747
rect 6362 11744 6368 11756
rect 6227 11716 6368 11744
rect 6227 11713 6239 11716
rect 6181 11707 6239 11713
rect 6362 11704 6368 11716
rect 6420 11704 6426 11756
rect 6457 11747 6515 11753
rect 6457 11713 6469 11747
rect 6503 11713 6515 11747
rect 6457 11707 6515 11713
rect 6270 11676 6276 11688
rect 5920 11648 6276 11676
rect 6270 11636 6276 11648
rect 6328 11676 6334 11688
rect 6472 11676 6500 11707
rect 6546 11704 6552 11756
rect 6604 11744 6610 11756
rect 6641 11747 6699 11753
rect 6641 11744 6653 11747
rect 6604 11716 6653 11744
rect 6604 11704 6610 11716
rect 6641 11713 6653 11716
rect 6687 11744 6699 11747
rect 7377 11747 7435 11753
rect 7377 11744 7389 11747
rect 6687 11716 7389 11744
rect 6687 11713 6699 11716
rect 6641 11707 6699 11713
rect 7377 11713 7389 11716
rect 7423 11713 7435 11747
rect 7377 11707 7435 11713
rect 7561 11747 7619 11753
rect 7561 11713 7573 11747
rect 7607 11713 7619 11747
rect 7561 11707 7619 11713
rect 7745 11747 7803 11753
rect 7745 11713 7757 11747
rect 7791 11744 7803 11747
rect 8018 11744 8024 11756
rect 7791 11716 8024 11744
rect 7791 11713 7803 11716
rect 7745 11707 7803 11713
rect 6328 11648 6500 11676
rect 6328 11636 6334 11648
rect 7006 11636 7012 11688
rect 7064 11676 7070 11688
rect 7576 11676 7604 11707
rect 8018 11704 8024 11716
rect 8076 11704 8082 11756
rect 10962 11747 10968 11756
rect 10888 11719 10968 11747
rect 7834 11676 7840 11688
rect 7064 11648 7840 11676
rect 7064 11636 7070 11648
rect 7834 11636 7840 11648
rect 7892 11636 7898 11688
rect 9585 11679 9643 11685
rect 9585 11645 9597 11679
rect 9631 11645 9643 11679
rect 9585 11639 9643 11645
rect 5166 11500 5172 11552
rect 5224 11500 5230 11552
rect 5718 11500 5724 11552
rect 5776 11540 5782 11552
rect 5905 11543 5963 11549
rect 5905 11540 5917 11543
rect 5776 11512 5917 11540
rect 5776 11500 5782 11512
rect 5905 11509 5917 11512
rect 5951 11509 5963 11543
rect 5905 11503 5963 11509
rect 6549 11543 6607 11549
rect 6549 11509 6561 11543
rect 6595 11540 6607 11543
rect 7098 11540 7104 11552
rect 6595 11512 7104 11540
rect 6595 11509 6607 11512
rect 6549 11503 6607 11509
rect 7098 11500 7104 11512
rect 7156 11500 7162 11552
rect 8294 11500 8300 11552
rect 8352 11500 8358 11552
rect 8938 11500 8944 11552
rect 8996 11540 9002 11552
rect 9600 11540 9628 11639
rect 9858 11636 9864 11688
rect 9916 11636 9922 11688
rect 10410 11636 10416 11688
rect 10468 11676 10474 11688
rect 10888 11676 10916 11719
rect 10962 11704 10968 11719
rect 11020 11704 11026 11756
rect 12820 11676 12848 11775
rect 13814 11772 13820 11784
rect 13872 11772 13878 11824
rect 18690 11772 18696 11824
rect 18748 11772 18754 11824
rect 18800 11821 18828 11852
rect 18874 11840 18880 11892
rect 18932 11880 18938 11892
rect 19061 11883 19119 11889
rect 19061 11880 19073 11883
rect 18932 11852 19073 11880
rect 18932 11840 18938 11852
rect 19061 11849 19073 11852
rect 19107 11849 19119 11883
rect 19061 11843 19119 11849
rect 19153 11883 19211 11889
rect 19153 11849 19165 11883
rect 19199 11880 19211 11883
rect 19702 11880 19708 11892
rect 19199 11852 19708 11880
rect 19199 11849 19211 11852
rect 19153 11843 19211 11849
rect 18785 11815 18843 11821
rect 18785 11781 18797 11815
rect 18831 11781 18843 11815
rect 18785 11775 18843 11781
rect 12986 11704 12992 11756
rect 13044 11704 13050 11756
rect 13170 11704 13176 11756
rect 13228 11704 13234 11756
rect 13262 11704 13268 11756
rect 13320 11704 13326 11756
rect 13357 11747 13415 11753
rect 13357 11713 13369 11747
rect 13403 11744 13415 11747
rect 14366 11744 14372 11756
rect 13403 11716 14372 11744
rect 13403 11713 13415 11716
rect 13357 11707 13415 11713
rect 14366 11704 14372 11716
rect 14424 11704 14430 11756
rect 18414 11704 18420 11756
rect 18472 11704 18478 11756
rect 18598 11753 18604 11756
rect 18565 11747 18604 11753
rect 18565 11713 18577 11747
rect 18565 11707 18604 11713
rect 18598 11704 18604 11707
rect 18656 11704 18662 11756
rect 18923 11747 18981 11753
rect 18923 11713 18935 11747
rect 18969 11744 18981 11747
rect 19168 11744 19196 11843
rect 19702 11840 19708 11852
rect 19760 11840 19766 11892
rect 20254 11840 20260 11892
rect 20312 11880 20318 11892
rect 21450 11880 21456 11892
rect 20312 11852 21456 11880
rect 20312 11840 20318 11852
rect 21450 11840 21456 11852
rect 21508 11840 21514 11892
rect 22646 11840 22652 11892
rect 22704 11840 22710 11892
rect 25498 11840 25504 11892
rect 25556 11880 25562 11892
rect 25556 11852 26924 11880
rect 25556 11840 25562 11852
rect 20272 11812 20300 11840
rect 20194 11784 20300 11812
rect 20625 11815 20683 11821
rect 20625 11781 20637 11815
rect 20671 11812 20683 11815
rect 20714 11812 20720 11824
rect 20671 11784 20720 11812
rect 20671 11781 20683 11784
rect 20625 11775 20683 11781
rect 20714 11772 20720 11784
rect 20772 11772 20778 11824
rect 23382 11772 23388 11824
rect 23440 11772 23446 11824
rect 26160 11812 26188 11852
rect 26082 11784 26188 11812
rect 26234 11772 26240 11824
rect 26292 11812 26298 11824
rect 26896 11812 26924 11852
rect 27338 11840 27344 11892
rect 27396 11840 27402 11892
rect 27890 11812 27896 11824
rect 26292 11784 26832 11812
rect 26896 11784 27896 11812
rect 26292 11772 26298 11784
rect 18969 11716 19196 11744
rect 22097 11747 22155 11753
rect 18969 11713 18981 11716
rect 18923 11707 18981 11713
rect 22097 11713 22109 11747
rect 22143 11744 22155 11747
rect 22278 11744 22284 11756
rect 22143 11716 22284 11744
rect 22143 11713 22155 11716
rect 22097 11707 22155 11713
rect 22278 11704 22284 11716
rect 22336 11704 22342 11756
rect 22370 11704 22376 11756
rect 22428 11704 22434 11756
rect 24394 11704 24400 11756
rect 24452 11704 24458 11756
rect 26804 11753 26832 11784
rect 27890 11772 27896 11784
rect 27948 11772 27954 11824
rect 26789 11747 26847 11753
rect 26789 11713 26801 11747
rect 26835 11713 26847 11747
rect 26789 11707 26847 11713
rect 26878 11704 26884 11756
rect 26936 11744 26942 11756
rect 26973 11747 27031 11753
rect 26973 11744 26985 11747
rect 26936 11716 26985 11744
rect 26936 11704 26942 11716
rect 26973 11713 26985 11716
rect 27019 11713 27031 11747
rect 26973 11707 27031 11713
rect 27154 11704 27160 11756
rect 27212 11704 27218 11756
rect 28350 11704 28356 11756
rect 28408 11704 28414 11756
rect 10468 11648 10916 11676
rect 10980 11648 12848 11676
rect 10468 11636 10474 11648
rect 10980 11540 11008 11648
rect 13078 11636 13084 11688
rect 13136 11676 13142 11688
rect 13722 11676 13728 11688
rect 13136 11648 13728 11676
rect 13136 11636 13142 11648
rect 13722 11636 13728 11648
rect 13780 11636 13786 11688
rect 17862 11636 17868 11688
rect 17920 11676 17926 11688
rect 20254 11676 20260 11688
rect 17920 11648 20260 11676
rect 17920 11636 17926 11648
rect 20254 11636 20260 11648
rect 20312 11636 20318 11688
rect 20901 11679 20959 11685
rect 20901 11645 20913 11679
rect 20947 11676 20959 11679
rect 20990 11676 20996 11688
rect 20947 11648 20996 11676
rect 20947 11645 20959 11648
rect 20901 11639 20959 11645
rect 11054 11568 11060 11620
rect 11112 11608 11118 11620
rect 13262 11608 13268 11620
rect 11112 11580 13268 11608
rect 11112 11568 11118 11580
rect 13262 11568 13268 11580
rect 13320 11568 13326 11620
rect 15194 11608 15200 11620
rect 13372 11580 15200 11608
rect 8996 11512 11008 11540
rect 11333 11543 11391 11549
rect 8996 11500 9002 11512
rect 11333 11509 11345 11543
rect 11379 11540 11391 11543
rect 11698 11540 11704 11552
rect 11379 11512 11704 11540
rect 11379 11509 11391 11512
rect 11333 11503 11391 11509
rect 11698 11500 11704 11512
rect 11756 11540 11762 11552
rect 11974 11540 11980 11552
rect 11756 11512 11980 11540
rect 11756 11500 11762 11512
rect 11974 11500 11980 11512
rect 12032 11500 12038 11552
rect 12526 11500 12532 11552
rect 12584 11540 12590 11552
rect 13372 11540 13400 11580
rect 15194 11568 15200 11580
rect 15252 11568 15258 11620
rect 12584 11512 13400 11540
rect 12584 11500 12590 11512
rect 13538 11500 13544 11552
rect 13596 11540 13602 11552
rect 13633 11543 13691 11549
rect 13633 11540 13645 11543
rect 13596 11512 13645 11540
rect 13596 11500 13602 11512
rect 13633 11509 13645 11512
rect 13679 11509 13691 11543
rect 13633 11503 13691 11509
rect 19242 11500 19248 11552
rect 19300 11540 19306 11552
rect 20916 11540 20944 11639
rect 20990 11636 20996 11648
rect 21048 11636 21054 11688
rect 22557 11679 22615 11685
rect 22557 11645 22569 11679
rect 22603 11676 22615 11679
rect 24121 11679 24179 11685
rect 24121 11676 24133 11679
rect 22603 11648 24133 11676
rect 22603 11645 22615 11648
rect 22557 11639 22615 11645
rect 24121 11645 24133 11648
rect 24167 11645 24179 11679
rect 24121 11639 24179 11645
rect 26513 11679 26571 11685
rect 26513 11645 26525 11679
rect 26559 11676 26571 11679
rect 27430 11676 27436 11688
rect 26559 11648 27436 11676
rect 26559 11645 26571 11648
rect 26513 11639 26571 11645
rect 27430 11636 27436 11648
rect 27488 11636 27494 11688
rect 21542 11568 21548 11620
rect 21600 11608 21606 11620
rect 22646 11608 22652 11620
rect 21600 11580 22652 11608
rect 21600 11568 21606 11580
rect 22646 11568 22652 11580
rect 22704 11568 22710 11620
rect 19300 11512 20944 11540
rect 22189 11543 22247 11549
rect 19300 11500 19306 11512
rect 22189 11509 22201 11543
rect 22235 11540 22247 11543
rect 22554 11540 22560 11552
rect 22235 11512 22560 11540
rect 22235 11509 22247 11512
rect 22189 11503 22247 11509
rect 22554 11500 22560 11512
rect 22612 11500 22618 11552
rect 25038 11500 25044 11552
rect 25096 11500 25102 11552
rect 26510 11500 26516 11552
rect 26568 11540 26574 11552
rect 26973 11543 27031 11549
rect 26973 11540 26985 11543
rect 26568 11512 26985 11540
rect 26568 11500 26574 11512
rect 26973 11509 26985 11512
rect 27019 11509 27031 11543
rect 26973 11503 27031 11509
rect 27062 11500 27068 11552
rect 27120 11540 27126 11552
rect 27338 11540 27344 11552
rect 27120 11512 27344 11540
rect 27120 11500 27126 11512
rect 27338 11500 27344 11512
rect 27396 11540 27402 11552
rect 28169 11543 28227 11549
rect 28169 11540 28181 11543
rect 27396 11512 28181 11540
rect 27396 11500 27402 11512
rect 28169 11509 28181 11512
rect 28215 11509 28227 11543
rect 28169 11503 28227 11509
rect 1104 11450 28704 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 28704 11450
rect 1104 11376 28704 11398
rect 3602 11296 3608 11348
rect 3660 11336 3666 11348
rect 4341 11339 4399 11345
rect 4341 11336 4353 11339
rect 3660 11308 4353 11336
rect 3660 11296 3666 11308
rect 4341 11305 4353 11308
rect 4387 11305 4399 11339
rect 4341 11299 4399 11305
rect 5353 11339 5411 11345
rect 5353 11305 5365 11339
rect 5399 11336 5411 11339
rect 5442 11336 5448 11348
rect 5399 11308 5448 11336
rect 5399 11305 5411 11308
rect 5353 11299 5411 11305
rect 5442 11296 5448 11308
rect 5500 11296 5506 11348
rect 8018 11296 8024 11348
rect 8076 11336 8082 11348
rect 8076 11308 10272 11336
rect 8076 11296 8082 11308
rect 6638 11268 6644 11280
rect 5000 11240 6644 11268
rect 5000 11209 5028 11240
rect 6638 11228 6644 11240
rect 6696 11228 6702 11280
rect 7929 11271 7987 11277
rect 7929 11268 7941 11271
rect 6748 11240 7941 11268
rect 6748 11212 6776 11240
rect 7929 11237 7941 11240
rect 7975 11237 7987 11271
rect 7929 11231 7987 11237
rect 4985 11203 5043 11209
rect 4985 11169 4997 11203
rect 5031 11169 5043 11203
rect 4985 11163 5043 11169
rect 5718 11160 5724 11212
rect 5776 11160 5782 11212
rect 5810 11160 5816 11212
rect 5868 11200 5874 11212
rect 5905 11203 5963 11209
rect 5905 11200 5917 11203
rect 5868 11172 5917 11200
rect 5868 11160 5874 11172
rect 5905 11169 5917 11172
rect 5951 11169 5963 11203
rect 5905 11163 5963 11169
rect 6730 11160 6736 11212
rect 6788 11160 6794 11212
rect 6914 11160 6920 11212
rect 6972 11160 6978 11212
rect 4709 11135 4767 11141
rect 4709 11101 4721 11135
rect 4755 11132 4767 11135
rect 5166 11132 5172 11144
rect 4755 11104 5172 11132
rect 4755 11101 4767 11104
rect 4709 11095 4767 11101
rect 5166 11092 5172 11104
rect 5224 11092 5230 11144
rect 5629 11135 5687 11141
rect 5629 11101 5641 11135
rect 5675 11101 5687 11135
rect 5629 11095 5687 11101
rect 6089 11135 6147 11141
rect 6089 11101 6101 11135
rect 6135 11132 6147 11135
rect 6178 11132 6184 11144
rect 6135 11104 6184 11132
rect 6135 11101 6147 11104
rect 6089 11095 6147 11101
rect 5644 11064 5672 11095
rect 6178 11092 6184 11104
rect 6236 11092 6242 11144
rect 6270 11092 6276 11144
rect 6328 11092 6334 11144
rect 6546 11092 6552 11144
rect 6604 11092 6610 11144
rect 7834 11092 7840 11144
rect 7892 11092 7898 11144
rect 8036 11141 8064 11296
rect 10244 11268 10272 11308
rect 10778 11296 10784 11348
rect 10836 11296 10842 11348
rect 12066 11296 12072 11348
rect 12124 11336 12130 11348
rect 12618 11336 12624 11348
rect 12124 11308 12624 11336
rect 12124 11296 12130 11308
rect 12618 11296 12624 11308
rect 12676 11296 12682 11348
rect 12802 11296 12808 11348
rect 12860 11336 12866 11348
rect 12897 11339 12955 11345
rect 12897 11336 12909 11339
rect 12860 11308 12909 11336
rect 12860 11296 12866 11308
rect 12897 11305 12909 11308
rect 12943 11305 12955 11339
rect 12897 11299 12955 11305
rect 13081 11339 13139 11345
rect 13081 11305 13093 11339
rect 13127 11305 13139 11339
rect 13081 11299 13139 11305
rect 11054 11268 11060 11280
rect 10244 11240 11060 11268
rect 11054 11228 11060 11240
rect 11112 11228 11118 11280
rect 12250 11228 12256 11280
rect 12308 11268 12314 11280
rect 12526 11268 12532 11280
rect 12308 11240 12532 11268
rect 12308 11228 12314 11240
rect 12526 11228 12532 11240
rect 12584 11228 12590 11280
rect 12986 11268 12992 11280
rect 12728 11240 12992 11268
rect 8938 11160 8944 11212
rect 8996 11160 9002 11212
rect 9214 11160 9220 11212
rect 9272 11160 9278 11212
rect 10689 11203 10747 11209
rect 10689 11169 10701 11203
rect 10735 11200 10747 11203
rect 11333 11203 11391 11209
rect 11333 11200 11345 11203
rect 10735 11172 11345 11200
rect 10735 11169 10747 11172
rect 10689 11163 10747 11169
rect 11333 11169 11345 11172
rect 11379 11169 11391 11203
rect 11333 11163 11391 11169
rect 8021 11135 8079 11141
rect 8021 11101 8033 11135
rect 8067 11101 8079 11135
rect 11348 11132 11376 11163
rect 11514 11160 11520 11212
rect 11572 11200 11578 11212
rect 12728 11200 12756 11240
rect 12986 11228 12992 11240
rect 13044 11228 13050 11280
rect 11572 11172 11928 11200
rect 11572 11160 11578 11172
rect 11900 11141 11928 11172
rect 12360 11172 12756 11200
rect 11655 11135 11713 11141
rect 11655 11132 11667 11135
rect 11348 11104 11667 11132
rect 8021 11095 8079 11101
rect 11655 11101 11667 11104
rect 11701 11101 11713 11135
rect 11655 11095 11713 11101
rect 11885 11135 11943 11141
rect 11885 11101 11897 11135
rect 11931 11101 11943 11135
rect 11885 11095 11943 11101
rect 12068 11135 12126 11141
rect 12068 11101 12080 11135
rect 12114 11101 12126 11135
rect 12068 11095 12126 11101
rect 6365 11067 6423 11073
rect 6365 11064 6377 11067
rect 5644 11036 6377 11064
rect 6365 11033 6377 11036
rect 6411 11064 6423 11067
rect 6454 11064 6460 11076
rect 6411 11036 6460 11064
rect 6411 11033 6423 11036
rect 6365 11027 6423 11033
rect 6454 11024 6460 11036
rect 6512 11024 6518 11076
rect 7006 11024 7012 11076
rect 7064 11064 7070 11076
rect 7742 11064 7748 11076
rect 7064 11036 7748 11064
rect 7064 11024 7070 11036
rect 7742 11024 7748 11036
rect 7800 11024 7806 11076
rect 10870 11064 10876 11076
rect 10442 11036 10876 11064
rect 10870 11024 10876 11036
rect 10928 11024 10934 11076
rect 11422 11064 11428 11076
rect 10980 11036 11428 11064
rect 10980 11008 11008 11036
rect 11422 11024 11428 11036
rect 11480 11064 11486 11076
rect 11793 11067 11851 11073
rect 11793 11064 11805 11067
rect 11480 11036 11805 11064
rect 11480 11024 11486 11036
rect 11793 11033 11805 11036
rect 11839 11033 11851 11067
rect 12084 11064 12112 11095
rect 12158 11092 12164 11144
rect 12216 11092 12222 11144
rect 12250 11092 12256 11144
rect 12308 11092 12314 11144
rect 12360 11141 12388 11172
rect 12802 11160 12808 11212
rect 12860 11200 12866 11212
rect 13096 11200 13124 11299
rect 13354 11296 13360 11348
rect 13412 11296 13418 11348
rect 13541 11339 13599 11345
rect 13541 11305 13553 11339
rect 13587 11305 13599 11339
rect 13541 11299 13599 11305
rect 13556 11268 13584 11299
rect 13630 11296 13636 11348
rect 13688 11336 13694 11348
rect 16390 11336 16396 11348
rect 13688 11308 16396 11336
rect 13688 11296 13694 11308
rect 16390 11296 16396 11308
rect 16448 11336 16454 11348
rect 20438 11336 20444 11348
rect 16448 11308 20444 11336
rect 16448 11296 16454 11308
rect 20438 11296 20444 11308
rect 20496 11296 20502 11348
rect 20622 11296 20628 11348
rect 20680 11336 20686 11348
rect 20680 11308 21128 11336
rect 20680 11296 20686 11308
rect 14366 11268 14372 11280
rect 13556 11240 14372 11268
rect 14366 11228 14372 11240
rect 14424 11228 14430 11280
rect 15286 11268 15292 11280
rect 14476 11240 15292 11268
rect 12860 11172 13124 11200
rect 12860 11160 12866 11172
rect 13262 11160 13268 11212
rect 13320 11200 13326 11212
rect 14476 11200 14504 11240
rect 15286 11228 15292 11240
rect 15344 11228 15350 11280
rect 16758 11228 16764 11280
rect 16816 11268 16822 11280
rect 17221 11271 17279 11277
rect 17221 11268 17233 11271
rect 16816 11240 17233 11268
rect 16816 11228 16822 11240
rect 17221 11237 17233 11240
rect 17267 11237 17279 11271
rect 17221 11231 17279 11237
rect 18506 11228 18512 11280
rect 18564 11268 18570 11280
rect 18564 11240 20944 11268
rect 18564 11228 18570 11240
rect 15378 11200 15384 11212
rect 13320 11172 14504 11200
rect 14568 11172 15384 11200
rect 13320 11160 13326 11172
rect 12345 11135 12403 11141
rect 12345 11101 12357 11135
rect 12391 11101 12403 11135
rect 12621 11135 12679 11141
rect 12621 11132 12633 11135
rect 12345 11095 12403 11101
rect 12452 11104 12633 11132
rect 12268 11064 12296 11092
rect 12452 11064 12480 11104
rect 12621 11101 12633 11104
rect 12667 11101 12679 11135
rect 12621 11095 12679 11101
rect 12710 11092 12716 11144
rect 12768 11132 12774 11144
rect 13998 11132 14004 11144
rect 12768 11104 13492 11132
rect 12768 11092 12774 11104
rect 12084 11036 12296 11064
rect 12406 11036 12480 11064
rect 11793 11027 11851 11033
rect 4798 10956 4804 11008
rect 4856 10956 4862 11008
rect 10962 10956 10968 11008
rect 11020 10956 11026 11008
rect 11514 10956 11520 11008
rect 11572 10956 11578 11008
rect 12066 10956 12072 11008
rect 12124 10996 12130 11008
rect 12406 10996 12434 11036
rect 12526 11024 12532 11076
rect 12584 11024 12590 11076
rect 13262 11024 13268 11076
rect 13320 11024 13326 11076
rect 13078 11005 13084 11008
rect 12124 10968 12434 10996
rect 13065 10999 13084 11005
rect 12124 10956 12130 10968
rect 13065 10965 13077 10999
rect 13065 10959 13084 10965
rect 13078 10956 13084 10959
rect 13136 10956 13142 11008
rect 13464 10996 13492 11104
rect 13648 11104 14004 11132
rect 13525 11067 13583 11073
rect 13525 11033 13537 11067
rect 13571 11064 13583 11067
rect 13648 11064 13676 11104
rect 13998 11092 14004 11104
rect 14056 11092 14062 11144
rect 14292 11141 14320 11172
rect 14277 11135 14335 11141
rect 14277 11101 14289 11135
rect 14323 11101 14335 11135
rect 14277 11095 14335 11101
rect 14366 11092 14372 11144
rect 14424 11132 14430 11144
rect 14568 11132 14596 11172
rect 15378 11160 15384 11172
rect 15436 11160 15442 11212
rect 15473 11203 15531 11209
rect 15473 11169 15485 11203
rect 15519 11200 15531 11203
rect 18138 11200 18144 11212
rect 15519 11172 18144 11200
rect 15519 11169 15531 11172
rect 15473 11163 15531 11169
rect 18138 11160 18144 11172
rect 18196 11160 18202 11212
rect 19306 11172 20669 11200
rect 14424 11104 14596 11132
rect 14424 11092 14430 11104
rect 14642 11092 14648 11144
rect 14700 11092 14706 11144
rect 17034 11092 17040 11144
rect 17092 11132 17098 11144
rect 17770 11132 17776 11144
rect 17092 11104 17776 11132
rect 17092 11092 17098 11104
rect 17770 11092 17776 11104
rect 17828 11132 17834 11144
rect 19306 11132 19334 11172
rect 17828 11104 19334 11132
rect 17828 11092 17834 11104
rect 19518 11092 19524 11144
rect 19576 11092 19582 11144
rect 20530 11092 20536 11144
rect 20588 11092 20594 11144
rect 20641 11141 20669 11172
rect 20916 11141 20944 11240
rect 21100 11200 21128 11308
rect 21174 11296 21180 11348
rect 21232 11296 21238 11348
rect 22370 11296 22376 11348
rect 22428 11296 22434 11348
rect 22186 11268 22192 11280
rect 21744 11240 22192 11268
rect 21744 11200 21772 11240
rect 22186 11228 22192 11240
rect 22244 11228 22250 11280
rect 21910 11200 21916 11212
rect 21100 11172 21772 11200
rect 20626 11135 20684 11141
rect 20626 11101 20638 11135
rect 20672 11101 20684 11135
rect 20626 11095 20684 11101
rect 20901 11135 20959 11141
rect 20901 11101 20913 11135
rect 20947 11101 20959 11135
rect 20901 11095 20959 11101
rect 21039 11135 21097 11141
rect 21039 11101 21051 11135
rect 21085 11132 21097 11135
rect 21542 11132 21548 11144
rect 21085 11104 21548 11132
rect 21085 11101 21097 11104
rect 21039 11095 21097 11101
rect 13571 11036 13676 11064
rect 13725 11067 13783 11073
rect 13571 11033 13583 11036
rect 13525 11027 13583 11033
rect 13725 11033 13737 11067
rect 13771 11064 13783 11067
rect 13814 11064 13820 11076
rect 13771 11036 13820 11064
rect 13771 11033 13783 11036
rect 13725 11027 13783 11033
rect 13814 11024 13820 11036
rect 13872 11064 13878 11076
rect 14461 11067 14519 11073
rect 13872 11036 14412 11064
rect 13872 11024 13878 11036
rect 13906 10996 13912 11008
rect 13464 10968 13912 10996
rect 13906 10956 13912 10968
rect 13964 10956 13970 11008
rect 14090 10956 14096 11008
rect 14148 10956 14154 11008
rect 14384 10996 14412 11036
rect 14461 11033 14473 11067
rect 14507 11064 14519 11067
rect 15194 11064 15200 11076
rect 14507 11036 15200 11064
rect 14507 11033 14519 11036
rect 14461 11027 14519 11033
rect 15194 11024 15200 11036
rect 15252 11064 15258 11076
rect 15252 11036 15608 11064
rect 15252 11024 15258 11036
rect 15580 11008 15608 11036
rect 15746 11024 15752 11076
rect 15804 11024 15810 11076
rect 17126 11064 17132 11076
rect 16974 11036 17132 11064
rect 17126 11024 17132 11036
rect 17184 11064 17190 11076
rect 17402 11064 17408 11076
rect 17184 11036 17408 11064
rect 17184 11024 17190 11036
rect 17402 11024 17408 11036
rect 17460 11064 17466 11076
rect 17862 11064 17868 11076
rect 17460 11036 17868 11064
rect 17460 11024 17466 11036
rect 17862 11024 17868 11036
rect 17920 11024 17926 11076
rect 18690 11024 18696 11076
rect 18748 11064 18754 11076
rect 20809 11067 20867 11073
rect 20809 11064 20821 11067
rect 18748 11036 20821 11064
rect 18748 11024 18754 11036
rect 20809 11033 20821 11036
rect 20855 11033 20867 11067
rect 20916 11064 20944 11095
rect 21542 11092 21548 11104
rect 21600 11092 21606 11144
rect 21744 11141 21772 11172
rect 21836 11172 21916 11200
rect 21836 11141 21864 11172
rect 21910 11160 21916 11172
rect 21968 11160 21974 11212
rect 22462 11200 22468 11212
rect 22112 11172 22468 11200
rect 22112 11141 22140 11172
rect 22462 11160 22468 11172
rect 22520 11160 22526 11212
rect 24213 11203 24271 11209
rect 24213 11169 24225 11203
rect 24259 11200 24271 11203
rect 24394 11200 24400 11212
rect 24259 11172 24400 11200
rect 24259 11169 24271 11172
rect 24213 11163 24271 11169
rect 24394 11160 24400 11172
rect 24452 11160 24458 11212
rect 26234 11160 26240 11212
rect 26292 11200 26298 11212
rect 26329 11203 26387 11209
rect 26329 11200 26341 11203
rect 26292 11172 26341 11200
rect 26292 11160 26298 11172
rect 26329 11169 26341 11172
rect 26375 11169 26387 11203
rect 26329 11163 26387 11169
rect 26602 11160 26608 11212
rect 26660 11160 26666 11212
rect 28074 11160 28080 11212
rect 28132 11160 28138 11212
rect 21729 11135 21787 11141
rect 21729 11101 21741 11135
rect 21775 11101 21787 11135
rect 21729 11095 21787 11101
rect 21822 11135 21880 11141
rect 21822 11101 21834 11135
rect 21868 11101 21880 11135
rect 22097 11135 22155 11141
rect 22097 11132 22109 11135
rect 21822 11095 21880 11101
rect 21928 11104 22109 11132
rect 21928 11064 21956 11104
rect 22097 11101 22109 11104
rect 22143 11101 22155 11135
rect 22097 11095 22155 11101
rect 22235 11135 22293 11141
rect 22235 11101 22247 11135
rect 22281 11132 22293 11135
rect 22281 11104 22508 11132
rect 22281 11101 22293 11104
rect 22235 11095 22293 11101
rect 20916 11036 21956 11064
rect 22005 11067 22063 11073
rect 20809 11027 20867 11033
rect 22005 11033 22017 11067
rect 22051 11033 22063 11067
rect 22005 11027 22063 11033
rect 14642 10996 14648 11008
rect 14384 10968 14648 10996
rect 14642 10956 14648 10968
rect 14700 10956 14706 11008
rect 15562 10956 15568 11008
rect 15620 10956 15626 11008
rect 22020 10996 22048 11027
rect 22278 10996 22284 11008
rect 22020 10968 22284 10996
rect 22278 10956 22284 10968
rect 22336 10956 22342 11008
rect 22480 11005 22508 11104
rect 23382 11024 23388 11076
rect 23440 11024 23446 11076
rect 23934 11024 23940 11076
rect 23992 11024 23998 11076
rect 27890 11064 27896 11076
rect 27830 11036 27896 11064
rect 27890 11024 27896 11036
rect 27948 11024 27954 11076
rect 22465 10999 22523 11005
rect 22465 10965 22477 10999
rect 22511 10996 22523 10999
rect 23106 10996 23112 11008
rect 22511 10968 23112 10996
rect 22511 10965 22523 10968
rect 22465 10959 22523 10965
rect 23106 10956 23112 10968
rect 23164 10956 23170 11008
rect 1104 10906 28704 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 28704 10906
rect 1104 10832 28704 10854
rect 4798 10752 4804 10804
rect 4856 10792 4862 10804
rect 5445 10795 5503 10801
rect 5445 10792 5457 10795
rect 4856 10764 5457 10792
rect 4856 10752 4862 10764
rect 5445 10761 5457 10764
rect 5491 10761 5503 10795
rect 5445 10755 5503 10761
rect 6546 10752 6552 10804
rect 6604 10752 6610 10804
rect 12161 10795 12219 10801
rect 12161 10761 12173 10795
rect 12207 10792 12219 10795
rect 13078 10792 13084 10804
rect 12207 10764 13084 10792
rect 12207 10761 12219 10764
rect 12161 10755 12219 10761
rect 13078 10752 13084 10764
rect 13136 10752 13142 10804
rect 15473 10795 15531 10801
rect 15473 10761 15485 10795
rect 15519 10792 15531 10795
rect 15746 10792 15752 10804
rect 15519 10764 15752 10792
rect 15519 10761 15531 10764
rect 15473 10755 15531 10761
rect 15746 10752 15752 10764
rect 15804 10752 15810 10804
rect 16285 10795 16343 10801
rect 16285 10761 16297 10795
rect 16331 10792 16343 10795
rect 16666 10792 16672 10804
rect 16331 10764 16672 10792
rect 16331 10761 16343 10764
rect 16285 10755 16343 10761
rect 16666 10752 16672 10764
rect 16724 10752 16730 10804
rect 18598 10792 18604 10804
rect 16960 10764 18604 10792
rect 5000 10696 6132 10724
rect 5000 10665 5028 10696
rect 6104 10668 6132 10696
rect 7006 10684 7012 10736
rect 7064 10684 7070 10736
rect 8202 10724 8208 10736
rect 8036 10696 8208 10724
rect 4985 10659 5043 10665
rect 4985 10625 4997 10659
rect 5031 10625 5043 10659
rect 4985 10619 5043 10625
rect 5626 10616 5632 10668
rect 5684 10616 5690 10668
rect 5718 10616 5724 10668
rect 5776 10616 5782 10668
rect 5813 10659 5871 10665
rect 5813 10625 5825 10659
rect 5859 10625 5871 10659
rect 5813 10619 5871 10625
rect 5077 10591 5135 10597
rect 5077 10557 5089 10591
rect 5123 10557 5135 10591
rect 5077 10551 5135 10557
rect 5353 10591 5411 10597
rect 5353 10557 5365 10591
rect 5399 10588 5411 10591
rect 5828 10588 5856 10619
rect 5902 10616 5908 10668
rect 5960 10656 5966 10668
rect 5997 10659 6055 10665
rect 5997 10656 6009 10659
rect 5960 10628 6009 10656
rect 5960 10616 5966 10628
rect 5997 10625 6009 10628
rect 6043 10625 6055 10659
rect 5997 10619 6055 10625
rect 6086 10616 6092 10668
rect 6144 10656 6150 10668
rect 6365 10659 6423 10665
rect 6365 10656 6377 10659
rect 6144 10628 6377 10656
rect 6144 10616 6150 10628
rect 6365 10625 6377 10628
rect 6411 10625 6423 10659
rect 6365 10619 6423 10625
rect 6454 10616 6460 10668
rect 6512 10656 6518 10668
rect 8036 10665 8064 10696
rect 8202 10684 8208 10696
rect 8260 10684 8266 10736
rect 8294 10684 8300 10736
rect 8352 10684 8358 10736
rect 8754 10684 8760 10736
rect 8812 10684 8818 10736
rect 13262 10724 13268 10736
rect 12544 10696 13268 10724
rect 6549 10659 6607 10665
rect 6549 10656 6561 10659
rect 6512 10628 6561 10656
rect 6512 10616 6518 10628
rect 6549 10625 6561 10628
rect 6595 10625 6607 10659
rect 6549 10619 6607 10625
rect 6917 10659 6975 10665
rect 6917 10625 6929 10659
rect 6963 10625 6975 10659
rect 6917 10619 6975 10625
rect 8021 10659 8079 10665
rect 8021 10625 8033 10659
rect 8067 10625 8079 10659
rect 8021 10619 8079 10625
rect 10137 10659 10195 10665
rect 10137 10625 10149 10659
rect 10183 10656 10195 10659
rect 11514 10656 11520 10668
rect 10183 10628 11520 10656
rect 10183 10625 10195 10628
rect 10137 10619 10195 10625
rect 5399 10560 5856 10588
rect 6932 10588 6960 10619
rect 11514 10616 11520 10628
rect 11572 10616 11578 10668
rect 11793 10659 11851 10665
rect 11793 10625 11805 10659
rect 11839 10656 11851 10659
rect 12066 10656 12072 10668
rect 11839 10628 12072 10656
rect 11839 10625 11851 10628
rect 11793 10619 11851 10625
rect 12066 10616 12072 10628
rect 12124 10616 12130 10668
rect 12544 10665 12572 10696
rect 13262 10684 13268 10696
rect 13320 10724 13326 10736
rect 13449 10727 13507 10733
rect 13449 10724 13461 10727
rect 13320 10696 13461 10724
rect 13320 10684 13326 10696
rect 13449 10693 13461 10696
rect 13495 10693 13507 10727
rect 15657 10727 15715 10733
rect 15657 10724 15669 10727
rect 13449 10687 13507 10693
rect 15488 10696 15669 10724
rect 15488 10668 15516 10696
rect 15657 10693 15669 10696
rect 15703 10693 15715 10727
rect 15657 10687 15715 10693
rect 16390 10684 16396 10736
rect 16448 10724 16454 10736
rect 16485 10727 16543 10733
rect 16485 10724 16497 10727
rect 16448 10696 16497 10724
rect 16448 10684 16454 10696
rect 16485 10693 16497 10696
rect 16531 10724 16543 10727
rect 16960 10724 16988 10764
rect 18598 10752 18604 10764
rect 18656 10752 18662 10804
rect 22462 10752 22468 10804
rect 22520 10792 22526 10804
rect 22520 10764 22784 10792
rect 22520 10752 22526 10764
rect 16531 10696 16988 10724
rect 16531 10693 16543 10696
rect 16485 10687 16543 10693
rect 17862 10684 17868 10736
rect 17920 10684 17926 10736
rect 18230 10684 18236 10736
rect 18288 10724 18294 10736
rect 21450 10724 21456 10736
rect 18288 10696 18828 10724
rect 21298 10696 21456 10724
rect 18288 10684 18294 10696
rect 12529 10659 12587 10665
rect 12529 10625 12541 10659
rect 12575 10625 12587 10659
rect 12529 10619 12587 10625
rect 12621 10659 12679 10665
rect 12621 10625 12633 10659
rect 12667 10656 12679 10659
rect 12802 10656 12808 10668
rect 12667 10628 12808 10656
rect 12667 10625 12679 10628
rect 12621 10619 12679 10625
rect 12802 10616 12808 10628
rect 12860 10616 12866 10668
rect 13725 10659 13783 10665
rect 13725 10625 13737 10659
rect 13771 10656 13783 10659
rect 14642 10656 14648 10668
rect 13771 10628 14648 10656
rect 13771 10625 13783 10628
rect 13725 10619 13783 10625
rect 14642 10616 14648 10628
rect 14700 10616 14706 10668
rect 15470 10616 15476 10668
rect 15528 10616 15534 10668
rect 18800 10665 18828 10696
rect 21450 10684 21456 10696
rect 21508 10684 21514 10736
rect 22278 10684 22284 10736
rect 22336 10724 22342 10736
rect 22756 10733 22784 10764
rect 23934 10752 23940 10804
rect 23992 10792 23998 10804
rect 24305 10795 24363 10801
rect 24305 10792 24317 10795
rect 23992 10764 24317 10792
rect 23992 10752 23998 10764
rect 24305 10761 24317 10764
rect 24351 10761 24363 10795
rect 24305 10755 24363 10761
rect 26786 10752 26792 10804
rect 26844 10792 26850 10804
rect 26844 10764 27844 10792
rect 26844 10752 26850 10764
rect 22649 10727 22707 10733
rect 22649 10724 22661 10727
rect 22336 10696 22661 10724
rect 22336 10684 22342 10696
rect 22649 10693 22661 10696
rect 22695 10693 22707 10727
rect 22649 10687 22707 10693
rect 22741 10727 22799 10733
rect 22741 10693 22753 10727
rect 22787 10693 22799 10727
rect 24210 10724 24216 10736
rect 22741 10687 22799 10693
rect 23032 10696 24216 10724
rect 18785 10659 18843 10665
rect 18785 10625 18797 10659
rect 18831 10656 18843 10659
rect 19242 10656 19248 10668
rect 18831 10628 19248 10656
rect 18831 10625 18843 10628
rect 18785 10619 18843 10625
rect 19242 10616 19248 10628
rect 19300 10656 19306 10668
rect 19518 10656 19524 10668
rect 19300 10628 19524 10656
rect 19300 10616 19306 10628
rect 19518 10616 19524 10628
rect 19576 10656 19582 10668
rect 19797 10659 19855 10665
rect 19797 10656 19809 10659
rect 19576 10628 19809 10656
rect 19576 10616 19582 10628
rect 19797 10625 19809 10628
rect 19843 10625 19855 10659
rect 19797 10619 19855 10625
rect 22186 10616 22192 10668
rect 22244 10656 22250 10668
rect 22554 10665 22560 10668
rect 22373 10659 22431 10665
rect 22373 10656 22385 10659
rect 22244 10628 22385 10656
rect 22244 10616 22250 10628
rect 22373 10625 22385 10628
rect 22419 10625 22431 10659
rect 22373 10619 22431 10625
rect 22521 10659 22560 10665
rect 22521 10625 22533 10659
rect 22521 10619 22560 10625
rect 22554 10616 22560 10619
rect 22612 10616 22618 10668
rect 22879 10659 22937 10665
rect 22879 10625 22891 10659
rect 22925 10656 22937 10659
rect 23032 10656 23060 10696
rect 24210 10684 24216 10696
rect 24268 10684 24274 10736
rect 26053 10727 26111 10733
rect 26053 10693 26065 10727
rect 26099 10724 26111 10727
rect 26234 10724 26240 10736
rect 26099 10696 26240 10724
rect 26099 10693 26111 10696
rect 26053 10687 26111 10693
rect 26234 10684 26240 10696
rect 26292 10684 26298 10736
rect 26418 10684 26424 10736
rect 26476 10724 26482 10736
rect 26970 10724 26976 10736
rect 26476 10696 26976 10724
rect 26476 10684 26482 10696
rect 26970 10684 26976 10696
rect 27028 10724 27034 10736
rect 27249 10727 27307 10733
rect 27249 10724 27261 10727
rect 27028 10696 27261 10724
rect 27028 10684 27034 10696
rect 27249 10693 27261 10696
rect 27295 10693 27307 10727
rect 27249 10687 27307 10693
rect 22925 10628 23060 10656
rect 22925 10625 22937 10628
rect 22879 10619 22937 10625
rect 23106 10616 23112 10668
rect 23164 10616 23170 10668
rect 23474 10616 23480 10668
rect 23532 10656 23538 10668
rect 23937 10659 23995 10665
rect 23937 10656 23949 10659
rect 23532 10628 23949 10656
rect 23532 10616 23538 10628
rect 23937 10625 23949 10628
rect 23983 10625 23995 10659
rect 23937 10619 23995 10625
rect 24121 10659 24179 10665
rect 24121 10625 24133 10659
rect 24167 10625 24179 10659
rect 24121 10619 24179 10625
rect 7837 10591 7895 10597
rect 7837 10588 7849 10591
rect 6932 10560 7849 10588
rect 5399 10557 5411 10560
rect 5353 10551 5411 10557
rect 7837 10557 7849 10560
rect 7883 10557 7895 10591
rect 7837 10551 7895 10557
rect 5092 10520 5120 10551
rect 6362 10520 6368 10532
rect 5092 10492 6368 10520
rect 6362 10480 6368 10492
rect 6420 10480 6426 10532
rect 6546 10480 6552 10532
rect 6604 10520 6610 10532
rect 7190 10520 7196 10532
rect 6604 10492 7196 10520
rect 6604 10480 6610 10492
rect 7190 10480 7196 10492
rect 7248 10480 7254 10532
rect 7852 10452 7880 10551
rect 10318 10548 10324 10600
rect 10376 10548 10382 10600
rect 10413 10591 10471 10597
rect 10413 10557 10425 10591
rect 10459 10588 10471 10591
rect 10597 10591 10655 10597
rect 10597 10588 10609 10591
rect 10459 10560 10609 10588
rect 10459 10557 10471 10560
rect 10413 10551 10471 10557
rect 10597 10557 10609 10560
rect 10643 10557 10655 10591
rect 10597 10551 10655 10557
rect 10686 10548 10692 10600
rect 10744 10588 10750 10600
rect 11149 10591 11207 10597
rect 11149 10588 11161 10591
rect 10744 10560 11161 10588
rect 10744 10548 10750 10560
rect 11149 10557 11161 10560
rect 11195 10557 11207 10591
rect 11149 10551 11207 10557
rect 11882 10548 11888 10600
rect 11940 10548 11946 10600
rect 13449 10591 13507 10597
rect 13449 10557 13461 10591
rect 13495 10588 13507 10591
rect 13538 10588 13544 10600
rect 13495 10560 13544 10588
rect 13495 10557 13507 10560
rect 13449 10551 13507 10557
rect 13538 10548 13544 10560
rect 13596 10548 13602 10600
rect 13633 10591 13691 10597
rect 13633 10557 13645 10591
rect 13679 10588 13691 10591
rect 14090 10588 14096 10600
rect 13679 10560 14096 10588
rect 13679 10557 13691 10560
rect 13633 10551 13691 10557
rect 14090 10548 14096 10560
rect 14148 10548 14154 10600
rect 14200 10560 16988 10588
rect 9769 10523 9827 10529
rect 9769 10489 9781 10523
rect 9815 10520 9827 10523
rect 12250 10520 12256 10532
rect 9815 10492 12256 10520
rect 9815 10489 9827 10492
rect 9769 10483 9827 10489
rect 12250 10480 12256 10492
rect 12308 10480 12314 10532
rect 12805 10523 12863 10529
rect 12805 10489 12817 10523
rect 12851 10520 12863 10523
rect 12894 10520 12900 10532
rect 12851 10492 12900 10520
rect 12851 10489 12863 10492
rect 12805 10483 12863 10489
rect 12894 10480 12900 10492
rect 12952 10520 12958 10532
rect 14200 10520 14228 10560
rect 12952 10492 14228 10520
rect 12952 10480 12958 10492
rect 14274 10480 14280 10532
rect 14332 10520 14338 10532
rect 16025 10523 16083 10529
rect 16025 10520 16037 10523
rect 14332 10492 16037 10520
rect 14332 10480 14338 10492
rect 16025 10489 16037 10492
rect 16071 10520 16083 10523
rect 16117 10523 16175 10529
rect 16117 10520 16129 10523
rect 16071 10492 16129 10520
rect 16071 10489 16083 10492
rect 16025 10483 16083 10489
rect 16117 10489 16129 10492
rect 16163 10489 16175 10523
rect 16117 10483 16175 10489
rect 8754 10452 8760 10464
rect 7852 10424 8760 10452
rect 8754 10412 8760 10424
rect 8812 10412 8818 10464
rect 9950 10412 9956 10464
rect 10008 10412 10014 10464
rect 15654 10412 15660 10464
rect 15712 10412 15718 10464
rect 16301 10455 16359 10461
rect 16301 10421 16313 10455
rect 16347 10452 16359 10455
rect 16482 10452 16488 10464
rect 16347 10424 16488 10452
rect 16347 10421 16359 10424
rect 16301 10415 16359 10421
rect 16482 10412 16488 10424
rect 16540 10412 16546 10464
rect 16960 10452 16988 10560
rect 17034 10548 17040 10600
rect 17092 10548 17098 10600
rect 18506 10548 18512 10600
rect 18564 10548 18570 10600
rect 20070 10548 20076 10600
rect 20128 10548 20134 10600
rect 23753 10591 23811 10597
rect 23753 10557 23765 10591
rect 23799 10588 23811 10591
rect 23845 10591 23903 10597
rect 23845 10588 23857 10591
rect 23799 10560 23857 10588
rect 23799 10557 23811 10560
rect 23753 10551 23811 10557
rect 23845 10557 23857 10560
rect 23891 10557 23903 10591
rect 23845 10551 23903 10557
rect 23017 10523 23075 10529
rect 23017 10489 23029 10523
rect 23063 10520 23075 10523
rect 24136 10520 24164 10619
rect 24578 10616 24584 10668
rect 24636 10656 24642 10668
rect 25225 10659 25283 10665
rect 25225 10656 25237 10659
rect 24636 10628 25237 10656
rect 24636 10616 24642 10628
rect 25225 10625 25237 10628
rect 25271 10625 25283 10659
rect 25225 10619 25283 10625
rect 27246 10548 27252 10600
rect 27304 10588 27310 10600
rect 27356 10588 27384 10764
rect 27816 10733 27844 10764
rect 27801 10727 27859 10733
rect 27801 10693 27813 10727
rect 27847 10693 27859 10727
rect 27801 10687 27859 10693
rect 27433 10659 27491 10665
rect 27433 10625 27445 10659
rect 27479 10656 27491 10659
rect 27522 10656 27528 10668
rect 27479 10628 27528 10656
rect 27479 10625 27491 10628
rect 27433 10619 27491 10625
rect 27522 10616 27528 10628
rect 27580 10616 27586 10668
rect 27304 10560 27384 10588
rect 27304 10548 27310 10560
rect 23063 10492 24164 10520
rect 23063 10489 23075 10492
rect 23017 10483 23075 10489
rect 18322 10452 18328 10464
rect 16960 10424 18328 10452
rect 18322 10412 18328 10424
rect 18380 10412 18386 10464
rect 21542 10412 21548 10464
rect 21600 10452 21606 10464
rect 21910 10452 21916 10464
rect 21600 10424 21916 10452
rect 21600 10412 21606 10424
rect 21910 10412 21916 10424
rect 21968 10412 21974 10464
rect 27065 10455 27123 10461
rect 27065 10421 27077 10455
rect 27111 10452 27123 10455
rect 27430 10452 27436 10464
rect 27111 10424 27436 10452
rect 27111 10421 27123 10424
rect 27065 10415 27123 10421
rect 27430 10412 27436 10424
rect 27488 10412 27494 10464
rect 27890 10412 27896 10464
rect 27948 10412 27954 10464
rect 1104 10362 28704 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 28704 10362
rect 1104 10288 28704 10310
rect 5445 10251 5503 10257
rect 5445 10217 5457 10251
rect 5491 10248 5503 10251
rect 6086 10248 6092 10260
rect 5491 10220 6092 10248
rect 5491 10217 5503 10220
rect 5445 10211 5503 10217
rect 6086 10208 6092 10220
rect 6144 10208 6150 10260
rect 13998 10208 14004 10260
rect 14056 10248 14062 10260
rect 14093 10251 14151 10257
rect 14093 10248 14105 10251
rect 14056 10220 14105 10248
rect 14056 10208 14062 10220
rect 14093 10217 14105 10220
rect 14139 10217 14151 10251
rect 14093 10211 14151 10217
rect 15654 10208 15660 10260
rect 15712 10208 15718 10260
rect 15930 10208 15936 10260
rect 15988 10248 15994 10260
rect 16390 10248 16396 10260
rect 15988 10220 16396 10248
rect 15988 10208 15994 10220
rect 16390 10208 16396 10220
rect 16448 10208 16454 10260
rect 16666 10208 16672 10260
rect 16724 10248 16730 10260
rect 18417 10251 18475 10257
rect 18417 10248 18429 10251
rect 16724 10220 18429 10248
rect 16724 10208 16730 10220
rect 18417 10217 18429 10220
rect 18463 10217 18475 10251
rect 18417 10211 18475 10217
rect 7650 10140 7656 10192
rect 7708 10140 7714 10192
rect 6270 10112 6276 10124
rect 5276 10084 6276 10112
rect 5276 10053 5304 10084
rect 6270 10072 6276 10084
rect 6328 10072 6334 10124
rect 6549 10115 6607 10121
rect 6549 10081 6561 10115
rect 6595 10112 6607 10115
rect 7009 10115 7067 10121
rect 7009 10112 7021 10115
rect 6595 10084 7021 10112
rect 6595 10081 6607 10084
rect 6549 10075 6607 10081
rect 7009 10081 7021 10084
rect 7055 10081 7067 10115
rect 7009 10075 7067 10081
rect 7101 10115 7159 10121
rect 7101 10081 7113 10115
rect 7147 10112 7159 10115
rect 7282 10112 7288 10124
rect 7147 10084 7288 10112
rect 7147 10081 7159 10084
rect 7101 10075 7159 10081
rect 7282 10072 7288 10084
rect 7340 10072 7346 10124
rect 9217 10115 9275 10121
rect 9217 10081 9229 10115
rect 9263 10112 9275 10115
rect 9950 10112 9956 10124
rect 9263 10084 9956 10112
rect 9263 10081 9275 10084
rect 9217 10075 9275 10081
rect 9950 10072 9956 10084
rect 10008 10072 10014 10124
rect 14182 10072 14188 10124
rect 14240 10112 14246 10124
rect 14461 10115 14519 10121
rect 14461 10112 14473 10115
rect 14240 10084 14473 10112
rect 14240 10072 14246 10084
rect 14461 10081 14473 10084
rect 14507 10112 14519 10115
rect 14550 10112 14556 10124
rect 14507 10084 14556 10112
rect 14507 10081 14519 10084
rect 14461 10075 14519 10081
rect 14550 10072 14556 10084
rect 14608 10072 14614 10124
rect 15841 10115 15899 10121
rect 15841 10081 15853 10115
rect 15887 10112 15899 10115
rect 16850 10112 16856 10124
rect 15887 10084 16856 10112
rect 15887 10081 15899 10084
rect 15841 10075 15899 10081
rect 16850 10072 16856 10084
rect 16908 10072 16914 10124
rect 18138 10072 18144 10124
rect 18196 10072 18202 10124
rect 18233 10115 18291 10121
rect 18233 10081 18245 10115
rect 18279 10112 18291 10115
rect 18322 10112 18328 10124
rect 18279 10084 18328 10112
rect 18279 10081 18291 10084
rect 18233 10075 18291 10081
rect 18322 10072 18328 10084
rect 18380 10072 18386 10124
rect 18432 10112 18460 10211
rect 18506 10208 18512 10260
rect 18564 10248 18570 10260
rect 18601 10251 18659 10257
rect 18601 10248 18613 10251
rect 18564 10220 18613 10248
rect 18564 10208 18570 10220
rect 18601 10217 18613 10220
rect 18647 10217 18659 10251
rect 18601 10211 18659 10217
rect 18432 10084 18828 10112
rect 5261 10047 5319 10053
rect 5261 10013 5273 10047
rect 5307 10013 5319 10047
rect 5261 10007 5319 10013
rect 5445 10047 5503 10053
rect 5445 10013 5457 10047
rect 5491 10044 5503 10047
rect 5994 10044 6000 10056
rect 5491 10016 6000 10044
rect 5491 10013 5503 10016
rect 5445 10007 5503 10013
rect 5994 10004 6000 10016
rect 6052 10004 6058 10056
rect 6638 10004 6644 10056
rect 6696 10004 6702 10056
rect 6730 10004 6736 10056
rect 6788 10004 6794 10056
rect 6914 10004 6920 10056
rect 6972 10004 6978 10056
rect 7190 10004 7196 10056
rect 7248 10004 7254 10056
rect 7653 10047 7711 10053
rect 7653 10044 7665 10047
rect 7300 10016 7665 10044
rect 6822 9936 6828 9988
rect 6880 9976 6886 9988
rect 7300 9976 7328 10016
rect 7653 10013 7665 10016
rect 7699 10013 7711 10047
rect 7653 10007 7711 10013
rect 7834 10004 7840 10056
rect 7892 10004 7898 10056
rect 8754 10004 8760 10056
rect 8812 10044 8818 10056
rect 8941 10047 8999 10053
rect 8941 10044 8953 10047
rect 8812 10016 8953 10044
rect 8812 10004 8818 10016
rect 8941 10013 8953 10016
rect 8987 10013 8999 10047
rect 8941 10007 8999 10013
rect 12529 10047 12587 10053
rect 12529 10013 12541 10047
rect 12575 10044 12587 10047
rect 13630 10044 13636 10056
rect 12575 10016 13636 10044
rect 12575 10013 12587 10016
rect 12529 10007 12587 10013
rect 13630 10004 13636 10016
rect 13688 10004 13694 10056
rect 14274 10004 14280 10056
rect 14332 10004 14338 10056
rect 15930 10004 15936 10056
rect 15988 10004 15994 10056
rect 16025 10047 16083 10053
rect 16025 10013 16037 10047
rect 16071 10013 16083 10047
rect 16025 10007 16083 10013
rect 16117 10047 16175 10053
rect 16117 10013 16129 10047
rect 16163 10044 16175 10047
rect 16482 10044 16488 10056
rect 16163 10016 16488 10044
rect 16163 10013 16175 10016
rect 16117 10007 16175 10013
rect 6880 9948 7328 9976
rect 7377 9979 7435 9985
rect 6880 9936 6886 9948
rect 7377 9945 7389 9979
rect 7423 9976 7435 9979
rect 7469 9979 7527 9985
rect 7469 9976 7481 9979
rect 7423 9948 7481 9976
rect 7423 9945 7435 9948
rect 7377 9939 7435 9945
rect 7469 9945 7481 9948
rect 7515 9945 7527 9979
rect 11793 9979 11851 9985
rect 10442 9948 10916 9976
rect 7469 9939 7527 9945
rect 10888 9920 10916 9948
rect 11793 9945 11805 9979
rect 11839 9976 11851 9979
rect 11882 9976 11888 9988
rect 11839 9948 11888 9976
rect 11839 9945 11851 9948
rect 11793 9939 11851 9945
rect 11882 9936 11888 9948
rect 11940 9936 11946 9988
rect 16040 9976 16068 10007
rect 16482 10004 16488 10016
rect 16540 10004 16546 10056
rect 18506 10004 18512 10056
rect 18564 10004 18570 10056
rect 18598 10004 18604 10056
rect 18656 10004 18662 10056
rect 18800 10053 18828 10084
rect 19518 10072 19524 10124
rect 19576 10112 19582 10124
rect 19613 10115 19671 10121
rect 19613 10112 19625 10115
rect 19576 10084 19625 10112
rect 19576 10072 19582 10084
rect 19613 10081 19625 10084
rect 19659 10081 19671 10115
rect 19613 10075 19671 10081
rect 26234 10072 26240 10124
rect 26292 10112 26298 10124
rect 26513 10115 26571 10121
rect 26513 10112 26525 10115
rect 26292 10084 26525 10112
rect 26292 10072 26298 10084
rect 26513 10081 26525 10084
rect 26559 10081 26571 10115
rect 26513 10075 26571 10081
rect 26789 10115 26847 10121
rect 26789 10081 26801 10115
rect 26835 10112 26847 10115
rect 27338 10112 27344 10124
rect 26835 10084 27344 10112
rect 26835 10081 26847 10084
rect 26789 10075 26847 10081
rect 27338 10072 27344 10084
rect 27396 10072 27402 10124
rect 18785 10047 18843 10053
rect 18785 10013 18797 10047
rect 18831 10013 18843 10047
rect 18785 10007 18843 10013
rect 20438 10004 20444 10056
rect 20496 10044 20502 10056
rect 22738 10044 22744 10056
rect 20496 10016 22744 10044
rect 20496 10004 20502 10016
rect 22738 10004 22744 10016
rect 22796 10044 22802 10056
rect 24578 10044 24584 10056
rect 22796 10016 24584 10044
rect 22796 10004 22802 10016
rect 24578 10004 24584 10016
rect 24636 10004 24642 10056
rect 26418 10004 26424 10056
rect 26476 10004 26482 10056
rect 27890 10004 27896 10056
rect 27948 10004 27954 10056
rect 16040 9948 16160 9976
rect 9950 9868 9956 9920
rect 10008 9908 10014 9920
rect 10686 9908 10692 9920
rect 10008 9880 10692 9908
rect 10008 9868 10014 9880
rect 10686 9868 10692 9880
rect 10744 9868 10750 9920
rect 10870 9868 10876 9920
rect 10928 9908 10934 9920
rect 14458 9908 14464 9920
rect 10928 9880 14464 9908
rect 10928 9868 10934 9880
rect 14458 9868 14464 9880
rect 14516 9868 14522 9920
rect 16132 9908 16160 9948
rect 17402 9936 17408 9988
rect 17460 9936 17466 9988
rect 17862 9936 17868 9988
rect 17920 9936 17926 9988
rect 20346 9936 20352 9988
rect 20404 9976 20410 9988
rect 20533 9979 20591 9985
rect 20533 9976 20545 9979
rect 20404 9948 20545 9976
rect 20404 9936 20410 9948
rect 20533 9945 20545 9948
rect 20579 9945 20591 9979
rect 20533 9939 20591 9945
rect 20714 9936 20720 9988
rect 20772 9976 20778 9988
rect 21818 9976 21824 9988
rect 20772 9948 21824 9976
rect 20772 9936 20778 9948
rect 21818 9936 21824 9948
rect 21876 9936 21882 9988
rect 24762 9936 24768 9988
rect 24820 9976 24826 9988
rect 25317 9979 25375 9985
rect 25317 9976 25329 9979
rect 24820 9948 25329 9976
rect 24820 9936 24826 9948
rect 25317 9945 25329 9948
rect 25363 9945 25375 9979
rect 25317 9939 25375 9945
rect 17034 9908 17040 9920
rect 16132 9880 17040 9908
rect 17034 9868 17040 9880
rect 17092 9868 17098 9920
rect 18230 9868 18236 9920
rect 18288 9868 18294 9920
rect 20898 9868 20904 9920
rect 20956 9868 20962 9920
rect 26326 9868 26332 9920
rect 26384 9868 26390 9920
rect 27522 9868 27528 9920
rect 27580 9908 27586 9920
rect 28261 9911 28319 9917
rect 28261 9908 28273 9911
rect 27580 9880 28273 9908
rect 27580 9868 27586 9880
rect 28261 9877 28273 9880
rect 28307 9877 28319 9911
rect 28261 9871 28319 9877
rect 1104 9818 28704 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 28704 9818
rect 1104 9744 28704 9766
rect 6362 9664 6368 9716
rect 6420 9664 6426 9716
rect 7561 9707 7619 9713
rect 7561 9673 7573 9707
rect 7607 9704 7619 9707
rect 7834 9704 7840 9716
rect 7607 9676 7840 9704
rect 7607 9673 7619 9676
rect 7561 9667 7619 9673
rect 7834 9664 7840 9676
rect 7892 9664 7898 9716
rect 14016 9676 14688 9704
rect 14016 9648 14044 9676
rect 6638 9596 6644 9648
rect 6696 9636 6702 9648
rect 6696 9608 7052 9636
rect 6696 9596 6702 9608
rect 6549 9571 6607 9577
rect 6549 9537 6561 9571
rect 6595 9537 6607 9571
rect 6549 9531 6607 9537
rect 6825 9571 6883 9577
rect 6825 9537 6837 9571
rect 6871 9568 6883 9571
rect 6914 9568 6920 9580
rect 6871 9540 6920 9568
rect 6871 9537 6883 9540
rect 6825 9531 6883 9537
rect 6564 9432 6592 9531
rect 6914 9528 6920 9540
rect 6972 9528 6978 9580
rect 7024 9577 7052 9608
rect 7190 9596 7196 9648
rect 7248 9596 7254 9648
rect 12713 9639 12771 9645
rect 12713 9605 12725 9639
rect 12759 9636 12771 9639
rect 13081 9639 13139 9645
rect 13081 9636 13093 9639
rect 12759 9608 13093 9636
rect 12759 9605 12771 9608
rect 12713 9599 12771 9605
rect 13081 9605 13093 9608
rect 13127 9605 13139 9639
rect 13998 9636 14004 9648
rect 13081 9599 13139 9605
rect 13280 9608 14004 9636
rect 7009 9571 7067 9577
rect 7009 9537 7021 9571
rect 7055 9537 7067 9571
rect 7009 9531 7067 9537
rect 7098 9528 7104 9580
rect 7156 9528 7162 9580
rect 7208 9568 7236 9596
rect 7377 9571 7435 9577
rect 7377 9568 7389 9571
rect 7208 9540 7389 9568
rect 7377 9537 7389 9540
rect 7423 9537 7435 9571
rect 7377 9531 7435 9537
rect 10594 9528 10600 9580
rect 10652 9568 10658 9580
rect 10870 9568 10876 9580
rect 10652 9540 10876 9568
rect 10652 9528 10658 9540
rect 10870 9528 10876 9540
rect 10928 9528 10934 9580
rect 11882 9528 11888 9580
rect 11940 9528 11946 9580
rect 13280 9577 13308 9608
rect 13998 9596 14004 9608
rect 14056 9596 14062 9648
rect 14461 9639 14519 9645
rect 14461 9605 14473 9639
rect 14507 9605 14519 9639
rect 14461 9599 14519 9605
rect 12897 9571 12955 9577
rect 12897 9537 12909 9571
rect 12943 9537 12955 9571
rect 12897 9531 12955 9537
rect 12989 9571 13047 9577
rect 12989 9537 13001 9571
rect 13035 9568 13047 9571
rect 13265 9571 13323 9577
rect 13265 9568 13277 9571
rect 13035 9540 13277 9568
rect 13035 9537 13047 9540
rect 12989 9531 13047 9537
rect 13265 9537 13277 9540
rect 13311 9537 13323 9571
rect 13265 9531 13323 9537
rect 13357 9571 13415 9577
rect 13357 9537 13369 9571
rect 13403 9537 13415 9571
rect 13357 9531 13415 9537
rect 7190 9460 7196 9512
rect 7248 9460 7254 9512
rect 12912 9500 12940 9531
rect 12912 9472 13032 9500
rect 7006 9432 7012 9444
rect 6564 9404 7012 9432
rect 7006 9392 7012 9404
rect 7064 9432 7070 9444
rect 13004 9432 13032 9472
rect 13078 9460 13084 9512
rect 13136 9460 13142 9512
rect 13372 9500 13400 9531
rect 14182 9528 14188 9580
rect 14240 9528 14246 9580
rect 14274 9528 14280 9580
rect 14332 9528 14338 9580
rect 14476 9568 14504 9599
rect 14553 9571 14611 9577
rect 14553 9568 14565 9571
rect 14476 9540 14565 9568
rect 14553 9537 14565 9540
rect 14599 9537 14611 9571
rect 14660 9568 14688 9676
rect 18322 9664 18328 9716
rect 18380 9704 18386 9716
rect 18380 9676 19196 9704
rect 18380 9664 18386 9676
rect 17497 9639 17555 9645
rect 17497 9605 17509 9639
rect 17543 9636 17555 9639
rect 17681 9639 17739 9645
rect 17681 9636 17693 9639
rect 17543 9608 17693 9636
rect 17543 9605 17555 9608
rect 17497 9599 17555 9605
rect 17681 9605 17693 9608
rect 17727 9605 17739 9639
rect 17681 9599 17739 9605
rect 17865 9639 17923 9645
rect 17865 9605 17877 9639
rect 17911 9636 17923 9639
rect 18230 9636 18236 9648
rect 17911 9608 18236 9636
rect 17911 9605 17923 9608
rect 17865 9599 17923 9605
rect 18230 9596 18236 9608
rect 18288 9596 18294 9648
rect 18782 9596 18788 9648
rect 18840 9636 18846 9648
rect 19061 9639 19119 9645
rect 19061 9636 19073 9639
rect 18840 9608 19073 9636
rect 18840 9596 18846 9608
rect 19061 9605 19073 9608
rect 19107 9605 19119 9639
rect 19061 9599 19119 9605
rect 14737 9571 14795 9577
rect 14737 9568 14749 9571
rect 14660 9540 14749 9568
rect 14553 9531 14611 9537
rect 14737 9537 14749 9540
rect 14783 9537 14795 9571
rect 14737 9531 14795 9537
rect 16666 9528 16672 9580
rect 16724 9568 16730 9580
rect 17589 9571 17647 9577
rect 17589 9568 17601 9571
rect 16724 9540 17601 9568
rect 16724 9528 16730 9540
rect 17589 9537 17601 9540
rect 17635 9537 17647 9571
rect 17589 9531 17647 9537
rect 17770 9528 17776 9580
rect 17828 9568 17834 9580
rect 17957 9571 18015 9577
rect 17957 9568 17969 9571
rect 17828 9540 17969 9568
rect 17828 9528 17834 9540
rect 17957 9537 17969 9540
rect 18003 9537 18015 9571
rect 17957 9531 18015 9537
rect 13814 9500 13820 9512
rect 13372 9472 13820 9500
rect 13814 9460 13820 9472
rect 13872 9500 13878 9512
rect 14090 9500 14096 9512
rect 13872 9472 14096 9500
rect 13872 9460 13878 9472
rect 14090 9460 14096 9472
rect 14148 9460 14154 9512
rect 14461 9503 14519 9509
rect 14461 9469 14473 9503
rect 14507 9500 14519 9503
rect 15470 9500 15476 9512
rect 14507 9472 15476 9500
rect 14507 9469 14519 9472
rect 14461 9463 14519 9469
rect 13449 9435 13507 9441
rect 13449 9432 13461 9435
rect 7064 9404 7328 9432
rect 13004 9404 13461 9432
rect 7064 9392 7070 9404
rect 7300 9376 7328 9404
rect 13449 9401 13461 9404
rect 13495 9401 13507 9435
rect 13449 9395 13507 9401
rect 7282 9324 7288 9376
rect 7340 9324 7346 9376
rect 9858 9324 9864 9376
rect 9916 9364 9922 9376
rect 10962 9364 10968 9376
rect 9916 9336 10968 9364
rect 9916 9324 9922 9336
rect 10962 9324 10968 9336
rect 11020 9324 11026 9376
rect 12342 9324 12348 9376
rect 12400 9364 12406 9376
rect 12713 9367 12771 9373
rect 12713 9364 12725 9367
rect 12400 9336 12725 9364
rect 12400 9324 12406 9336
rect 12713 9333 12725 9336
rect 12759 9333 12771 9367
rect 12713 9327 12771 9333
rect 13078 9324 13084 9376
rect 13136 9364 13142 9376
rect 14476 9364 14504 9463
rect 15470 9460 15476 9472
rect 15528 9460 15534 9512
rect 16390 9460 16396 9512
rect 16448 9500 16454 9512
rect 16853 9503 16911 9509
rect 16853 9500 16865 9503
rect 16448 9472 16865 9500
rect 16448 9460 16454 9472
rect 16853 9469 16865 9472
rect 16899 9469 16911 9503
rect 16853 9463 16911 9469
rect 18233 9503 18291 9509
rect 18233 9469 18245 9503
rect 18279 9500 18291 9503
rect 18322 9500 18328 9512
rect 18279 9472 18328 9500
rect 18279 9469 18291 9472
rect 18233 9463 18291 9469
rect 18322 9460 18328 9472
rect 18380 9460 18386 9512
rect 19076 9500 19104 9599
rect 19168 9568 19196 9676
rect 20070 9664 20076 9716
rect 20128 9664 20134 9716
rect 27430 9704 27436 9716
rect 26252 9676 27436 9704
rect 19277 9639 19335 9645
rect 19277 9605 19289 9639
rect 19323 9636 19335 9639
rect 19794 9636 19800 9648
rect 19323 9608 19800 9636
rect 19323 9605 19335 9608
rect 19277 9599 19335 9605
rect 19794 9596 19800 9608
rect 19852 9596 19858 9648
rect 19889 9639 19947 9645
rect 19889 9605 19901 9639
rect 19935 9605 19947 9639
rect 22646 9636 22652 9648
rect 19889 9599 19947 9605
rect 20456 9608 22652 9636
rect 19904 9568 19932 9599
rect 20254 9568 20260 9580
rect 19168 9540 20260 9568
rect 20254 9528 20260 9540
rect 20312 9528 20318 9580
rect 20346 9528 20352 9580
rect 20404 9528 20410 9580
rect 20456 9512 20484 9608
rect 22646 9596 22652 9608
rect 22704 9596 22710 9648
rect 22738 9596 22744 9648
rect 22796 9596 22802 9648
rect 26252 9636 26280 9676
rect 27430 9664 27436 9676
rect 27488 9664 27494 9716
rect 26068 9608 26280 9636
rect 26482 9608 27476 9636
rect 20533 9571 20591 9577
rect 20533 9537 20545 9571
rect 20579 9568 20591 9571
rect 20714 9568 20720 9580
rect 20579 9540 20720 9568
rect 20579 9537 20591 9540
rect 20533 9531 20591 9537
rect 20714 9528 20720 9540
rect 20772 9528 20778 9580
rect 21174 9528 21180 9580
rect 21232 9568 21238 9580
rect 21453 9571 21511 9577
rect 21453 9568 21465 9571
rect 21232 9540 21465 9568
rect 21232 9528 21238 9540
rect 21453 9537 21465 9540
rect 21499 9568 21511 9571
rect 21913 9571 21971 9577
rect 21913 9568 21925 9571
rect 21499 9540 21925 9568
rect 21499 9537 21511 9540
rect 21453 9531 21511 9537
rect 21913 9537 21925 9540
rect 21959 9537 21971 9571
rect 21913 9531 21971 9537
rect 23658 9528 23664 9580
rect 23716 9568 23722 9580
rect 24581 9571 24639 9577
rect 24581 9568 24593 9571
rect 23716 9540 24593 9568
rect 23716 9528 23722 9540
rect 24581 9537 24593 9540
rect 24627 9568 24639 9571
rect 24762 9568 24768 9580
rect 24627 9540 24768 9568
rect 24627 9537 24639 9540
rect 24581 9531 24639 9537
rect 24762 9528 24768 9540
rect 24820 9528 24826 9580
rect 26068 9577 26096 9608
rect 26053 9571 26111 9577
rect 26053 9537 26065 9571
rect 26099 9537 26111 9571
rect 26053 9531 26111 9537
rect 26234 9528 26240 9580
rect 26292 9528 26298 9580
rect 26326 9528 26332 9580
rect 26384 9528 26390 9580
rect 26482 9577 26510 9608
rect 26467 9571 26525 9577
rect 26467 9537 26479 9571
rect 26513 9537 26525 9571
rect 26467 9531 26525 9537
rect 26786 9528 26792 9580
rect 26844 9568 26850 9580
rect 27448 9568 27476 9608
rect 27522 9568 27528 9580
rect 26844 9540 27384 9568
rect 27448 9540 27528 9568
rect 26844 9528 26850 9540
rect 20438 9500 20444 9512
rect 19076 9472 20444 9500
rect 20438 9460 20444 9472
rect 20496 9460 20502 9512
rect 20625 9503 20683 9509
rect 20625 9469 20637 9503
rect 20671 9469 20683 9503
rect 20625 9463 20683 9469
rect 26605 9503 26663 9509
rect 26605 9469 26617 9503
rect 26651 9500 26663 9503
rect 26878 9500 26884 9512
rect 26651 9472 26884 9500
rect 26651 9469 26663 9472
rect 26605 9463 26663 9469
rect 17862 9392 17868 9444
rect 17920 9392 17926 9444
rect 18141 9435 18199 9441
rect 18141 9401 18153 9435
rect 18187 9432 18199 9435
rect 18598 9432 18604 9444
rect 18187 9404 18604 9432
rect 18187 9401 18199 9404
rect 18141 9395 18199 9401
rect 18598 9392 18604 9404
rect 18656 9392 18662 9444
rect 19429 9435 19487 9441
rect 19429 9432 19441 9435
rect 18800 9404 19441 9432
rect 13136 9336 14504 9364
rect 13136 9324 13142 9336
rect 14550 9324 14556 9376
rect 14608 9324 14614 9376
rect 16850 9324 16856 9376
rect 16908 9364 16914 9376
rect 18049 9367 18107 9373
rect 18049 9364 18061 9367
rect 16908 9336 18061 9364
rect 16908 9324 16914 9336
rect 18049 9333 18061 9336
rect 18095 9364 18107 9367
rect 18800 9364 18828 9404
rect 19429 9401 19441 9404
rect 19475 9432 19487 9435
rect 19521 9435 19579 9441
rect 19521 9432 19533 9435
rect 19475 9404 19533 9432
rect 19475 9401 19487 9404
rect 19429 9395 19487 9401
rect 19521 9401 19533 9404
rect 19567 9401 19579 9435
rect 19521 9395 19579 9401
rect 19812 9404 20392 9432
rect 18095 9336 18828 9364
rect 18095 9333 18107 9336
rect 18049 9327 18107 9333
rect 19242 9324 19248 9376
rect 19300 9364 19306 9376
rect 19812 9364 19840 9404
rect 19300 9336 19840 9364
rect 19889 9367 19947 9373
rect 19300 9324 19306 9336
rect 19889 9333 19901 9367
rect 19935 9364 19947 9367
rect 20165 9367 20223 9373
rect 20165 9364 20177 9367
rect 19935 9336 20177 9364
rect 19935 9333 19947 9336
rect 19889 9327 19947 9333
rect 20165 9333 20177 9336
rect 20211 9333 20223 9367
rect 20364 9364 20392 9404
rect 20640 9364 20668 9463
rect 26878 9460 26884 9472
rect 26936 9500 26942 9512
rect 27249 9503 27307 9509
rect 27249 9500 27261 9503
rect 26936 9472 27261 9500
rect 26936 9460 26942 9472
rect 27249 9469 27261 9472
rect 27295 9469 27307 9503
rect 27356 9500 27384 9540
rect 27522 9528 27528 9540
rect 27580 9528 27586 9580
rect 27893 9571 27951 9577
rect 27893 9537 27905 9571
rect 27939 9568 27951 9571
rect 28074 9568 28080 9580
rect 27939 9540 28080 9568
rect 27939 9537 27951 9540
rect 27893 9531 27951 9537
rect 28074 9528 28080 9540
rect 28132 9528 28138 9580
rect 28166 9528 28172 9580
rect 28224 9528 28230 9580
rect 27356 9472 27660 9500
rect 27249 9463 27307 9469
rect 25682 9392 25688 9444
rect 25740 9432 25746 9444
rect 27632 9441 27660 9472
rect 26697 9435 26755 9441
rect 26697 9432 26709 9435
rect 25740 9404 26709 9432
rect 25740 9392 25746 9404
rect 26697 9401 26709 9404
rect 26743 9401 26755 9435
rect 26697 9395 26755 9401
rect 27617 9435 27675 9441
rect 27617 9401 27629 9435
rect 27663 9401 27675 9435
rect 27617 9395 27675 9401
rect 21542 9364 21548 9376
rect 20364 9336 21548 9364
rect 20165 9327 20223 9333
rect 21542 9324 21548 9336
rect 21600 9324 21606 9376
rect 25866 9324 25872 9376
rect 25924 9364 25930 9376
rect 26053 9367 26111 9373
rect 26053 9364 26065 9367
rect 25924 9336 26065 9364
rect 25924 9324 25930 9336
rect 26053 9333 26065 9336
rect 26099 9333 26111 9367
rect 26053 9327 26111 9333
rect 26970 9324 26976 9376
rect 27028 9324 27034 9376
rect 27062 9324 27068 9376
rect 27120 9364 27126 9376
rect 27157 9367 27215 9373
rect 27157 9364 27169 9367
rect 27120 9336 27169 9364
rect 27120 9324 27126 9336
rect 27157 9333 27169 9336
rect 27203 9333 27215 9367
rect 27157 9327 27215 9333
rect 27430 9324 27436 9376
rect 27488 9364 27494 9376
rect 27801 9367 27859 9373
rect 27801 9364 27813 9367
rect 27488 9336 27813 9364
rect 27488 9324 27494 9336
rect 27801 9333 27813 9336
rect 27847 9333 27859 9367
rect 27801 9327 27859 9333
rect 1104 9274 28704 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 28704 9274
rect 1104 9200 28704 9222
rect 6638 9120 6644 9172
rect 6696 9160 6702 9172
rect 6733 9163 6791 9169
rect 6733 9160 6745 9163
rect 6696 9132 6745 9160
rect 6696 9120 6702 9132
rect 6733 9129 6745 9132
rect 6779 9129 6791 9163
rect 6733 9123 6791 9129
rect 7282 9120 7288 9172
rect 7340 9160 7346 9172
rect 7340 9132 14596 9160
rect 7340 9120 7346 9132
rect 6454 9052 6460 9104
rect 6512 9092 6518 9104
rect 10137 9095 10195 9101
rect 6512 9064 7236 9092
rect 6512 9052 6518 9064
rect 6549 9027 6607 9033
rect 6549 9024 6561 9027
rect 6380 8996 6561 9024
rect 5626 8916 5632 8968
rect 5684 8916 5690 8968
rect 6380 8965 6408 8996
rect 6549 8993 6561 8996
rect 6595 9024 6607 9027
rect 7006 9024 7012 9036
rect 6595 8996 7012 9024
rect 6595 8993 6607 8996
rect 6549 8987 6607 8993
rect 7006 8984 7012 8996
rect 7064 8984 7070 9036
rect 7208 9033 7236 9064
rect 10137 9061 10149 9095
rect 10183 9061 10195 9095
rect 14568 9092 14596 9132
rect 14642 9120 14648 9172
rect 14700 9120 14706 9172
rect 16666 9120 16672 9172
rect 16724 9120 16730 9172
rect 17586 9120 17592 9172
rect 17644 9160 17650 9172
rect 19242 9160 19248 9172
rect 17644 9132 19248 9160
rect 17644 9120 17650 9132
rect 19242 9120 19248 9132
rect 19300 9120 19306 9172
rect 19794 9120 19800 9172
rect 19852 9160 19858 9172
rect 20165 9163 20223 9169
rect 20165 9160 20177 9163
rect 19852 9132 20177 9160
rect 19852 9120 19858 9132
rect 20165 9129 20177 9132
rect 20211 9160 20223 9163
rect 20625 9163 20683 9169
rect 20211 9132 20300 9160
rect 20211 9129 20223 9132
rect 20165 9123 20223 9129
rect 15562 9092 15568 9104
rect 14568 9064 15568 9092
rect 10137 9055 10195 9061
rect 7193 9027 7251 9033
rect 7193 8993 7205 9027
rect 7239 8993 7251 9027
rect 10042 9024 10048 9036
rect 7193 8987 7251 8993
rect 9784 8996 10048 9024
rect 6181 8959 6239 8965
rect 6181 8925 6193 8959
rect 6227 8925 6239 8959
rect 6181 8919 6239 8925
rect 6365 8959 6423 8965
rect 6365 8925 6377 8959
rect 6411 8925 6423 8959
rect 6365 8919 6423 8925
rect 6196 8888 6224 8919
rect 6454 8916 6460 8968
rect 6512 8916 6518 8968
rect 6641 8959 6699 8965
rect 6641 8925 6653 8959
rect 6687 8956 6699 8959
rect 7377 8959 7435 8965
rect 7377 8956 7389 8959
rect 6687 8928 7389 8956
rect 6687 8925 6699 8928
rect 6641 8919 6699 8925
rect 7377 8925 7389 8928
rect 7423 8956 7435 8959
rect 9398 8956 9404 8968
rect 7423 8928 9404 8956
rect 7423 8925 7435 8928
rect 7377 8919 7435 8925
rect 9398 8916 9404 8928
rect 9456 8916 9462 8968
rect 9784 8965 9812 8996
rect 10042 8984 10048 8996
rect 10100 8984 10106 9036
rect 9585 8959 9643 8965
rect 9585 8925 9597 8959
rect 9631 8925 9643 8959
rect 9585 8919 9643 8925
rect 9769 8959 9827 8965
rect 9769 8925 9781 8959
rect 9815 8925 9827 8959
rect 9769 8919 9827 8925
rect 6917 8891 6975 8897
rect 6917 8888 6929 8891
rect 6196 8860 6929 8888
rect 6917 8857 6929 8860
rect 6963 8857 6975 8891
rect 6917 8851 6975 8857
rect 5077 8823 5135 8829
rect 5077 8789 5089 8823
rect 5123 8820 5135 8823
rect 5258 8820 5264 8832
rect 5123 8792 5264 8820
rect 5123 8789 5135 8792
rect 5077 8783 5135 8789
rect 5258 8780 5264 8792
rect 5316 8780 5322 8832
rect 6273 8823 6331 8829
rect 6273 8789 6285 8823
rect 6319 8820 6331 8823
rect 6362 8820 6368 8832
rect 6319 8792 6368 8820
rect 6319 8789 6331 8792
rect 6273 8783 6331 8789
rect 6362 8780 6368 8792
rect 6420 8780 6426 8832
rect 6932 8820 6960 8851
rect 7006 8848 7012 8900
rect 7064 8888 7070 8900
rect 7101 8891 7159 8897
rect 7101 8888 7113 8891
rect 7064 8860 7113 8888
rect 7064 8848 7070 8860
rect 7101 8857 7113 8860
rect 7147 8857 7159 8891
rect 7101 8851 7159 8857
rect 8294 8848 8300 8900
rect 8352 8888 8358 8900
rect 9600 8888 9628 8919
rect 9858 8916 9864 8968
rect 9916 8916 9922 8968
rect 9950 8916 9956 8968
rect 10008 8916 10014 8968
rect 10152 8956 10180 9055
rect 15562 9052 15568 9064
rect 15620 9052 15626 9104
rect 20272 9101 20300 9132
rect 20625 9129 20637 9163
rect 20671 9160 20683 9163
rect 20898 9160 20904 9172
rect 20671 9132 20904 9160
rect 20671 9129 20683 9132
rect 20625 9123 20683 9129
rect 20898 9120 20904 9132
rect 20956 9120 20962 9172
rect 26421 9163 26479 9169
rect 26421 9129 26433 9163
rect 26467 9160 26479 9163
rect 26694 9160 26700 9172
rect 26467 9132 26700 9160
rect 26467 9129 26479 9132
rect 26421 9123 26479 9129
rect 26694 9120 26700 9132
rect 26752 9120 26758 9172
rect 26878 9120 26884 9172
rect 26936 9120 26942 9172
rect 20257 9095 20315 9101
rect 20257 9061 20269 9095
rect 20303 9061 20315 9095
rect 20257 9055 20315 9061
rect 24397 9095 24455 9101
rect 24397 9061 24409 9095
rect 24443 9092 24455 9095
rect 25314 9092 25320 9104
rect 24443 9064 25320 9092
rect 24443 9061 24455 9064
rect 24397 9055 24455 9061
rect 25314 9052 25320 9064
rect 25372 9052 25378 9104
rect 26234 9052 26240 9104
rect 26292 9092 26298 9104
rect 27062 9092 27068 9104
rect 26292 9064 27068 9092
rect 26292 9052 26298 9064
rect 27062 9052 27068 9064
rect 27120 9092 27126 9104
rect 28166 9092 28172 9104
rect 27120 9064 28172 9092
rect 27120 9052 27126 9064
rect 28166 9052 28172 9064
rect 28224 9052 28230 9104
rect 10226 8984 10232 9036
rect 10284 9024 10290 9036
rect 10284 8996 10548 9024
rect 10284 8984 10290 8996
rect 10520 8965 10548 8996
rect 12342 8984 12348 9036
rect 12400 8984 12406 9036
rect 15105 9027 15163 9033
rect 15105 8993 15117 9027
rect 15151 9024 15163 9027
rect 15930 9024 15936 9036
rect 15151 8996 15936 9024
rect 15151 8993 15163 8996
rect 15105 8987 15163 8993
rect 15930 8984 15936 8996
rect 15988 8984 15994 9036
rect 17037 9027 17095 9033
rect 17037 8993 17049 9027
rect 17083 9024 17095 9027
rect 17218 9024 17224 9036
rect 17083 8996 17224 9024
rect 17083 8993 17095 8996
rect 17037 8987 17095 8993
rect 17218 8984 17224 8996
rect 17276 9024 17282 9036
rect 17770 9024 17776 9036
rect 17276 8996 17776 9024
rect 17276 8984 17282 8996
rect 17770 8984 17776 8996
rect 17828 8984 17834 9036
rect 18874 8984 18880 9036
rect 18932 9024 18938 9036
rect 19797 9027 19855 9033
rect 19797 9024 19809 9027
rect 18932 8996 19809 9024
rect 18932 8984 18938 8996
rect 19797 8993 19809 8996
rect 19843 9024 19855 9027
rect 20714 9024 20720 9036
rect 19843 8996 20720 9024
rect 19843 8993 19855 8996
rect 19797 8987 19855 8993
rect 20714 8984 20720 8996
rect 20772 8984 20778 9036
rect 20901 9027 20959 9033
rect 20901 8993 20913 9027
rect 20947 9024 20959 9027
rect 21174 9024 21180 9036
rect 20947 8996 21180 9024
rect 20947 8993 20959 8996
rect 20901 8987 20959 8993
rect 21174 8984 21180 8996
rect 21232 8984 21238 9036
rect 22646 8984 22652 9036
rect 22704 9024 22710 9036
rect 23385 9027 23443 9033
rect 23385 9024 23397 9027
rect 22704 8996 23397 9024
rect 22704 8984 22710 8996
rect 23385 8993 23397 8996
rect 23431 8993 23443 9027
rect 23385 8987 23443 8993
rect 24026 8984 24032 9036
rect 24084 9024 24090 9036
rect 25593 9027 25651 9033
rect 25593 9024 25605 9027
rect 24084 8996 25605 9024
rect 24084 8984 24090 8996
rect 25593 8993 25605 8996
rect 25639 8993 25651 9027
rect 25593 8987 25651 8993
rect 25866 8984 25872 9036
rect 25924 8984 25930 9036
rect 25961 9027 26019 9033
rect 25961 8993 25973 9027
rect 26007 9024 26019 9027
rect 26786 9024 26792 9036
rect 26007 8996 26556 9024
rect 26007 8993 26019 8996
rect 25961 8987 26019 8993
rect 10413 8959 10471 8965
rect 10413 8956 10425 8959
rect 10152 8928 10425 8956
rect 10413 8925 10425 8928
rect 10459 8925 10471 8959
rect 10413 8919 10471 8925
rect 10505 8959 10563 8965
rect 10505 8925 10517 8959
rect 10551 8925 10563 8959
rect 10505 8919 10563 8925
rect 10781 8959 10839 8965
rect 10781 8925 10793 8959
rect 10827 8956 10839 8959
rect 10873 8959 10931 8965
rect 10873 8956 10885 8959
rect 10827 8928 10885 8956
rect 10827 8925 10839 8928
rect 10781 8919 10839 8925
rect 10873 8925 10885 8928
rect 10919 8925 10931 8959
rect 10873 8919 10931 8925
rect 10962 8916 10968 8968
rect 11020 8956 11026 8968
rect 11425 8959 11483 8965
rect 11425 8956 11437 8959
rect 11020 8928 11437 8956
rect 11020 8916 11026 8928
rect 11425 8925 11437 8928
rect 11471 8925 11483 8959
rect 11425 8919 11483 8925
rect 11882 8916 11888 8968
rect 11940 8956 11946 8968
rect 12069 8959 12127 8965
rect 12069 8956 12081 8959
rect 11940 8928 12081 8956
rect 11940 8916 11946 8928
rect 12069 8925 12081 8928
rect 12115 8925 12127 8959
rect 12069 8919 12127 8925
rect 14826 8916 14832 8968
rect 14884 8916 14890 8968
rect 15010 8916 15016 8968
rect 15068 8916 15074 8968
rect 15197 8959 15255 8965
rect 15197 8925 15209 8959
rect 15243 8925 15255 8959
rect 15197 8919 15255 8925
rect 15381 8959 15439 8965
rect 15381 8925 15393 8959
rect 15427 8956 15439 8959
rect 15562 8956 15568 8968
rect 15427 8928 15568 8956
rect 15427 8925 15439 8928
rect 15381 8919 15439 8925
rect 9674 8888 9680 8900
rect 8352 8860 9680 8888
rect 8352 8848 8358 8860
rect 9674 8848 9680 8860
rect 9732 8848 9738 8900
rect 10594 8848 10600 8900
rect 10652 8848 10658 8900
rect 12802 8848 12808 8900
rect 12860 8848 12866 8900
rect 15212 8888 15240 8919
rect 15562 8916 15568 8928
rect 15620 8916 15626 8968
rect 16850 8916 16856 8968
rect 16908 8916 16914 8968
rect 19981 8959 20039 8965
rect 19981 8925 19993 8959
rect 20027 8956 20039 8959
rect 20070 8956 20076 8968
rect 20027 8928 20076 8956
rect 20027 8925 20039 8928
rect 19981 8919 20039 8925
rect 20070 8916 20076 8928
rect 20128 8956 20134 8968
rect 20346 8956 20352 8968
rect 20128 8928 20352 8956
rect 20128 8916 20134 8928
rect 20346 8916 20352 8928
rect 20404 8956 20410 8968
rect 20530 8956 20536 8968
rect 20404 8928 20536 8956
rect 20404 8916 20410 8928
rect 20530 8916 20536 8928
rect 20588 8916 20594 8968
rect 22278 8916 22284 8968
rect 22336 8916 22342 8968
rect 24213 8959 24271 8965
rect 24213 8925 24225 8959
rect 24259 8956 24271 8959
rect 24302 8956 24308 8968
rect 24259 8928 24308 8956
rect 24259 8925 24271 8928
rect 24213 8919 24271 8925
rect 24302 8916 24308 8928
rect 24360 8956 24366 8968
rect 24670 8956 24676 8968
rect 24360 8928 24676 8956
rect 24360 8916 24366 8928
rect 24670 8916 24676 8928
rect 24728 8916 24734 8968
rect 25038 8916 25044 8968
rect 25096 8916 25102 8968
rect 25777 8959 25835 8965
rect 25777 8925 25789 8959
rect 25823 8925 25835 8959
rect 25777 8919 25835 8925
rect 15286 8888 15292 8900
rect 15212 8860 15292 8888
rect 15286 8848 15292 8860
rect 15344 8888 15350 8900
rect 16482 8888 16488 8900
rect 15344 8860 16488 8888
rect 15344 8848 15350 8860
rect 16482 8848 16488 8860
rect 16540 8848 16546 8900
rect 21082 8848 21088 8900
rect 21140 8888 21146 8900
rect 21177 8891 21235 8897
rect 21177 8888 21189 8891
rect 21140 8860 21189 8888
rect 21140 8848 21146 8860
rect 21177 8857 21189 8860
rect 21223 8857 21235 8891
rect 21177 8851 21235 8857
rect 24121 8891 24179 8897
rect 24121 8857 24133 8891
rect 24167 8888 24179 8891
rect 24486 8888 24492 8900
rect 24167 8860 24492 8888
rect 24167 8857 24179 8860
rect 24121 8851 24179 8857
rect 24486 8848 24492 8860
rect 24544 8888 24550 8900
rect 24765 8891 24823 8897
rect 24765 8888 24777 8891
rect 24544 8860 24777 8888
rect 24544 8848 24550 8860
rect 24765 8857 24777 8860
rect 24811 8857 24823 8891
rect 24765 8851 24823 8857
rect 24949 8891 25007 8897
rect 24949 8857 24961 8891
rect 24995 8888 25007 8891
rect 25133 8891 25191 8897
rect 25133 8888 25145 8891
rect 24995 8860 25145 8888
rect 24995 8857 25007 8860
rect 24949 8851 25007 8857
rect 25133 8857 25145 8860
rect 25179 8888 25191 8891
rect 25222 8888 25228 8900
rect 25179 8860 25228 8888
rect 25179 8857 25191 8860
rect 25133 8851 25191 8857
rect 25222 8848 25228 8860
rect 25280 8848 25286 8900
rect 25792 8888 25820 8919
rect 26050 8916 26056 8968
rect 26108 8916 26114 8968
rect 26237 8959 26295 8965
rect 26237 8925 26249 8959
rect 26283 8956 26295 8959
rect 26326 8956 26332 8968
rect 26283 8928 26332 8956
rect 26283 8925 26295 8928
rect 26237 8919 26295 8925
rect 26252 8888 26280 8919
rect 26326 8916 26332 8928
rect 26384 8916 26390 8968
rect 25792 8860 26280 8888
rect 26528 8888 26556 8996
rect 26620 8996 26792 9024
rect 26620 8965 26648 8996
rect 26786 8984 26792 8996
rect 26844 8984 26850 9036
rect 26878 8984 26884 9036
rect 26936 9024 26942 9036
rect 26936 8996 27384 9024
rect 26936 8984 26942 8996
rect 26605 8959 26663 8965
rect 26605 8925 26617 8959
rect 26651 8925 26663 8959
rect 26605 8919 26663 8925
rect 26697 8959 26755 8965
rect 26697 8925 26709 8959
rect 26743 8956 26755 8959
rect 26970 8956 26976 8968
rect 26743 8928 26976 8956
rect 26743 8925 26755 8928
rect 26697 8919 26755 8925
rect 26970 8916 26976 8928
rect 27028 8916 27034 8968
rect 27062 8916 27068 8968
rect 27120 8916 27126 8968
rect 27356 8965 27384 8996
rect 27341 8959 27399 8965
rect 27341 8925 27353 8959
rect 27387 8925 27399 8959
rect 27341 8919 27399 8925
rect 27430 8916 27436 8968
rect 27488 8956 27494 8968
rect 27525 8959 27583 8965
rect 27525 8956 27537 8959
rect 27488 8928 27537 8956
rect 27488 8916 27494 8928
rect 27525 8925 27537 8928
rect 27571 8925 27583 8959
rect 27525 8919 27583 8925
rect 27249 8891 27307 8897
rect 27249 8888 27261 8891
rect 26528 8860 27261 8888
rect 27249 8857 27261 8860
rect 27295 8888 27307 8891
rect 28074 8888 28080 8900
rect 27295 8860 28080 8888
rect 27295 8857 27307 8860
rect 27249 8851 27307 8857
rect 28074 8848 28080 8860
rect 28132 8848 28138 8900
rect 7190 8820 7196 8832
rect 6932 8792 7196 8820
rect 7190 8780 7196 8792
rect 7248 8820 7254 8832
rect 7561 8823 7619 8829
rect 7561 8820 7573 8823
rect 7248 8792 7573 8820
rect 7248 8780 7254 8792
rect 7561 8789 7573 8792
rect 7607 8789 7619 8823
rect 7561 8783 7619 8789
rect 9306 8780 9312 8832
rect 9364 8820 9370 8832
rect 10229 8823 10287 8829
rect 10229 8820 10241 8823
rect 9364 8792 10241 8820
rect 9364 8780 9370 8792
rect 10229 8789 10241 8792
rect 10275 8789 10287 8823
rect 10229 8783 10287 8789
rect 13817 8823 13875 8829
rect 13817 8789 13829 8823
rect 13863 8820 13875 8823
rect 14090 8820 14096 8832
rect 13863 8792 14096 8820
rect 13863 8789 13875 8792
rect 13817 8783 13875 8789
rect 14090 8780 14096 8792
rect 14148 8820 14154 8832
rect 15102 8820 15108 8832
rect 14148 8792 15108 8820
rect 14148 8780 14154 8792
rect 15102 8780 15108 8792
rect 15160 8780 15166 8832
rect 15194 8780 15200 8832
rect 15252 8780 15258 8832
rect 15470 8780 15476 8832
rect 15528 8820 15534 8832
rect 19886 8820 19892 8832
rect 15528 8792 19892 8820
rect 15528 8780 15534 8792
rect 19886 8780 19892 8792
rect 19944 8820 19950 8832
rect 20625 8823 20683 8829
rect 20625 8820 20637 8823
rect 19944 8792 20637 8820
rect 19944 8780 19950 8792
rect 20625 8789 20637 8792
rect 20671 8789 20683 8823
rect 20625 8783 20683 8789
rect 20806 8780 20812 8832
rect 20864 8780 20870 8832
rect 22738 8780 22744 8832
rect 22796 8820 22802 8832
rect 22833 8823 22891 8829
rect 22833 8820 22845 8823
rect 22796 8792 22845 8820
rect 22796 8780 22802 8792
rect 22833 8789 22845 8792
rect 22879 8789 22891 8823
rect 22833 8783 22891 8789
rect 24578 8780 24584 8832
rect 24636 8780 24642 8832
rect 24670 8780 24676 8832
rect 24728 8780 24734 8832
rect 26602 8780 26608 8832
rect 26660 8820 26666 8832
rect 27709 8823 27767 8829
rect 27709 8820 27721 8823
rect 26660 8792 27721 8820
rect 26660 8780 26666 8792
rect 27709 8789 27721 8792
rect 27755 8789 27767 8823
rect 27709 8783 27767 8789
rect 1104 8730 28704 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 28704 8730
rect 1104 8656 28704 8678
rect 4801 8619 4859 8625
rect 4801 8585 4813 8619
rect 4847 8585 4859 8619
rect 4801 8579 4859 8585
rect 3234 8548 3240 8560
rect 3068 8520 3240 8548
rect 3068 8489 3096 8520
rect 3234 8508 3240 8520
rect 3292 8508 3298 8560
rect 4614 8548 4620 8560
rect 4554 8520 4620 8548
rect 4614 8508 4620 8520
rect 4672 8508 4678 8560
rect 4816 8548 4844 8579
rect 5258 8576 5264 8628
rect 5316 8576 5322 8628
rect 6733 8619 6791 8625
rect 6733 8585 6745 8619
rect 6779 8616 6791 8619
rect 7006 8616 7012 8628
rect 6779 8588 7012 8616
rect 6779 8585 6791 8588
rect 6733 8579 6791 8585
rect 7006 8576 7012 8588
rect 7064 8616 7070 8628
rect 7374 8616 7380 8628
rect 7064 8588 7380 8616
rect 7064 8576 7070 8588
rect 7374 8576 7380 8588
rect 7432 8576 7438 8628
rect 8386 8576 8392 8628
rect 8444 8616 8450 8628
rect 10686 8616 10692 8628
rect 8444 8588 10692 8616
rect 8444 8576 8450 8588
rect 10686 8576 10692 8588
rect 10744 8576 10750 8628
rect 10781 8619 10839 8625
rect 10781 8585 10793 8619
rect 10827 8616 10839 8619
rect 10962 8616 10968 8628
rect 10827 8588 10968 8616
rect 10827 8585 10839 8588
rect 10781 8579 10839 8585
rect 10962 8576 10968 8588
rect 11020 8576 11026 8628
rect 14550 8616 14556 8628
rect 12728 8588 14556 8616
rect 5626 8548 5632 8560
rect 4816 8520 5632 8548
rect 5626 8508 5632 8520
rect 5684 8548 5690 8560
rect 6454 8548 6460 8560
rect 5684 8520 6460 8548
rect 5684 8508 5690 8520
rect 6454 8508 6460 8520
rect 6512 8508 6518 8560
rect 9306 8508 9312 8560
rect 9364 8508 9370 8560
rect 10318 8508 10324 8560
rect 10376 8508 10382 8560
rect 12728 8557 12756 8588
rect 14550 8576 14556 8588
rect 14608 8576 14614 8628
rect 14737 8619 14795 8625
rect 14737 8585 14749 8619
rect 14783 8616 14795 8619
rect 15010 8616 15016 8628
rect 14783 8588 15016 8616
rect 14783 8585 14795 8588
rect 14737 8579 14795 8585
rect 15010 8576 15016 8588
rect 15068 8576 15074 8628
rect 15562 8616 15568 8628
rect 15120 8588 15568 8616
rect 12713 8551 12771 8557
rect 12713 8517 12725 8551
rect 12759 8517 12771 8551
rect 12713 8511 12771 8517
rect 12802 8508 12808 8560
rect 12860 8548 12866 8560
rect 12860 8520 13202 8548
rect 12860 8508 12866 8520
rect 14182 8508 14188 8560
rect 14240 8548 14246 8560
rect 15120 8557 15148 8588
rect 15562 8576 15568 8588
rect 15620 8576 15626 8628
rect 20530 8576 20536 8628
rect 20588 8576 20594 8628
rect 21082 8576 21088 8628
rect 21140 8625 21146 8628
rect 21140 8616 21149 8625
rect 21140 8588 21185 8616
rect 21140 8579 21149 8588
rect 21140 8576 21146 8579
rect 21818 8576 21824 8628
rect 21876 8616 21882 8628
rect 21913 8619 21971 8625
rect 21913 8616 21925 8619
rect 21876 8588 21925 8616
rect 21876 8576 21882 8588
rect 21913 8585 21925 8588
rect 21959 8585 21971 8619
rect 22738 8616 22744 8628
rect 21913 8579 21971 8585
rect 22066 8588 22744 8616
rect 14461 8551 14519 8557
rect 14461 8548 14473 8551
rect 14240 8520 14473 8548
rect 14240 8508 14246 8520
rect 14461 8517 14473 8520
rect 14507 8548 14519 8551
rect 15105 8551 15163 8557
rect 14507 8520 15056 8548
rect 14507 8517 14519 8520
rect 14461 8511 14519 8517
rect 3053 8483 3111 8489
rect 3053 8449 3065 8483
rect 3099 8449 3111 8483
rect 3053 8443 3111 8449
rect 6546 8440 6552 8492
rect 6604 8440 6610 8492
rect 6822 8440 6828 8492
rect 6880 8440 6886 8492
rect 6914 8440 6920 8492
rect 6972 8440 6978 8492
rect 7006 8440 7012 8492
rect 7064 8440 7070 8492
rect 7101 8483 7159 8489
rect 7101 8449 7113 8483
rect 7147 8470 7159 8483
rect 7147 8449 7236 8470
rect 7101 8443 7236 8449
rect 7116 8442 7236 8443
rect 3329 8415 3387 8421
rect 3329 8381 3341 8415
rect 3375 8412 3387 8415
rect 3375 8384 4936 8412
rect 3375 8381 3387 8384
rect 3329 8375 3387 8381
rect 4908 8353 4936 8384
rect 5350 8372 5356 8424
rect 5408 8372 5414 8424
rect 5442 8372 5448 8424
rect 5500 8372 5506 8424
rect 5902 8372 5908 8424
rect 5960 8412 5966 8424
rect 6365 8415 6423 8421
rect 6365 8412 6377 8415
rect 5960 8384 6377 8412
rect 5960 8372 5966 8384
rect 6365 8381 6377 8384
rect 6411 8381 6423 8415
rect 7208 8412 7236 8442
rect 7282 8440 7288 8492
rect 7340 8440 7346 8492
rect 8294 8440 8300 8492
rect 8352 8440 8358 8492
rect 14277 8483 14335 8489
rect 14277 8480 14289 8483
rect 13924 8452 14289 8480
rect 6365 8375 6423 8381
rect 7116 8384 7236 8412
rect 4893 8347 4951 8353
rect 4893 8313 4905 8347
rect 4939 8313 4951 8347
rect 6380 8344 6408 8375
rect 7116 8344 7144 8384
rect 8312 8344 8340 8440
rect 8754 8372 8760 8424
rect 8812 8412 8818 8424
rect 9033 8415 9091 8421
rect 9033 8412 9045 8415
rect 8812 8384 9045 8412
rect 8812 8372 8818 8384
rect 9033 8381 9045 8384
rect 9079 8381 9091 8415
rect 9033 8375 9091 8381
rect 9398 8372 9404 8424
rect 9456 8412 9462 8424
rect 9456 8384 11836 8412
rect 9456 8372 9462 8384
rect 6380 8316 7144 8344
rect 7208 8316 8340 8344
rect 11808 8344 11836 8384
rect 11882 8372 11888 8424
rect 11940 8412 11946 8424
rect 12437 8415 12495 8421
rect 12437 8412 12449 8415
rect 11940 8384 12449 8412
rect 11940 8372 11946 8384
rect 12437 8381 12449 8384
rect 12483 8381 12495 8415
rect 13924 8412 13952 8452
rect 14277 8449 14289 8452
rect 14323 8480 14335 8483
rect 14918 8480 14924 8492
rect 14323 8452 14924 8480
rect 14323 8449 14335 8452
rect 14277 8443 14335 8449
rect 14918 8440 14924 8452
rect 14976 8440 14982 8492
rect 15028 8489 15056 8520
rect 15105 8517 15117 8551
rect 15151 8517 15163 8551
rect 15105 8511 15163 8517
rect 15304 8520 15700 8548
rect 15304 8492 15332 8520
rect 15013 8483 15071 8489
rect 15013 8449 15025 8483
rect 15059 8449 15071 8483
rect 15013 8443 15071 8449
rect 15286 8440 15292 8492
rect 15344 8440 15350 8492
rect 15381 8483 15439 8489
rect 15381 8449 15393 8483
rect 15427 8449 15439 8483
rect 15381 8443 15439 8449
rect 12437 8375 12495 8381
rect 12544 8384 13952 8412
rect 12544 8344 12572 8384
rect 14182 8372 14188 8424
rect 14240 8372 14246 8424
rect 15396 8412 15424 8443
rect 15562 8440 15568 8492
rect 15620 8440 15626 8492
rect 15672 8489 15700 8520
rect 16390 8508 16396 8560
rect 16448 8548 16454 8560
rect 16945 8551 17003 8557
rect 16945 8548 16957 8551
rect 16448 8520 16957 8548
rect 16448 8508 16454 8520
rect 16945 8517 16957 8520
rect 16991 8517 17003 8551
rect 16945 8511 17003 8517
rect 17037 8551 17095 8557
rect 17037 8517 17049 8551
rect 17083 8548 17095 8551
rect 17402 8548 17408 8560
rect 17083 8520 17408 8548
rect 17083 8517 17095 8520
rect 17037 8511 17095 8517
rect 17402 8508 17408 8520
rect 17460 8508 17466 8560
rect 19702 8508 19708 8560
rect 19760 8508 19766 8560
rect 20162 8508 20168 8560
rect 20220 8508 20226 8560
rect 20346 8508 20352 8560
rect 20404 8557 20410 8560
rect 20404 8551 20423 8557
rect 20411 8517 20423 8551
rect 20404 8511 20423 8517
rect 20625 8551 20683 8557
rect 20625 8517 20637 8551
rect 20671 8548 20683 8551
rect 20993 8551 21051 8557
rect 20993 8548 21005 8551
rect 20671 8520 21005 8548
rect 20671 8517 20683 8520
rect 20625 8511 20683 8517
rect 20993 8517 21005 8520
rect 21039 8517 21051 8551
rect 20993 8511 21051 8517
rect 21177 8551 21235 8557
rect 21177 8517 21189 8551
rect 21223 8548 21235 8551
rect 22066 8548 22094 8588
rect 22738 8576 22744 8588
rect 22796 8576 22802 8628
rect 23937 8619 23995 8625
rect 23937 8585 23949 8619
rect 23983 8616 23995 8619
rect 24118 8616 24124 8628
rect 23983 8588 24124 8616
rect 23983 8585 23995 8588
rect 23937 8579 23995 8585
rect 24118 8576 24124 8588
rect 24176 8616 24182 8628
rect 24578 8616 24584 8628
rect 24176 8588 24584 8616
rect 24176 8576 24182 8588
rect 24578 8576 24584 8588
rect 24636 8576 24642 8628
rect 24670 8548 24676 8560
rect 21223 8520 22094 8548
rect 23952 8520 24164 8548
rect 21223 8517 21235 8520
rect 21177 8511 21235 8517
rect 20404 8508 20410 8511
rect 15657 8483 15715 8489
rect 15657 8449 15669 8483
rect 15703 8449 15715 8483
rect 15657 8443 15715 8449
rect 15933 8483 15991 8489
rect 15933 8449 15945 8483
rect 15979 8480 15991 8483
rect 16408 8480 16436 8508
rect 23952 8492 23980 8520
rect 16853 8483 16911 8489
rect 16853 8480 16865 8483
rect 15979 8452 16436 8480
rect 16500 8452 16865 8480
rect 15979 8449 15991 8452
rect 15933 8443 15991 8449
rect 14936 8384 15424 8412
rect 11808 8316 12572 8344
rect 4893 8307 4951 8313
rect 5718 8236 5724 8288
rect 5776 8276 5782 8288
rect 7208 8276 7236 8316
rect 14936 8288 14964 8384
rect 15746 8372 15752 8424
rect 15804 8412 15810 8424
rect 16500 8412 16528 8452
rect 16853 8449 16865 8452
rect 16899 8449 16911 8483
rect 16853 8443 16911 8449
rect 17218 8440 17224 8492
rect 17276 8440 17282 8492
rect 17494 8440 17500 8492
rect 17552 8440 17558 8492
rect 17586 8440 17592 8492
rect 17644 8440 17650 8492
rect 17678 8440 17684 8492
rect 17736 8440 17742 8492
rect 17862 8440 17868 8492
rect 17920 8440 17926 8492
rect 20070 8440 20076 8492
rect 20128 8440 20134 8492
rect 20530 8440 20536 8492
rect 20588 8480 20594 8492
rect 20901 8483 20959 8489
rect 20901 8480 20913 8483
rect 20588 8452 20913 8480
rect 20588 8440 20594 8452
rect 20901 8449 20913 8452
rect 20947 8449 20959 8483
rect 21269 8483 21327 8489
rect 21269 8480 21281 8483
rect 20901 8443 20959 8449
rect 21008 8452 21281 8480
rect 15804 8384 16528 8412
rect 15804 8372 15810 8384
rect 16758 8372 16764 8424
rect 16816 8412 16822 8424
rect 17604 8412 17632 8440
rect 16816 8384 17632 8412
rect 16816 8372 16822 8384
rect 19426 8372 19432 8424
rect 19484 8412 19490 8424
rect 20162 8412 20168 8424
rect 19484 8384 20168 8412
rect 19484 8372 19490 8384
rect 20162 8372 20168 8384
rect 20220 8372 20226 8424
rect 20254 8372 20260 8424
rect 20312 8412 20318 8424
rect 20625 8415 20683 8421
rect 20625 8412 20637 8415
rect 20312 8384 20637 8412
rect 20312 8372 20318 8384
rect 20625 8381 20637 8384
rect 20671 8381 20683 8415
rect 21008 8412 21036 8452
rect 21269 8449 21281 8452
rect 21315 8449 21327 8483
rect 21269 8443 21327 8449
rect 22278 8440 22284 8492
rect 22336 8440 22342 8492
rect 23845 8483 23903 8489
rect 23845 8449 23857 8483
rect 23891 8480 23903 8483
rect 23934 8480 23940 8492
rect 23891 8452 23940 8480
rect 23891 8449 23903 8452
rect 23845 8443 23903 8449
rect 23934 8440 23940 8452
rect 23992 8440 23998 8492
rect 24136 8489 24164 8520
rect 24412 8520 24676 8548
rect 24029 8483 24087 8489
rect 24029 8449 24041 8483
rect 24075 8449 24087 8483
rect 24029 8443 24087 8449
rect 24121 8483 24179 8489
rect 24121 8449 24133 8483
rect 24167 8449 24179 8483
rect 24121 8443 24179 8449
rect 20625 8375 20683 8381
rect 20824 8384 21036 8412
rect 19794 8304 19800 8356
rect 19852 8344 19858 8356
rect 20824 8353 20852 8384
rect 21082 8372 21088 8424
rect 21140 8412 21146 8424
rect 23385 8415 23443 8421
rect 23385 8412 23397 8415
rect 21140 8384 23397 8412
rect 21140 8372 21146 8384
rect 23385 8381 23397 8384
rect 23431 8381 23443 8415
rect 23385 8375 23443 8381
rect 23658 8372 23664 8424
rect 23716 8372 23722 8424
rect 20809 8347 20867 8353
rect 20809 8344 20821 8347
rect 19852 8316 20821 8344
rect 19852 8304 19858 8316
rect 20809 8313 20821 8316
rect 20855 8313 20867 8347
rect 24044 8344 24072 8443
rect 24210 8372 24216 8424
rect 24268 8412 24274 8424
rect 24412 8421 24440 8520
rect 24670 8508 24676 8520
rect 24728 8508 24734 8560
rect 25038 8508 25044 8560
rect 25096 8508 25102 8560
rect 25332 8520 26004 8548
rect 24581 8483 24639 8489
rect 24581 8449 24593 8483
rect 24627 8480 24639 8483
rect 25056 8480 25084 8508
rect 25332 8492 25360 8520
rect 24627 8452 25084 8480
rect 24627 8449 24639 8452
rect 24581 8443 24639 8449
rect 25222 8440 25228 8492
rect 25280 8440 25286 8492
rect 25314 8440 25320 8492
rect 25372 8440 25378 8492
rect 25682 8440 25688 8492
rect 25740 8440 25746 8492
rect 25976 8489 26004 8520
rect 25777 8483 25835 8489
rect 25777 8449 25789 8483
rect 25823 8449 25835 8483
rect 25777 8443 25835 8449
rect 25961 8483 26019 8489
rect 25961 8449 25973 8483
rect 26007 8449 26019 8483
rect 25961 8443 26019 8449
rect 24397 8415 24455 8421
rect 24397 8412 24409 8415
rect 24268 8384 24409 8412
rect 24268 8372 24274 8384
rect 24397 8381 24409 8384
rect 24443 8381 24455 8415
rect 24397 8375 24455 8381
rect 24762 8372 24768 8424
rect 24820 8412 24826 8424
rect 24857 8415 24915 8421
rect 24857 8412 24869 8415
rect 24820 8384 24869 8412
rect 24820 8372 24826 8384
rect 24857 8381 24869 8384
rect 24903 8381 24915 8415
rect 24857 8375 24915 8381
rect 25038 8372 25044 8424
rect 25096 8372 25102 8424
rect 25133 8415 25191 8421
rect 25133 8381 25145 8415
rect 25179 8412 25191 8415
rect 25406 8412 25412 8424
rect 25179 8384 25412 8412
rect 25179 8381 25191 8384
rect 25133 8375 25191 8381
rect 25406 8372 25412 8384
rect 25464 8372 25470 8424
rect 25792 8412 25820 8443
rect 26050 8440 26056 8492
rect 26108 8440 26114 8492
rect 26326 8412 26332 8424
rect 25792 8384 26332 8412
rect 26326 8372 26332 8384
rect 26384 8372 26390 8424
rect 24670 8344 24676 8356
rect 24044 8316 24676 8344
rect 20809 8307 20867 8313
rect 24670 8304 24676 8316
rect 24728 8304 24734 8356
rect 24946 8304 24952 8356
rect 25004 8344 25010 8356
rect 25501 8347 25559 8353
rect 25501 8344 25513 8347
rect 25004 8316 25513 8344
rect 25004 8304 25010 8316
rect 25501 8313 25513 8316
rect 25547 8313 25559 8347
rect 25501 8307 25559 8313
rect 5776 8248 7236 8276
rect 5776 8236 5782 8248
rect 7282 8236 7288 8288
rect 7340 8236 7346 8288
rect 9490 8236 9496 8288
rect 9548 8276 9554 8288
rect 9858 8276 9864 8288
rect 9548 8248 9864 8276
rect 9548 8236 9554 8248
rect 9858 8236 9864 8248
rect 9916 8236 9922 8288
rect 14645 8279 14703 8285
rect 14645 8245 14657 8279
rect 14691 8276 14703 8279
rect 14918 8276 14924 8288
rect 14691 8248 14924 8276
rect 14691 8245 14703 8248
rect 14645 8239 14703 8245
rect 14918 8236 14924 8248
rect 14976 8236 14982 8288
rect 16114 8236 16120 8288
rect 16172 8236 16178 8288
rect 16666 8236 16672 8288
rect 16724 8236 16730 8288
rect 17310 8236 17316 8288
rect 17368 8236 17374 8288
rect 19518 8236 19524 8288
rect 19576 8236 19582 8288
rect 19705 8279 19763 8285
rect 19705 8245 19717 8279
rect 19751 8276 19763 8279
rect 19886 8276 19892 8288
rect 19751 8248 19892 8276
rect 19751 8245 19763 8248
rect 19705 8239 19763 8245
rect 19886 8236 19892 8248
rect 19944 8236 19950 8288
rect 20254 8236 20260 8288
rect 20312 8276 20318 8288
rect 20349 8279 20407 8285
rect 20349 8276 20361 8279
rect 20312 8248 20361 8276
rect 20312 8236 20318 8248
rect 20349 8245 20361 8248
rect 20395 8245 20407 8279
rect 20349 8239 20407 8245
rect 24302 8236 24308 8288
rect 24360 8236 24366 8288
rect 24394 8236 24400 8288
rect 24452 8276 24458 8288
rect 24765 8279 24823 8285
rect 24765 8276 24777 8279
rect 24452 8248 24777 8276
rect 24452 8236 24458 8248
rect 24765 8245 24777 8248
rect 24811 8245 24823 8279
rect 24765 8239 24823 8245
rect 1104 8186 28704 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 28704 8186
rect 1104 8112 28704 8134
rect 5169 8075 5227 8081
rect 5169 8041 5181 8075
rect 5215 8072 5227 8075
rect 5350 8072 5356 8084
rect 5215 8044 5356 8072
rect 5215 8041 5227 8044
rect 5169 8035 5227 8041
rect 5350 8032 5356 8044
rect 5408 8032 5414 8084
rect 7098 8032 7104 8084
rect 7156 8072 7162 8084
rect 7193 8075 7251 8081
rect 7193 8072 7205 8075
rect 7156 8044 7205 8072
rect 7156 8032 7162 8044
rect 7193 8041 7205 8044
rect 7239 8041 7251 8075
rect 9950 8072 9956 8084
rect 7193 8035 7251 8041
rect 9140 8044 9956 8072
rect 5718 8004 5724 8016
rect 4632 7976 5724 8004
rect 4632 7877 4660 7976
rect 5718 7964 5724 7976
rect 5776 7964 5782 8016
rect 5997 8007 6055 8013
rect 5997 7973 6009 8007
rect 6043 7973 6055 8007
rect 8386 8004 8392 8016
rect 5997 7967 6055 7973
rect 6840 7976 8392 8004
rect 6012 7936 6040 7967
rect 4816 7908 6040 7936
rect 4816 7877 4844 7908
rect 6454 7896 6460 7948
rect 6512 7896 6518 7948
rect 4617 7871 4675 7877
rect 4617 7837 4629 7871
rect 4663 7837 4675 7871
rect 4617 7831 4675 7837
rect 4801 7871 4859 7877
rect 4801 7837 4813 7871
rect 4847 7837 4859 7871
rect 4801 7831 4859 7837
rect 4985 7871 5043 7877
rect 4985 7837 4997 7871
rect 5031 7868 5043 7871
rect 5902 7868 5908 7880
rect 5031 7840 5908 7868
rect 5031 7837 5043 7840
rect 4985 7831 5043 7837
rect 5902 7828 5908 7840
rect 5960 7828 5966 7880
rect 6362 7828 6368 7880
rect 6420 7828 6426 7880
rect 6840 7877 6868 7976
rect 8386 7964 8392 7976
rect 8444 7964 8450 8016
rect 7190 7936 7196 7948
rect 7024 7908 7196 7936
rect 7024 7877 7052 7908
rect 7190 7896 7196 7908
rect 7248 7896 7254 7948
rect 9140 7945 9168 8044
rect 9950 8032 9956 8044
rect 10008 8032 10014 8084
rect 10045 8075 10103 8081
rect 10045 8041 10057 8075
rect 10091 8072 10103 8075
rect 10594 8072 10600 8084
rect 10091 8044 10600 8072
rect 10091 8041 10103 8044
rect 10045 8035 10103 8041
rect 10594 8032 10600 8044
rect 10652 8032 10658 8084
rect 14737 8075 14795 8081
rect 14737 8041 14749 8075
rect 14783 8072 14795 8075
rect 14826 8072 14832 8084
rect 14783 8044 14832 8072
rect 14783 8041 14795 8044
rect 14737 8035 14795 8041
rect 14826 8032 14832 8044
rect 14884 8032 14890 8084
rect 15930 8032 15936 8084
rect 15988 8032 15994 8084
rect 16301 8075 16359 8081
rect 16301 8041 16313 8075
rect 16347 8072 16359 8075
rect 16666 8072 16672 8084
rect 16347 8044 16672 8072
rect 16347 8041 16359 8044
rect 16301 8035 16359 8041
rect 16666 8032 16672 8044
rect 16724 8032 16730 8084
rect 19702 8032 19708 8084
rect 19760 8072 19766 8084
rect 19797 8075 19855 8081
rect 19797 8072 19809 8075
rect 19760 8044 19809 8072
rect 19760 8032 19766 8044
rect 19797 8041 19809 8044
rect 19843 8041 19855 8075
rect 19797 8035 19855 8041
rect 24302 8032 24308 8084
rect 24360 8072 24366 8084
rect 25041 8075 25099 8081
rect 25041 8072 25053 8075
rect 24360 8044 25053 8072
rect 24360 8032 24366 8044
rect 25041 8041 25053 8044
rect 25087 8072 25099 8075
rect 25406 8072 25412 8084
rect 25087 8044 25412 8072
rect 25087 8041 25099 8044
rect 25041 8035 25099 8041
rect 25406 8032 25412 8044
rect 25464 8032 25470 8084
rect 26145 8075 26203 8081
rect 26145 8041 26157 8075
rect 26191 8041 26203 8075
rect 26145 8035 26203 8041
rect 9646 7976 9809 8004
rect 9125 7939 9183 7945
rect 9125 7905 9137 7939
rect 9171 7905 9183 7939
rect 9646 7936 9674 7976
rect 9125 7899 9183 7905
rect 9324 7908 9674 7936
rect 9781 7936 9809 7976
rect 10134 7964 10140 8016
rect 10192 8004 10198 8016
rect 10873 8007 10931 8013
rect 10873 8004 10885 8007
rect 10192 7976 10885 8004
rect 10192 7964 10198 7976
rect 10873 7973 10885 7976
rect 10919 7973 10931 8007
rect 17494 8004 17500 8016
rect 10873 7967 10931 7973
rect 16960 7976 17500 8004
rect 9781 7908 10364 7936
rect 9324 7880 9352 7908
rect 6825 7871 6883 7877
rect 6825 7837 6837 7871
rect 6871 7837 6883 7871
rect 6825 7831 6883 7837
rect 7009 7871 7067 7877
rect 7009 7837 7021 7871
rect 7055 7837 7067 7871
rect 7009 7831 7067 7837
rect 7098 7828 7104 7880
rect 7156 7828 7162 7880
rect 7282 7828 7288 7880
rect 7340 7868 7346 7880
rect 7561 7871 7619 7877
rect 7561 7868 7573 7871
rect 7340 7840 7573 7868
rect 7340 7828 7346 7840
rect 7561 7837 7573 7840
rect 7607 7837 7619 7871
rect 7561 7831 7619 7837
rect 9306 7828 9312 7880
rect 9364 7828 9370 7880
rect 9582 7828 9588 7880
rect 9640 7828 9646 7880
rect 9858 7828 9864 7880
rect 9916 7828 9922 7880
rect 10336 7877 10364 7908
rect 10410 7896 10416 7948
rect 10468 7936 10474 7948
rect 11333 7939 11391 7945
rect 11333 7936 11345 7939
rect 10468 7908 11345 7936
rect 10468 7896 10474 7908
rect 11333 7905 11345 7908
rect 11379 7905 11391 7939
rect 11333 7899 11391 7905
rect 15197 7939 15255 7945
rect 15197 7905 15209 7939
rect 15243 7936 15255 7939
rect 15470 7936 15476 7948
rect 15243 7908 15476 7936
rect 15243 7905 15255 7908
rect 15197 7899 15255 7905
rect 15470 7896 15476 7908
rect 15528 7936 15534 7948
rect 15654 7936 15660 7948
rect 15528 7908 15660 7936
rect 15528 7896 15534 7908
rect 15654 7896 15660 7908
rect 15712 7896 15718 7948
rect 16960 7880 16988 7976
rect 17494 7964 17500 7976
rect 17552 7964 17558 8016
rect 24118 7964 24124 8016
rect 24176 7964 24182 8016
rect 24670 7964 24676 8016
rect 24728 8004 24734 8016
rect 25777 8007 25835 8013
rect 25777 8004 25789 8007
rect 24728 7976 25789 8004
rect 24728 7964 24734 7976
rect 25777 7973 25789 7976
rect 25823 7973 25835 8007
rect 26160 8004 26188 8035
rect 26326 8032 26332 8084
rect 26384 8032 26390 8084
rect 26510 8032 26516 8084
rect 26568 8072 26574 8084
rect 26878 8072 26884 8084
rect 26568 8044 26884 8072
rect 26568 8032 26574 8044
rect 26878 8032 26884 8044
rect 26936 8032 26942 8084
rect 26421 8007 26479 8013
rect 26421 8004 26433 8007
rect 26160 7976 26433 8004
rect 25777 7967 25835 7973
rect 26421 7973 26433 7976
rect 26467 8004 26479 8007
rect 26786 8004 26792 8016
rect 26467 7976 26792 8004
rect 26467 7973 26479 7976
rect 26421 7967 26479 7973
rect 26786 7964 26792 7976
rect 26844 7964 26850 8016
rect 17037 7939 17095 7945
rect 17037 7905 17049 7939
rect 17083 7936 17095 7939
rect 17218 7936 17224 7948
rect 17083 7908 17224 7936
rect 17083 7905 17095 7908
rect 17037 7899 17095 7905
rect 17218 7896 17224 7908
rect 17276 7896 17282 7948
rect 18414 7936 18420 7948
rect 18064 7908 18420 7936
rect 10321 7871 10379 7877
rect 10321 7837 10333 7871
rect 10367 7837 10379 7871
rect 10321 7831 10379 7837
rect 10597 7871 10655 7877
rect 10597 7837 10609 7871
rect 10643 7837 10655 7871
rect 10597 7831 10655 7837
rect 10781 7871 10839 7877
rect 10781 7837 10793 7871
rect 10827 7868 10839 7871
rect 10962 7868 10968 7880
rect 10827 7840 10968 7868
rect 10827 7837 10839 7840
rect 10781 7831 10839 7837
rect 4893 7803 4951 7809
rect 4893 7769 4905 7803
rect 4939 7800 4951 7803
rect 5534 7800 5540 7812
rect 4939 7772 5540 7800
rect 4939 7769 4951 7772
rect 4893 7763 4951 7769
rect 5534 7760 5540 7772
rect 5592 7800 5598 7812
rect 7190 7800 7196 7812
rect 5592 7772 7196 7800
rect 5592 7760 5598 7772
rect 7190 7760 7196 7772
rect 7248 7760 7254 7812
rect 7374 7760 7380 7812
rect 7432 7760 7438 7812
rect 10612 7800 10640 7831
rect 10962 7828 10968 7840
rect 11020 7868 11026 7880
rect 11149 7871 11207 7877
rect 11149 7868 11161 7871
rect 11020 7840 11161 7868
rect 11020 7828 11026 7840
rect 11149 7837 11161 7840
rect 11195 7868 11207 7871
rect 11241 7871 11299 7877
rect 11241 7868 11253 7871
rect 11195 7840 11253 7868
rect 11195 7837 11207 7840
rect 11149 7831 11207 7837
rect 11241 7837 11253 7840
rect 11287 7837 11299 7871
rect 11241 7831 11299 7837
rect 11425 7871 11483 7877
rect 11425 7837 11437 7871
rect 11471 7868 11483 7871
rect 12802 7868 12808 7880
rect 11471 7840 12808 7868
rect 11471 7837 11483 7840
rect 11425 7831 11483 7837
rect 9968 7772 10640 7800
rect 5261 7735 5319 7741
rect 5261 7701 5273 7735
rect 5307 7732 5319 7735
rect 5442 7732 5448 7744
rect 5307 7704 5448 7732
rect 5307 7701 5319 7704
rect 5261 7695 5319 7701
rect 5442 7692 5448 7704
rect 5500 7692 5506 7744
rect 6638 7692 6644 7744
rect 6696 7692 6702 7744
rect 9493 7735 9551 7741
rect 9493 7701 9505 7735
rect 9539 7732 9551 7735
rect 9582 7732 9588 7744
rect 9539 7704 9588 7732
rect 9539 7701 9551 7704
rect 9493 7695 9551 7701
rect 9582 7692 9588 7704
rect 9640 7692 9646 7744
rect 9674 7692 9680 7744
rect 9732 7692 9738 7744
rect 9766 7692 9772 7744
rect 9824 7732 9830 7744
rect 9968 7732 9996 7772
rect 9824 7704 9996 7732
rect 10137 7735 10195 7741
rect 9824 7692 9830 7704
rect 10137 7701 10149 7735
rect 10183 7732 10195 7735
rect 10502 7732 10508 7744
rect 10183 7704 10508 7732
rect 10183 7701 10195 7704
rect 10137 7695 10195 7701
rect 10502 7692 10508 7704
rect 10560 7692 10566 7744
rect 10612 7732 10640 7772
rect 10870 7760 10876 7812
rect 10928 7760 10934 7812
rect 11440 7800 11468 7831
rect 12802 7828 12808 7840
rect 12860 7828 12866 7880
rect 14918 7828 14924 7880
rect 14976 7828 14982 7880
rect 15013 7871 15071 7877
rect 15013 7837 15025 7871
rect 15059 7837 15071 7871
rect 15013 7831 15071 7837
rect 10980 7772 11468 7800
rect 15028 7800 15056 7831
rect 15102 7828 15108 7880
rect 15160 7868 15166 7880
rect 15289 7871 15347 7877
rect 15289 7868 15301 7871
rect 15160 7840 15301 7868
rect 15160 7828 15166 7840
rect 15289 7837 15301 7840
rect 15335 7837 15347 7871
rect 15289 7831 15347 7837
rect 16114 7828 16120 7880
rect 16172 7828 16178 7880
rect 16393 7871 16451 7877
rect 16393 7837 16405 7871
rect 16439 7868 16451 7871
rect 16577 7871 16635 7877
rect 16577 7868 16589 7871
rect 16439 7840 16589 7868
rect 16439 7837 16451 7840
rect 16393 7831 16451 7837
rect 16577 7837 16589 7840
rect 16623 7837 16635 7871
rect 16577 7831 16635 7837
rect 16758 7828 16764 7880
rect 16816 7828 16822 7880
rect 16942 7828 16948 7880
rect 17000 7828 17006 7880
rect 17129 7871 17187 7877
rect 17129 7837 17141 7871
rect 17175 7837 17187 7871
rect 17129 7831 17187 7837
rect 15194 7800 15200 7812
rect 15028 7772 15200 7800
rect 10980 7732 11008 7772
rect 15194 7760 15200 7772
rect 15252 7760 15258 7812
rect 10612 7704 11008 7732
rect 11057 7735 11115 7741
rect 11057 7701 11069 7735
rect 11103 7732 11115 7735
rect 11606 7732 11612 7744
rect 11103 7704 11612 7732
rect 11103 7701 11115 7704
rect 11057 7695 11115 7701
rect 11606 7692 11612 7704
rect 11664 7692 11670 7744
rect 17144 7732 17172 7831
rect 17310 7828 17316 7880
rect 17368 7828 17374 7880
rect 18064 7877 18092 7908
rect 18414 7896 18420 7908
rect 18472 7936 18478 7948
rect 20254 7936 20260 7948
rect 18472 7908 19104 7936
rect 18472 7896 18478 7908
rect 19076 7880 19104 7908
rect 19352 7908 20260 7936
rect 18049 7871 18107 7877
rect 18049 7837 18061 7871
rect 18095 7837 18107 7871
rect 18049 7831 18107 7837
rect 18322 7828 18328 7880
rect 18380 7868 18386 7880
rect 18509 7871 18567 7877
rect 18509 7868 18521 7871
rect 18380 7840 18521 7868
rect 18380 7828 18386 7840
rect 18509 7837 18521 7840
rect 18555 7837 18567 7871
rect 18509 7831 18567 7837
rect 18601 7871 18659 7877
rect 18601 7837 18613 7871
rect 18647 7868 18659 7871
rect 18782 7868 18788 7880
rect 18647 7840 18788 7868
rect 18647 7837 18659 7840
rect 18601 7831 18659 7837
rect 18782 7828 18788 7840
rect 18840 7828 18846 7880
rect 18874 7828 18880 7880
rect 18932 7828 18938 7880
rect 19058 7828 19064 7880
rect 19116 7868 19122 7880
rect 19352 7877 19380 7908
rect 20254 7896 20260 7908
rect 20312 7896 20318 7948
rect 24213 7939 24271 7945
rect 24213 7905 24225 7939
rect 24259 7936 24271 7939
rect 24578 7936 24584 7948
rect 24259 7908 24584 7936
rect 24259 7905 24271 7908
rect 24213 7899 24271 7905
rect 24578 7896 24584 7908
rect 24636 7896 24642 7948
rect 24854 7896 24860 7948
rect 24912 7936 24918 7948
rect 24912 7908 24957 7936
rect 24912 7896 24918 7908
rect 25222 7896 25228 7948
rect 25280 7896 25286 7948
rect 26053 7939 26111 7945
rect 26053 7905 26065 7939
rect 26099 7936 26111 7939
rect 26326 7936 26332 7948
rect 26099 7908 26332 7936
rect 26099 7905 26111 7908
rect 26053 7899 26111 7905
rect 26326 7896 26332 7908
rect 26384 7936 26390 7948
rect 26602 7936 26608 7948
rect 26384 7908 26608 7936
rect 26384 7896 26390 7908
rect 26602 7896 26608 7908
rect 26660 7896 26666 7948
rect 19337 7871 19395 7877
rect 19337 7868 19349 7871
rect 19116 7840 19349 7868
rect 19116 7828 19122 7840
rect 19337 7837 19349 7840
rect 19383 7837 19395 7871
rect 19337 7831 19395 7837
rect 19426 7828 19432 7880
rect 19484 7828 19490 7880
rect 19613 7871 19671 7877
rect 19613 7837 19625 7871
rect 19659 7868 19671 7871
rect 20346 7868 20352 7880
rect 19659 7840 20352 7868
rect 19659 7837 19671 7840
rect 19613 7831 19671 7837
rect 17770 7760 17776 7812
rect 17828 7800 17834 7812
rect 17865 7803 17923 7809
rect 17865 7800 17877 7803
rect 17828 7772 17877 7800
rect 17828 7760 17834 7772
rect 17865 7769 17877 7772
rect 17911 7769 17923 7803
rect 17865 7763 17923 7769
rect 18233 7803 18291 7809
rect 18233 7769 18245 7803
rect 18279 7800 18291 7803
rect 18693 7803 18751 7809
rect 18279 7772 18552 7800
rect 18279 7769 18291 7772
rect 18233 7763 18291 7769
rect 17402 7732 17408 7744
rect 17144 7704 17408 7732
rect 17402 7692 17408 7704
rect 17460 7692 17466 7744
rect 18322 7692 18328 7744
rect 18380 7692 18386 7744
rect 18524 7732 18552 7772
rect 18693 7769 18705 7803
rect 18739 7800 18751 7803
rect 18966 7800 18972 7812
rect 18739 7772 18972 7800
rect 18739 7769 18751 7772
rect 18693 7763 18751 7769
rect 18966 7760 18972 7772
rect 19024 7760 19030 7812
rect 19150 7760 19156 7812
rect 19208 7800 19214 7812
rect 19628 7800 19656 7831
rect 20346 7828 20352 7840
rect 20404 7868 20410 7880
rect 22094 7868 22100 7880
rect 20404 7840 22100 7868
rect 20404 7828 20410 7840
rect 22094 7828 22100 7840
rect 22152 7828 22158 7880
rect 23753 7871 23811 7877
rect 23753 7837 23765 7871
rect 23799 7868 23811 7871
rect 24302 7868 24308 7880
rect 23799 7840 24308 7868
rect 23799 7837 23811 7840
rect 23753 7831 23811 7837
rect 24302 7828 24308 7840
rect 24360 7828 24366 7880
rect 24486 7828 24492 7880
rect 24544 7868 24550 7880
rect 24673 7871 24731 7877
rect 24673 7868 24685 7871
rect 24544 7840 24685 7868
rect 24544 7828 24550 7840
rect 24673 7837 24685 7840
rect 24719 7837 24731 7871
rect 24673 7831 24731 7837
rect 24765 7871 24823 7877
rect 24765 7837 24777 7871
rect 24811 7868 24823 7871
rect 25130 7868 25136 7880
rect 24811 7864 24900 7868
rect 24964 7864 25136 7868
rect 24811 7840 25136 7864
rect 24811 7837 24823 7840
rect 24765 7831 24823 7837
rect 24872 7836 24992 7840
rect 25130 7828 25136 7840
rect 25188 7868 25194 7880
rect 25317 7871 25375 7877
rect 25317 7868 25329 7871
rect 25188 7840 25329 7868
rect 25188 7828 25194 7840
rect 25317 7837 25329 7840
rect 25363 7837 25375 7871
rect 25317 7831 25375 7837
rect 26145 7871 26203 7877
rect 26145 7837 26157 7871
rect 26191 7868 26203 7871
rect 26510 7868 26516 7880
rect 26191 7840 26516 7868
rect 26191 7837 26203 7840
rect 26145 7831 26203 7837
rect 26510 7828 26516 7840
rect 26568 7828 26574 7880
rect 28350 7828 28356 7880
rect 28408 7828 28414 7880
rect 19208 7772 19656 7800
rect 19208 7760 19214 7772
rect 23934 7760 23940 7812
rect 23992 7800 23998 7812
rect 25041 7803 25099 7809
rect 25041 7800 25053 7803
rect 23992 7772 25053 7800
rect 23992 7760 23998 7772
rect 25041 7769 25053 7772
rect 25087 7769 25099 7803
rect 25682 7800 25688 7812
rect 25041 7763 25099 7769
rect 25516 7772 25688 7800
rect 19242 7732 19248 7744
rect 18524 7704 19248 7732
rect 19242 7692 19248 7704
rect 19300 7692 19306 7744
rect 23842 7692 23848 7744
rect 23900 7732 23906 7744
rect 25516 7741 25544 7772
rect 25682 7760 25688 7772
rect 25740 7800 25746 7812
rect 26237 7803 26295 7809
rect 26237 7800 26249 7803
rect 25740 7772 26249 7800
rect 25740 7760 25746 7772
rect 26237 7769 26249 7772
rect 26283 7769 26295 7803
rect 26237 7763 26295 7769
rect 24397 7735 24455 7741
rect 24397 7732 24409 7735
rect 23900 7704 24409 7732
rect 23900 7692 23906 7704
rect 24397 7701 24409 7704
rect 24443 7701 24455 7735
rect 24397 7695 24455 7701
rect 25501 7735 25559 7741
rect 25501 7701 25513 7735
rect 25547 7701 25559 7735
rect 25501 7695 25559 7701
rect 27522 7692 27528 7744
rect 27580 7732 27586 7744
rect 28169 7735 28227 7741
rect 28169 7732 28181 7735
rect 27580 7704 28181 7732
rect 27580 7692 27586 7704
rect 28169 7701 28181 7704
rect 28215 7701 28227 7735
rect 28169 7695 28227 7701
rect 1104 7642 28704 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 28704 7642
rect 1104 7568 28704 7590
rect 4985 7531 5043 7537
rect 4985 7497 4997 7531
rect 5031 7497 5043 7531
rect 4985 7491 5043 7497
rect 5000 7460 5028 7491
rect 5442 7488 5448 7540
rect 5500 7488 5506 7540
rect 5537 7531 5595 7537
rect 5537 7497 5549 7531
rect 5583 7528 5595 7531
rect 6365 7531 6423 7537
rect 6365 7528 6377 7531
rect 5583 7500 6377 7528
rect 5583 7497 5595 7500
rect 5537 7491 5595 7497
rect 6365 7497 6377 7500
rect 6411 7497 6423 7531
rect 6365 7491 6423 7497
rect 6454 7488 6460 7540
rect 6512 7528 6518 7540
rect 7193 7531 7251 7537
rect 7193 7528 7205 7531
rect 6512 7500 7205 7528
rect 6512 7488 6518 7500
rect 7193 7497 7205 7500
rect 7239 7497 7251 7531
rect 7193 7491 7251 7497
rect 9306 7488 9312 7540
rect 9364 7528 9370 7540
rect 10597 7531 10655 7537
rect 10597 7528 10609 7531
rect 9364 7500 10609 7528
rect 9364 7488 9370 7500
rect 10597 7497 10609 7500
rect 10643 7497 10655 7531
rect 10597 7491 10655 7497
rect 11790 7488 11796 7540
rect 11848 7528 11854 7540
rect 17589 7531 17647 7537
rect 11848 7500 12388 7528
rect 11848 7488 11854 7500
rect 5902 7460 5908 7472
rect 5000 7432 5908 7460
rect 5902 7420 5908 7432
rect 5960 7420 5966 7472
rect 6914 7460 6920 7472
rect 6564 7432 6920 7460
rect 4614 7352 4620 7404
rect 4672 7392 4678 7404
rect 5258 7392 5264 7404
rect 4672 7364 5264 7392
rect 4672 7352 4678 7364
rect 5258 7352 5264 7364
rect 5316 7352 5322 7404
rect 6564 7401 6592 7432
rect 6914 7420 6920 7432
rect 6972 7460 6978 7472
rect 10410 7460 10416 7472
rect 6972 7432 7144 7460
rect 10258 7432 10416 7460
rect 6972 7420 6978 7432
rect 6549 7395 6607 7401
rect 6549 7361 6561 7395
rect 6595 7361 6607 7395
rect 6549 7355 6607 7361
rect 6638 7352 6644 7404
rect 6696 7352 6702 7404
rect 7116 7401 7144 7432
rect 10410 7420 10416 7432
rect 10468 7420 10474 7472
rect 11606 7420 11612 7472
rect 11664 7460 11670 7472
rect 12066 7460 12072 7472
rect 11664 7432 12072 7460
rect 11664 7420 11670 7432
rect 12066 7420 12072 7432
rect 12124 7469 12130 7472
rect 12360 7469 12388 7500
rect 17589 7497 17601 7531
rect 17635 7528 17647 7531
rect 17862 7528 17868 7540
rect 17635 7500 17868 7528
rect 17635 7497 17647 7500
rect 17589 7491 17647 7497
rect 17862 7488 17868 7500
rect 17920 7488 17926 7540
rect 18322 7488 18328 7540
rect 18380 7488 18386 7540
rect 19426 7528 19432 7540
rect 18800 7500 19432 7528
rect 12124 7463 12173 7469
rect 12124 7429 12127 7463
rect 12161 7429 12173 7463
rect 12124 7423 12173 7429
rect 12345 7463 12403 7469
rect 12345 7429 12357 7463
rect 12391 7429 12403 7463
rect 12345 7423 12403 7429
rect 12124 7420 12130 7423
rect 15010 7420 15016 7472
rect 15068 7460 15074 7472
rect 17126 7460 17132 7472
rect 15068 7432 17132 7460
rect 15068 7420 15074 7432
rect 17126 7420 17132 7432
rect 17184 7420 17190 7472
rect 18340 7460 18368 7488
rect 17788 7432 18368 7460
rect 7101 7395 7159 7401
rect 7101 7361 7113 7395
rect 7147 7361 7159 7395
rect 7101 7355 7159 7361
rect 7285 7395 7343 7401
rect 7285 7361 7297 7395
rect 7331 7392 7343 7395
rect 7374 7392 7380 7404
rect 7331 7364 7380 7392
rect 7331 7361 7343 7364
rect 7285 7355 7343 7361
rect 7374 7352 7380 7364
rect 7432 7352 7438 7404
rect 10962 7392 10968 7404
rect 10520 7364 10968 7392
rect 3234 7284 3240 7336
rect 3292 7284 3298 7336
rect 3513 7327 3571 7333
rect 3513 7293 3525 7327
rect 3559 7324 3571 7327
rect 3559 7296 5120 7324
rect 3559 7293 3571 7296
rect 3513 7287 3571 7293
rect 5092 7265 5120 7296
rect 5350 7284 5356 7336
rect 5408 7324 5414 7336
rect 5629 7327 5687 7333
rect 5629 7324 5641 7327
rect 5408 7296 5641 7324
rect 5408 7284 5414 7296
rect 5629 7293 5641 7296
rect 5675 7293 5687 7327
rect 5629 7287 5687 7293
rect 6454 7284 6460 7336
rect 6512 7324 6518 7336
rect 6917 7327 6975 7333
rect 6917 7324 6929 7327
rect 6512 7296 6929 7324
rect 6512 7284 6518 7296
rect 6917 7293 6929 7296
rect 6963 7293 6975 7327
rect 6917 7287 6975 7293
rect 7009 7327 7067 7333
rect 7009 7293 7021 7327
rect 7055 7324 7067 7327
rect 7190 7324 7196 7336
rect 7055 7296 7196 7324
rect 7055 7293 7067 7296
rect 7009 7287 7067 7293
rect 7190 7284 7196 7296
rect 7248 7324 7254 7336
rect 7248 7296 8248 7324
rect 7248 7284 7254 7296
rect 5077 7259 5135 7265
rect 5077 7225 5089 7259
rect 5123 7225 5135 7259
rect 5077 7219 5135 7225
rect 8220 7188 8248 7296
rect 8294 7284 8300 7336
rect 8352 7324 8358 7336
rect 8754 7324 8760 7336
rect 8352 7296 8760 7324
rect 8352 7284 8358 7296
rect 8754 7284 8760 7296
rect 8812 7284 8818 7336
rect 9030 7284 9036 7336
rect 9088 7284 9094 7336
rect 10520 7333 10548 7364
rect 10962 7352 10968 7364
rect 11020 7392 11026 7404
rect 11977 7395 12035 7401
rect 11977 7392 11989 7395
rect 11020 7364 11989 7392
rect 11020 7352 11026 7364
rect 11977 7361 11989 7364
rect 12023 7361 12035 7395
rect 11977 7355 12035 7361
rect 12253 7395 12311 7401
rect 12253 7361 12265 7395
rect 12299 7361 12311 7395
rect 12253 7355 12311 7361
rect 10505 7327 10563 7333
rect 10505 7293 10517 7327
rect 10551 7293 10563 7327
rect 10505 7287 10563 7293
rect 10873 7327 10931 7333
rect 10873 7293 10885 7327
rect 10919 7324 10931 7327
rect 11146 7324 11152 7336
rect 10919 7296 11152 7324
rect 10919 7293 10931 7296
rect 10873 7287 10931 7293
rect 11146 7284 11152 7296
rect 11204 7284 11210 7336
rect 12268 7324 12296 7355
rect 12434 7352 12440 7404
rect 12492 7352 12498 7404
rect 13081 7395 13139 7401
rect 13081 7361 13093 7395
rect 13127 7392 13139 7395
rect 13630 7392 13636 7404
rect 13127 7364 13636 7392
rect 13127 7361 13139 7364
rect 13081 7355 13139 7361
rect 13630 7352 13636 7364
rect 13688 7352 13694 7404
rect 17788 7401 17816 7432
rect 18414 7420 18420 7472
rect 18472 7420 18478 7472
rect 17773 7395 17831 7401
rect 17773 7361 17785 7395
rect 17819 7361 17831 7395
rect 17773 7355 17831 7361
rect 17954 7352 17960 7404
rect 18012 7352 18018 7404
rect 18046 7352 18052 7404
rect 18104 7352 18110 7404
rect 18279 7395 18337 7401
rect 18279 7392 18291 7395
rect 18156 7364 18291 7392
rect 12342 7324 12348 7336
rect 12268 7296 12348 7324
rect 12342 7284 12348 7296
rect 12400 7284 12406 7336
rect 12621 7327 12679 7333
rect 12621 7293 12633 7327
rect 12667 7324 12679 7327
rect 12710 7324 12716 7336
rect 12667 7296 12716 7324
rect 12667 7293 12679 7296
rect 12621 7287 12679 7293
rect 12710 7284 12716 7296
rect 12768 7284 12774 7336
rect 12986 7284 12992 7336
rect 13044 7284 13050 7336
rect 18156 7324 18184 7364
rect 18279 7361 18291 7364
rect 18325 7361 18337 7395
rect 18279 7355 18337 7361
rect 18506 7352 18512 7404
rect 18564 7352 18570 7404
rect 18690 7392 18696 7404
rect 18651 7364 18696 7392
rect 18690 7352 18696 7364
rect 18748 7352 18754 7404
rect 18800 7401 18828 7500
rect 19426 7488 19432 7500
rect 19484 7488 19490 7540
rect 21637 7531 21695 7537
rect 21637 7497 21649 7531
rect 21683 7528 21695 7531
rect 22094 7528 22100 7540
rect 21683 7500 22100 7528
rect 21683 7497 21695 7500
rect 21637 7491 21695 7497
rect 22094 7488 22100 7500
rect 22152 7488 22158 7540
rect 24302 7488 24308 7540
rect 24360 7528 24366 7540
rect 25222 7528 25228 7540
rect 24360 7500 25228 7528
rect 24360 7488 24366 7500
rect 25222 7488 25228 7500
rect 25280 7488 25286 7540
rect 26050 7528 26056 7540
rect 25608 7500 26056 7528
rect 19150 7420 19156 7472
rect 19208 7420 19214 7472
rect 19242 7420 19248 7472
rect 19300 7420 19306 7472
rect 19518 7420 19524 7472
rect 19576 7460 19582 7472
rect 20165 7463 20223 7469
rect 20165 7460 20177 7463
rect 19576 7432 20177 7460
rect 19576 7420 19582 7432
rect 20165 7429 20177 7432
rect 20211 7429 20223 7463
rect 21450 7460 21456 7472
rect 21390 7432 21456 7460
rect 20165 7423 20223 7429
rect 21450 7420 21456 7432
rect 21508 7420 21514 7472
rect 24670 7460 24676 7472
rect 24228 7432 24676 7460
rect 24228 7401 24256 7432
rect 24670 7420 24676 7432
rect 24728 7420 24734 7472
rect 18785 7395 18843 7401
rect 18785 7361 18797 7395
rect 18831 7361 18843 7395
rect 18785 7355 18843 7361
rect 19061 7395 19119 7401
rect 19061 7361 19073 7395
rect 19107 7361 19119 7395
rect 19061 7355 19119 7361
rect 19429 7395 19487 7401
rect 19429 7361 19441 7395
rect 19475 7361 19487 7395
rect 19429 7355 19487 7361
rect 24213 7395 24271 7401
rect 24213 7361 24225 7395
rect 24259 7361 24271 7395
rect 24213 7355 24271 7361
rect 17788 7296 18184 7324
rect 17788 7268 17816 7296
rect 18598 7284 18604 7336
rect 18656 7324 18662 7336
rect 19076 7324 19104 7355
rect 18656 7296 19104 7324
rect 18656 7284 18662 7296
rect 17770 7216 17776 7268
rect 17828 7216 17834 7268
rect 17954 7216 17960 7268
rect 18012 7256 18018 7268
rect 18877 7259 18935 7265
rect 18877 7256 18889 7259
rect 18012 7228 18889 7256
rect 18012 7216 18018 7228
rect 18877 7225 18889 7228
rect 18923 7225 18935 7259
rect 18877 7219 18935 7225
rect 9490 7188 9496 7200
rect 8220 7160 9496 7188
rect 9490 7148 9496 7160
rect 9548 7148 9554 7200
rect 9582 7148 9588 7200
rect 9640 7188 9646 7200
rect 10686 7188 10692 7200
rect 9640 7160 10692 7188
rect 9640 7148 9646 7160
rect 10686 7148 10692 7160
rect 10744 7148 10750 7200
rect 12526 7148 12532 7200
rect 12584 7188 12590 7200
rect 12713 7191 12771 7197
rect 12713 7188 12725 7191
rect 12584 7160 12725 7188
rect 12584 7148 12590 7160
rect 12713 7157 12725 7160
rect 12759 7157 12771 7191
rect 12713 7151 12771 7157
rect 18141 7191 18199 7197
rect 18141 7157 18153 7191
rect 18187 7188 18199 7191
rect 19444 7188 19472 7355
rect 24394 7352 24400 7404
rect 24452 7352 24458 7404
rect 25608 7392 25636 7500
rect 26050 7488 26056 7500
rect 26108 7528 26114 7540
rect 26513 7531 26571 7537
rect 26513 7528 26525 7531
rect 26108 7500 26525 7528
rect 26108 7488 26114 7500
rect 26513 7497 26525 7500
rect 26559 7497 26571 7531
rect 26513 7491 26571 7497
rect 25682 7420 25688 7472
rect 25740 7460 25746 7472
rect 25740 7432 26188 7460
rect 25740 7420 25746 7432
rect 26160 7401 26188 7432
rect 24688 7364 25636 7392
rect 25869 7395 25927 7401
rect 24688 7333 24716 7364
rect 25869 7361 25881 7395
rect 25915 7392 25927 7395
rect 26145 7395 26203 7401
rect 25915 7364 26004 7392
rect 25915 7361 25927 7364
rect 25869 7355 25927 7361
rect 19889 7327 19947 7333
rect 19889 7293 19901 7327
rect 19935 7324 19947 7327
rect 24673 7327 24731 7333
rect 19935 7296 20024 7324
rect 19935 7293 19947 7296
rect 19889 7287 19947 7293
rect 18187 7160 19472 7188
rect 19996 7188 20024 7296
rect 24673 7293 24685 7327
rect 24719 7293 24731 7327
rect 24673 7287 24731 7293
rect 25976 7256 26004 7364
rect 26145 7361 26157 7395
rect 26191 7361 26203 7395
rect 26145 7355 26203 7361
rect 26326 7352 26332 7404
rect 26384 7352 26390 7404
rect 26418 7352 26424 7404
rect 26476 7352 26482 7404
rect 26605 7395 26663 7401
rect 26605 7361 26617 7395
rect 26651 7361 26663 7395
rect 26605 7355 26663 7361
rect 26053 7327 26111 7333
rect 26053 7293 26065 7327
rect 26099 7324 26111 7327
rect 26234 7324 26240 7336
rect 26099 7296 26240 7324
rect 26099 7293 26111 7296
rect 26053 7287 26111 7293
rect 26234 7284 26240 7296
rect 26292 7324 26298 7336
rect 26620 7324 26648 7355
rect 28350 7352 28356 7404
rect 28408 7352 28414 7404
rect 26292 7296 26648 7324
rect 26292 7284 26298 7296
rect 26326 7256 26332 7268
rect 25976 7228 26332 7256
rect 26326 7216 26332 7228
rect 26384 7216 26390 7268
rect 21174 7188 21180 7200
rect 19996 7160 21180 7188
rect 18187 7157 18199 7160
rect 18141 7151 18199 7157
rect 21174 7148 21180 7160
rect 21232 7148 21238 7200
rect 24394 7148 24400 7200
rect 24452 7148 24458 7200
rect 25498 7148 25504 7200
rect 25556 7188 25562 7200
rect 26145 7191 26203 7197
rect 26145 7188 26157 7191
rect 25556 7160 26157 7188
rect 25556 7148 25562 7160
rect 26145 7157 26157 7160
rect 26191 7157 26203 7191
rect 26145 7151 26203 7157
rect 27890 7148 27896 7200
rect 27948 7188 27954 7200
rect 28169 7191 28227 7197
rect 28169 7188 28181 7191
rect 27948 7160 28181 7188
rect 27948 7148 27954 7160
rect 28169 7157 28181 7160
rect 28215 7157 28227 7191
rect 28169 7151 28227 7157
rect 1104 7098 28704 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 28704 7098
rect 1104 7024 28704 7046
rect 9030 6944 9036 6996
rect 9088 6984 9094 6996
rect 9585 6987 9643 6993
rect 9585 6984 9597 6987
rect 9088 6956 9597 6984
rect 9088 6944 9094 6956
rect 9585 6953 9597 6956
rect 9631 6953 9643 6987
rect 9585 6947 9643 6953
rect 10502 6944 10508 6996
rect 10560 6984 10566 6996
rect 11425 6987 11483 6993
rect 11425 6984 11437 6987
rect 10560 6956 11437 6984
rect 10560 6944 10566 6956
rect 11425 6953 11437 6956
rect 11471 6984 11483 6987
rect 11974 6984 11980 6996
rect 11471 6956 11980 6984
rect 11471 6953 11483 6956
rect 11425 6947 11483 6953
rect 11974 6944 11980 6956
rect 12032 6944 12038 6996
rect 12158 6993 12164 6996
rect 12148 6987 12164 6993
rect 12148 6953 12160 6987
rect 12148 6947 12164 6953
rect 12158 6944 12164 6947
rect 12216 6944 12222 6996
rect 12342 6944 12348 6996
rect 12400 6984 12406 6996
rect 14277 6987 14335 6993
rect 14277 6984 14289 6987
rect 12400 6956 14289 6984
rect 12400 6944 12406 6956
rect 14277 6953 14289 6956
rect 14323 6953 14335 6987
rect 14277 6947 14335 6953
rect 18046 6944 18052 6996
rect 18104 6984 18110 6996
rect 18417 6987 18475 6993
rect 18417 6984 18429 6987
rect 18104 6956 18429 6984
rect 18104 6944 18110 6956
rect 18417 6953 18429 6956
rect 18463 6953 18475 6987
rect 18417 6947 18475 6953
rect 18877 6987 18935 6993
rect 18877 6953 18889 6987
rect 18923 6984 18935 6987
rect 19058 6984 19064 6996
rect 18923 6956 19064 6984
rect 18923 6953 18935 6956
rect 18877 6947 18935 6953
rect 11333 6919 11391 6925
rect 11333 6885 11345 6919
rect 11379 6916 11391 6919
rect 11514 6916 11520 6928
rect 11379 6888 11520 6916
rect 11379 6885 11391 6888
rect 11333 6879 11391 6885
rect 11514 6876 11520 6888
rect 11572 6876 11578 6928
rect 18322 6876 18328 6928
rect 18380 6916 18386 6928
rect 18892 6916 18920 6947
rect 19058 6944 19064 6956
rect 19116 6944 19122 6996
rect 27522 6944 27528 6996
rect 27580 6984 27586 6996
rect 27997 6987 28055 6993
rect 27997 6984 28009 6987
rect 27580 6956 28009 6984
rect 27580 6944 27586 6956
rect 27997 6953 28009 6956
rect 28043 6953 28055 6987
rect 27997 6947 28055 6953
rect 18380 6888 18920 6916
rect 18380 6876 18386 6888
rect 10137 6851 10195 6857
rect 10137 6817 10149 6851
rect 10183 6848 10195 6851
rect 10962 6848 10968 6860
rect 10183 6820 10968 6848
rect 10183 6817 10195 6820
rect 10137 6811 10195 6817
rect 10962 6808 10968 6820
rect 11020 6808 11026 6860
rect 12526 6848 12532 6860
rect 11440 6820 12532 6848
rect 9766 6783 9824 6789
rect 9766 6749 9778 6783
rect 9812 6780 9824 6783
rect 10042 6780 10048 6792
rect 9812 6752 10048 6780
rect 9812 6749 9824 6752
rect 9766 6743 9824 6749
rect 10042 6740 10048 6752
rect 10100 6740 10106 6792
rect 10226 6740 10232 6792
rect 10284 6740 10290 6792
rect 10597 6783 10655 6789
rect 10597 6749 10609 6783
rect 10643 6749 10655 6783
rect 10597 6743 10655 6749
rect 10612 6712 10640 6743
rect 10686 6740 10692 6792
rect 10744 6740 10750 6792
rect 11146 6740 11152 6792
rect 11204 6740 11210 6792
rect 11440 6789 11468 6820
rect 12526 6808 12532 6820
rect 12584 6808 12590 6860
rect 17678 6808 17684 6860
rect 17736 6848 17742 6860
rect 17865 6851 17923 6857
rect 17865 6848 17877 6851
rect 17736 6820 17877 6848
rect 17736 6808 17742 6820
rect 17865 6817 17877 6820
rect 17911 6817 17923 6851
rect 18782 6848 18788 6860
rect 17865 6811 17923 6817
rect 18064 6820 18788 6848
rect 11425 6783 11483 6789
rect 11425 6749 11437 6783
rect 11471 6749 11483 6783
rect 11425 6743 11483 6749
rect 11514 6740 11520 6792
rect 11572 6740 11578 6792
rect 11882 6740 11888 6792
rect 11940 6740 11946 6792
rect 18064 6789 18092 6820
rect 18782 6808 18788 6820
rect 18840 6808 18846 6860
rect 14093 6783 14151 6789
rect 14093 6749 14105 6783
rect 14139 6749 14151 6783
rect 14093 6743 14151 6749
rect 18049 6783 18107 6789
rect 18049 6749 18061 6783
rect 18095 6749 18107 6783
rect 18598 6780 18604 6792
rect 18049 6743 18107 6749
rect 18156 6752 18604 6780
rect 10778 6712 10784 6724
rect 10612 6684 10784 6712
rect 10778 6672 10784 6684
rect 10836 6672 10842 6724
rect 11624 6684 12572 6712
rect 9769 6647 9827 6653
rect 9769 6613 9781 6647
rect 9815 6644 9827 6647
rect 10321 6647 10379 6653
rect 10321 6644 10333 6647
rect 9815 6616 10333 6644
rect 9815 6613 9827 6616
rect 9769 6607 9827 6613
rect 10321 6613 10333 6616
rect 10367 6613 10379 6647
rect 10321 6607 10379 6613
rect 11238 6604 11244 6656
rect 11296 6644 11302 6656
rect 11624 6644 11652 6684
rect 11296 6616 11652 6644
rect 11793 6647 11851 6653
rect 11296 6604 11302 6616
rect 11793 6613 11805 6647
rect 11839 6644 11851 6647
rect 12434 6644 12440 6656
rect 11839 6616 12440 6644
rect 11839 6613 11851 6616
rect 11793 6607 11851 6613
rect 12434 6604 12440 6616
rect 12492 6604 12498 6656
rect 12544 6644 12572 6684
rect 12618 6672 12624 6724
rect 12676 6672 12682 6724
rect 14108 6712 14136 6743
rect 13464 6684 14136 6712
rect 13464 6644 13492 6684
rect 17218 6672 17224 6724
rect 17276 6712 17282 6724
rect 18156 6712 18184 6752
rect 18598 6740 18604 6752
rect 18656 6740 18662 6792
rect 18693 6783 18751 6789
rect 18693 6749 18705 6783
rect 18739 6749 18751 6783
rect 18693 6743 18751 6749
rect 17276 6684 18184 6712
rect 17276 6672 17282 6684
rect 18230 6672 18236 6724
rect 18288 6672 18294 6724
rect 18708 6712 18736 6743
rect 18874 6740 18880 6792
rect 18932 6780 18938 6792
rect 18969 6783 19027 6789
rect 18969 6780 18981 6783
rect 18932 6752 18981 6780
rect 18932 6740 18938 6752
rect 18969 6749 18981 6752
rect 19015 6749 19027 6783
rect 18969 6743 19027 6749
rect 28258 6740 28264 6792
rect 28316 6740 28322 6792
rect 19150 6712 19156 6724
rect 18708 6684 19156 6712
rect 19150 6672 19156 6684
rect 19208 6672 19214 6724
rect 23566 6672 23572 6724
rect 23624 6712 23630 6724
rect 23845 6715 23903 6721
rect 23845 6712 23857 6715
rect 23624 6684 23857 6712
rect 23624 6672 23630 6684
rect 23845 6681 23857 6684
rect 23891 6681 23903 6715
rect 23845 6675 23903 6681
rect 24210 6672 24216 6724
rect 24268 6712 24274 6724
rect 26694 6712 26700 6724
rect 24268 6684 26700 6712
rect 24268 6672 24274 6684
rect 26694 6672 26700 6684
rect 26752 6672 26758 6724
rect 27246 6672 27252 6724
rect 27304 6672 27310 6724
rect 12544 6616 13492 6644
rect 13630 6604 13636 6656
rect 13688 6604 13694 6656
rect 19794 6604 19800 6656
rect 19852 6644 19858 6656
rect 23937 6647 23995 6653
rect 23937 6644 23949 6647
rect 19852 6616 23949 6644
rect 19852 6604 19858 6616
rect 23937 6613 23949 6616
rect 23983 6644 23995 6647
rect 24118 6644 24124 6656
rect 23983 6616 24124 6644
rect 23983 6613 23995 6616
rect 23937 6607 23995 6613
rect 24118 6604 24124 6616
rect 24176 6604 24182 6656
rect 26513 6647 26571 6653
rect 26513 6613 26525 6647
rect 26559 6644 26571 6647
rect 26602 6644 26608 6656
rect 26559 6616 26608 6644
rect 26559 6613 26571 6616
rect 26513 6607 26571 6613
rect 26602 6604 26608 6616
rect 26660 6604 26666 6656
rect 1104 6554 28704 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 28704 6554
rect 1104 6480 28704 6502
rect 12158 6400 12164 6452
rect 12216 6440 12222 6452
rect 12253 6443 12311 6449
rect 12253 6440 12265 6443
rect 12216 6412 12265 6440
rect 12216 6400 12222 6412
rect 12253 6409 12265 6412
rect 12299 6409 12311 6443
rect 12253 6403 12311 6409
rect 12710 6400 12716 6452
rect 12768 6400 12774 6452
rect 12802 6400 12808 6452
rect 12860 6440 12866 6452
rect 17957 6443 18015 6449
rect 17957 6440 17969 6443
rect 12860 6412 17969 6440
rect 12860 6400 12866 6412
rect 17957 6409 17969 6412
rect 18003 6409 18015 6443
rect 17957 6403 18015 6409
rect 22278 6400 22284 6452
rect 22336 6400 22342 6452
rect 23566 6400 23572 6452
rect 23624 6400 23630 6452
rect 24854 6400 24860 6452
rect 24912 6400 24918 6452
rect 27154 6400 27160 6452
rect 27212 6400 27218 6452
rect 13446 6332 13452 6384
rect 13504 6332 13510 6384
rect 14918 6332 14924 6384
rect 14976 6372 14982 6384
rect 15289 6375 15347 6381
rect 15289 6372 15301 6375
rect 14976 6344 15301 6372
rect 14976 6332 14982 6344
rect 15289 6341 15301 6344
rect 15335 6372 15347 6375
rect 16574 6372 16580 6384
rect 15335 6344 16580 6372
rect 15335 6341 15347 6344
rect 15289 6335 15347 6341
rect 16574 6332 16580 6344
rect 16632 6372 16638 6384
rect 16853 6375 16911 6381
rect 16853 6372 16865 6375
rect 16632 6344 16865 6372
rect 16632 6332 16638 6344
rect 16853 6341 16865 6344
rect 16899 6372 16911 6375
rect 17129 6375 17187 6381
rect 17129 6372 17141 6375
rect 16899 6344 17141 6372
rect 16899 6341 16911 6344
rect 16853 6335 16911 6341
rect 17129 6341 17141 6344
rect 17175 6341 17187 6375
rect 17129 6335 17187 6341
rect 17313 6375 17371 6381
rect 17313 6341 17325 6375
rect 17359 6372 17371 6375
rect 20438 6372 20444 6384
rect 17359 6344 20444 6372
rect 17359 6341 17371 6344
rect 17313 6335 17371 6341
rect 20438 6332 20444 6344
rect 20496 6332 20502 6384
rect 22296 6372 22324 6400
rect 22554 6372 22560 6384
rect 22296 6344 22560 6372
rect 22554 6332 22560 6344
rect 22612 6332 22618 6384
rect 24320 6344 24808 6372
rect 11514 6264 11520 6316
rect 11572 6304 11578 6316
rect 11885 6307 11943 6313
rect 11885 6304 11897 6307
rect 11572 6276 11897 6304
rect 11572 6264 11578 6276
rect 11885 6273 11897 6276
rect 11931 6273 11943 6307
rect 11885 6267 11943 6273
rect 11974 6264 11980 6316
rect 12032 6264 12038 6316
rect 12621 6307 12679 6313
rect 12621 6273 12633 6307
rect 12667 6304 12679 6307
rect 12710 6304 12716 6316
rect 12667 6276 12716 6304
rect 12667 6273 12679 6276
rect 12621 6267 12679 6273
rect 12710 6264 12716 6276
rect 12768 6304 12774 6316
rect 13630 6304 13636 6316
rect 12768 6276 13636 6304
rect 12768 6264 12774 6276
rect 13630 6264 13636 6276
rect 13688 6264 13694 6316
rect 13906 6264 13912 6316
rect 13964 6304 13970 6316
rect 14734 6304 14740 6316
rect 13964 6276 14740 6304
rect 13964 6264 13970 6276
rect 14734 6264 14740 6276
rect 14792 6304 14798 6316
rect 15930 6304 15936 6316
rect 14792 6276 15936 6304
rect 14792 6264 14798 6276
rect 15930 6264 15936 6276
rect 15988 6264 15994 6316
rect 16025 6307 16083 6313
rect 16025 6273 16037 6307
rect 16071 6273 16083 6307
rect 16025 6267 16083 6273
rect 16117 6307 16175 6313
rect 16117 6273 16129 6307
rect 16163 6273 16175 6307
rect 16117 6267 16175 6273
rect 12161 6239 12219 6245
rect 12161 6205 12173 6239
rect 12207 6236 12219 6239
rect 12526 6236 12532 6248
rect 12207 6208 12532 6236
rect 12207 6205 12219 6208
rect 12161 6199 12219 6205
rect 12526 6196 12532 6208
rect 12584 6196 12590 6248
rect 12897 6239 12955 6245
rect 12897 6205 12909 6239
rect 12943 6236 12955 6239
rect 12943 6208 13124 6236
rect 12943 6205 12955 6208
rect 12897 6199 12955 6205
rect 11790 6128 11796 6180
rect 11848 6168 11854 6180
rect 12069 6171 12127 6177
rect 12069 6168 12081 6171
rect 11848 6140 12081 6168
rect 11848 6128 11854 6140
rect 12069 6137 12081 6140
rect 12115 6137 12127 6171
rect 12069 6131 12127 6137
rect 13096 6112 13124 6208
rect 15378 6196 15384 6248
rect 15436 6236 15442 6248
rect 15436 6208 15884 6236
rect 15436 6196 15442 6208
rect 15194 6128 15200 6180
rect 15252 6168 15258 6180
rect 15856 6177 15884 6208
rect 16040 6180 16068 6267
rect 16132 6236 16160 6267
rect 16206 6264 16212 6316
rect 16264 6264 16270 6316
rect 16390 6264 16396 6316
rect 16448 6264 16454 6316
rect 17037 6307 17095 6313
rect 17037 6273 17049 6307
rect 17083 6273 17095 6307
rect 17037 6267 17095 6273
rect 18141 6307 18199 6313
rect 18141 6273 18153 6307
rect 18187 6273 18199 6307
rect 18141 6267 18199 6273
rect 18325 6307 18383 6313
rect 18325 6273 18337 6307
rect 18371 6304 18383 6307
rect 18506 6304 18512 6316
rect 18371 6276 18512 6304
rect 18371 6273 18383 6276
rect 18325 6267 18383 6273
rect 16850 6236 16856 6248
rect 16132 6208 16856 6236
rect 16850 6196 16856 6208
rect 16908 6236 16914 6248
rect 17052 6236 17080 6267
rect 16908 6208 17080 6236
rect 18156 6236 18184 6267
rect 18506 6264 18512 6276
rect 18564 6264 18570 6316
rect 23842 6264 23848 6316
rect 23900 6264 23906 6316
rect 24026 6264 24032 6316
rect 24084 6264 24090 6316
rect 24118 6264 24124 6316
rect 24176 6264 24182 6316
rect 24320 6313 24348 6344
rect 24305 6307 24363 6313
rect 24305 6273 24317 6307
rect 24351 6273 24363 6307
rect 24305 6267 24363 6273
rect 24578 6264 24584 6316
rect 24636 6264 24642 6316
rect 24780 6313 24808 6344
rect 24765 6307 24823 6313
rect 24765 6273 24777 6307
rect 24811 6304 24823 6307
rect 25038 6304 25044 6316
rect 24811 6276 25044 6304
rect 24811 6273 24823 6276
rect 24765 6267 24823 6273
rect 25038 6264 25044 6276
rect 25096 6304 25102 6316
rect 26145 6307 26203 6313
rect 25096 6276 26004 6304
rect 25096 6264 25102 6276
rect 18690 6236 18696 6248
rect 18156 6208 18696 6236
rect 16908 6196 16914 6208
rect 18690 6196 18696 6208
rect 18748 6236 18754 6248
rect 19058 6236 19064 6248
rect 18748 6208 19064 6236
rect 18748 6196 18754 6208
rect 19058 6196 19064 6208
rect 19116 6196 19122 6248
rect 21174 6196 21180 6248
rect 21232 6236 21238 6248
rect 21821 6239 21879 6245
rect 21821 6236 21833 6239
rect 21232 6208 21833 6236
rect 21232 6196 21238 6208
rect 21821 6205 21833 6208
rect 21867 6205 21879 6239
rect 21821 6199 21879 6205
rect 22097 6239 22155 6245
rect 22097 6205 22109 6239
rect 22143 6236 22155 6239
rect 23661 6239 23719 6245
rect 23661 6236 23673 6239
rect 22143 6208 23673 6236
rect 22143 6205 22155 6208
rect 22097 6199 22155 6205
rect 23661 6205 23673 6208
rect 23707 6205 23719 6239
rect 23661 6199 23719 6205
rect 15565 6171 15623 6177
rect 15565 6168 15577 6171
rect 15252 6140 15577 6168
rect 15252 6128 15258 6140
rect 15565 6137 15577 6140
rect 15611 6137 15623 6171
rect 15565 6131 15623 6137
rect 15841 6171 15899 6177
rect 15841 6137 15853 6171
rect 15887 6137 15899 6171
rect 15841 6131 15899 6137
rect 16022 6128 16028 6180
rect 16080 6128 16086 6180
rect 16666 6128 16672 6180
rect 16724 6168 16730 6180
rect 17310 6168 17316 6180
rect 16724 6140 17316 6168
rect 16724 6128 16730 6140
rect 17310 6128 17316 6140
rect 17368 6128 17374 6180
rect 23474 6128 23480 6180
rect 23532 6168 23538 6180
rect 23937 6171 23995 6177
rect 23937 6168 23949 6171
rect 23532 6140 23949 6168
rect 23532 6128 23538 6140
rect 23937 6137 23949 6140
rect 23983 6168 23995 6171
rect 24762 6168 24768 6180
rect 23983 6140 24768 6168
rect 23983 6137 23995 6140
rect 23937 6131 23995 6137
rect 24762 6128 24768 6140
rect 24820 6128 24826 6180
rect 25976 6177 26004 6276
rect 26145 6273 26157 6307
rect 26191 6273 26203 6307
rect 26145 6267 26203 6273
rect 25961 6171 26019 6177
rect 25961 6137 25973 6171
rect 26007 6137 26019 6171
rect 26160 6168 26188 6267
rect 26234 6264 26240 6316
rect 26292 6264 26298 6316
rect 26421 6307 26479 6313
rect 26421 6273 26433 6307
rect 26467 6304 26479 6307
rect 26786 6304 26792 6316
rect 26467 6276 26792 6304
rect 26467 6273 26479 6276
rect 26421 6267 26479 6273
rect 26786 6264 26792 6276
rect 26844 6264 26850 6316
rect 27341 6307 27399 6313
rect 27341 6273 27353 6307
rect 27387 6273 27399 6307
rect 27341 6267 27399 6273
rect 26234 6168 26240 6180
rect 26160 6140 26240 6168
rect 25961 6131 26019 6137
rect 26234 6128 26240 6140
rect 26292 6128 26298 6180
rect 27356 6168 27384 6267
rect 27614 6264 27620 6316
rect 27672 6264 27678 6316
rect 28350 6264 28356 6316
rect 28408 6264 28414 6316
rect 27525 6239 27583 6245
rect 27525 6205 27537 6239
rect 27571 6236 27583 6239
rect 27982 6236 27988 6248
rect 27571 6208 27988 6236
rect 27571 6205 27583 6208
rect 27525 6199 27583 6205
rect 27982 6196 27988 6208
rect 28040 6236 28046 6248
rect 28040 6208 28212 6236
rect 28040 6196 28046 6208
rect 27890 6168 27896 6180
rect 27356 6140 27896 6168
rect 27890 6128 27896 6140
rect 27948 6128 27954 6180
rect 28184 6177 28212 6208
rect 28169 6171 28227 6177
rect 28169 6137 28181 6171
rect 28215 6137 28227 6171
rect 28169 6131 28227 6137
rect 13078 6060 13084 6112
rect 13136 6100 13142 6112
rect 13173 6103 13231 6109
rect 13173 6100 13185 6103
rect 13136 6072 13185 6100
rect 13136 6060 13142 6072
rect 13173 6069 13185 6072
rect 13219 6069 13231 6103
rect 13173 6063 13231 6069
rect 13722 6060 13728 6112
rect 13780 6100 13786 6112
rect 15470 6100 15476 6112
rect 13780 6072 15476 6100
rect 13780 6060 13786 6072
rect 15470 6060 15476 6072
rect 15528 6060 15534 6112
rect 15746 6060 15752 6112
rect 15804 6060 15810 6112
rect 23750 6060 23756 6112
rect 23808 6100 23814 6112
rect 24489 6103 24547 6109
rect 24489 6100 24501 6103
rect 23808 6072 24501 6100
rect 23808 6060 23814 6072
rect 24489 6069 24501 6072
rect 24535 6069 24547 6103
rect 24489 6063 24547 6069
rect 26142 6060 26148 6112
rect 26200 6060 26206 6112
rect 27522 6060 27528 6112
rect 27580 6060 27586 6112
rect 1104 6010 28704 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 28704 6010
rect 1104 5936 28704 5958
rect 16942 5856 16948 5908
rect 17000 5896 17006 5908
rect 17037 5899 17095 5905
rect 17037 5896 17049 5899
rect 17000 5868 17049 5896
rect 17000 5856 17006 5868
rect 17037 5865 17049 5868
rect 17083 5865 17095 5899
rect 17037 5859 17095 5865
rect 17218 5856 17224 5908
rect 17276 5896 17282 5908
rect 17405 5899 17463 5905
rect 17405 5896 17417 5899
rect 17276 5868 17417 5896
rect 17276 5856 17282 5868
rect 17405 5865 17417 5868
rect 17451 5865 17463 5899
rect 17405 5859 17463 5865
rect 22925 5899 22983 5905
rect 22925 5865 22937 5899
rect 22971 5896 22983 5899
rect 24578 5896 24584 5908
rect 22971 5868 24584 5896
rect 22971 5865 22983 5868
rect 22925 5859 22983 5865
rect 24578 5856 24584 5868
rect 24636 5856 24642 5908
rect 25038 5896 25044 5908
rect 24688 5868 25044 5896
rect 6914 5828 6920 5840
rect 6288 5800 6920 5828
rect 6288 5701 6316 5800
rect 6914 5788 6920 5800
rect 6972 5788 6978 5840
rect 14734 5788 14740 5840
rect 14792 5788 14798 5840
rect 15470 5788 15476 5840
rect 15528 5788 15534 5840
rect 23569 5831 23627 5837
rect 23569 5797 23581 5831
rect 23615 5828 23627 5831
rect 24210 5828 24216 5840
rect 23615 5800 24216 5828
rect 23615 5797 23627 5800
rect 23569 5791 23627 5797
rect 24210 5788 24216 5800
rect 24268 5788 24274 5840
rect 24688 5828 24716 5868
rect 25038 5856 25044 5868
rect 25096 5856 25102 5908
rect 25869 5899 25927 5905
rect 25869 5865 25881 5899
rect 25915 5896 25927 5899
rect 26142 5896 26148 5908
rect 25915 5868 26148 5896
rect 25915 5865 25927 5868
rect 25869 5859 25927 5865
rect 26142 5856 26148 5868
rect 26200 5856 26206 5908
rect 26421 5899 26479 5905
rect 26421 5865 26433 5899
rect 26467 5896 26479 5899
rect 26510 5896 26516 5908
rect 26467 5868 26516 5896
rect 26467 5865 26479 5868
rect 26421 5859 26479 5865
rect 26510 5856 26516 5868
rect 26568 5896 26574 5908
rect 26694 5896 26700 5908
rect 26568 5868 26700 5896
rect 26568 5856 26574 5868
rect 26694 5856 26700 5868
rect 26752 5856 26758 5908
rect 24320 5800 24716 5828
rect 6733 5763 6791 5769
rect 6733 5760 6745 5763
rect 6564 5732 6745 5760
rect 5997 5695 6055 5701
rect 5997 5661 6009 5695
rect 6043 5661 6055 5695
rect 5997 5655 6055 5661
rect 6181 5695 6239 5701
rect 6181 5661 6193 5695
rect 6227 5692 6239 5695
rect 6273 5695 6331 5701
rect 6273 5692 6285 5695
rect 6227 5664 6285 5692
rect 6227 5661 6239 5664
rect 6181 5655 6239 5661
rect 6273 5661 6285 5664
rect 6319 5661 6331 5695
rect 6273 5655 6331 5661
rect 6012 5624 6040 5655
rect 6454 5652 6460 5704
rect 6512 5652 6518 5704
rect 6472 5624 6500 5652
rect 6012 5596 6500 5624
rect 6089 5559 6147 5565
rect 6089 5525 6101 5559
rect 6135 5556 6147 5559
rect 6564 5556 6592 5732
rect 6733 5729 6745 5732
rect 6779 5729 6791 5763
rect 16666 5760 16672 5772
rect 6733 5723 6791 5729
rect 15212 5732 16068 5760
rect 6917 5695 6975 5701
rect 6917 5692 6929 5695
rect 6656 5664 6929 5692
rect 6656 5568 6684 5664
rect 6917 5661 6929 5664
rect 6963 5661 6975 5695
rect 6917 5655 6975 5661
rect 14918 5652 14924 5704
rect 14976 5652 14982 5704
rect 15212 5701 15240 5732
rect 15197 5695 15255 5701
rect 15197 5661 15209 5695
rect 15243 5661 15255 5695
rect 15197 5655 15255 5661
rect 15289 5695 15347 5701
rect 15289 5661 15301 5695
rect 15335 5692 15347 5695
rect 15930 5692 15936 5704
rect 15335 5664 15936 5692
rect 15335 5661 15347 5664
rect 15289 5655 15347 5661
rect 15930 5652 15936 5664
rect 15988 5652 15994 5704
rect 11146 5584 11152 5636
rect 11204 5624 11210 5636
rect 16040 5624 16068 5732
rect 16224 5732 16672 5760
rect 16224 5704 16252 5732
rect 16666 5720 16672 5732
rect 16724 5720 16730 5772
rect 17494 5720 17500 5772
rect 17552 5720 17558 5772
rect 21453 5763 21511 5769
rect 21453 5729 21465 5763
rect 21499 5760 21511 5763
rect 23293 5763 23351 5769
rect 23293 5760 23305 5763
rect 21499 5732 23305 5760
rect 21499 5729 21511 5732
rect 21453 5723 21511 5729
rect 23293 5729 23305 5732
rect 23339 5729 23351 5763
rect 23293 5723 23351 5729
rect 16117 5695 16175 5701
rect 16117 5661 16129 5695
rect 16163 5692 16175 5695
rect 16206 5692 16212 5704
rect 16163 5664 16212 5692
rect 16163 5661 16175 5664
rect 16117 5655 16175 5661
rect 16206 5652 16212 5664
rect 16264 5652 16270 5704
rect 16577 5695 16635 5701
rect 16577 5661 16589 5695
rect 16623 5692 16635 5695
rect 16942 5692 16948 5704
rect 16623 5664 16948 5692
rect 16623 5661 16635 5664
rect 16577 5655 16635 5661
rect 16942 5652 16948 5664
rect 17000 5652 17006 5704
rect 17037 5695 17095 5701
rect 17037 5661 17049 5695
rect 17083 5661 17095 5695
rect 17037 5655 17095 5661
rect 16298 5624 16304 5636
rect 11204 5596 15976 5624
rect 16040 5596 16304 5624
rect 11204 5584 11210 5596
rect 6135 5528 6592 5556
rect 6135 5525 6147 5528
rect 6089 5519 6147 5525
rect 6638 5516 6644 5568
rect 6696 5516 6702 5568
rect 7101 5559 7159 5565
rect 7101 5525 7113 5559
rect 7147 5556 7159 5559
rect 7466 5556 7472 5568
rect 7147 5528 7472 5556
rect 7147 5525 7159 5528
rect 7101 5519 7159 5525
rect 7466 5516 7472 5528
rect 7524 5516 7530 5568
rect 10226 5516 10232 5568
rect 10284 5556 10290 5568
rect 13078 5556 13084 5568
rect 10284 5528 13084 5556
rect 10284 5516 10290 5528
rect 13078 5516 13084 5528
rect 13136 5516 13142 5568
rect 15105 5559 15163 5565
rect 15105 5525 15117 5559
rect 15151 5556 15163 5559
rect 15286 5556 15292 5568
rect 15151 5528 15292 5556
rect 15151 5525 15163 5528
rect 15105 5519 15163 5525
rect 15286 5516 15292 5528
rect 15344 5516 15350 5568
rect 15948 5556 15976 5596
rect 16298 5584 16304 5596
rect 16356 5624 16362 5636
rect 17052 5624 17080 5655
rect 17310 5652 17316 5704
rect 17368 5652 17374 5704
rect 17678 5652 17684 5704
rect 17736 5652 17742 5704
rect 21174 5652 21180 5704
rect 21232 5652 21238 5704
rect 22554 5652 22560 5704
rect 22612 5652 22618 5704
rect 23474 5652 23480 5704
rect 23532 5652 23538 5704
rect 23661 5695 23719 5701
rect 23661 5661 23673 5695
rect 23707 5661 23719 5695
rect 23661 5655 23719 5661
rect 16356 5596 17080 5624
rect 23676 5624 23704 5655
rect 23750 5652 23756 5704
rect 23808 5652 23814 5704
rect 23937 5695 23995 5701
rect 23937 5661 23949 5695
rect 23983 5692 23995 5695
rect 24320 5692 24348 5800
rect 24854 5788 24860 5840
rect 24912 5788 24918 5840
rect 24394 5720 24400 5772
rect 24452 5760 24458 5772
rect 24765 5763 24823 5769
rect 24765 5760 24777 5763
rect 24452 5732 24777 5760
rect 24452 5720 24458 5732
rect 24765 5729 24777 5732
rect 24811 5729 24823 5763
rect 24872 5760 24900 5788
rect 24872 5732 25360 5760
rect 24765 5723 24823 5729
rect 23983 5664 24348 5692
rect 24581 5695 24639 5701
rect 23983 5661 23995 5664
rect 23937 5655 23995 5661
rect 24581 5661 24593 5695
rect 24627 5661 24639 5695
rect 24581 5655 24639 5661
rect 24596 5624 24624 5655
rect 24670 5652 24676 5704
rect 24728 5652 24734 5704
rect 24854 5652 24860 5704
rect 24912 5652 24918 5704
rect 25038 5652 25044 5704
rect 25096 5652 25102 5704
rect 25332 5701 25360 5732
rect 27982 5720 27988 5772
rect 28040 5720 28046 5772
rect 25317 5695 25375 5701
rect 25317 5661 25329 5695
rect 25363 5661 25375 5695
rect 25317 5655 25375 5661
rect 25406 5652 25412 5704
rect 25464 5692 25470 5704
rect 25593 5695 25651 5701
rect 25593 5692 25605 5695
rect 25464 5664 25605 5692
rect 25464 5652 25470 5664
rect 25593 5661 25605 5664
rect 25639 5661 25651 5695
rect 25593 5655 25651 5661
rect 25961 5695 26019 5701
rect 25961 5661 25973 5695
rect 26007 5692 26019 5695
rect 26053 5695 26111 5701
rect 26053 5692 26065 5695
rect 26007 5664 26065 5692
rect 26007 5661 26019 5664
rect 25961 5655 26019 5661
rect 26053 5661 26065 5664
rect 26099 5692 26111 5695
rect 26099 5664 26556 5692
rect 26099 5661 26111 5664
rect 26053 5655 26111 5661
rect 25133 5627 25191 5633
rect 25133 5624 25145 5627
rect 23676 5596 24624 5624
rect 16356 5584 16362 5596
rect 16853 5559 16911 5565
rect 16853 5556 16865 5559
rect 15948 5528 16865 5556
rect 16853 5525 16865 5528
rect 16899 5556 16911 5559
rect 17770 5556 17776 5568
rect 16899 5528 17776 5556
rect 16899 5525 16911 5528
rect 16853 5519 16911 5525
rect 17770 5516 17776 5528
rect 17828 5516 17834 5568
rect 24394 5516 24400 5568
rect 24452 5516 24458 5568
rect 24596 5556 24624 5596
rect 24872 5596 25145 5624
rect 24872 5556 24900 5596
rect 25133 5593 25145 5596
rect 25179 5593 25191 5627
rect 25133 5587 25191 5593
rect 25498 5584 25504 5636
rect 25556 5584 25562 5636
rect 26234 5584 26240 5636
rect 26292 5584 26298 5636
rect 26528 5568 26556 5664
rect 28258 5652 28264 5704
rect 28316 5652 28322 5704
rect 27246 5584 27252 5636
rect 27304 5584 27310 5636
rect 24596 5528 24900 5556
rect 26510 5516 26516 5568
rect 26568 5516 26574 5568
rect 1104 5466 28704 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 28704 5466
rect 1104 5392 28704 5414
rect 6457 5355 6515 5361
rect 6457 5321 6469 5355
rect 6503 5352 6515 5355
rect 6638 5352 6644 5364
rect 6503 5324 6644 5352
rect 6503 5321 6515 5324
rect 6457 5315 6515 5321
rect 6638 5312 6644 5324
rect 6696 5312 6702 5364
rect 6730 5312 6736 5364
rect 6788 5352 6794 5364
rect 12342 5352 12348 5364
rect 6788 5324 12348 5352
rect 6788 5312 6794 5324
rect 5258 5284 5264 5296
rect 4830 5256 5264 5284
rect 5258 5244 5264 5256
rect 5316 5244 5322 5296
rect 6546 5284 6552 5296
rect 6012 5256 6552 5284
rect 5718 5176 5724 5228
rect 5776 5216 5782 5228
rect 6012 5225 6040 5256
rect 6546 5244 6552 5256
rect 6604 5244 6610 5296
rect 7377 5287 7435 5293
rect 7377 5284 7389 5287
rect 6656 5256 7389 5284
rect 5997 5219 6055 5225
rect 5997 5216 6009 5219
rect 5776 5188 6009 5216
rect 5776 5176 5782 5188
rect 5997 5185 6009 5188
rect 6043 5185 6055 5219
rect 5997 5179 6055 5185
rect 6178 5176 6184 5228
rect 6236 5216 6242 5228
rect 6656 5225 6684 5256
rect 7377 5253 7389 5256
rect 7423 5253 7435 5287
rect 7377 5247 7435 5253
rect 7466 5244 7472 5296
rect 7524 5284 7530 5296
rect 8205 5287 8263 5293
rect 8205 5284 8217 5287
rect 7524 5256 8217 5284
rect 7524 5244 7530 5256
rect 8205 5253 8217 5256
rect 8251 5253 8263 5287
rect 9214 5284 9220 5296
rect 8205 5247 8263 5253
rect 8312 5256 9220 5284
rect 6914 5225 6920 5228
rect 6365 5219 6423 5225
rect 6365 5216 6377 5219
rect 6236 5188 6377 5216
rect 6236 5176 6242 5188
rect 6365 5185 6377 5188
rect 6411 5185 6423 5219
rect 6365 5179 6423 5185
rect 6641 5219 6699 5225
rect 6641 5185 6653 5219
rect 6687 5185 6699 5219
rect 6641 5179 6699 5185
rect 6891 5219 6920 5225
rect 6891 5185 6903 5219
rect 6891 5179 6920 5185
rect 6914 5176 6920 5179
rect 6972 5176 6978 5228
rect 7009 5219 7067 5225
rect 7009 5185 7021 5219
rect 7055 5185 7067 5219
rect 7009 5179 7067 5185
rect 3326 5108 3332 5160
rect 3384 5108 3390 5160
rect 3602 5108 3608 5160
rect 3660 5108 3666 5160
rect 5813 5151 5871 5157
rect 5813 5117 5825 5151
rect 5859 5117 5871 5151
rect 5813 5111 5871 5117
rect 4982 5040 4988 5092
rect 5040 5080 5046 5092
rect 5629 5083 5687 5089
rect 5629 5080 5641 5083
rect 5040 5052 5641 5080
rect 5040 5040 5046 5052
rect 5629 5049 5641 5052
rect 5675 5049 5687 5083
rect 5828 5080 5856 5111
rect 5902 5108 5908 5160
rect 5960 5108 5966 5160
rect 6089 5151 6147 5157
rect 6089 5117 6101 5151
rect 6135 5148 6147 5151
rect 6270 5148 6276 5160
rect 6135 5120 6276 5148
rect 6135 5117 6147 5120
rect 6089 5111 6147 5117
rect 6270 5108 6276 5120
rect 6328 5108 6334 5160
rect 6454 5108 6460 5160
rect 6512 5148 6518 5160
rect 6733 5151 6791 5157
rect 6733 5148 6745 5151
rect 6512 5120 6745 5148
rect 6512 5108 6518 5120
rect 6733 5117 6745 5120
rect 6779 5117 6791 5151
rect 7024 5148 7052 5179
rect 7098 5176 7104 5228
rect 7156 5176 7162 5228
rect 7193 5219 7251 5225
rect 7193 5185 7205 5219
rect 7239 5216 7251 5219
rect 7558 5216 7564 5228
rect 7239 5188 7564 5216
rect 7239 5185 7251 5188
rect 7193 5179 7251 5185
rect 7558 5176 7564 5188
rect 7616 5176 7622 5228
rect 7653 5219 7711 5225
rect 7653 5185 7665 5219
rect 7699 5185 7711 5219
rect 7653 5179 7711 5185
rect 7466 5148 7472 5160
rect 7024 5120 7472 5148
rect 6733 5111 6791 5117
rect 7466 5108 7472 5120
rect 7524 5108 7530 5160
rect 6546 5080 6552 5092
rect 5828 5052 6552 5080
rect 5629 5043 5687 5049
rect 6546 5040 6552 5052
rect 6604 5040 6610 5092
rect 6641 5083 6699 5089
rect 6641 5049 6653 5083
rect 6687 5080 6699 5083
rect 7668 5080 7696 5179
rect 8018 5176 8024 5228
rect 8076 5176 8082 5228
rect 8312 5225 8340 5256
rect 9214 5244 9220 5256
rect 9272 5244 9278 5296
rect 9508 5293 9536 5324
rect 12342 5312 12348 5324
rect 12400 5312 12406 5364
rect 15194 5312 15200 5364
rect 15252 5352 15258 5364
rect 15381 5355 15439 5361
rect 15381 5352 15393 5355
rect 15252 5324 15393 5352
rect 15252 5312 15258 5324
rect 15381 5321 15393 5324
rect 15427 5321 15439 5355
rect 15381 5315 15439 5321
rect 15562 5312 15568 5364
rect 15620 5352 15626 5364
rect 15749 5355 15807 5361
rect 15749 5352 15761 5355
rect 15620 5324 15761 5352
rect 15620 5312 15626 5324
rect 15749 5321 15761 5324
rect 15795 5321 15807 5355
rect 15749 5315 15807 5321
rect 15930 5312 15936 5364
rect 15988 5352 15994 5364
rect 15988 5324 16988 5352
rect 15988 5312 15994 5324
rect 9493 5287 9551 5293
rect 9493 5253 9505 5287
rect 9539 5253 9551 5287
rect 9493 5247 9551 5253
rect 9582 5244 9588 5296
rect 9640 5293 9646 5296
rect 9640 5287 9669 5293
rect 9657 5253 9669 5287
rect 9640 5247 9669 5253
rect 9640 5244 9646 5247
rect 11790 5244 11796 5296
rect 11848 5284 11854 5296
rect 12434 5284 12440 5296
rect 11848 5256 12440 5284
rect 11848 5244 11854 5256
rect 12434 5244 12440 5256
rect 12492 5284 12498 5296
rect 13170 5284 13176 5296
rect 12492 5256 13176 5284
rect 12492 5244 12498 5256
rect 13170 5244 13176 5256
rect 13228 5244 13234 5296
rect 16393 5287 16451 5293
rect 16393 5284 16405 5287
rect 15304 5256 16405 5284
rect 15304 5228 15332 5256
rect 16393 5253 16405 5256
rect 16439 5284 16451 5287
rect 16482 5284 16488 5296
rect 16439 5256 16488 5284
rect 16439 5253 16451 5256
rect 16393 5247 16451 5253
rect 16482 5244 16488 5256
rect 16540 5244 16546 5296
rect 16850 5244 16856 5296
rect 16908 5244 16914 5296
rect 16960 5284 16988 5324
rect 17218 5312 17224 5364
rect 17276 5312 17282 5364
rect 18417 5355 18475 5361
rect 18417 5321 18429 5355
rect 18463 5352 18475 5355
rect 18506 5352 18512 5364
rect 18463 5324 18512 5352
rect 18463 5321 18475 5324
rect 18417 5315 18475 5321
rect 18506 5312 18512 5324
rect 18564 5312 18570 5364
rect 19058 5312 19064 5364
rect 19116 5312 19122 5364
rect 19426 5312 19432 5364
rect 19484 5352 19490 5364
rect 19889 5355 19947 5361
rect 19889 5352 19901 5355
rect 19484 5324 19901 5352
rect 19484 5312 19490 5324
rect 19889 5321 19901 5324
rect 19935 5321 19947 5355
rect 19889 5315 19947 5321
rect 20438 5312 20444 5364
rect 20496 5352 20502 5364
rect 21821 5355 21879 5361
rect 21821 5352 21833 5355
rect 20496 5324 21833 5352
rect 20496 5312 20502 5324
rect 21821 5321 21833 5324
rect 21867 5321 21879 5355
rect 21821 5315 21879 5321
rect 17865 5287 17923 5293
rect 17865 5284 17877 5287
rect 16960 5256 17877 5284
rect 17865 5253 17877 5256
rect 17911 5284 17923 5287
rect 17954 5284 17960 5296
rect 17911 5256 17960 5284
rect 17911 5253 17923 5256
rect 17865 5247 17923 5253
rect 17954 5244 17960 5256
rect 18012 5244 18018 5296
rect 18064 5256 18735 5284
rect 8297 5219 8355 5225
rect 8297 5185 8309 5219
rect 8343 5185 8355 5219
rect 8297 5179 8355 5185
rect 8389 5219 8447 5225
rect 8389 5185 8401 5219
rect 8435 5216 8447 5219
rect 8478 5216 8484 5228
rect 8435 5188 8484 5216
rect 8435 5185 8447 5188
rect 8389 5179 8447 5185
rect 8478 5176 8484 5188
rect 8536 5176 8542 5228
rect 8573 5219 8631 5225
rect 8573 5185 8585 5219
rect 8619 5216 8631 5219
rect 8619 5188 8800 5216
rect 8619 5185 8631 5188
rect 8573 5179 8631 5185
rect 7926 5108 7932 5160
rect 7984 5108 7990 5160
rect 8665 5151 8723 5157
rect 8665 5117 8677 5151
rect 8711 5117 8723 5151
rect 8772 5148 8800 5188
rect 8846 5176 8852 5228
rect 8904 5176 8910 5228
rect 9306 5176 9312 5228
rect 9364 5176 9370 5228
rect 9398 5176 9404 5228
rect 9456 5176 9462 5228
rect 9508 5188 10732 5216
rect 9508 5148 9536 5188
rect 8772 5120 9536 5148
rect 8665 5111 8723 5117
rect 6687 5052 7696 5080
rect 6687 5049 6699 5052
rect 6641 5043 6699 5049
rect 7742 5040 7748 5092
rect 7800 5080 7806 5092
rect 8481 5083 8539 5089
rect 8481 5080 8493 5083
rect 7800 5052 8493 5080
rect 7800 5040 7806 5052
rect 8481 5049 8493 5052
rect 8527 5080 8539 5083
rect 8680 5080 8708 5111
rect 9582 5108 9588 5160
rect 9640 5148 9646 5160
rect 9769 5151 9827 5157
rect 9769 5148 9781 5151
rect 9640 5120 9781 5148
rect 9640 5108 9646 5120
rect 9769 5117 9781 5120
rect 9815 5117 9827 5151
rect 9769 5111 9827 5117
rect 10704 5092 10732 5188
rect 12710 5176 12716 5228
rect 12768 5216 12774 5228
rect 12897 5219 12955 5225
rect 12897 5216 12909 5219
rect 12768 5188 12909 5216
rect 12768 5176 12774 5188
rect 12897 5185 12909 5188
rect 12943 5185 12955 5219
rect 12897 5179 12955 5185
rect 12986 5176 12992 5228
rect 13044 5216 13050 5228
rect 13081 5219 13139 5225
rect 13081 5216 13093 5219
rect 13044 5188 13093 5216
rect 13044 5176 13050 5188
rect 13081 5185 13093 5188
rect 13127 5185 13139 5219
rect 13081 5179 13139 5185
rect 15286 5176 15292 5228
rect 15344 5176 15350 5228
rect 15562 5176 15568 5228
rect 15620 5176 15626 5228
rect 15838 5176 15844 5228
rect 15896 5216 15902 5228
rect 16025 5219 16083 5225
rect 16025 5216 16037 5219
rect 15896 5188 16037 5216
rect 15896 5176 15902 5188
rect 16025 5185 16037 5188
rect 16071 5185 16083 5219
rect 16025 5179 16083 5185
rect 16301 5219 16359 5225
rect 16301 5185 16313 5219
rect 16347 5216 16359 5219
rect 16347 5214 16436 5216
rect 16347 5188 16528 5214
rect 16347 5185 16359 5188
rect 16408 5186 16528 5188
rect 16301 5179 16359 5185
rect 12250 5108 12256 5160
rect 12308 5148 12314 5160
rect 15657 5151 15715 5157
rect 12308 5120 15516 5148
rect 12308 5108 12314 5120
rect 8527 5052 8708 5080
rect 9033 5083 9091 5089
rect 8527 5049 8539 5052
rect 8481 5043 8539 5049
rect 9033 5049 9045 5083
rect 9079 5080 9091 5083
rect 9214 5080 9220 5092
rect 9079 5052 9220 5080
rect 9079 5049 9091 5052
rect 9033 5043 9091 5049
rect 9214 5040 9220 5052
rect 9272 5080 9278 5092
rect 10134 5080 10140 5092
rect 9272 5052 10140 5080
rect 9272 5040 9278 5052
rect 10134 5040 10140 5052
rect 10192 5040 10198 5092
rect 10686 5040 10692 5092
rect 10744 5080 10750 5092
rect 15378 5080 15384 5092
rect 10744 5052 15384 5080
rect 10744 5040 10750 5052
rect 15378 5040 15384 5052
rect 15436 5040 15442 5092
rect 5077 5015 5135 5021
rect 5077 4981 5089 5015
rect 5123 5012 5135 5015
rect 5534 5012 5540 5024
rect 5123 4984 5540 5012
rect 5123 4981 5135 4984
rect 5077 4975 5135 4981
rect 5534 4972 5540 4984
rect 5592 5012 5598 5024
rect 6454 5012 6460 5024
rect 5592 4984 6460 5012
rect 5592 4972 5598 4984
rect 6454 4972 6460 4984
rect 6512 4972 6518 5024
rect 7469 5015 7527 5021
rect 7469 4981 7481 5015
rect 7515 5012 7527 5015
rect 7650 5012 7656 5024
rect 7515 4984 7656 5012
rect 7515 4981 7527 4984
rect 7469 4975 7527 4981
rect 7650 4972 7656 4984
rect 7708 4972 7714 5024
rect 7837 5015 7895 5021
rect 7837 4981 7849 5015
rect 7883 5012 7895 5015
rect 8113 5015 8171 5021
rect 8113 5012 8125 5015
rect 7883 4984 8125 5012
rect 7883 4981 7895 4984
rect 7837 4975 7895 4981
rect 8113 4981 8125 4984
rect 8159 4981 8171 5015
rect 8113 4975 8171 4981
rect 9122 4972 9128 5024
rect 9180 4972 9186 5024
rect 12986 4972 12992 5024
rect 13044 4972 13050 5024
rect 15488 5012 15516 5120
rect 15657 5117 15669 5151
rect 15703 5117 15715 5151
rect 15657 5111 15715 5117
rect 16209 5151 16267 5157
rect 16209 5117 16221 5151
rect 16255 5117 16267 5151
rect 16500 5148 16528 5186
rect 16574 5176 16580 5228
rect 16632 5216 16638 5228
rect 16669 5219 16727 5225
rect 16669 5216 16681 5219
rect 16632 5188 16681 5216
rect 16632 5176 16638 5188
rect 16669 5185 16681 5188
rect 16715 5185 16727 5219
rect 16669 5179 16727 5185
rect 16868 5148 16896 5244
rect 18064 5228 18092 5256
rect 16942 5176 16948 5228
rect 17000 5176 17006 5228
rect 17037 5219 17095 5225
rect 17037 5185 17049 5219
rect 17083 5216 17095 5219
rect 17310 5216 17316 5228
rect 17083 5188 17316 5216
rect 17083 5185 17095 5188
rect 17037 5179 17095 5185
rect 17310 5176 17316 5188
rect 17368 5176 17374 5228
rect 18046 5176 18052 5228
rect 18104 5176 18110 5228
rect 18141 5219 18199 5225
rect 18141 5185 18153 5219
rect 18187 5216 18199 5219
rect 18601 5219 18659 5225
rect 18601 5216 18613 5219
rect 18187 5188 18613 5216
rect 18187 5185 18199 5188
rect 18141 5179 18199 5185
rect 18601 5185 18613 5188
rect 18647 5185 18659 5219
rect 18707 5216 18735 5256
rect 19518 5244 19524 5296
rect 19576 5244 19582 5296
rect 19794 5244 19800 5296
rect 19852 5244 19858 5296
rect 18707 5214 18736 5216
rect 18782 5214 18788 5228
rect 18707 5188 18788 5214
rect 18708 5186 18788 5188
rect 18601 5179 18659 5185
rect 17586 5148 17592 5160
rect 16500 5120 17592 5148
rect 16209 5111 16267 5117
rect 15565 5083 15623 5089
rect 15565 5049 15577 5083
rect 15611 5080 15623 5083
rect 15672 5080 15700 5111
rect 15611 5052 15700 5080
rect 16224 5080 16252 5111
rect 17586 5108 17592 5120
rect 17644 5108 17650 5160
rect 17678 5080 17684 5092
rect 16224 5052 17684 5080
rect 15611 5049 15623 5052
rect 15565 5043 15623 5049
rect 17678 5040 17684 5052
rect 17736 5080 17742 5092
rect 17865 5083 17923 5089
rect 17865 5080 17877 5083
rect 17736 5052 17877 5080
rect 17736 5040 17742 5052
rect 17865 5049 17877 5052
rect 17911 5049 17923 5083
rect 18616 5080 18644 5179
rect 18782 5176 18788 5186
rect 18840 5176 18846 5228
rect 18874 5176 18880 5228
rect 18932 5176 18938 5228
rect 19337 5219 19395 5225
rect 19337 5216 19349 5219
rect 18984 5188 19349 5216
rect 18682 5151 18740 5157
rect 18682 5117 18694 5151
rect 18728 5148 18740 5151
rect 18984 5148 19012 5188
rect 19337 5185 19349 5188
rect 19383 5216 19395 5219
rect 19536 5216 19564 5244
rect 19383 5188 19564 5216
rect 19383 5185 19395 5188
rect 19337 5179 19395 5185
rect 18728 5120 19012 5148
rect 19245 5151 19303 5157
rect 18728 5117 18740 5120
rect 18682 5111 18740 5117
rect 19245 5117 19257 5151
rect 19291 5117 19303 5151
rect 19245 5111 19303 5117
rect 19260 5080 19288 5111
rect 19426 5108 19432 5160
rect 19484 5108 19490 5160
rect 19521 5151 19579 5157
rect 19521 5117 19533 5151
rect 19567 5148 19579 5151
rect 21836 5148 21864 5315
rect 22278 5312 22284 5364
rect 22336 5352 22342 5364
rect 23750 5352 23756 5364
rect 22336 5324 23756 5352
rect 22336 5312 22342 5324
rect 23750 5312 23756 5324
rect 23808 5312 23814 5364
rect 24305 5355 24363 5361
rect 24305 5321 24317 5355
rect 24351 5352 24363 5355
rect 24854 5352 24860 5364
rect 24351 5324 24860 5352
rect 24351 5321 24363 5324
rect 24305 5315 24363 5321
rect 24854 5312 24860 5324
rect 24912 5312 24918 5364
rect 25685 5355 25743 5361
rect 25685 5321 25697 5355
rect 25731 5352 25743 5355
rect 25958 5352 25964 5364
rect 25731 5324 25964 5352
rect 25731 5321 25743 5324
rect 25685 5315 25743 5321
rect 22554 5244 22560 5296
rect 22612 5244 22618 5296
rect 23293 5287 23351 5293
rect 23293 5253 23305 5287
rect 23339 5284 23351 5287
rect 24394 5284 24400 5296
rect 23339 5256 24400 5284
rect 23339 5253 23351 5256
rect 23293 5247 23351 5253
rect 24394 5244 24400 5256
rect 24452 5244 24458 5296
rect 24670 5244 24676 5296
rect 24728 5284 24734 5296
rect 25700 5284 25728 5315
rect 25958 5312 25964 5324
rect 26016 5312 26022 5364
rect 27614 5312 27620 5364
rect 27672 5352 27678 5364
rect 27982 5352 27988 5364
rect 27672 5324 27988 5352
rect 27672 5312 27678 5324
rect 27982 5312 27988 5324
rect 28040 5352 28046 5364
rect 28169 5355 28227 5361
rect 28169 5352 28181 5355
rect 28040 5324 28181 5352
rect 28040 5312 28046 5324
rect 28169 5321 28181 5324
rect 28215 5321 28227 5355
rect 28169 5315 28227 5321
rect 24728 5256 25728 5284
rect 24728 5244 24734 5256
rect 26234 5244 26240 5296
rect 26292 5284 26298 5296
rect 26292 5256 26648 5284
rect 26292 5244 26298 5256
rect 23842 5176 23848 5228
rect 23900 5216 23906 5228
rect 24581 5219 24639 5225
rect 24581 5216 24593 5219
rect 23900 5188 24593 5216
rect 23900 5176 23906 5188
rect 24581 5185 24593 5188
rect 24627 5185 24639 5219
rect 24581 5179 24639 5185
rect 24765 5219 24823 5225
rect 24765 5185 24777 5219
rect 24811 5216 24823 5219
rect 24946 5216 24952 5228
rect 24811 5188 24952 5216
rect 24811 5185 24823 5188
rect 24765 5179 24823 5185
rect 24946 5176 24952 5188
rect 25004 5176 25010 5228
rect 25038 5176 25044 5228
rect 25096 5176 25102 5228
rect 25317 5219 25375 5225
rect 25317 5185 25329 5219
rect 25363 5216 25375 5219
rect 25498 5216 25504 5228
rect 25363 5188 25504 5216
rect 25363 5185 25375 5188
rect 25317 5179 25375 5185
rect 25498 5176 25504 5188
rect 25556 5216 25562 5228
rect 25869 5219 25927 5225
rect 25869 5216 25881 5219
rect 25556 5188 25881 5216
rect 25556 5176 25562 5188
rect 25869 5185 25881 5188
rect 25915 5185 25927 5219
rect 25869 5179 25927 5185
rect 26510 5176 26516 5228
rect 26568 5176 26574 5228
rect 26620 5225 26648 5256
rect 26605 5219 26663 5225
rect 26605 5185 26617 5219
rect 26651 5185 26663 5219
rect 26605 5179 26663 5185
rect 28350 5176 28356 5228
rect 28408 5176 28414 5228
rect 19567 5120 19748 5148
rect 21836 5120 22324 5148
rect 19567 5117 19579 5120
rect 19521 5111 19579 5117
rect 19610 5080 19616 5092
rect 18616 5052 19616 5080
rect 17865 5043 17923 5049
rect 19610 5040 19616 5052
rect 19668 5040 19674 5092
rect 16666 5012 16672 5024
rect 15488 4984 16672 5012
rect 16666 4972 16672 4984
rect 16724 5012 16730 5024
rect 18874 5012 18880 5024
rect 16724 4984 18880 5012
rect 16724 4972 16730 4984
rect 18874 4972 18880 4984
rect 18932 4972 18938 5024
rect 18966 4972 18972 5024
rect 19024 5012 19030 5024
rect 19720 5012 19748 5120
rect 20162 5040 20168 5092
rect 20220 5080 20226 5092
rect 22186 5080 22192 5092
rect 20220 5052 22192 5080
rect 20220 5040 20226 5052
rect 22186 5040 22192 5052
rect 22244 5040 22250 5092
rect 19024 4984 19748 5012
rect 22296 5012 22324 5120
rect 23566 5108 23572 5160
rect 23624 5108 23630 5160
rect 23661 5151 23719 5157
rect 23661 5117 23673 5151
rect 23707 5117 23719 5151
rect 23661 5111 23719 5117
rect 23676 5012 23704 5111
rect 24854 5108 24860 5160
rect 24912 5108 24918 5160
rect 25593 5151 25651 5157
rect 25593 5117 25605 5151
rect 25639 5148 25651 5151
rect 26145 5151 26203 5157
rect 26145 5148 26157 5151
rect 25639 5120 26157 5148
rect 25639 5117 25651 5120
rect 25593 5111 25651 5117
rect 26145 5117 26157 5120
rect 26191 5148 26203 5151
rect 26237 5151 26295 5157
rect 26237 5148 26249 5151
rect 26191 5120 26249 5148
rect 26191 5117 26203 5120
rect 26145 5111 26203 5117
rect 26237 5117 26249 5120
rect 26283 5117 26295 5151
rect 26237 5111 26295 5117
rect 26421 5151 26479 5157
rect 26421 5117 26433 5151
rect 26467 5148 26479 5151
rect 26786 5148 26792 5160
rect 26467 5120 26792 5148
rect 26467 5117 26479 5120
rect 26421 5111 26479 5117
rect 26786 5108 26792 5120
rect 26844 5108 26850 5160
rect 24673 5083 24731 5089
rect 24673 5049 24685 5083
rect 24719 5080 24731 5083
rect 25133 5083 25191 5089
rect 25133 5080 25145 5083
rect 24719 5052 25145 5080
rect 24719 5049 24731 5052
rect 24673 5043 24731 5049
rect 25133 5049 25145 5052
rect 25179 5049 25191 5083
rect 25133 5043 25191 5049
rect 22296 4984 23704 5012
rect 19024 4972 19030 4984
rect 24394 4972 24400 5024
rect 24452 4972 24458 5024
rect 25498 4972 25504 5024
rect 25556 4972 25562 5024
rect 26053 5015 26111 5021
rect 26053 4981 26065 5015
rect 26099 5012 26111 5015
rect 26326 5012 26332 5024
rect 26099 4984 26332 5012
rect 26099 4981 26111 4984
rect 26053 4975 26111 4981
rect 26326 4972 26332 4984
rect 26384 4972 26390 5024
rect 1104 4922 28704 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 28704 4922
rect 1104 4848 28704 4870
rect 3602 4768 3608 4820
rect 3660 4808 3666 4820
rect 4709 4811 4767 4817
rect 4709 4808 4721 4811
rect 3660 4780 4721 4808
rect 3660 4768 3666 4780
rect 4709 4777 4721 4780
rect 4755 4777 4767 4811
rect 4709 4771 4767 4777
rect 5169 4811 5227 4817
rect 5169 4777 5181 4811
rect 5215 4808 5227 4811
rect 5350 4808 5356 4820
rect 5215 4780 5356 4808
rect 5215 4777 5227 4780
rect 5169 4771 5227 4777
rect 5350 4768 5356 4780
rect 5408 4768 5414 4820
rect 5902 4768 5908 4820
rect 5960 4808 5966 4820
rect 6089 4811 6147 4817
rect 6089 4808 6101 4811
rect 5960 4780 6101 4808
rect 5960 4768 5966 4780
rect 6089 4777 6101 4780
rect 6135 4777 6147 4811
rect 6089 4771 6147 4777
rect 6178 4768 6184 4820
rect 6236 4808 6242 4820
rect 6273 4811 6331 4817
rect 6273 4808 6285 4811
rect 6236 4780 6285 4808
rect 6236 4768 6242 4780
rect 6273 4777 6285 4780
rect 6319 4777 6331 4811
rect 6273 4771 6331 4777
rect 5721 4675 5779 4681
rect 5721 4641 5733 4675
rect 5767 4672 5779 4675
rect 6086 4672 6092 4684
rect 5767 4644 6092 4672
rect 5767 4641 5779 4644
rect 5721 4635 5779 4641
rect 6086 4632 6092 4644
rect 6144 4632 6150 4684
rect 6288 4672 6316 4771
rect 6546 4768 6552 4820
rect 6604 4808 6610 4820
rect 6733 4811 6791 4817
rect 6733 4808 6745 4811
rect 6604 4780 6745 4808
rect 6604 4768 6610 4780
rect 6733 4777 6745 4780
rect 6779 4777 6791 4811
rect 6733 4771 6791 4777
rect 7006 4768 7012 4820
rect 7064 4808 7070 4820
rect 7745 4811 7803 4817
rect 7745 4808 7757 4811
rect 7064 4780 7757 4808
rect 7064 4768 7070 4780
rect 7745 4777 7757 4780
rect 7791 4808 7803 4811
rect 8018 4808 8024 4820
rect 7791 4780 8024 4808
rect 7791 4777 7803 4780
rect 7745 4771 7803 4777
rect 8018 4768 8024 4780
rect 8076 4768 8082 4820
rect 9125 4811 9183 4817
rect 9125 4777 9137 4811
rect 9171 4808 9183 4811
rect 9306 4808 9312 4820
rect 9171 4780 9312 4808
rect 9171 4777 9183 4780
rect 9125 4771 9183 4777
rect 9306 4768 9312 4780
rect 9364 4768 9370 4820
rect 9398 4768 9404 4820
rect 9456 4808 9462 4820
rect 10413 4811 10471 4817
rect 10413 4808 10425 4811
rect 9456 4780 10425 4808
rect 9456 4768 9462 4780
rect 10413 4777 10425 4780
rect 10459 4777 10471 4811
rect 13541 4811 13599 4817
rect 13541 4808 13553 4811
rect 10413 4771 10471 4777
rect 11992 4780 13553 4808
rect 6454 4700 6460 4752
rect 6512 4740 6518 4752
rect 6641 4743 6699 4749
rect 6641 4740 6653 4743
rect 6512 4712 6653 4740
rect 6512 4700 6518 4712
rect 6641 4709 6653 4712
rect 6687 4740 6699 4743
rect 7193 4743 7251 4749
rect 7193 4740 7205 4743
rect 6687 4712 7205 4740
rect 6687 4709 6699 4712
rect 6641 4703 6699 4709
rect 7193 4709 7205 4712
rect 7239 4709 7251 4743
rect 7466 4740 7472 4752
rect 7193 4703 7251 4709
rect 7300 4712 7472 4740
rect 6825 4675 6883 4681
rect 6288 4644 6592 4672
rect 4893 4607 4951 4613
rect 4893 4573 4905 4607
rect 4939 4573 4951 4607
rect 4893 4567 4951 4573
rect 4908 4536 4936 4567
rect 4982 4564 4988 4616
rect 5040 4564 5046 4616
rect 5261 4607 5319 4613
rect 5261 4573 5273 4607
rect 5307 4604 5319 4607
rect 5442 4604 5448 4616
rect 5307 4576 5448 4604
rect 5307 4573 5319 4576
rect 5261 4567 5319 4573
rect 5442 4564 5448 4576
rect 5500 4564 5506 4616
rect 5537 4607 5595 4613
rect 5537 4573 5549 4607
rect 5583 4573 5595 4607
rect 5537 4567 5595 4573
rect 6365 4607 6423 4613
rect 6365 4573 6377 4607
rect 6411 4573 6423 4607
rect 6365 4567 6423 4573
rect 5353 4539 5411 4545
rect 5353 4536 5365 4539
rect 4908 4508 5365 4536
rect 5353 4505 5365 4508
rect 5399 4505 5411 4539
rect 5552 4536 5580 4567
rect 5810 4536 5816 4548
rect 5552 4508 5816 4536
rect 5353 4499 5411 4505
rect 5810 4496 5816 4508
rect 5868 4496 5874 4548
rect 6380 4468 6408 4567
rect 6454 4564 6460 4616
rect 6512 4564 6518 4616
rect 6564 4613 6592 4644
rect 6825 4641 6837 4675
rect 6871 4672 6883 4675
rect 7300 4672 7328 4712
rect 7466 4700 7472 4712
rect 7524 4700 7530 4752
rect 7558 4700 7564 4752
rect 7616 4740 7622 4752
rect 8205 4743 8263 4749
rect 8205 4740 8217 4743
rect 7616 4712 8217 4740
rect 7616 4700 7622 4712
rect 8205 4709 8217 4712
rect 8251 4709 8263 4743
rect 9582 4740 9588 4752
rect 8205 4703 8263 4709
rect 8588 4712 9588 4740
rect 6871 4644 7328 4672
rect 7484 4644 8156 4672
rect 6871 4641 6883 4644
rect 6825 4635 6883 4641
rect 6549 4607 6607 4613
rect 6549 4573 6561 4607
rect 6595 4573 6607 4607
rect 6549 4567 6607 4573
rect 6840 4468 6868 4635
rect 7006 4564 7012 4616
rect 7064 4564 7070 4616
rect 7484 4613 7512 4644
rect 8128 4613 8156 4644
rect 8478 4632 8484 4684
rect 8536 4632 8542 4684
rect 8588 4681 8616 4712
rect 9582 4700 9588 4712
rect 9640 4700 9646 4752
rect 8573 4675 8631 4681
rect 8573 4641 8585 4675
rect 8619 4641 8631 4675
rect 8573 4635 8631 4641
rect 9858 4632 9864 4684
rect 9916 4672 9922 4684
rect 10505 4675 10563 4681
rect 10505 4672 10517 4675
rect 9916 4644 10517 4672
rect 9916 4632 9922 4644
rect 10505 4641 10517 4644
rect 10551 4641 10563 4675
rect 10505 4635 10563 4641
rect 7469 4607 7527 4613
rect 7469 4573 7481 4607
rect 7515 4573 7527 4607
rect 7469 4567 7527 4573
rect 7837 4607 7895 4613
rect 7837 4573 7849 4607
rect 7883 4573 7895 4607
rect 7837 4567 7895 4573
rect 8113 4607 8171 4613
rect 8113 4573 8125 4607
rect 8159 4604 8171 4607
rect 8294 4604 8300 4616
rect 8159 4576 8300 4604
rect 8159 4573 8171 4576
rect 8113 4567 8171 4573
rect 7377 4539 7435 4545
rect 7377 4505 7389 4539
rect 7423 4536 7435 4539
rect 7742 4536 7748 4548
rect 7423 4508 7748 4536
rect 7423 4505 7435 4508
rect 7377 4499 7435 4505
rect 7742 4496 7748 4508
rect 7800 4496 7806 4548
rect 7852 4536 7880 4567
rect 8294 4564 8300 4576
rect 8352 4564 8358 4616
rect 8386 4564 8392 4616
rect 8444 4564 8450 4616
rect 8662 4564 8668 4616
rect 8720 4564 8726 4616
rect 8754 4564 8760 4616
rect 8812 4604 8818 4616
rect 9039 4607 9097 4613
rect 9039 4604 9051 4607
rect 8812 4576 9051 4604
rect 8812 4564 8818 4576
rect 9039 4573 9051 4576
rect 9085 4604 9097 4607
rect 9085 4576 9168 4604
rect 9085 4573 9097 4576
rect 9039 4567 9097 4573
rect 8680 4536 8708 4564
rect 7852 4508 8708 4536
rect 9140 4536 9168 4576
rect 9214 4564 9220 4616
rect 9272 4564 9278 4616
rect 9490 4564 9496 4616
rect 9548 4564 9554 4616
rect 9582 4564 9588 4616
rect 9640 4564 9646 4616
rect 10134 4564 10140 4616
rect 10192 4604 10198 4616
rect 10229 4607 10287 4613
rect 10229 4604 10241 4607
rect 10192 4576 10241 4604
rect 10192 4564 10198 4576
rect 10229 4573 10241 4576
rect 10275 4573 10287 4607
rect 10229 4567 10287 4573
rect 10686 4564 10692 4616
rect 10744 4564 10750 4616
rect 11992 4613 12020 4780
rect 13541 4777 13553 4780
rect 13587 4808 13599 4811
rect 13906 4808 13912 4820
rect 13587 4780 13912 4808
rect 13587 4777 13599 4780
rect 13541 4771 13599 4777
rect 13906 4768 13912 4780
rect 13964 4768 13970 4820
rect 16114 4768 16120 4820
rect 16172 4768 16178 4820
rect 16390 4768 16396 4820
rect 16448 4768 16454 4820
rect 16669 4811 16727 4817
rect 16669 4777 16681 4811
rect 16715 4808 16727 4811
rect 18046 4808 18052 4820
rect 16715 4780 18052 4808
rect 16715 4777 16727 4780
rect 16669 4771 16727 4777
rect 18046 4768 18052 4780
rect 18104 4808 18110 4820
rect 18325 4811 18383 4817
rect 18325 4808 18337 4811
rect 18104 4780 18337 4808
rect 18104 4768 18110 4780
rect 18325 4777 18337 4780
rect 18371 4777 18383 4811
rect 18325 4771 18383 4777
rect 18506 4768 18512 4820
rect 18564 4768 18570 4820
rect 23569 4811 23627 4817
rect 23569 4777 23581 4811
rect 23615 4808 23627 4811
rect 24854 4808 24860 4820
rect 23615 4780 24860 4808
rect 23615 4777 23627 4780
rect 23569 4771 23627 4777
rect 24854 4768 24860 4780
rect 24912 4768 24918 4820
rect 25498 4768 25504 4820
rect 25556 4808 25562 4820
rect 25866 4808 25872 4820
rect 25556 4780 25872 4808
rect 25556 4768 25562 4780
rect 25866 4768 25872 4780
rect 25924 4808 25930 4820
rect 25961 4811 26019 4817
rect 25961 4808 25973 4811
rect 25924 4780 25973 4808
rect 25924 4768 25930 4780
rect 25961 4777 25973 4780
rect 26007 4777 26019 4811
rect 25961 4771 26019 4777
rect 26234 4768 26240 4820
rect 26292 4808 26298 4820
rect 26513 4811 26571 4817
rect 26513 4808 26525 4811
rect 26292 4780 26525 4808
rect 26292 4768 26298 4780
rect 26513 4777 26525 4780
rect 26559 4777 26571 4811
rect 26513 4771 26571 4777
rect 12618 4700 12624 4752
rect 12676 4740 12682 4752
rect 12676 4712 13676 4740
rect 12676 4700 12682 4712
rect 12434 4632 12440 4684
rect 12492 4632 12498 4684
rect 12986 4672 12992 4684
rect 12544 4644 12992 4672
rect 10781 4607 10839 4613
rect 10781 4573 10793 4607
rect 10827 4573 10839 4607
rect 10781 4567 10839 4573
rect 11977 4607 12035 4613
rect 11977 4573 11989 4607
rect 12023 4573 12035 4607
rect 11977 4567 12035 4573
rect 9309 4539 9367 4545
rect 9309 4536 9321 4539
rect 9140 4508 9321 4536
rect 9309 4505 9321 4508
rect 9355 4536 9367 4539
rect 10045 4539 10103 4545
rect 10045 4536 10057 4539
rect 9355 4508 10057 4536
rect 9355 4505 9367 4508
rect 9309 4499 9367 4505
rect 10045 4505 10057 4508
rect 10091 4505 10103 4539
rect 10045 4499 10103 4505
rect 10502 4496 10508 4548
rect 10560 4536 10566 4548
rect 10796 4536 10824 4567
rect 12158 4564 12164 4616
rect 12216 4564 12222 4616
rect 12452 4591 12480 4632
rect 12544 4613 12572 4644
rect 12986 4632 12992 4644
rect 13044 4632 13050 4684
rect 13648 4616 13676 4712
rect 15562 4700 15568 4752
rect 15620 4740 15626 4752
rect 16942 4740 16948 4752
rect 15620 4712 16948 4740
rect 15620 4700 15626 4712
rect 16942 4700 16948 4712
rect 17000 4740 17006 4752
rect 18690 4740 18696 4752
rect 17000 4712 18696 4740
rect 17000 4700 17006 4712
rect 18690 4700 18696 4712
rect 18748 4700 18754 4752
rect 19426 4740 19432 4752
rect 18800 4712 19432 4740
rect 15746 4632 15752 4684
rect 15804 4632 15810 4684
rect 16482 4632 16488 4684
rect 16540 4632 16546 4684
rect 17310 4672 17316 4684
rect 16684 4644 17316 4672
rect 12529 4607 12587 4613
rect 12437 4585 12495 4591
rect 12437 4551 12449 4585
rect 12483 4551 12495 4585
rect 12529 4573 12541 4607
rect 12575 4573 12587 4607
rect 12529 4567 12587 4573
rect 12618 4564 12624 4616
rect 12676 4564 12682 4616
rect 12802 4564 12808 4616
rect 12860 4564 12866 4616
rect 12894 4564 12900 4616
rect 12952 4564 12958 4616
rect 13170 4564 13176 4616
rect 13228 4564 13234 4616
rect 13446 4564 13452 4616
rect 13504 4564 13510 4616
rect 13630 4564 13636 4616
rect 13688 4564 13694 4616
rect 13722 4564 13728 4616
rect 13780 4564 13786 4616
rect 13909 4607 13967 4613
rect 13909 4573 13921 4607
rect 13955 4604 13967 4607
rect 14550 4604 14556 4616
rect 13955 4576 14556 4604
rect 13955 4573 13967 4576
rect 13909 4567 13967 4573
rect 14550 4564 14556 4576
rect 14608 4564 14614 4616
rect 15838 4564 15844 4616
rect 15896 4564 15902 4616
rect 16206 4564 16212 4616
rect 16264 4564 16270 4616
rect 16393 4607 16451 4613
rect 16393 4573 16405 4607
rect 16439 4604 16451 4607
rect 16574 4604 16580 4616
rect 16439 4576 16580 4604
rect 16439 4573 16451 4576
rect 16393 4567 16451 4573
rect 16574 4564 16580 4576
rect 16632 4564 16638 4616
rect 12437 4545 12495 4551
rect 10560 4508 10824 4536
rect 12069 4539 12127 4545
rect 10560 4496 10566 4508
rect 12069 4505 12081 4539
rect 12115 4536 12127 4539
rect 12820 4536 12848 4564
rect 12115 4508 12388 4536
rect 12820 4508 13216 4536
rect 12115 4505 12127 4508
rect 12069 4499 12127 4505
rect 6380 4440 6868 4468
rect 7558 4428 7564 4480
rect 7616 4428 7622 4480
rect 7926 4428 7932 4480
rect 7984 4468 7990 4480
rect 9953 4471 10011 4477
rect 9953 4468 9965 4471
rect 7984 4440 9965 4468
rect 7984 4428 7990 4440
rect 9953 4437 9965 4440
rect 9999 4468 10011 4471
rect 11974 4468 11980 4480
rect 9999 4440 11980 4468
rect 9999 4437 10011 4440
rect 9953 4431 10011 4437
rect 11974 4428 11980 4440
rect 12032 4468 12038 4480
rect 12253 4471 12311 4477
rect 12253 4468 12265 4471
rect 12032 4440 12265 4468
rect 12032 4428 12038 4440
rect 12253 4437 12265 4440
rect 12299 4437 12311 4471
rect 12360 4468 12388 4508
rect 12986 4468 12992 4480
rect 12360 4440 12992 4468
rect 12253 4431 12311 4437
rect 12986 4428 12992 4440
rect 13044 4428 13050 4480
rect 13188 4468 13216 4508
rect 13354 4496 13360 4548
rect 13412 4496 13418 4548
rect 15194 4496 15200 4548
rect 15252 4536 15258 4548
rect 16684 4536 16712 4644
rect 17310 4632 17316 4644
rect 17368 4672 17374 4684
rect 18800 4672 18828 4712
rect 19426 4700 19432 4712
rect 19484 4700 19490 4752
rect 24394 4740 24400 4752
rect 22756 4712 24400 4740
rect 19794 4672 19800 4684
rect 17368 4644 18828 4672
rect 18892 4644 19800 4672
rect 17368 4632 17374 4644
rect 16761 4607 16819 4613
rect 16761 4573 16773 4607
rect 16807 4604 16819 4607
rect 16850 4604 16856 4616
rect 16807 4576 16856 4604
rect 16807 4573 16819 4576
rect 16761 4567 16819 4573
rect 16850 4564 16856 4576
rect 16908 4564 16914 4616
rect 17034 4564 17040 4616
rect 17092 4564 17098 4616
rect 17218 4564 17224 4616
rect 17276 4564 17282 4616
rect 18892 4613 18920 4644
rect 19794 4632 19800 4644
rect 19852 4632 19858 4684
rect 22557 4675 22615 4681
rect 22557 4641 22569 4675
rect 22603 4672 22615 4675
rect 22756 4672 22784 4712
rect 24394 4700 24400 4712
rect 24452 4700 24458 4752
rect 22603 4644 22784 4672
rect 22833 4675 22891 4681
rect 22603 4641 22615 4644
rect 22557 4635 22615 4641
rect 22833 4641 22845 4675
rect 22879 4672 22891 4675
rect 23566 4672 23572 4684
rect 22879 4644 23572 4672
rect 22879 4641 22891 4644
rect 22833 4635 22891 4641
rect 23566 4632 23572 4644
rect 23624 4632 23630 4684
rect 26694 4672 26700 4684
rect 26252 4644 26700 4672
rect 18417 4607 18475 4613
rect 18417 4573 18429 4607
rect 18463 4604 18475 4607
rect 18877 4607 18935 4613
rect 18877 4604 18889 4607
rect 18463 4576 18889 4604
rect 18463 4573 18475 4576
rect 18417 4567 18475 4573
rect 18877 4573 18889 4576
rect 18923 4573 18935 4607
rect 18877 4567 18935 4573
rect 19058 4564 19064 4616
rect 19116 4604 19122 4616
rect 19116 4576 19380 4604
rect 19116 4564 19122 4576
rect 15252 4508 16712 4536
rect 16868 4536 16896 4564
rect 18693 4539 18751 4545
rect 16868 4508 18276 4536
rect 15252 4496 15258 4508
rect 13814 4468 13820 4480
rect 13188 4440 13820 4468
rect 13814 4428 13820 4440
rect 13872 4428 13878 4480
rect 16853 4471 16911 4477
rect 16853 4437 16865 4471
rect 16899 4468 16911 4471
rect 17126 4468 17132 4480
rect 16899 4440 17132 4468
rect 16899 4437 16911 4440
rect 16853 4431 16911 4437
rect 17126 4428 17132 4440
rect 17184 4428 17190 4480
rect 18248 4468 18276 4508
rect 18693 4505 18705 4539
rect 18739 4505 18751 4539
rect 18693 4499 18751 4505
rect 18708 4468 18736 4499
rect 19242 4496 19248 4548
rect 19300 4496 19306 4548
rect 19352 4536 19380 4576
rect 19610 4564 19616 4616
rect 19668 4564 19674 4616
rect 20162 4564 20168 4616
rect 20220 4564 20226 4616
rect 20438 4564 20444 4616
rect 20496 4564 20502 4616
rect 22925 4607 22983 4613
rect 22925 4573 22937 4607
rect 22971 4573 22983 4607
rect 22925 4567 22983 4573
rect 19797 4539 19855 4545
rect 19797 4536 19809 4539
rect 19352 4508 19809 4536
rect 19797 4505 19809 4508
rect 19843 4505 19855 4539
rect 22554 4536 22560 4548
rect 22126 4508 22560 4536
rect 19797 4499 19855 4505
rect 22554 4496 22560 4508
rect 22612 4496 22618 4548
rect 18248 4440 18736 4468
rect 18782 4428 18788 4480
rect 18840 4468 18846 4480
rect 19429 4471 19487 4477
rect 19429 4468 19441 4471
rect 18840 4440 19441 4468
rect 18840 4428 18846 4440
rect 19429 4437 19441 4440
rect 19475 4437 19487 4471
rect 19429 4431 19487 4437
rect 19518 4428 19524 4480
rect 19576 4428 19582 4480
rect 19978 4428 19984 4480
rect 20036 4428 20042 4480
rect 20254 4428 20260 4480
rect 20312 4428 20318 4480
rect 20990 4428 20996 4480
rect 21048 4468 21054 4480
rect 21085 4471 21143 4477
rect 21085 4468 21097 4471
rect 21048 4440 21097 4468
rect 21048 4428 21054 4440
rect 21085 4437 21097 4440
rect 21131 4468 21143 4471
rect 22940 4468 22968 4567
rect 25958 4564 25964 4616
rect 26016 4564 26022 4616
rect 26252 4613 26280 4644
rect 26694 4632 26700 4644
rect 26752 4632 26758 4684
rect 27982 4632 27988 4684
rect 28040 4632 28046 4684
rect 26145 4607 26203 4613
rect 26145 4573 26157 4607
rect 26191 4604 26203 4607
rect 26237 4607 26295 4613
rect 26237 4604 26249 4607
rect 26191 4576 26249 4604
rect 26191 4573 26203 4576
rect 26145 4567 26203 4573
rect 26237 4573 26249 4576
rect 26283 4573 26295 4607
rect 26237 4567 26295 4573
rect 26421 4607 26479 4613
rect 26421 4573 26433 4607
rect 26467 4604 26479 4607
rect 26602 4604 26608 4616
rect 26467 4576 26608 4604
rect 26467 4573 26479 4576
rect 26421 4567 26479 4573
rect 26602 4564 26608 4576
rect 26660 4564 26666 4616
rect 28258 4564 28264 4616
rect 28316 4564 28322 4616
rect 27246 4496 27252 4548
rect 27304 4496 27310 4548
rect 21131 4440 22968 4468
rect 21131 4437 21143 4440
rect 21085 4431 21143 4437
rect 26234 4428 26240 4480
rect 26292 4468 26298 4480
rect 26329 4471 26387 4477
rect 26329 4468 26341 4471
rect 26292 4440 26341 4468
rect 26292 4428 26298 4440
rect 26329 4437 26341 4440
rect 26375 4437 26387 4471
rect 26329 4431 26387 4437
rect 1104 4378 28704 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 28704 4378
rect 1104 4304 28704 4326
rect 6178 4224 6184 4276
rect 6236 4224 6242 4276
rect 6270 4224 6276 4276
rect 6328 4264 6334 4276
rect 6328 4236 7328 4264
rect 6328 4224 6334 4236
rect 5350 4156 5356 4208
rect 5408 4196 5414 4208
rect 5408 4168 6684 4196
rect 5408 4156 5414 4168
rect 5994 4088 6000 4140
rect 6052 4088 6058 4140
rect 6365 4131 6423 4137
rect 6365 4097 6377 4131
rect 6411 4128 6423 4131
rect 6454 4128 6460 4140
rect 6411 4100 6460 4128
rect 6411 4097 6423 4100
rect 6365 4091 6423 4097
rect 6454 4088 6460 4100
rect 6512 4088 6518 4140
rect 6656 4128 6684 4168
rect 6730 4156 6736 4208
rect 6788 4156 6794 4208
rect 7190 4196 7196 4208
rect 6840 4168 7196 4196
rect 6840 4128 6868 4168
rect 7190 4156 7196 4168
rect 7248 4156 7254 4208
rect 7300 4140 7328 4236
rect 8294 4224 8300 4276
rect 8352 4264 8358 4276
rect 8481 4267 8539 4273
rect 8481 4264 8493 4267
rect 8352 4236 8493 4264
rect 8352 4224 8358 4236
rect 8481 4233 8493 4236
rect 8527 4233 8539 4267
rect 8481 4227 8539 4233
rect 9122 4224 9128 4276
rect 9180 4264 9186 4276
rect 9217 4267 9275 4273
rect 9217 4264 9229 4267
rect 9180 4236 9229 4264
rect 9180 4224 9186 4236
rect 9217 4233 9229 4236
rect 9263 4233 9275 4267
rect 9217 4227 9275 4233
rect 12066 4224 12072 4276
rect 12124 4224 12130 4276
rect 12342 4224 12348 4276
rect 12400 4264 12406 4276
rect 12400 4236 12940 4264
rect 12400 4224 12406 4236
rect 8386 4156 8392 4208
rect 8444 4196 8450 4208
rect 8846 4196 8852 4208
rect 8444 4168 8852 4196
rect 8444 4156 8450 4168
rect 6656 4100 6868 4128
rect 7009 4131 7067 4137
rect 7009 4097 7021 4131
rect 7055 4097 7067 4131
rect 7009 4091 7067 4097
rect 5810 4020 5816 4072
rect 5868 4060 5874 4072
rect 6638 4060 6644 4072
rect 5868 4032 6644 4060
rect 5868 4020 5874 4032
rect 6638 4020 6644 4032
rect 6696 4020 6702 4072
rect 7024 4060 7052 4091
rect 7098 4088 7104 4140
rect 7156 4088 7162 4140
rect 7282 4088 7288 4140
rect 7340 4088 7346 4140
rect 8496 4137 8524 4168
rect 8846 4156 8852 4168
rect 8904 4196 8910 4208
rect 9585 4199 9643 4205
rect 9585 4196 9597 4199
rect 8904 4168 9597 4196
rect 8904 4156 8910 4168
rect 9585 4165 9597 4168
rect 9631 4165 9643 4199
rect 9585 4159 9643 4165
rect 9953 4199 10011 4205
rect 9953 4165 9965 4199
rect 9999 4196 10011 4199
rect 10594 4196 10600 4208
rect 9999 4168 10600 4196
rect 9999 4165 10011 4168
rect 9953 4159 10011 4165
rect 10594 4156 10600 4168
rect 10652 4156 10658 4208
rect 11974 4156 11980 4208
rect 12032 4156 12038 4208
rect 12084 4196 12112 4224
rect 12912 4205 12940 4236
rect 13722 4224 13728 4276
rect 13780 4264 13786 4276
rect 16485 4267 16543 4273
rect 13780 4236 14228 4264
rect 13780 4224 13786 4236
rect 12187 4199 12245 4205
rect 12187 4196 12199 4199
rect 12084 4168 12199 4196
rect 12187 4165 12199 4168
rect 12233 4196 12245 4199
rect 12759 4199 12817 4205
rect 12759 4196 12771 4199
rect 12233 4168 12771 4196
rect 12233 4165 12245 4168
rect 12187 4159 12245 4165
rect 12759 4165 12771 4168
rect 12805 4165 12817 4199
rect 12759 4159 12817 4165
rect 12897 4199 12955 4205
rect 12897 4165 12909 4199
rect 12943 4165 12955 4199
rect 12897 4159 12955 4165
rect 8481 4131 8539 4137
rect 8481 4097 8493 4131
rect 8527 4097 8539 4131
rect 8481 4091 8539 4097
rect 8665 4131 8723 4137
rect 8665 4097 8677 4131
rect 8711 4128 8723 4131
rect 8754 4128 8760 4140
rect 8711 4100 8760 4128
rect 8711 4097 8723 4100
rect 8665 4091 8723 4097
rect 8754 4088 8760 4100
rect 8812 4088 8818 4140
rect 9125 4131 9183 4137
rect 9125 4097 9137 4131
rect 9171 4128 9183 4131
rect 9769 4131 9827 4137
rect 9769 4128 9781 4131
rect 9171 4100 9781 4128
rect 9171 4097 9183 4100
rect 9125 4091 9183 4097
rect 9769 4097 9781 4100
rect 9815 4128 9827 4131
rect 9858 4128 9864 4140
rect 9815 4100 9864 4128
rect 9815 4097 9827 4100
rect 9769 4091 9827 4097
rect 8570 4060 8576 4072
rect 7024 4032 8576 4060
rect 8570 4020 8576 4032
rect 8628 4060 8634 4072
rect 9140 4060 9168 4091
rect 9858 4088 9864 4100
rect 9916 4128 9922 4140
rect 10502 4128 10508 4140
rect 9916 4100 10508 4128
rect 9916 4088 9922 4100
rect 10502 4088 10508 4100
rect 10560 4088 10566 4140
rect 10689 4131 10747 4137
rect 10689 4097 10701 4131
rect 10735 4128 10747 4131
rect 11422 4128 11428 4140
rect 10735 4100 11428 4128
rect 10735 4097 10747 4100
rect 10689 4091 10747 4097
rect 11422 4088 11428 4100
rect 11480 4088 11486 4140
rect 11885 4131 11943 4137
rect 11885 4097 11897 4131
rect 11931 4097 11943 4131
rect 11885 4091 11943 4097
rect 12069 4131 12127 4137
rect 12069 4097 12081 4131
rect 12115 4128 12127 4131
rect 12912 4128 12940 4159
rect 12986 4156 12992 4208
rect 13044 4156 13050 4208
rect 13354 4156 13360 4208
rect 13412 4196 13418 4208
rect 14093 4199 14151 4205
rect 14093 4196 14105 4199
rect 13412 4168 14105 4196
rect 13412 4156 13418 4168
rect 13740 4137 13768 4168
rect 14093 4165 14105 4168
rect 14139 4165 14151 4199
rect 14093 4159 14151 4165
rect 12115 4100 12940 4128
rect 13081 4131 13139 4137
rect 12115 4097 12127 4100
rect 12069 4091 12127 4097
rect 13081 4097 13093 4131
rect 13127 4128 13139 4131
rect 13725 4131 13783 4137
rect 13127 4100 13676 4128
rect 13127 4097 13139 4100
rect 13081 4091 13139 4097
rect 8628 4032 9168 4060
rect 9309 4063 9367 4069
rect 8628 4020 8634 4032
rect 9309 4029 9321 4063
rect 9355 4060 9367 4063
rect 10226 4060 10232 4072
rect 9355 4032 10232 4060
rect 9355 4029 9367 4032
rect 9309 4023 9367 4029
rect 7558 3992 7564 4004
rect 6748 3964 7564 3992
rect 6748 3933 6776 3964
rect 7558 3952 7564 3964
rect 7616 3952 7622 4004
rect 7834 3952 7840 4004
rect 7892 3992 7898 4004
rect 9324 3992 9352 4023
rect 10226 4020 10232 4032
rect 10284 4060 10290 4072
rect 10413 4063 10471 4069
rect 10413 4060 10425 4063
rect 10284 4032 10425 4060
rect 10284 4020 10290 4032
rect 10413 4029 10425 4032
rect 10459 4029 10471 4063
rect 10413 4023 10471 4029
rect 10597 4063 10655 4069
rect 10597 4029 10609 4063
rect 10643 4060 10655 4063
rect 11701 4063 11759 4069
rect 11701 4060 11713 4063
rect 10643 4032 11713 4060
rect 10643 4029 10655 4032
rect 10597 4023 10655 4029
rect 11701 4029 11713 4032
rect 11747 4029 11759 4063
rect 11900 4060 11928 4091
rect 11974 4060 11980 4072
rect 11900 4032 11980 4060
rect 11701 4023 11759 4029
rect 11974 4020 11980 4032
rect 12032 4020 12038 4072
rect 12342 4020 12348 4072
rect 12400 4020 12406 4072
rect 12621 4063 12679 4069
rect 12621 4029 12633 4063
rect 12667 4029 12679 4063
rect 12621 4023 12679 4029
rect 13449 4063 13507 4069
rect 13449 4029 13461 4063
rect 13495 4029 13507 4063
rect 13449 4023 13507 4029
rect 7892 3964 9352 3992
rect 7892 3952 7898 3964
rect 6733 3927 6791 3933
rect 6733 3893 6745 3927
rect 6779 3893 6791 3927
rect 6733 3887 6791 3893
rect 6914 3884 6920 3936
rect 6972 3884 6978 3936
rect 7469 3927 7527 3933
rect 7469 3893 7481 3927
rect 7515 3924 7527 3927
rect 7650 3924 7656 3936
rect 7515 3896 7656 3924
rect 7515 3893 7527 3896
rect 7469 3887 7527 3893
rect 7650 3884 7656 3896
rect 7708 3884 7714 3936
rect 8754 3884 8760 3936
rect 8812 3884 8818 3936
rect 10870 3884 10876 3936
rect 10928 3924 10934 3936
rect 11057 3927 11115 3933
rect 11057 3924 11069 3927
rect 10928 3896 11069 3924
rect 10928 3884 10934 3896
rect 11057 3893 11069 3896
rect 11103 3893 11115 3927
rect 12636 3924 12664 4023
rect 13354 3952 13360 4004
rect 13412 3952 13418 4004
rect 13464 3992 13492 4023
rect 13538 4020 13544 4072
rect 13596 4020 13602 4072
rect 13648 4060 13676 4100
rect 13725 4097 13737 4131
rect 13771 4097 13783 4131
rect 13725 4091 13783 4097
rect 13814 4088 13820 4140
rect 13872 4088 13878 4140
rect 13906 4088 13912 4140
rect 13964 4088 13970 4140
rect 14200 4128 14228 4236
rect 16485 4233 16497 4267
rect 16531 4264 16543 4267
rect 17034 4264 17040 4276
rect 16531 4236 17040 4264
rect 16531 4233 16543 4236
rect 16485 4227 16543 4233
rect 17034 4224 17040 4236
rect 17092 4224 17098 4276
rect 17218 4224 17224 4276
rect 17276 4264 17282 4276
rect 17681 4267 17739 4273
rect 17681 4264 17693 4267
rect 17276 4236 17693 4264
rect 17276 4224 17282 4236
rect 17681 4233 17693 4236
rect 17727 4233 17739 4267
rect 19518 4264 19524 4276
rect 17681 4227 17739 4233
rect 18340 4236 19524 4264
rect 15838 4156 15844 4208
rect 15896 4196 15902 4208
rect 16025 4199 16083 4205
rect 16025 4196 16037 4199
rect 15896 4168 16037 4196
rect 15896 4156 15902 4168
rect 16025 4165 16037 4168
rect 16071 4196 16083 4199
rect 16390 4196 16396 4208
rect 16071 4168 16396 4196
rect 16071 4165 16083 4168
rect 16025 4159 16083 4165
rect 16390 4156 16396 4168
rect 16448 4196 16454 4208
rect 18340 4205 18368 4236
rect 19518 4224 19524 4236
rect 19576 4264 19582 4276
rect 20533 4267 20591 4273
rect 20533 4264 20545 4267
rect 19576 4236 20545 4264
rect 19576 4224 19582 4236
rect 20533 4233 20545 4236
rect 20579 4233 20591 4267
rect 20533 4227 20591 4233
rect 22554 4224 22560 4276
rect 22612 4264 22618 4276
rect 22612 4236 23704 4264
rect 22612 4224 22618 4236
rect 18325 4199 18383 4205
rect 16448 4168 16804 4196
rect 16448 4156 16454 4168
rect 14369 4131 14427 4137
rect 14369 4128 14381 4131
rect 14200 4100 14381 4128
rect 14369 4097 14381 4100
rect 14415 4097 14427 4131
rect 14369 4091 14427 4097
rect 14550 4088 14556 4140
rect 14608 4088 14614 4140
rect 16301 4131 16359 4137
rect 16301 4097 16313 4131
rect 16347 4128 16359 4131
rect 16574 4128 16580 4140
rect 16347 4100 16580 4128
rect 16347 4097 16359 4100
rect 16301 4091 16359 4097
rect 16574 4088 16580 4100
rect 16632 4088 16638 4140
rect 16666 4088 16672 4140
rect 16724 4088 16730 4140
rect 16776 4128 16804 4168
rect 18325 4165 18337 4199
rect 18371 4165 18383 4199
rect 18325 4159 18383 4165
rect 18874 4156 18880 4208
rect 18932 4196 18938 4208
rect 19245 4199 19303 4205
rect 19245 4196 19257 4199
rect 18932 4168 19257 4196
rect 18932 4156 18938 4168
rect 19245 4165 19257 4168
rect 19291 4165 19303 4199
rect 19702 4196 19708 4208
rect 19245 4159 19303 4165
rect 19352 4168 19708 4196
rect 16945 4131 17003 4137
rect 16945 4128 16957 4131
rect 16776 4100 16957 4128
rect 16945 4097 16957 4100
rect 16991 4097 17003 4131
rect 16945 4091 17003 4097
rect 17313 4131 17371 4137
rect 17313 4097 17325 4131
rect 17359 4128 17371 4131
rect 17494 4128 17500 4140
rect 17359 4100 17500 4128
rect 17359 4097 17371 4100
rect 17313 4091 17371 4097
rect 17494 4088 17500 4100
rect 17552 4088 17558 4140
rect 17954 4088 17960 4140
rect 18012 4088 18018 4140
rect 18785 4131 18843 4137
rect 18785 4128 18797 4131
rect 18156 4100 18797 4128
rect 14277 4063 14335 4069
rect 14277 4060 14289 4063
rect 13648 4032 14289 4060
rect 14277 4029 14289 4032
rect 14323 4029 14335 4063
rect 14277 4023 14335 4029
rect 15746 4020 15752 4072
rect 15804 4060 15810 4072
rect 15930 4060 15936 4072
rect 15804 4032 15936 4060
rect 15804 4020 15810 4032
rect 15930 4020 15936 4032
rect 15988 4060 15994 4072
rect 16117 4063 16175 4069
rect 16117 4060 16129 4063
rect 15988 4032 16129 4060
rect 15988 4020 15994 4032
rect 16117 4029 16129 4032
rect 16163 4029 16175 4063
rect 16117 4023 16175 4029
rect 16758 4020 16764 4072
rect 16816 4060 16822 4072
rect 16853 4063 16911 4069
rect 16853 4060 16865 4063
rect 16816 4032 16865 4060
rect 16816 4020 16822 4032
rect 16853 4029 16865 4032
rect 16899 4029 16911 4063
rect 16853 4023 16911 4029
rect 17037 4063 17095 4069
rect 17037 4029 17049 4063
rect 17083 4029 17095 4063
rect 17037 4023 17095 4029
rect 17129 4063 17187 4069
rect 17129 4029 17141 4063
rect 17175 4029 17187 4063
rect 17129 4023 17187 4029
rect 17865 4063 17923 4069
rect 17865 4029 17877 4063
rect 17911 4060 17923 4063
rect 18156 4060 18184 4100
rect 18785 4097 18797 4100
rect 18831 4128 18843 4131
rect 19153 4131 19211 4137
rect 19153 4128 19165 4131
rect 18831 4100 19165 4128
rect 18831 4097 18843 4100
rect 18785 4091 18843 4097
rect 19153 4097 19165 4100
rect 19199 4128 19211 4131
rect 19352 4128 19380 4168
rect 19702 4156 19708 4168
rect 19760 4196 19766 4208
rect 23566 4196 23572 4208
rect 19760 4168 20300 4196
rect 19760 4156 19766 4168
rect 20272 4140 20300 4168
rect 23032 4168 23572 4196
rect 19199 4100 19380 4128
rect 19199 4097 19211 4100
rect 19153 4091 19211 4097
rect 19886 4088 19892 4140
rect 19944 4128 19950 4140
rect 19981 4131 20039 4137
rect 19981 4128 19993 4131
rect 19944 4100 19993 4128
rect 19944 4088 19950 4100
rect 19981 4097 19993 4100
rect 20027 4097 20039 4131
rect 19981 4091 20039 4097
rect 20073 4131 20131 4137
rect 20073 4097 20085 4131
rect 20119 4128 20131 4131
rect 20162 4128 20168 4140
rect 20119 4100 20168 4128
rect 20119 4097 20131 4100
rect 20073 4091 20131 4097
rect 20162 4088 20168 4100
rect 20220 4088 20226 4140
rect 20254 4088 20260 4140
rect 20312 4088 20318 4140
rect 20622 4088 20628 4140
rect 20680 4088 20686 4140
rect 20990 4088 20996 4140
rect 21048 4088 21054 4140
rect 23032 4137 23060 4168
rect 23566 4156 23572 4168
rect 23624 4156 23630 4208
rect 23676 4196 23704 4236
rect 25958 4224 25964 4276
rect 26016 4264 26022 4276
rect 26053 4267 26111 4273
rect 26053 4264 26065 4267
rect 26016 4236 26065 4264
rect 26016 4224 26022 4236
rect 26053 4233 26065 4236
rect 26099 4233 26111 4267
rect 26053 4227 26111 4233
rect 26234 4224 26240 4276
rect 26292 4224 26298 4276
rect 26786 4224 26792 4276
rect 26844 4264 26850 4276
rect 27433 4267 27491 4273
rect 27433 4264 27445 4267
rect 26844 4236 27445 4264
rect 26844 4224 26850 4236
rect 27433 4233 27445 4236
rect 27479 4233 27491 4267
rect 27433 4227 27491 4233
rect 26252 4196 26280 4224
rect 23676 4168 23782 4196
rect 25792 4168 26280 4196
rect 23017 4131 23075 4137
rect 23017 4097 23029 4131
rect 23063 4097 23075 4131
rect 23017 4091 23075 4097
rect 25593 4131 25651 4137
rect 25593 4097 25605 4131
rect 25639 4128 25651 4131
rect 25792 4128 25820 4168
rect 26602 4156 26608 4208
rect 26660 4196 26666 4208
rect 26697 4199 26755 4205
rect 26697 4196 26709 4199
rect 26660 4168 26709 4196
rect 26660 4156 26666 4168
rect 26697 4165 26709 4168
rect 26743 4196 26755 4199
rect 26973 4199 27031 4205
rect 26973 4196 26985 4199
rect 26743 4168 26985 4196
rect 26743 4165 26755 4168
rect 26697 4159 26755 4165
rect 26973 4165 26985 4168
rect 27019 4165 27031 4199
rect 26973 4159 27031 4165
rect 25639 4100 25820 4128
rect 25639 4097 25651 4100
rect 25593 4091 25651 4097
rect 25866 4088 25872 4140
rect 25924 4088 25930 4140
rect 25958 4088 25964 4140
rect 26016 4128 26022 4140
rect 26237 4131 26295 4137
rect 26237 4128 26249 4131
rect 26016 4100 26249 4128
rect 26016 4088 26022 4100
rect 26237 4097 26249 4100
rect 26283 4128 26295 4131
rect 27249 4131 27307 4137
rect 27249 4128 27261 4131
rect 26283 4100 27261 4128
rect 26283 4097 26295 4100
rect 26237 4091 26295 4097
rect 27249 4097 27261 4100
rect 27295 4097 27307 4131
rect 27249 4091 27307 4097
rect 27525 4131 27583 4137
rect 27525 4097 27537 4131
rect 27571 4128 27583 4131
rect 27614 4128 27620 4140
rect 27571 4100 27620 4128
rect 27571 4097 27583 4100
rect 27525 4091 27583 4097
rect 27614 4088 27620 4100
rect 27672 4088 27678 4140
rect 27706 4088 27712 4140
rect 27764 4128 27770 4140
rect 27893 4131 27951 4137
rect 27893 4128 27905 4131
rect 27764 4100 27905 4128
rect 27764 4088 27770 4100
rect 27893 4097 27905 4100
rect 27939 4097 27951 4131
rect 27893 4091 27951 4097
rect 17911 4032 18184 4060
rect 18233 4063 18291 4069
rect 17911 4029 17923 4032
rect 17865 4023 17923 4029
rect 18233 4029 18245 4063
rect 18279 4060 18291 4063
rect 18506 4060 18512 4072
rect 18279 4032 18512 4060
rect 18279 4029 18291 4032
rect 18233 4023 18291 4029
rect 13630 3992 13636 4004
rect 13464 3964 13636 3992
rect 13630 3952 13636 3964
rect 13688 3992 13694 4004
rect 14461 3995 14519 4001
rect 14461 3992 14473 3995
rect 13688 3964 14473 3992
rect 13688 3952 13694 3964
rect 14461 3961 14473 3964
rect 14507 3961 14519 3995
rect 17052 3992 17080 4023
rect 14461 3955 14519 3961
rect 16316 3964 17080 3992
rect 16316 3936 16344 3964
rect 12710 3924 12716 3936
rect 12636 3896 12716 3924
rect 11057 3887 11115 3893
rect 12710 3884 12716 3896
rect 12768 3884 12774 3936
rect 12894 3884 12900 3936
rect 12952 3924 12958 3936
rect 13265 3927 13323 3933
rect 13265 3924 13277 3927
rect 12952 3896 13277 3924
rect 12952 3884 12958 3896
rect 13265 3893 13277 3896
rect 13311 3893 13323 3927
rect 13265 3887 13323 3893
rect 15194 3884 15200 3936
rect 15252 3924 15258 3936
rect 16298 3924 16304 3936
rect 15252 3896 16304 3924
rect 15252 3884 15258 3896
rect 16298 3884 16304 3896
rect 16356 3884 16362 3936
rect 16574 3884 16580 3936
rect 16632 3924 16638 3936
rect 17144 3924 17172 4023
rect 18506 4020 18512 4032
rect 18564 4060 18570 4072
rect 18601 4063 18659 4069
rect 18601 4060 18613 4063
rect 18564 4032 18613 4060
rect 18564 4020 18570 4032
rect 18601 4029 18613 4032
rect 18647 4029 18659 4063
rect 18601 4023 18659 4029
rect 18693 4063 18751 4069
rect 18693 4029 18705 4063
rect 18739 4029 18751 4063
rect 18693 4023 18751 4029
rect 18877 4063 18935 4069
rect 18877 4029 18889 4063
rect 18923 4029 18935 4063
rect 18877 4023 18935 4029
rect 17586 3952 17592 4004
rect 17644 3992 17650 4004
rect 18708 3992 18736 4023
rect 17644 3964 18736 3992
rect 18892 3992 18920 4023
rect 19426 4020 19432 4072
rect 19484 4060 19490 4072
rect 20441 4063 20499 4069
rect 20441 4060 20453 4063
rect 19484 4032 20453 4060
rect 19484 4020 19490 4032
rect 20441 4029 20453 4032
rect 20487 4029 20499 4063
rect 20441 4023 20499 4029
rect 23290 4020 23296 4072
rect 23348 4020 23354 4072
rect 25406 4020 25412 4072
rect 25464 4020 25470 4072
rect 25685 4063 25743 4069
rect 25685 4029 25697 4063
rect 25731 4029 25743 4063
rect 25685 4023 25743 4029
rect 25777 4063 25835 4069
rect 25777 4029 25789 4063
rect 25823 4029 25835 4063
rect 25777 4023 25835 4029
rect 26421 4063 26479 4069
rect 26421 4029 26433 4063
rect 26467 4060 26479 4063
rect 26510 4060 26516 4072
rect 26467 4032 26516 4060
rect 26467 4029 26479 4032
rect 26421 4023 26479 4029
rect 20257 3995 20315 4001
rect 20257 3992 20269 3995
rect 18892 3964 20269 3992
rect 17644 3952 17650 3964
rect 16632 3896 17172 3924
rect 16632 3884 16638 3896
rect 18322 3884 18328 3936
rect 18380 3924 18386 3936
rect 18417 3927 18475 3933
rect 18417 3924 18429 3927
rect 18380 3896 18429 3924
rect 18380 3884 18386 3896
rect 18417 3893 18429 3896
rect 18463 3893 18475 3927
rect 18708 3924 18736 3964
rect 20257 3961 20269 3964
rect 20303 3961 20315 3995
rect 20257 3955 20315 3961
rect 25590 3952 25596 4004
rect 25648 3992 25654 4004
rect 25700 3992 25728 4023
rect 25648 3964 25728 3992
rect 25648 3952 25654 3964
rect 19978 3924 19984 3936
rect 18708 3896 19984 3924
rect 18417 3887 18475 3893
rect 19978 3884 19984 3896
rect 20036 3884 20042 3936
rect 20530 3884 20536 3936
rect 20588 3924 20594 3936
rect 20809 3927 20867 3933
rect 20809 3924 20821 3927
rect 20588 3896 20821 3924
rect 20588 3884 20594 3896
rect 20809 3893 20821 3896
rect 20855 3893 20867 3927
rect 20809 3887 20867 3893
rect 24765 3927 24823 3933
rect 24765 3893 24777 3927
rect 24811 3924 24823 3927
rect 25682 3924 25688 3936
rect 24811 3896 25688 3924
rect 24811 3893 24823 3896
rect 24765 3887 24823 3893
rect 25682 3884 25688 3896
rect 25740 3924 25746 3936
rect 25792 3924 25820 4023
rect 26510 4020 26516 4032
rect 26568 4060 26574 4072
rect 27065 4063 27123 4069
rect 27065 4060 27077 4063
rect 26568 4032 27077 4060
rect 26568 4020 26574 4032
rect 27065 4029 27077 4032
rect 27111 4029 27123 4063
rect 27065 4023 27123 4029
rect 27246 3952 27252 4004
rect 27304 3992 27310 4004
rect 27430 3992 27436 4004
rect 27304 3964 27436 3992
rect 27304 3952 27310 3964
rect 27430 3952 27436 3964
rect 27488 3992 27494 4004
rect 27709 3995 27767 4001
rect 27709 3992 27721 3995
rect 27488 3964 27721 3992
rect 27488 3952 27494 3964
rect 27709 3961 27721 3964
rect 27755 3961 27767 3995
rect 27709 3955 27767 3961
rect 28077 3995 28135 4001
rect 28077 3961 28089 3995
rect 28123 3992 28135 3995
rect 28166 3992 28172 4004
rect 28123 3964 28172 3992
rect 28123 3961 28135 3964
rect 28077 3955 28135 3961
rect 28166 3952 28172 3964
rect 28224 3952 28230 4004
rect 26237 3927 26295 3933
rect 26237 3924 26249 3927
rect 25740 3896 26249 3924
rect 25740 3884 25746 3896
rect 26237 3893 26249 3896
rect 26283 3924 26295 3927
rect 26973 3927 27031 3933
rect 26973 3924 26985 3927
rect 26283 3896 26985 3924
rect 26283 3893 26295 3896
rect 26237 3887 26295 3893
rect 26973 3893 26985 3896
rect 27019 3893 27031 3927
rect 26973 3887 27031 3893
rect 1104 3834 28704 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 28704 3834
rect 1104 3760 28704 3782
rect 4801 3723 4859 3729
rect 4801 3689 4813 3723
rect 4847 3720 4859 3723
rect 5810 3720 5816 3732
rect 4847 3692 5816 3720
rect 4847 3689 4859 3692
rect 4801 3683 4859 3689
rect 5810 3680 5816 3692
rect 5868 3680 5874 3732
rect 6291 3723 6349 3729
rect 6291 3689 6303 3723
rect 6337 3720 6349 3723
rect 7377 3723 7435 3729
rect 7377 3720 7389 3723
rect 6337 3692 7389 3720
rect 6337 3689 6349 3692
rect 6291 3683 6349 3689
rect 7377 3689 7389 3692
rect 7423 3689 7435 3723
rect 7377 3683 7435 3689
rect 9401 3723 9459 3729
rect 9401 3689 9413 3723
rect 9447 3720 9459 3723
rect 9582 3720 9588 3732
rect 9447 3692 9588 3720
rect 9447 3689 9459 3692
rect 9401 3683 9459 3689
rect 9582 3680 9588 3692
rect 9640 3720 9646 3732
rect 11422 3720 11428 3732
rect 9640 3692 11428 3720
rect 9640 3680 9646 3692
rect 11422 3680 11428 3692
rect 11480 3680 11486 3732
rect 11606 3680 11612 3732
rect 11664 3720 11670 3732
rect 11664 3692 13308 3720
rect 11664 3680 11670 3692
rect 7190 3612 7196 3664
rect 7248 3652 7254 3664
rect 7834 3652 7840 3664
rect 7248 3624 7840 3652
rect 7248 3612 7254 3624
rect 7834 3612 7840 3624
rect 7892 3612 7898 3664
rect 11790 3652 11796 3664
rect 11164 3624 11796 3652
rect 3326 3544 3332 3596
rect 3384 3584 3390 3596
rect 3384 3556 6592 3584
rect 3384 3544 3390 3556
rect 6564 3525 6592 3556
rect 6638 3544 6644 3596
rect 6696 3544 6702 3596
rect 7285 3587 7343 3593
rect 7285 3553 7297 3587
rect 7331 3584 7343 3587
rect 7331 3556 7788 3584
rect 7331 3553 7343 3556
rect 7285 3547 7343 3553
rect 6549 3519 6607 3525
rect 6549 3485 6561 3519
rect 6595 3485 6607 3519
rect 6549 3479 6607 3485
rect 6564 3448 6592 3479
rect 6914 3476 6920 3528
rect 6972 3516 6978 3528
rect 7561 3519 7619 3525
rect 7561 3516 7573 3519
rect 6972 3488 7573 3516
rect 6972 3476 6978 3488
rect 7561 3485 7573 3488
rect 7607 3485 7619 3519
rect 7561 3479 7619 3485
rect 7650 3476 7656 3528
rect 7708 3476 7714 3528
rect 7760 3516 7788 3556
rect 10870 3544 10876 3596
rect 10928 3544 10934 3596
rect 11164 3593 11192 3624
rect 11790 3612 11796 3624
rect 11848 3612 11854 3664
rect 13280 3652 13308 3692
rect 13722 3680 13728 3732
rect 13780 3720 13786 3732
rect 13780 3692 14688 3720
rect 13780 3680 13786 3692
rect 11900 3624 12112 3652
rect 13280 3624 13676 3652
rect 11149 3587 11207 3593
rect 11149 3553 11161 3587
rect 11195 3553 11207 3587
rect 11149 3547 11207 3553
rect 11514 3544 11520 3596
rect 11572 3544 11578 3596
rect 7929 3519 7987 3525
rect 7929 3516 7941 3519
rect 7760 3488 7941 3516
rect 7929 3485 7941 3488
rect 7975 3485 7987 3519
rect 7929 3479 7987 3485
rect 11422 3476 11428 3528
rect 11480 3476 11486 3528
rect 8202 3448 8208 3460
rect 5842 3420 6408 3448
rect 6564 3420 8208 3448
rect 5258 3340 5264 3392
rect 5316 3380 5322 3392
rect 5920 3380 5948 3420
rect 5316 3352 5948 3380
rect 6380 3380 6408 3420
rect 8202 3408 8208 3420
rect 8260 3408 8266 3460
rect 10410 3408 10416 3460
rect 10468 3448 10474 3460
rect 11900 3448 11928 3624
rect 11974 3544 11980 3596
rect 12032 3544 12038 3596
rect 12084 3584 12112 3624
rect 12618 3584 12624 3596
rect 12084 3556 12624 3584
rect 12618 3544 12624 3556
rect 12676 3584 12682 3596
rect 12676 3556 13400 3584
rect 12676 3544 12682 3556
rect 13372 3528 13400 3556
rect 13354 3476 13360 3528
rect 13412 3476 13418 3528
rect 13648 3516 13676 3624
rect 14660 3593 14688 3692
rect 15470 3680 15476 3732
rect 15528 3720 15534 3732
rect 16945 3723 17003 3729
rect 16945 3720 16957 3723
rect 15528 3692 16957 3720
rect 15528 3680 15534 3692
rect 16945 3689 16957 3692
rect 16991 3720 17003 3723
rect 17129 3723 17187 3729
rect 17129 3720 17141 3723
rect 16991 3692 17141 3720
rect 16991 3689 17003 3692
rect 16945 3683 17003 3689
rect 17129 3689 17141 3692
rect 17175 3689 17187 3723
rect 17129 3683 17187 3689
rect 17497 3723 17555 3729
rect 17497 3689 17509 3723
rect 17543 3720 17555 3723
rect 17586 3720 17592 3732
rect 17543 3692 17592 3720
rect 17543 3689 17555 3692
rect 17497 3683 17555 3689
rect 17586 3680 17592 3692
rect 17644 3680 17650 3732
rect 17954 3680 17960 3732
rect 18012 3720 18018 3732
rect 18601 3723 18659 3729
rect 18601 3720 18613 3723
rect 18012 3692 18613 3720
rect 18012 3680 18018 3692
rect 18601 3689 18613 3692
rect 18647 3689 18659 3723
rect 18601 3683 18659 3689
rect 19242 3680 19248 3732
rect 19300 3680 19306 3732
rect 19794 3680 19800 3732
rect 19852 3720 19858 3732
rect 20165 3723 20223 3729
rect 20165 3720 20177 3723
rect 19852 3692 20177 3720
rect 19852 3680 19858 3692
rect 20165 3689 20177 3692
rect 20211 3720 20223 3723
rect 20622 3720 20628 3732
rect 20211 3692 20628 3720
rect 20211 3689 20223 3692
rect 20165 3683 20223 3689
rect 20622 3680 20628 3692
rect 20680 3680 20686 3732
rect 23109 3723 23167 3729
rect 23109 3689 23121 3723
rect 23155 3689 23167 3723
rect 23109 3683 23167 3689
rect 23569 3723 23627 3729
rect 23569 3689 23581 3723
rect 23615 3720 23627 3723
rect 23615 3692 26096 3720
rect 23615 3689 23627 3692
rect 23569 3683 23627 3689
rect 16206 3652 16212 3664
rect 15120 3624 16212 3652
rect 14645 3587 14703 3593
rect 14645 3553 14657 3587
rect 14691 3553 14703 3587
rect 14645 3547 14703 3553
rect 15120 3516 15148 3624
rect 16206 3612 16212 3624
rect 16264 3612 16270 3664
rect 17034 3612 17040 3664
rect 17092 3652 17098 3664
rect 17604 3652 17632 3680
rect 20990 3652 20996 3664
rect 17092 3624 17908 3652
rect 17092 3612 17098 3624
rect 17773 3587 17831 3593
rect 17773 3584 17785 3587
rect 15396 3556 17785 3584
rect 13648 3488 15148 3516
rect 15194 3476 15200 3528
rect 15252 3476 15258 3528
rect 15396 3525 15424 3556
rect 17773 3553 17785 3556
rect 17819 3553 17831 3587
rect 17773 3547 17831 3553
rect 15381 3519 15439 3525
rect 15381 3485 15393 3519
rect 15427 3485 15439 3519
rect 15381 3479 15439 3485
rect 15470 3476 15476 3528
rect 15528 3476 15534 3528
rect 15933 3519 15991 3525
rect 15933 3516 15945 3519
rect 15580 3488 15945 3516
rect 10468 3420 11928 3448
rect 10468 3408 10474 3420
rect 12250 3408 12256 3460
rect 12308 3408 12314 3460
rect 15013 3451 15071 3457
rect 15013 3417 15025 3451
rect 15059 3448 15071 3451
rect 15580 3448 15608 3488
rect 15933 3485 15945 3488
rect 15979 3485 15991 3519
rect 15933 3479 15991 3485
rect 15059 3420 15608 3448
rect 15657 3451 15715 3457
rect 15059 3417 15071 3420
rect 15013 3411 15071 3417
rect 15657 3417 15669 3451
rect 15703 3448 15715 3451
rect 15948 3448 15976 3479
rect 16022 3476 16028 3528
rect 16080 3516 16086 3528
rect 16574 3516 16580 3528
rect 16080 3488 16580 3516
rect 16080 3476 16086 3488
rect 16574 3476 16580 3488
rect 16632 3476 16638 3528
rect 16942 3476 16948 3528
rect 17000 3516 17006 3528
rect 17037 3519 17095 3525
rect 17037 3516 17049 3519
rect 17000 3488 17049 3516
rect 17000 3476 17006 3488
rect 17037 3485 17049 3488
rect 17083 3485 17095 3519
rect 17037 3479 17095 3485
rect 17313 3519 17371 3525
rect 17313 3485 17325 3519
rect 17359 3485 17371 3519
rect 17313 3479 17371 3485
rect 15703 3420 15884 3448
rect 15948 3420 16620 3448
rect 15703 3417 15715 3420
rect 15657 3411 15715 3417
rect 10502 3380 10508 3392
rect 6380 3352 10508 3380
rect 5316 3340 5322 3352
rect 10502 3340 10508 3352
rect 10560 3340 10566 3392
rect 11793 3383 11851 3389
rect 11793 3349 11805 3383
rect 11839 3380 11851 3383
rect 12986 3380 12992 3392
rect 11839 3352 12992 3380
rect 11839 3349 11851 3352
rect 11793 3343 11851 3349
rect 12986 3340 12992 3352
rect 13044 3380 13050 3392
rect 13538 3380 13544 3392
rect 13044 3352 13544 3380
rect 13044 3340 13050 3352
rect 13538 3340 13544 3352
rect 13596 3340 13602 3392
rect 14090 3340 14096 3392
rect 14148 3340 14154 3392
rect 15746 3340 15752 3392
rect 15804 3340 15810 3392
rect 15856 3380 15884 3420
rect 16022 3380 16028 3392
rect 15856 3352 16028 3380
rect 16022 3340 16028 3352
rect 16080 3340 16086 3392
rect 16114 3340 16120 3392
rect 16172 3380 16178 3392
rect 16592 3389 16620 3420
rect 16850 3408 16856 3460
rect 16908 3448 16914 3460
rect 17126 3448 17132 3460
rect 16908 3420 17132 3448
rect 16908 3408 16914 3420
rect 17126 3408 17132 3420
rect 17184 3448 17190 3460
rect 17328 3448 17356 3479
rect 17402 3476 17408 3528
rect 17460 3516 17466 3528
rect 17880 3525 17908 3624
rect 19076 3624 20996 3652
rect 19076 3593 19104 3624
rect 20990 3612 20996 3624
rect 21048 3612 21054 3664
rect 19061 3587 19119 3593
rect 19061 3553 19073 3587
rect 19107 3553 19119 3587
rect 19061 3547 19119 3553
rect 19702 3544 19708 3596
rect 19760 3544 19766 3596
rect 19794 3544 19800 3596
rect 19852 3544 19858 3596
rect 21542 3544 21548 3596
rect 21600 3584 21606 3596
rect 23124 3584 23152 3683
rect 25314 3612 25320 3664
rect 25372 3652 25378 3664
rect 25685 3655 25743 3661
rect 25685 3652 25697 3655
rect 25372 3624 25697 3652
rect 25372 3612 25378 3624
rect 25685 3621 25697 3624
rect 25731 3652 25743 3655
rect 25958 3652 25964 3664
rect 25731 3624 25964 3652
rect 25731 3621 25743 3624
rect 25685 3615 25743 3621
rect 25958 3612 25964 3624
rect 26016 3612 26022 3664
rect 26068 3652 26096 3692
rect 26326 3680 26332 3732
rect 26384 3720 26390 3732
rect 26421 3723 26479 3729
rect 26421 3720 26433 3723
rect 26384 3692 26433 3720
rect 26384 3680 26390 3692
rect 26421 3689 26433 3692
rect 26467 3689 26479 3723
rect 26421 3683 26479 3689
rect 26510 3680 26516 3732
rect 26568 3680 26574 3732
rect 26878 3652 26884 3664
rect 26068 3624 26884 3652
rect 26878 3612 26884 3624
rect 26936 3612 26942 3664
rect 21600 3556 23152 3584
rect 21600 3544 21606 3556
rect 23566 3544 23572 3596
rect 23624 3584 23630 3596
rect 28258 3584 28264 3596
rect 23624 3556 28264 3584
rect 23624 3544 23630 3556
rect 28258 3544 28264 3556
rect 28316 3544 28322 3596
rect 17589 3519 17647 3525
rect 17589 3516 17601 3519
rect 17460 3488 17601 3516
rect 17460 3476 17466 3488
rect 17589 3485 17601 3488
rect 17635 3516 17647 3519
rect 17681 3519 17739 3525
rect 17681 3516 17693 3519
rect 17635 3488 17693 3516
rect 17635 3485 17647 3488
rect 17589 3479 17647 3485
rect 17681 3485 17693 3488
rect 17727 3485 17739 3519
rect 17681 3479 17739 3485
rect 17865 3519 17923 3525
rect 17865 3485 17877 3519
rect 17911 3485 17923 3519
rect 17865 3479 17923 3485
rect 18785 3519 18843 3525
rect 18785 3485 18797 3519
rect 18831 3485 18843 3519
rect 18785 3479 18843 3485
rect 18969 3519 19027 3525
rect 18969 3485 18981 3519
rect 19015 3516 19027 3519
rect 20162 3516 20168 3528
rect 19015 3488 20168 3516
rect 19015 3485 19027 3488
rect 18969 3479 19027 3485
rect 17184 3420 17356 3448
rect 17184 3408 17190 3420
rect 16393 3383 16451 3389
rect 16393 3380 16405 3383
rect 16172 3352 16405 3380
rect 16172 3340 16178 3352
rect 16393 3349 16405 3352
rect 16439 3349 16451 3383
rect 16393 3343 16451 3349
rect 16577 3383 16635 3389
rect 16577 3349 16589 3383
rect 16623 3349 16635 3383
rect 16577 3343 16635 3349
rect 16942 3340 16948 3392
rect 17000 3380 17006 3392
rect 17420 3380 17448 3476
rect 18800 3448 18828 3479
rect 20162 3476 20168 3488
rect 20220 3476 20226 3528
rect 20530 3476 20536 3528
rect 20588 3476 20594 3528
rect 21266 3476 21272 3528
rect 21324 3476 21330 3528
rect 22830 3476 22836 3528
rect 22888 3516 22894 3528
rect 23290 3516 23296 3528
rect 22888 3488 23296 3516
rect 22888 3476 22894 3488
rect 23290 3476 23296 3488
rect 23348 3476 23354 3528
rect 23382 3476 23388 3528
rect 23440 3476 23446 3528
rect 25314 3476 25320 3528
rect 25372 3476 25378 3528
rect 25501 3519 25559 3525
rect 25501 3485 25513 3519
rect 25547 3516 25559 3519
rect 25547 3488 26188 3516
rect 25547 3485 25559 3488
rect 25501 3479 25559 3485
rect 19334 3448 19340 3460
rect 18800 3420 19340 3448
rect 19334 3408 19340 3420
rect 19392 3448 19398 3460
rect 19886 3448 19892 3460
rect 19392 3420 19892 3448
rect 19392 3408 19398 3420
rect 19886 3408 19892 3420
rect 19944 3408 19950 3460
rect 21542 3408 21548 3460
rect 21600 3408 21606 3460
rect 22554 3408 22560 3460
rect 22612 3408 22618 3460
rect 23109 3451 23167 3457
rect 23109 3417 23121 3451
rect 23155 3448 23167 3451
rect 23934 3448 23940 3460
rect 23155 3420 23940 3448
rect 23155 3417 23167 3420
rect 23109 3411 23167 3417
rect 23934 3408 23940 3420
rect 23992 3408 23998 3460
rect 24857 3451 24915 3457
rect 24857 3417 24869 3451
rect 24903 3417 24915 3451
rect 24857 3411 24915 3417
rect 25409 3451 25467 3457
rect 25409 3417 25421 3451
rect 25455 3448 25467 3451
rect 25590 3448 25596 3460
rect 25455 3420 25596 3448
rect 25455 3417 25467 3420
rect 25409 3411 25467 3417
rect 17000 3352 17448 3380
rect 17000 3340 17006 3352
rect 19426 3340 19432 3392
rect 19484 3380 19490 3392
rect 19613 3383 19671 3389
rect 19613 3380 19625 3383
rect 19484 3352 19625 3380
rect 19484 3340 19490 3352
rect 19613 3349 19625 3352
rect 19659 3349 19671 3383
rect 19613 3343 19671 3349
rect 23017 3383 23075 3389
rect 23017 3349 23029 3383
rect 23063 3380 23075 3383
rect 24302 3380 24308 3392
rect 23063 3352 24308 3380
rect 23063 3349 23075 3352
rect 23017 3343 23075 3349
rect 24302 3340 24308 3352
rect 24360 3340 24366 3392
rect 24394 3340 24400 3392
rect 24452 3380 24458 3392
rect 24581 3383 24639 3389
rect 24581 3380 24593 3383
rect 24452 3352 24593 3380
rect 24452 3340 24458 3352
rect 24581 3349 24593 3352
rect 24627 3349 24639 3383
rect 24872 3380 24900 3411
rect 25590 3408 25596 3420
rect 25648 3408 25654 3460
rect 25682 3408 25688 3460
rect 25740 3408 25746 3460
rect 26160 3457 26188 3488
rect 26234 3476 26240 3528
rect 26292 3476 26298 3528
rect 26145 3451 26203 3457
rect 26145 3417 26157 3451
rect 26191 3448 26203 3451
rect 26510 3448 26516 3460
rect 26191 3420 26516 3448
rect 26191 3417 26203 3420
rect 26145 3411 26203 3417
rect 26510 3408 26516 3420
rect 26568 3408 26574 3460
rect 27430 3408 27436 3460
rect 27488 3408 27494 3460
rect 27890 3408 27896 3460
rect 27948 3448 27954 3460
rect 27985 3451 28043 3457
rect 27985 3448 27997 3451
rect 27948 3420 27997 3448
rect 27948 3408 27954 3420
rect 27985 3417 27997 3420
rect 28031 3417 28043 3451
rect 27985 3411 28043 3417
rect 27154 3380 27160 3392
rect 24872 3352 27160 3380
rect 24581 3343 24639 3349
rect 27154 3340 27160 3352
rect 27212 3340 27218 3392
rect 1104 3290 28704 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 28704 3290
rect 1104 3216 28704 3238
rect 5994 3136 6000 3188
rect 6052 3176 6058 3188
rect 11606 3176 11612 3188
rect 6052 3148 11612 3176
rect 6052 3136 6058 3148
rect 6638 3068 6644 3120
rect 6696 3068 6702 3120
rect 6549 3043 6607 3049
rect 6549 3009 6561 3043
rect 6595 3040 6607 3043
rect 6656 3040 6684 3068
rect 6595 3012 6684 3040
rect 6595 3009 6607 3012
rect 6549 3003 6607 3009
rect 6641 2975 6699 2981
rect 6641 2941 6653 2975
rect 6687 2972 6699 2975
rect 6840 2972 6868 3148
rect 11606 3136 11612 3148
rect 11664 3136 11670 3188
rect 12250 3136 12256 3188
rect 12308 3176 12314 3188
rect 12437 3179 12495 3185
rect 12437 3176 12449 3179
rect 12308 3148 12449 3176
rect 12308 3136 12314 3148
rect 12437 3145 12449 3148
rect 12483 3145 12495 3179
rect 12437 3139 12495 3145
rect 12894 3136 12900 3188
rect 12952 3136 12958 3188
rect 13354 3136 13360 3188
rect 13412 3136 13418 3188
rect 16390 3136 16396 3188
rect 16448 3136 16454 3188
rect 16758 3136 16764 3188
rect 16816 3136 16822 3188
rect 18966 3136 18972 3188
rect 19024 3176 19030 3188
rect 19245 3179 19303 3185
rect 19245 3176 19257 3179
rect 19024 3148 19257 3176
rect 19024 3136 19030 3148
rect 19245 3145 19257 3148
rect 19291 3145 19303 3179
rect 19245 3139 19303 3145
rect 19518 3136 19524 3188
rect 19576 3136 19582 3188
rect 23569 3179 23627 3185
rect 22480 3148 23428 3176
rect 8481 3111 8539 3117
rect 8481 3077 8493 3111
rect 8527 3108 8539 3111
rect 8754 3108 8760 3120
rect 8527 3080 8760 3108
rect 8527 3077 8539 3080
rect 8481 3071 8539 3077
rect 8754 3068 8760 3080
rect 8812 3068 8818 3120
rect 10410 3108 10416 3120
rect 9706 3080 10416 3108
rect 10410 3068 10416 3080
rect 10468 3068 10474 3120
rect 10502 3068 10508 3120
rect 10560 3108 10566 3120
rect 12805 3111 12863 3117
rect 10560 3080 12756 3108
rect 10560 3068 10566 3080
rect 8202 3000 8208 3052
rect 8260 3000 8266 3052
rect 12345 3043 12403 3049
rect 12345 3009 12357 3043
rect 12391 3009 12403 3043
rect 12728 3040 12756 3080
rect 12805 3077 12817 3111
rect 12851 3108 12863 3111
rect 14090 3108 14096 3120
rect 12851 3080 14096 3108
rect 12851 3077 12863 3080
rect 12805 3071 12863 3077
rect 14090 3068 14096 3080
rect 14148 3068 14154 3120
rect 14458 3068 14464 3120
rect 14516 3068 14522 3120
rect 16298 3068 16304 3120
rect 16356 3108 16362 3120
rect 17037 3111 17095 3117
rect 17037 3108 17049 3111
rect 16356 3080 17049 3108
rect 16356 3068 16362 3080
rect 17037 3077 17049 3080
rect 17083 3077 17095 3111
rect 20530 3108 20536 3120
rect 17037 3071 17095 3077
rect 18984 3080 20536 3108
rect 13633 3043 13691 3049
rect 13633 3040 13645 3043
rect 12728 3012 13645 3040
rect 12345 3003 12403 3009
rect 13633 3009 13645 3012
rect 13679 3009 13691 3043
rect 13633 3003 13691 3009
rect 16669 3043 16727 3049
rect 16669 3009 16681 3043
rect 16715 3040 16727 3043
rect 16758 3040 16764 3052
rect 16715 3012 16764 3040
rect 16715 3009 16727 3012
rect 16669 3003 16727 3009
rect 6687 2944 6868 2972
rect 6917 2975 6975 2981
rect 6687 2941 6699 2944
rect 6641 2935 6699 2941
rect 6917 2941 6929 2975
rect 6963 2972 6975 2975
rect 7006 2972 7012 2984
rect 6963 2944 7012 2972
rect 6963 2941 6975 2944
rect 6917 2935 6975 2941
rect 7006 2932 7012 2944
rect 7064 2932 7070 2984
rect 9858 2932 9864 2984
rect 9916 2972 9922 2984
rect 9953 2975 10011 2981
rect 9953 2972 9965 2975
rect 9916 2944 9965 2972
rect 9916 2932 9922 2944
rect 9953 2941 9965 2944
rect 9999 2941 10011 2975
rect 12360 2972 12388 3003
rect 12802 2972 12808 2984
rect 12360 2944 12808 2972
rect 9953 2935 10011 2941
rect 12802 2932 12808 2944
rect 12860 2932 12866 2984
rect 13078 2932 13084 2984
rect 13136 2932 13142 2984
rect 13648 2972 13676 3003
rect 16758 3000 16764 3012
rect 16816 3000 16822 3052
rect 16853 3043 16911 3049
rect 16853 3009 16865 3043
rect 16899 3009 16911 3043
rect 16853 3003 16911 3009
rect 14185 2975 14243 2981
rect 14185 2972 14197 2975
rect 13648 2944 14197 2972
rect 14185 2941 14197 2944
rect 14231 2941 14243 2975
rect 14185 2935 14243 2941
rect 15933 2975 15991 2981
rect 15933 2941 15945 2975
rect 15979 2972 15991 2975
rect 16868 2972 16896 3003
rect 16942 3000 16948 3052
rect 17000 3000 17006 3052
rect 17126 3000 17132 3052
rect 17184 3040 17190 3052
rect 18984 3049 19012 3080
rect 18969 3043 19027 3049
rect 18969 3040 18981 3043
rect 17184 3012 18981 3040
rect 17184 3000 17190 3012
rect 18969 3009 18981 3012
rect 19015 3009 19027 3043
rect 18969 3003 19027 3009
rect 19153 3043 19211 3049
rect 19153 3009 19165 3043
rect 19199 3040 19211 3043
rect 19334 3040 19340 3052
rect 19199 3012 19340 3040
rect 19199 3009 19211 3012
rect 19153 3003 19211 3009
rect 19334 3000 19340 3012
rect 19392 3000 19398 3052
rect 19429 3043 19487 3049
rect 19429 3009 19441 3043
rect 19475 3040 19487 3043
rect 19610 3040 19616 3052
rect 19475 3012 19616 3040
rect 19475 3009 19487 3012
rect 19429 3003 19487 3009
rect 19610 3000 19616 3012
rect 19668 3000 19674 3052
rect 19720 3049 19748 3080
rect 20530 3068 20536 3080
rect 20588 3068 20594 3120
rect 22480 3108 22508 3148
rect 22554 3108 22560 3120
rect 22480 3080 22560 3108
rect 22554 3068 22560 3080
rect 22612 3068 22618 3120
rect 23400 3108 23428 3148
rect 23569 3145 23581 3179
rect 23615 3176 23627 3179
rect 23842 3176 23848 3188
rect 23615 3148 23848 3176
rect 23615 3145 23627 3148
rect 23569 3139 23627 3145
rect 23842 3136 23848 3148
rect 23900 3136 23906 3188
rect 23952 3148 24072 3176
rect 23952 3108 23980 3148
rect 23400 3080 23980 3108
rect 24044 3108 24072 3148
rect 25314 3136 25320 3188
rect 25372 3176 25378 3188
rect 25409 3179 25467 3185
rect 25409 3176 25421 3179
rect 25372 3148 25421 3176
rect 25372 3136 25378 3148
rect 25409 3145 25421 3148
rect 25455 3145 25467 3179
rect 25409 3139 25467 3145
rect 26234 3136 26240 3188
rect 26292 3136 26298 3188
rect 26418 3136 26424 3188
rect 26476 3136 26482 3188
rect 27706 3136 27712 3188
rect 27764 3136 27770 3188
rect 24394 3108 24400 3120
rect 24044 3080 24400 3108
rect 24394 3068 24400 3080
rect 24452 3068 24458 3120
rect 26252 3108 26280 3136
rect 25792 3080 26280 3108
rect 19720 3043 19793 3049
rect 19720 3012 19747 3043
rect 19735 3009 19747 3012
rect 19781 3009 19793 3043
rect 19735 3003 19793 3009
rect 19889 3043 19947 3049
rect 19889 3009 19901 3043
rect 19935 3040 19947 3043
rect 19978 3040 19984 3052
rect 19935 3012 19984 3040
rect 19935 3009 19947 3012
rect 19889 3003 19947 3009
rect 19978 3000 19984 3012
rect 20036 3000 20042 3052
rect 21266 3000 21272 3052
rect 21324 3040 21330 3052
rect 21821 3043 21879 3049
rect 21821 3040 21833 3043
rect 21324 3012 21833 3040
rect 21324 3000 21330 3012
rect 21821 3009 21833 3012
rect 21867 3009 21879 3043
rect 21821 3003 21879 3009
rect 23566 3000 23572 3052
rect 23624 3040 23630 3052
rect 25792 3049 25820 3080
rect 28166 3068 28172 3120
rect 28224 3068 28230 3120
rect 23661 3043 23719 3049
rect 23661 3040 23673 3043
rect 23624 3012 23673 3040
rect 23624 3000 23630 3012
rect 23661 3009 23673 3012
rect 23707 3009 23719 3043
rect 23661 3003 23719 3009
rect 25777 3043 25835 3049
rect 25777 3009 25789 3043
rect 25823 3009 25835 3043
rect 25777 3003 25835 3009
rect 25869 3043 25927 3049
rect 25869 3009 25881 3043
rect 25915 3040 25927 3043
rect 25958 3040 25964 3052
rect 25915 3012 25964 3040
rect 25915 3009 25927 3012
rect 25869 3003 25927 3009
rect 25958 3000 25964 3012
rect 26016 3000 26022 3052
rect 26237 3043 26295 3049
rect 26237 3009 26249 3043
rect 26283 3009 26295 3043
rect 26237 3003 26295 3009
rect 17034 2972 17040 2984
rect 15979 2944 17040 2972
rect 15979 2941 15991 2944
rect 15933 2935 15991 2941
rect 17034 2932 17040 2944
rect 17092 2932 17098 2984
rect 12253 2907 12311 2913
rect 12253 2873 12265 2907
rect 12299 2904 12311 2907
rect 13446 2904 13452 2916
rect 12299 2876 13452 2904
rect 12299 2873 12311 2876
rect 12253 2867 12311 2873
rect 13446 2864 13452 2876
rect 13504 2864 13510 2916
rect 16301 2907 16359 2913
rect 16301 2873 16313 2907
rect 16347 2904 16359 2907
rect 17144 2904 17172 3000
rect 22097 2975 22155 2981
rect 22097 2941 22109 2975
rect 22143 2972 22155 2975
rect 22186 2972 22192 2984
rect 22143 2944 22192 2972
rect 22143 2941 22155 2944
rect 22097 2935 22155 2941
rect 22186 2932 22192 2944
rect 22244 2972 22250 2984
rect 23382 2972 23388 2984
rect 22244 2944 23388 2972
rect 22244 2932 22250 2944
rect 23382 2932 23388 2944
rect 23440 2932 23446 2984
rect 23492 2944 25636 2972
rect 16347 2876 17172 2904
rect 16347 2873 16359 2876
rect 16301 2867 16359 2873
rect 14550 2796 14556 2848
rect 14608 2836 14614 2848
rect 18322 2836 18328 2848
rect 14608 2808 18328 2836
rect 14608 2796 14614 2808
rect 18322 2796 18328 2808
rect 18380 2796 18386 2848
rect 21450 2796 21456 2848
rect 21508 2836 21514 2848
rect 23492 2836 23520 2944
rect 25608 2904 25636 2944
rect 25682 2932 25688 2984
rect 25740 2972 25746 2984
rect 26252 2972 26280 3003
rect 27522 3000 27528 3052
rect 27580 3000 27586 3052
rect 25740 2944 26280 2972
rect 25740 2932 25746 2944
rect 27614 2904 27620 2916
rect 25608 2876 27620 2904
rect 27614 2864 27620 2876
rect 27672 2904 27678 2916
rect 27893 2907 27951 2913
rect 27893 2904 27905 2907
rect 27672 2876 27905 2904
rect 27672 2864 27678 2876
rect 27893 2873 27905 2876
rect 27939 2873 27951 2907
rect 27893 2867 27951 2873
rect 23934 2845 23940 2848
rect 21508 2808 23520 2836
rect 23924 2839 23940 2845
rect 21508 2796 21514 2808
rect 23924 2805 23936 2839
rect 23924 2799 23940 2805
rect 23934 2796 23940 2799
rect 23992 2796 23998 2848
rect 26237 2839 26295 2845
rect 26237 2805 26249 2839
rect 26283 2836 26295 2839
rect 26510 2836 26516 2848
rect 26283 2808 26516 2836
rect 26283 2805 26295 2808
rect 26237 2799 26295 2805
rect 26510 2796 26516 2808
rect 26568 2796 26574 2848
rect 1104 2746 28704 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 28704 2746
rect 1104 2672 28704 2694
rect 21542 2592 21548 2644
rect 21600 2592 21606 2644
rect 22186 2592 22192 2644
rect 22244 2592 22250 2644
rect 22830 2592 22836 2644
rect 22888 2592 22894 2644
rect 23477 2635 23535 2641
rect 23477 2601 23489 2635
rect 23523 2632 23535 2635
rect 23934 2632 23940 2644
rect 23523 2604 23940 2632
rect 23523 2601 23535 2604
rect 23477 2595 23535 2601
rect 23934 2592 23940 2604
rect 23992 2592 23998 2644
rect 21266 2388 21272 2440
rect 21324 2428 21330 2440
rect 21361 2431 21419 2437
rect 21361 2428 21373 2431
rect 21324 2400 21373 2428
rect 21324 2388 21330 2400
rect 21361 2397 21373 2400
rect 21407 2397 21419 2431
rect 21361 2391 21419 2397
rect 21910 2388 21916 2440
rect 21968 2428 21974 2440
rect 22005 2431 22063 2437
rect 22005 2428 22017 2431
rect 21968 2400 22017 2428
rect 21968 2388 21974 2400
rect 22005 2397 22017 2400
rect 22051 2397 22063 2431
rect 22005 2391 22063 2397
rect 22554 2388 22560 2440
rect 22612 2428 22618 2440
rect 22649 2431 22707 2437
rect 22649 2428 22661 2431
rect 22612 2400 22661 2428
rect 22612 2388 22618 2400
rect 22649 2397 22661 2400
rect 22695 2397 22707 2431
rect 22649 2391 22707 2397
rect 23198 2388 23204 2440
rect 23256 2428 23262 2440
rect 23293 2431 23351 2437
rect 23293 2428 23305 2431
rect 23256 2400 23305 2428
rect 23256 2388 23262 2400
rect 23293 2397 23305 2400
rect 23339 2397 23351 2431
rect 23293 2391 23351 2397
rect 1104 2202 28704 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 28704 2202
rect 1104 2128 28704 2150
<< via1 >>
rect 4874 29350 4926 29402
rect 4938 29350 4990 29402
rect 5002 29350 5054 29402
rect 5066 29350 5118 29402
rect 5130 29350 5182 29402
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 4874 28262 4926 28314
rect 4938 28262 4990 28314
rect 5002 28262 5054 28314
rect 5066 28262 5118 28314
rect 5130 28262 5182 28314
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 4874 27174 4926 27226
rect 4938 27174 4990 27226
rect 5002 27174 5054 27226
rect 5066 27174 5118 27226
rect 5130 27174 5182 27226
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 4874 26086 4926 26138
rect 4938 26086 4990 26138
rect 5002 26086 5054 26138
rect 5066 26086 5118 26138
rect 5130 26086 5182 26138
rect 7840 25848 7892 25900
rect 8576 25848 8628 25900
rect 17776 25916 17828 25968
rect 22836 25916 22888 25968
rect 9588 25891 9640 25900
rect 9588 25857 9597 25891
rect 9597 25857 9631 25891
rect 9631 25857 9640 25891
rect 9588 25848 9640 25857
rect 10324 25848 10376 25900
rect 15292 25891 15344 25900
rect 15292 25857 15301 25891
rect 15301 25857 15335 25891
rect 15335 25857 15344 25891
rect 15292 25848 15344 25857
rect 17684 25848 17736 25900
rect 8944 25780 8996 25832
rect 11980 25780 12032 25832
rect 16948 25780 17000 25832
rect 21180 25823 21232 25832
rect 21180 25789 21189 25823
rect 21189 25789 21223 25823
rect 21223 25789 21232 25823
rect 21180 25780 21232 25789
rect 23296 25823 23348 25832
rect 23296 25789 23305 25823
rect 23305 25789 23339 25823
rect 23339 25789 23348 25823
rect 23296 25780 23348 25789
rect 24032 25823 24084 25832
rect 24032 25789 24041 25823
rect 24041 25789 24075 25823
rect 24075 25789 24084 25823
rect 24032 25780 24084 25789
rect 24308 25823 24360 25832
rect 24308 25789 24317 25823
rect 24317 25789 24351 25823
rect 24351 25789 24360 25823
rect 24308 25780 24360 25789
rect 21456 25712 21508 25764
rect 5540 25687 5592 25696
rect 5540 25653 5549 25687
rect 5549 25653 5583 25687
rect 5583 25653 5592 25687
rect 5540 25644 5592 25653
rect 8392 25687 8444 25696
rect 8392 25653 8401 25687
rect 8401 25653 8435 25687
rect 8435 25653 8444 25687
rect 8392 25644 8444 25653
rect 9772 25687 9824 25696
rect 9772 25653 9781 25687
rect 9781 25653 9815 25687
rect 9815 25653 9824 25687
rect 9772 25644 9824 25653
rect 11060 25644 11112 25696
rect 15476 25644 15528 25696
rect 19524 25644 19576 25696
rect 22928 25644 22980 25696
rect 25780 25687 25832 25696
rect 25780 25653 25789 25687
rect 25789 25653 25823 25687
rect 25823 25653 25832 25687
rect 25780 25644 25832 25653
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 8576 25483 8628 25492
rect 8576 25449 8585 25483
rect 8585 25449 8619 25483
rect 8619 25449 8628 25483
rect 8576 25440 8628 25449
rect 8944 25483 8996 25492
rect 8944 25449 8953 25483
rect 8953 25449 8987 25483
rect 8987 25449 8996 25483
rect 8944 25440 8996 25449
rect 5448 25304 5500 25356
rect 8392 25347 8444 25356
rect 8392 25313 8401 25347
rect 8401 25313 8435 25347
rect 8435 25313 8444 25347
rect 8392 25304 8444 25313
rect 9956 25372 10008 25424
rect 11980 25440 12032 25492
rect 21180 25440 21232 25492
rect 21548 25440 21600 25492
rect 24308 25440 24360 25492
rect 12992 25372 13044 25424
rect 4712 25236 4764 25288
rect 7840 25236 7892 25288
rect 15476 25347 15528 25356
rect 15476 25313 15485 25347
rect 15485 25313 15519 25347
rect 15519 25313 15528 25347
rect 15476 25304 15528 25313
rect 19524 25347 19576 25356
rect 19524 25313 19533 25347
rect 19533 25313 19567 25347
rect 19567 25313 19576 25347
rect 19524 25304 19576 25313
rect 8760 25279 8812 25288
rect 8760 25245 8769 25279
rect 8769 25245 8803 25279
rect 8803 25245 8812 25279
rect 8760 25236 8812 25245
rect 9588 25236 9640 25288
rect 5540 25168 5592 25220
rect 5908 25168 5960 25220
rect 10692 25279 10744 25288
rect 10692 25245 10701 25279
rect 10701 25245 10735 25279
rect 10735 25245 10744 25279
rect 10692 25236 10744 25245
rect 6920 25143 6972 25152
rect 6920 25109 6929 25143
rect 6929 25109 6963 25143
rect 6963 25109 6972 25143
rect 6920 25100 6972 25109
rect 7196 25100 7248 25152
rect 9680 25143 9732 25152
rect 9680 25109 9689 25143
rect 9689 25109 9723 25143
rect 9723 25109 9732 25143
rect 9680 25100 9732 25109
rect 9864 25100 9916 25152
rect 10416 25143 10468 25152
rect 10968 25211 11020 25220
rect 10968 25177 10977 25211
rect 10977 25177 11011 25211
rect 11011 25177 11020 25211
rect 10968 25168 11020 25177
rect 12624 25168 12676 25220
rect 13820 25279 13872 25288
rect 13820 25245 13829 25279
rect 13829 25245 13863 25279
rect 13863 25245 13872 25279
rect 13820 25236 13872 25245
rect 14372 25236 14424 25288
rect 15200 25279 15252 25288
rect 15200 25245 15209 25279
rect 15209 25245 15243 25279
rect 15243 25245 15252 25279
rect 15200 25236 15252 25245
rect 17592 25236 17644 25288
rect 19248 25279 19300 25288
rect 19248 25245 19257 25279
rect 19257 25245 19291 25279
rect 19291 25245 19300 25279
rect 19248 25236 19300 25245
rect 21272 25279 21324 25288
rect 21272 25245 21281 25279
rect 21281 25245 21315 25279
rect 21315 25245 21324 25279
rect 21272 25236 21324 25245
rect 22100 25279 22152 25288
rect 22100 25245 22109 25279
rect 22109 25245 22143 25279
rect 22143 25245 22152 25279
rect 22100 25236 22152 25245
rect 22928 25279 22980 25288
rect 22928 25245 22937 25279
rect 22937 25245 22971 25279
rect 22971 25245 22980 25279
rect 23756 25347 23808 25356
rect 23756 25313 23765 25347
rect 23765 25313 23799 25347
rect 23799 25313 23808 25347
rect 23756 25304 23808 25313
rect 24860 25304 24912 25356
rect 22928 25236 22980 25245
rect 26148 25279 26200 25288
rect 26148 25245 26157 25279
rect 26157 25245 26191 25279
rect 26191 25245 26200 25279
rect 26148 25236 26200 25245
rect 26332 25279 26384 25288
rect 26332 25245 26341 25279
rect 26341 25245 26375 25279
rect 26375 25245 26384 25279
rect 26332 25236 26384 25245
rect 27160 25279 27212 25288
rect 27160 25245 27169 25279
rect 27169 25245 27203 25279
rect 27203 25245 27212 25279
rect 27160 25236 27212 25245
rect 13636 25168 13688 25220
rect 16028 25168 16080 25220
rect 20536 25168 20588 25220
rect 10416 25109 10441 25143
rect 10441 25109 10468 25143
rect 10416 25100 10468 25109
rect 12532 25143 12584 25152
rect 12532 25109 12541 25143
rect 12541 25109 12575 25143
rect 12575 25109 12584 25143
rect 12532 25100 12584 25109
rect 14556 25100 14608 25152
rect 16948 25143 17000 25152
rect 16948 25109 16957 25143
rect 16957 25109 16991 25143
rect 16991 25109 17000 25143
rect 16948 25100 17000 25109
rect 21364 25143 21416 25152
rect 21364 25109 21373 25143
rect 21373 25109 21407 25143
rect 21407 25109 21416 25143
rect 21364 25100 21416 25109
rect 23020 25100 23072 25152
rect 25136 25100 25188 25152
rect 27804 25100 27856 25152
rect 4874 24998 4926 25050
rect 4938 24998 4990 25050
rect 5002 24998 5054 25050
rect 5066 24998 5118 25050
rect 5130 24998 5182 25050
rect 7840 24939 7892 24948
rect 7840 24905 7849 24939
rect 7849 24905 7883 24939
rect 7883 24905 7892 24939
rect 7840 24896 7892 24905
rect 10968 24896 11020 24948
rect 4712 24871 4764 24880
rect 4712 24837 4721 24871
rect 4721 24837 4755 24871
rect 4755 24837 4764 24871
rect 4712 24828 4764 24837
rect 6920 24828 6972 24880
rect 10324 24871 10376 24880
rect 10324 24837 10333 24871
rect 10333 24837 10367 24871
rect 10367 24837 10376 24871
rect 10324 24828 10376 24837
rect 13360 24828 13412 24880
rect 4804 24692 4856 24744
rect 5908 24692 5960 24744
rect 10048 24803 10100 24812
rect 10048 24769 10057 24803
rect 10057 24769 10091 24803
rect 10091 24769 10100 24803
rect 10048 24760 10100 24769
rect 10416 24760 10468 24812
rect 11520 24803 11572 24812
rect 11520 24769 11529 24803
rect 11529 24769 11563 24803
rect 11563 24769 11572 24803
rect 11520 24760 11572 24769
rect 9588 24735 9640 24744
rect 9588 24701 9597 24735
rect 9597 24701 9631 24735
rect 9631 24701 9640 24735
rect 9588 24692 9640 24701
rect 11060 24692 11112 24744
rect 9680 24624 9732 24676
rect 9956 24624 10008 24676
rect 5448 24556 5500 24608
rect 9128 24556 9180 24608
rect 9864 24599 9916 24608
rect 9864 24565 9873 24599
rect 9873 24565 9907 24599
rect 9907 24565 9916 24599
rect 9864 24556 9916 24565
rect 10968 24556 11020 24608
rect 13452 24760 13504 24812
rect 13820 24803 13872 24812
rect 13820 24769 13829 24803
rect 13829 24769 13863 24803
rect 13863 24769 13872 24803
rect 13820 24760 13872 24769
rect 11796 24735 11848 24744
rect 11796 24701 11805 24735
rect 11805 24701 11839 24735
rect 11839 24701 11848 24735
rect 11796 24692 11848 24701
rect 12532 24692 12584 24744
rect 13084 24692 13136 24744
rect 14096 24803 14148 24812
rect 14096 24769 14105 24803
rect 14105 24769 14139 24803
rect 14139 24769 14148 24803
rect 14096 24760 14148 24769
rect 14188 24803 14240 24812
rect 14188 24769 14197 24803
rect 14197 24769 14231 24803
rect 14231 24769 14240 24803
rect 14188 24760 14240 24769
rect 15384 24896 15436 24948
rect 16028 24828 16080 24880
rect 17868 24896 17920 24948
rect 22100 24896 22152 24948
rect 23296 24896 23348 24948
rect 23756 24896 23808 24948
rect 17776 24871 17828 24880
rect 17776 24837 17785 24871
rect 17785 24837 17819 24871
rect 17819 24837 17828 24871
rect 17776 24828 17828 24837
rect 16212 24760 16264 24812
rect 16764 24760 16816 24812
rect 17040 24760 17092 24812
rect 13636 24667 13688 24676
rect 13636 24633 13645 24667
rect 13645 24633 13679 24667
rect 13679 24633 13688 24667
rect 13636 24624 13688 24633
rect 14372 24667 14424 24676
rect 14372 24633 14381 24667
rect 14381 24633 14415 24667
rect 14415 24633 14424 24667
rect 14372 24624 14424 24633
rect 12808 24556 12860 24608
rect 13820 24556 13872 24608
rect 16304 24624 16356 24676
rect 17132 24692 17184 24744
rect 19248 24760 19300 24812
rect 22468 24760 22520 24812
rect 15200 24556 15252 24608
rect 15384 24556 15436 24608
rect 16856 24556 16908 24608
rect 17408 24556 17460 24608
rect 19156 24735 19208 24744
rect 19156 24701 19165 24735
rect 19165 24701 19199 24735
rect 19199 24701 19208 24735
rect 19156 24692 19208 24701
rect 21364 24692 21416 24744
rect 22284 24692 22336 24744
rect 17684 24624 17736 24676
rect 21548 24624 21600 24676
rect 17868 24556 17920 24608
rect 21732 24556 21784 24608
rect 22008 24624 22060 24676
rect 23020 24803 23072 24812
rect 23020 24769 23029 24803
rect 23029 24769 23063 24803
rect 23063 24769 23072 24803
rect 23020 24760 23072 24769
rect 25688 24828 25740 24880
rect 26424 24896 26476 24948
rect 27160 24896 27212 24948
rect 24860 24760 24912 24812
rect 25136 24803 25188 24812
rect 25136 24769 25145 24803
rect 25145 24769 25179 24803
rect 25179 24769 25188 24803
rect 25136 24760 25188 24769
rect 26976 24803 27028 24812
rect 26976 24769 26985 24803
rect 26985 24769 27019 24803
rect 27019 24769 27028 24803
rect 26976 24760 27028 24769
rect 27160 24803 27212 24812
rect 27160 24769 27169 24803
rect 27169 24769 27203 24803
rect 27203 24769 27212 24803
rect 27160 24760 27212 24769
rect 27896 24760 27948 24812
rect 25780 24556 25832 24608
rect 26332 24667 26384 24676
rect 26332 24633 26341 24667
rect 26341 24633 26375 24667
rect 26375 24633 26384 24667
rect 26332 24624 26384 24633
rect 26792 24556 26844 24608
rect 27988 24556 28040 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 8760 24352 8812 24404
rect 10416 24352 10468 24404
rect 11060 24352 11112 24404
rect 13820 24352 13872 24404
rect 14096 24352 14148 24404
rect 15292 24352 15344 24404
rect 16212 24352 16264 24404
rect 16948 24352 17000 24404
rect 12808 24327 12860 24336
rect 12808 24293 12817 24327
rect 12817 24293 12851 24327
rect 12851 24293 12860 24327
rect 12808 24284 12860 24293
rect 15844 24284 15896 24336
rect 5448 24216 5500 24268
rect 6920 24259 6972 24268
rect 6920 24225 6929 24259
rect 6929 24225 6963 24259
rect 6963 24225 6972 24259
rect 6920 24216 6972 24225
rect 9588 24216 9640 24268
rect 10692 24216 10744 24268
rect 11796 24216 11848 24268
rect 13084 24216 13136 24268
rect 13268 24216 13320 24268
rect 15200 24216 15252 24268
rect 16028 24259 16080 24268
rect 16028 24225 16037 24259
rect 16037 24225 16071 24259
rect 16071 24225 16080 24259
rect 17040 24284 17092 24336
rect 16028 24216 16080 24225
rect 7196 24123 7248 24132
rect 7196 24089 7205 24123
rect 7205 24089 7239 24123
rect 7239 24089 7248 24123
rect 7196 24080 7248 24089
rect 5908 24012 5960 24064
rect 9220 24123 9272 24132
rect 9220 24089 9229 24123
rect 9229 24089 9263 24123
rect 9263 24089 9272 24123
rect 9220 24080 9272 24089
rect 11244 24123 11296 24132
rect 11244 24089 11253 24123
rect 11253 24089 11287 24123
rect 11287 24089 11296 24123
rect 11244 24080 11296 24089
rect 11704 24080 11756 24132
rect 11612 24012 11664 24064
rect 12992 24123 13044 24132
rect 12992 24089 13019 24123
rect 13019 24089 13044 24123
rect 12992 24080 13044 24089
rect 15660 24148 15712 24200
rect 16212 24148 16264 24200
rect 17408 24352 17460 24404
rect 19156 24352 19208 24404
rect 21272 24352 21324 24404
rect 26976 24352 27028 24404
rect 21456 24284 21508 24336
rect 22008 24284 22060 24336
rect 26240 24284 26292 24336
rect 17592 24216 17644 24268
rect 19524 24216 19576 24268
rect 21180 24216 21232 24268
rect 24032 24216 24084 24268
rect 20168 24148 20220 24200
rect 14556 24123 14608 24132
rect 14556 24089 14565 24123
rect 14565 24089 14599 24123
rect 14599 24089 14608 24123
rect 14556 24080 14608 24089
rect 13360 24012 13412 24064
rect 16304 24123 16356 24132
rect 16304 24089 16313 24123
rect 16313 24089 16347 24123
rect 16347 24089 16356 24123
rect 16304 24080 16356 24089
rect 18052 24080 18104 24132
rect 21088 24191 21140 24200
rect 21088 24157 21097 24191
rect 21097 24157 21131 24191
rect 21131 24157 21140 24191
rect 21088 24148 21140 24157
rect 19432 24012 19484 24064
rect 19616 24055 19668 24064
rect 19616 24021 19625 24055
rect 19625 24021 19659 24055
rect 19659 24021 19668 24055
rect 19616 24012 19668 24021
rect 19708 24055 19760 24064
rect 19708 24021 19717 24055
rect 19717 24021 19751 24055
rect 19751 24021 19760 24055
rect 21272 24080 21324 24132
rect 21456 24191 21508 24200
rect 21456 24157 21465 24191
rect 21465 24157 21499 24191
rect 21499 24157 21508 24191
rect 21456 24148 21508 24157
rect 21548 24191 21600 24200
rect 21548 24157 21557 24191
rect 21557 24157 21591 24191
rect 21591 24157 21600 24191
rect 21548 24148 21600 24157
rect 21732 24191 21784 24200
rect 21732 24157 21741 24191
rect 21741 24157 21775 24191
rect 21775 24157 21784 24191
rect 21732 24148 21784 24157
rect 22284 24191 22336 24200
rect 22284 24157 22293 24191
rect 22293 24157 22327 24191
rect 22327 24157 22336 24191
rect 22284 24148 22336 24157
rect 25596 24216 25648 24268
rect 26516 24259 26568 24268
rect 26516 24225 26525 24259
rect 26525 24225 26559 24259
rect 26559 24225 26568 24259
rect 26516 24216 26568 24225
rect 26792 24259 26844 24268
rect 26792 24225 26801 24259
rect 26801 24225 26835 24259
rect 26835 24225 26844 24259
rect 26792 24216 26844 24225
rect 22836 24080 22888 24132
rect 19708 24012 19760 24021
rect 20996 24012 21048 24064
rect 21640 24012 21692 24064
rect 25872 24191 25924 24200
rect 25872 24157 25881 24191
rect 25881 24157 25915 24191
rect 25915 24157 25924 24191
rect 25872 24148 25924 24157
rect 26424 24191 26476 24200
rect 26424 24157 26433 24191
rect 26433 24157 26467 24191
rect 26467 24157 26476 24191
rect 26424 24148 26476 24157
rect 26148 24012 26200 24064
rect 27804 24080 27856 24132
rect 26424 24012 26476 24064
rect 4874 23910 4926 23962
rect 4938 23910 4990 23962
rect 5002 23910 5054 23962
rect 5066 23910 5118 23962
rect 5130 23910 5182 23962
rect 9220 23851 9272 23860
rect 9220 23817 9229 23851
rect 9229 23817 9263 23851
rect 9263 23817 9272 23851
rect 9220 23808 9272 23817
rect 10048 23808 10100 23860
rect 14188 23808 14240 23860
rect 16212 23808 16264 23860
rect 16764 23851 16816 23860
rect 16764 23817 16773 23851
rect 16773 23817 16807 23851
rect 16807 23817 16816 23851
rect 16764 23808 16816 23817
rect 19708 23808 19760 23860
rect 20168 23851 20220 23860
rect 20168 23817 20177 23851
rect 20177 23817 20211 23851
rect 20211 23817 20220 23851
rect 20168 23808 20220 23817
rect 21088 23808 21140 23860
rect 25596 23808 25648 23860
rect 25872 23808 25924 23860
rect 9864 23740 9916 23792
rect 9128 23715 9180 23724
rect 9128 23681 9137 23715
rect 9137 23681 9171 23715
rect 9171 23681 9180 23715
rect 9128 23672 9180 23681
rect 9772 23672 9824 23724
rect 11060 23715 11112 23724
rect 11060 23681 11069 23715
rect 11069 23681 11103 23715
rect 11103 23681 11112 23715
rect 11060 23672 11112 23681
rect 11612 23672 11664 23724
rect 13452 23740 13504 23792
rect 17868 23783 17920 23792
rect 17868 23749 17877 23783
rect 17877 23749 17911 23783
rect 17911 23749 17920 23783
rect 17868 23740 17920 23749
rect 17960 23740 18012 23792
rect 19616 23740 19668 23792
rect 21272 23783 21324 23792
rect 12164 23715 12216 23724
rect 12164 23681 12173 23715
rect 12173 23681 12207 23715
rect 12207 23681 12216 23715
rect 12164 23672 12216 23681
rect 11980 23604 12032 23656
rect 12992 23672 13044 23724
rect 16028 23672 16080 23724
rect 16120 23715 16172 23724
rect 16120 23681 16129 23715
rect 16129 23681 16163 23715
rect 16163 23681 16172 23715
rect 16120 23672 16172 23681
rect 16304 23715 16356 23724
rect 16304 23681 16313 23715
rect 16313 23681 16347 23715
rect 16347 23681 16356 23715
rect 16304 23672 16356 23681
rect 16856 23715 16908 23724
rect 16856 23681 16865 23715
rect 16865 23681 16899 23715
rect 16899 23681 16908 23715
rect 16856 23672 16908 23681
rect 19432 23672 19484 23724
rect 17592 23647 17644 23656
rect 17592 23613 17601 23647
rect 17601 23613 17635 23647
rect 17635 23613 17644 23647
rect 17592 23604 17644 23613
rect 11520 23536 11572 23588
rect 12164 23536 12216 23588
rect 17132 23536 17184 23588
rect 19616 23604 19668 23656
rect 19800 23715 19852 23724
rect 19800 23681 19809 23715
rect 19809 23681 19843 23715
rect 19843 23681 19852 23715
rect 19800 23672 19852 23681
rect 21272 23749 21281 23783
rect 21281 23749 21315 23783
rect 21315 23749 21324 23783
rect 21272 23740 21324 23749
rect 20996 23715 21048 23724
rect 20996 23681 21005 23715
rect 21005 23681 21039 23715
rect 21039 23681 21048 23715
rect 20996 23672 21048 23681
rect 21180 23715 21232 23724
rect 21180 23681 21187 23715
rect 21187 23681 21232 23715
rect 21180 23672 21232 23681
rect 21364 23715 21416 23724
rect 21364 23681 21373 23715
rect 21373 23681 21407 23715
rect 21407 23681 21416 23715
rect 21364 23672 21416 23681
rect 21640 23672 21692 23724
rect 22928 23740 22980 23792
rect 26332 23740 26384 23792
rect 20812 23647 20864 23656
rect 20812 23613 20821 23647
rect 20821 23613 20855 23647
rect 20855 23613 20864 23647
rect 20812 23604 20864 23613
rect 22008 23604 22060 23656
rect 25688 23715 25740 23724
rect 25688 23681 25697 23715
rect 25697 23681 25731 23715
rect 25731 23681 25740 23715
rect 25688 23672 25740 23681
rect 26424 23715 26476 23724
rect 26424 23681 26433 23715
rect 26433 23681 26467 23715
rect 26467 23681 26476 23715
rect 26424 23672 26476 23681
rect 27988 23740 28040 23792
rect 27160 23672 27212 23724
rect 27896 23604 27948 23656
rect 26884 23536 26936 23588
rect 11152 23468 11204 23520
rect 21640 23511 21692 23520
rect 21640 23477 21649 23511
rect 21649 23477 21683 23511
rect 21683 23477 21692 23511
rect 21640 23468 21692 23477
rect 22100 23468 22152 23520
rect 25044 23468 25096 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 11244 23264 11296 23316
rect 19800 23264 19852 23316
rect 27896 23264 27948 23316
rect 15384 23196 15436 23248
rect 20812 23196 20864 23248
rect 10968 23171 11020 23180
rect 10968 23137 10977 23171
rect 10977 23137 11011 23171
rect 11011 23137 11020 23171
rect 10968 23128 11020 23137
rect 15752 23128 15804 23180
rect 17132 23128 17184 23180
rect 17592 23128 17644 23180
rect 21732 23128 21784 23180
rect 26516 23171 26568 23180
rect 26516 23137 26525 23171
rect 26525 23137 26559 23171
rect 26559 23137 26568 23171
rect 26516 23128 26568 23137
rect 26884 23128 26936 23180
rect 11152 23103 11204 23112
rect 11152 23069 11161 23103
rect 11161 23069 11195 23103
rect 11195 23069 11204 23103
rect 11152 23060 11204 23069
rect 15108 23060 15160 23112
rect 15844 23103 15896 23112
rect 15844 23069 15853 23103
rect 15853 23069 15887 23103
rect 15887 23069 15896 23103
rect 15844 23060 15896 23069
rect 16120 23103 16172 23112
rect 16120 23069 16129 23103
rect 16129 23069 16163 23103
rect 16163 23069 16172 23103
rect 16120 23060 16172 23069
rect 19340 23060 19392 23112
rect 21640 23103 21692 23112
rect 21640 23069 21649 23103
rect 21649 23069 21683 23103
rect 21683 23069 21692 23103
rect 21640 23060 21692 23069
rect 15292 23035 15344 23044
rect 15292 23001 15301 23035
rect 15301 23001 15335 23035
rect 15335 23001 15344 23035
rect 15292 22992 15344 23001
rect 17500 23035 17552 23044
rect 17500 23001 17509 23035
rect 17509 23001 17543 23035
rect 17543 23001 17552 23035
rect 17500 22992 17552 23001
rect 17960 22992 18012 23044
rect 20996 22992 21048 23044
rect 21364 22992 21416 23044
rect 22100 23060 22152 23112
rect 22836 23060 22888 23112
rect 26424 23060 26476 23112
rect 27804 22992 27856 23044
rect 15568 22924 15620 22976
rect 23940 22924 23992 22976
rect 26332 22967 26384 22976
rect 26332 22933 26341 22967
rect 26341 22933 26375 22967
rect 26375 22933 26384 22967
rect 26332 22924 26384 22933
rect 4874 22822 4926 22874
rect 4938 22822 4990 22874
rect 5002 22822 5054 22874
rect 5066 22822 5118 22874
rect 5130 22822 5182 22874
rect 15292 22720 15344 22772
rect 17960 22720 18012 22772
rect 18880 22720 18932 22772
rect 8116 22652 8168 22704
rect 13268 22695 13320 22704
rect 13268 22661 13277 22695
rect 13277 22661 13311 22695
rect 13311 22661 13320 22695
rect 13268 22652 13320 22661
rect 15844 22652 15896 22704
rect 22100 22652 22152 22704
rect 7748 22627 7800 22636
rect 7748 22593 7757 22627
rect 7757 22593 7791 22627
rect 7791 22593 7800 22627
rect 7748 22584 7800 22593
rect 9680 22584 9732 22636
rect 13084 22584 13136 22636
rect 14096 22627 14148 22636
rect 14096 22593 14105 22627
rect 14105 22593 14139 22627
rect 14139 22593 14148 22627
rect 14096 22584 14148 22593
rect 15016 22516 15068 22568
rect 7840 22448 7892 22500
rect 15292 22627 15344 22636
rect 15292 22593 15301 22627
rect 15301 22593 15335 22627
rect 15335 22593 15344 22627
rect 15292 22584 15344 22593
rect 15384 22584 15436 22636
rect 23940 22627 23992 22636
rect 23940 22593 23949 22627
rect 23949 22593 23983 22627
rect 23983 22593 23992 22627
rect 23940 22584 23992 22593
rect 24584 22652 24636 22704
rect 28356 22652 28408 22704
rect 15936 22516 15988 22568
rect 20352 22559 20404 22568
rect 20352 22525 20361 22559
rect 20361 22525 20395 22559
rect 20395 22525 20404 22559
rect 20352 22516 20404 22525
rect 22376 22559 22428 22568
rect 22376 22525 22385 22559
rect 22385 22525 22419 22559
rect 22419 22525 22428 22559
rect 22376 22516 22428 22525
rect 23480 22516 23532 22568
rect 15568 22448 15620 22500
rect 16488 22448 16540 22500
rect 22836 22448 22888 22500
rect 9036 22380 9088 22432
rect 12072 22380 12124 22432
rect 14372 22380 14424 22432
rect 15200 22423 15252 22432
rect 15200 22389 15209 22423
rect 15209 22389 15243 22423
rect 15243 22389 15252 22423
rect 15200 22380 15252 22389
rect 15476 22423 15528 22432
rect 15476 22389 15485 22423
rect 15485 22389 15519 22423
rect 15519 22389 15528 22423
rect 15476 22380 15528 22389
rect 16672 22423 16724 22432
rect 16672 22389 16681 22423
rect 16681 22389 16715 22423
rect 16715 22389 16724 22423
rect 16672 22380 16724 22389
rect 19524 22380 19576 22432
rect 21824 22423 21876 22432
rect 21824 22389 21833 22423
rect 21833 22389 21867 22423
rect 21867 22389 21876 22423
rect 21824 22380 21876 22389
rect 23020 22380 23072 22432
rect 24952 22627 25004 22636
rect 24952 22593 24961 22627
rect 24961 22593 24995 22627
rect 24995 22593 25004 22627
rect 24952 22584 25004 22593
rect 25228 22627 25280 22636
rect 25228 22593 25237 22627
rect 25237 22593 25271 22627
rect 25271 22593 25280 22627
rect 25228 22584 25280 22593
rect 26424 22627 26476 22636
rect 26424 22593 26433 22627
rect 26433 22593 26467 22627
rect 26467 22593 26476 22627
rect 26424 22584 26476 22593
rect 25044 22559 25096 22568
rect 25044 22525 25053 22559
rect 25053 22525 25087 22559
rect 25087 22525 25096 22559
rect 25044 22516 25096 22525
rect 25596 22559 25648 22568
rect 25596 22525 25605 22559
rect 25605 22525 25639 22559
rect 25639 22525 25648 22559
rect 25596 22516 25648 22525
rect 26332 22516 26384 22568
rect 27896 22584 27948 22636
rect 27436 22516 27488 22568
rect 27620 22559 27672 22568
rect 27620 22525 27629 22559
rect 27629 22525 27663 22559
rect 27663 22525 27672 22559
rect 27620 22516 27672 22525
rect 26608 22448 26660 22500
rect 27988 22448 28040 22500
rect 24860 22380 24912 22432
rect 26148 22423 26200 22432
rect 26148 22389 26157 22423
rect 26157 22389 26191 22423
rect 26191 22389 26200 22423
rect 26148 22380 26200 22389
rect 26976 22423 27028 22432
rect 26976 22389 26985 22423
rect 26985 22389 27019 22423
rect 27019 22389 27028 22423
rect 26976 22380 27028 22389
rect 28080 22380 28132 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 15936 22219 15988 22228
rect 15936 22185 15945 22219
rect 15945 22185 15979 22219
rect 15979 22185 15988 22219
rect 15936 22176 15988 22185
rect 16488 22176 16540 22228
rect 19524 22219 19576 22228
rect 19524 22185 19554 22219
rect 19554 22185 19576 22219
rect 19524 22176 19576 22185
rect 21824 22176 21876 22228
rect 22836 22219 22888 22228
rect 22836 22185 22845 22219
rect 22845 22185 22879 22219
rect 22879 22185 22888 22219
rect 22836 22176 22888 22185
rect 26148 22176 26200 22228
rect 26976 22176 27028 22228
rect 16120 22108 16172 22160
rect 6920 22040 6972 22092
rect 7932 22040 7984 22092
rect 8116 22040 8168 22092
rect 8576 21972 8628 22024
rect 10968 21972 11020 22024
rect 4804 21904 4856 21956
rect 5540 21947 5592 21956
rect 5540 21913 5549 21947
rect 5549 21913 5583 21947
rect 5583 21913 5592 21947
rect 5540 21904 5592 21913
rect 6276 21947 6328 21956
rect 6276 21913 6285 21947
rect 6285 21913 6319 21947
rect 6319 21913 6328 21947
rect 6276 21904 6328 21913
rect 7840 21947 7892 21956
rect 7840 21913 7849 21947
rect 7849 21913 7883 21947
rect 7883 21913 7892 21947
rect 7840 21904 7892 21913
rect 7932 21904 7984 21956
rect 9588 21904 9640 21956
rect 13176 22040 13228 22092
rect 17592 22040 17644 22092
rect 19248 22083 19300 22092
rect 19248 22049 19257 22083
rect 19257 22049 19291 22083
rect 19291 22049 19300 22083
rect 19248 22040 19300 22049
rect 11428 22015 11480 22024
rect 11428 21981 11437 22015
rect 11437 21981 11471 22015
rect 11471 21981 11480 22015
rect 11428 21972 11480 21981
rect 12072 22015 12124 22024
rect 12072 21981 12081 22015
rect 12081 21981 12115 22015
rect 12115 21981 12124 22015
rect 12072 21972 12124 21981
rect 16120 21972 16172 22024
rect 16672 22015 16724 22024
rect 16672 21981 16681 22015
rect 16681 21981 16715 22015
rect 16715 21981 16724 22015
rect 16672 21972 16724 21981
rect 24032 22040 24084 22092
rect 24216 21972 24268 22024
rect 4068 21879 4120 21888
rect 4068 21845 4077 21879
rect 4077 21845 4111 21879
rect 4111 21845 4120 21879
rect 4068 21836 4120 21845
rect 7012 21836 7064 21888
rect 9128 21836 9180 21888
rect 11796 21836 11848 21888
rect 11888 21879 11940 21888
rect 11888 21845 11897 21879
rect 11897 21845 11931 21879
rect 11931 21845 11940 21879
rect 11888 21836 11940 21845
rect 12440 21947 12492 21956
rect 12440 21913 12449 21947
rect 12449 21913 12483 21947
rect 12483 21913 12492 21947
rect 12440 21904 12492 21913
rect 12900 21904 12952 21956
rect 15476 21904 15528 21956
rect 15936 21904 15988 21956
rect 17592 21947 17644 21956
rect 17592 21913 17601 21947
rect 17601 21913 17635 21947
rect 17635 21913 17644 21947
rect 17592 21904 17644 21913
rect 18880 21904 18932 21956
rect 19800 21904 19852 21956
rect 20536 21904 20588 21956
rect 24584 21904 24636 21956
rect 25504 21904 25556 21956
rect 26516 21904 26568 21956
rect 28448 21904 28500 21956
rect 12716 21836 12768 21888
rect 15108 21836 15160 21888
rect 19340 21836 19392 21888
rect 20996 21879 21048 21888
rect 20996 21845 21005 21879
rect 21005 21845 21039 21879
rect 21039 21845 21048 21879
rect 20996 21836 21048 21845
rect 22744 21836 22796 21888
rect 23112 21836 23164 21888
rect 23480 21836 23532 21888
rect 23664 21879 23716 21888
rect 23664 21845 23673 21879
rect 23673 21845 23707 21879
rect 23707 21845 23716 21879
rect 23664 21836 23716 21845
rect 25228 21836 25280 21888
rect 27344 21836 27396 21888
rect 4874 21734 4926 21786
rect 4938 21734 4990 21786
rect 5002 21734 5054 21786
rect 5066 21734 5118 21786
rect 5130 21734 5182 21786
rect 5540 21632 5592 21684
rect 4988 21564 5040 21616
rect 7840 21632 7892 21684
rect 14096 21632 14148 21684
rect 16488 21675 16540 21684
rect 4068 21496 4120 21548
rect 5080 21539 5132 21548
rect 5080 21505 5089 21539
rect 5089 21505 5123 21539
rect 5123 21505 5132 21539
rect 5080 21496 5132 21505
rect 5356 21496 5408 21548
rect 5816 21539 5868 21548
rect 5816 21505 5825 21539
rect 5825 21505 5859 21539
rect 5859 21505 5868 21539
rect 5816 21496 5868 21505
rect 11704 21564 11756 21616
rect 11796 21607 11848 21616
rect 11796 21573 11805 21607
rect 11805 21573 11839 21607
rect 11839 21573 11848 21607
rect 11796 21564 11848 21573
rect 6092 21496 6144 21548
rect 6920 21496 6972 21548
rect 7564 21496 7616 21548
rect 9220 21496 9272 21548
rect 5356 21360 5408 21412
rect 5724 21428 5776 21480
rect 8668 21428 8720 21480
rect 6092 21292 6144 21344
rect 6184 21335 6236 21344
rect 6184 21301 6193 21335
rect 6193 21301 6227 21335
rect 6227 21301 6236 21335
rect 6184 21292 6236 21301
rect 7196 21360 7248 21412
rect 9588 21539 9640 21548
rect 9588 21505 9597 21539
rect 9597 21505 9631 21539
rect 9631 21505 9640 21539
rect 9588 21496 9640 21505
rect 12900 21496 12952 21548
rect 13268 21496 13320 21548
rect 9864 21471 9916 21480
rect 9864 21437 9873 21471
rect 9873 21437 9907 21471
rect 9907 21437 9916 21471
rect 9864 21428 9916 21437
rect 16488 21641 16497 21675
rect 16497 21641 16531 21675
rect 16531 21641 16540 21675
rect 16488 21632 16540 21641
rect 20352 21632 20404 21684
rect 20996 21632 21048 21684
rect 22376 21632 22428 21684
rect 16304 21564 16356 21616
rect 18880 21564 18932 21616
rect 19248 21564 19300 21616
rect 22652 21564 22704 21616
rect 19340 21496 19392 21548
rect 22192 21539 22244 21548
rect 22192 21505 22201 21539
rect 22201 21505 22235 21539
rect 22235 21505 22244 21539
rect 22192 21496 22244 21505
rect 24032 21632 24084 21684
rect 24584 21632 24636 21684
rect 23020 21607 23072 21616
rect 23020 21573 23029 21607
rect 23029 21573 23063 21607
rect 23063 21573 23072 21607
rect 23020 21564 23072 21573
rect 25504 21632 25556 21684
rect 25596 21632 25648 21684
rect 26424 21632 26476 21684
rect 25044 21564 25096 21616
rect 27344 21607 27396 21616
rect 26608 21496 26660 21548
rect 27344 21573 27353 21607
rect 27353 21573 27387 21607
rect 27387 21573 27396 21607
rect 27344 21564 27396 21573
rect 10968 21360 11020 21412
rect 6920 21292 6972 21344
rect 13084 21360 13136 21412
rect 14372 21471 14424 21480
rect 14372 21437 14381 21471
rect 14381 21437 14415 21471
rect 14415 21437 14424 21471
rect 14372 21428 14424 21437
rect 15476 21428 15528 21480
rect 19616 21428 19668 21480
rect 21456 21471 21508 21480
rect 21456 21437 21465 21471
rect 21465 21437 21499 21471
rect 21499 21437 21508 21471
rect 21456 21428 21508 21437
rect 22744 21471 22796 21480
rect 22744 21437 22753 21471
rect 22753 21437 22787 21471
rect 22787 21437 22796 21471
rect 22744 21428 22796 21437
rect 24216 21428 24268 21480
rect 12900 21292 12952 21344
rect 14832 21292 14884 21344
rect 25228 21471 25280 21480
rect 25228 21437 25237 21471
rect 25237 21437 25271 21471
rect 25271 21437 25280 21471
rect 25228 21428 25280 21437
rect 26332 21471 26384 21480
rect 26332 21437 26341 21471
rect 26341 21437 26375 21471
rect 26375 21437 26384 21471
rect 26332 21428 26384 21437
rect 27436 21539 27488 21548
rect 27436 21505 27450 21539
rect 27450 21505 27484 21539
rect 27484 21505 27488 21539
rect 27436 21496 27488 21505
rect 28264 21471 28316 21480
rect 28264 21437 28273 21471
rect 28273 21437 28307 21471
rect 28307 21437 28316 21471
rect 28264 21428 28316 21437
rect 26792 21360 26844 21412
rect 27160 21292 27212 21344
rect 28172 21292 28224 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 5724 21088 5776 21140
rect 6276 21088 6328 21140
rect 11428 21088 11480 21140
rect 5080 20952 5132 21004
rect 5172 20927 5224 20936
rect 5172 20893 5181 20927
rect 5181 20893 5215 20927
rect 5215 20893 5224 20927
rect 5172 20884 5224 20893
rect 5356 20927 5408 20936
rect 5356 20893 5365 20927
rect 5365 20893 5399 20927
rect 5399 20893 5408 20927
rect 5356 20884 5408 20893
rect 5540 20927 5592 20936
rect 5540 20893 5549 20927
rect 5549 20893 5583 20927
rect 5583 20893 5592 20927
rect 5540 20884 5592 20893
rect 5816 20884 5868 20936
rect 6184 20927 6236 20936
rect 6184 20893 6193 20927
rect 6193 20893 6227 20927
rect 6227 20893 6236 20927
rect 6184 20884 6236 20893
rect 4712 20816 4764 20868
rect 4988 20816 5040 20868
rect 5908 20816 5960 20868
rect 7840 20884 7892 20936
rect 8392 20884 8444 20936
rect 9220 20952 9272 21004
rect 12440 21088 12492 21140
rect 15476 21131 15528 21140
rect 15476 21097 15485 21131
rect 15485 21097 15519 21131
rect 15519 21097 15528 21131
rect 15476 21088 15528 21097
rect 17500 21131 17552 21140
rect 17500 21097 17509 21131
rect 17509 21097 17543 21131
rect 17543 21097 17552 21131
rect 17500 21088 17552 21097
rect 23664 21088 23716 21140
rect 6368 20859 6420 20868
rect 6368 20825 6377 20859
rect 6377 20825 6411 20859
rect 6411 20825 6420 20859
rect 6368 20816 6420 20825
rect 7012 20816 7064 20868
rect 7564 20816 7616 20868
rect 8208 20748 8260 20800
rect 9128 20927 9180 20936
rect 9128 20893 9137 20927
rect 9137 20893 9171 20927
rect 9171 20893 9180 20927
rect 9128 20884 9180 20893
rect 9312 20927 9364 20936
rect 9312 20893 9321 20927
rect 9321 20893 9355 20927
rect 9355 20893 9364 20927
rect 9312 20884 9364 20893
rect 11152 20884 11204 20936
rect 11888 20884 11940 20936
rect 14832 20995 14884 21004
rect 14832 20961 14841 20995
rect 14841 20961 14875 20995
rect 14875 20961 14884 20995
rect 14832 20952 14884 20961
rect 19248 20952 19300 21004
rect 9956 20816 10008 20868
rect 12716 20927 12768 20936
rect 12716 20893 12725 20927
rect 12725 20893 12759 20927
rect 12759 20893 12768 20927
rect 12716 20884 12768 20893
rect 12900 20927 12952 20936
rect 12900 20893 12909 20927
rect 12909 20893 12943 20927
rect 12943 20893 12952 20927
rect 12900 20884 12952 20893
rect 15200 20884 15252 20936
rect 15844 20927 15896 20936
rect 15844 20893 15853 20927
rect 15853 20893 15887 20927
rect 15887 20893 15896 20927
rect 15844 20884 15896 20893
rect 9312 20748 9364 20800
rect 9772 20748 9824 20800
rect 14372 20816 14424 20868
rect 17960 20927 18012 20936
rect 17960 20893 17969 20927
rect 17969 20893 18003 20927
rect 18003 20893 18012 20927
rect 17960 20884 18012 20893
rect 22744 20952 22796 21004
rect 24032 20952 24084 21004
rect 24768 20952 24820 21004
rect 26792 20995 26844 21004
rect 26792 20961 26801 20995
rect 26801 20961 26835 20995
rect 26835 20961 26844 20995
rect 26792 20952 26844 20961
rect 23112 20884 23164 20936
rect 25504 20884 25556 20936
rect 18420 20816 18472 20868
rect 20168 20859 20220 20868
rect 20168 20825 20177 20859
rect 20177 20825 20211 20859
rect 20211 20825 20220 20859
rect 20168 20816 20220 20825
rect 20628 20816 20680 20868
rect 22284 20816 22336 20868
rect 24400 20859 24452 20868
rect 24400 20825 24409 20859
rect 24409 20825 24443 20859
rect 24443 20825 24452 20859
rect 24400 20816 24452 20825
rect 26792 20816 26844 20868
rect 12716 20748 12768 20800
rect 12992 20748 13044 20800
rect 15936 20748 15988 20800
rect 17408 20748 17460 20800
rect 21640 20791 21692 20800
rect 21640 20757 21649 20791
rect 21649 20757 21683 20791
rect 21683 20757 21692 20791
rect 21640 20748 21692 20757
rect 27804 20748 27856 20800
rect 4874 20646 4926 20698
rect 4938 20646 4990 20698
rect 5002 20646 5054 20698
rect 5066 20646 5118 20698
rect 5130 20646 5182 20698
rect 4804 20544 4856 20596
rect 5448 20476 5500 20528
rect 5908 20544 5960 20596
rect 8116 20544 8168 20596
rect 9404 20544 9456 20596
rect 9864 20544 9916 20596
rect 5816 20519 5868 20528
rect 5816 20485 5825 20519
rect 5825 20485 5859 20519
rect 5859 20485 5868 20519
rect 5816 20476 5868 20485
rect 6368 20476 6420 20528
rect 5724 20451 5776 20460
rect 5724 20417 5733 20451
rect 5733 20417 5767 20451
rect 5767 20417 5776 20451
rect 5724 20408 5776 20417
rect 6920 20476 6972 20528
rect 8392 20476 8444 20528
rect 8576 20476 8628 20528
rect 10968 20476 11020 20528
rect 14096 20544 14148 20596
rect 16396 20544 16448 20596
rect 16304 20476 16356 20528
rect 3608 20383 3660 20392
rect 3608 20349 3617 20383
rect 3617 20349 3651 20383
rect 3651 20349 3660 20383
rect 3608 20340 3660 20349
rect 5540 20340 5592 20392
rect 5264 20204 5316 20256
rect 5632 20204 5684 20256
rect 7012 20247 7064 20256
rect 7012 20213 7021 20247
rect 7021 20213 7055 20247
rect 7055 20213 7064 20247
rect 7012 20204 7064 20213
rect 7196 20451 7248 20460
rect 7196 20417 7205 20451
rect 7205 20417 7239 20451
rect 7239 20417 7248 20451
rect 7196 20408 7248 20417
rect 7288 20451 7340 20460
rect 7288 20417 7297 20451
rect 7297 20417 7331 20451
rect 7331 20417 7340 20451
rect 7288 20408 7340 20417
rect 9772 20451 9824 20460
rect 9772 20417 9781 20451
rect 9781 20417 9815 20451
rect 9815 20417 9824 20451
rect 9772 20408 9824 20417
rect 7564 20340 7616 20392
rect 8116 20383 8168 20392
rect 8116 20349 8125 20383
rect 8125 20349 8159 20383
rect 8159 20349 8168 20383
rect 8116 20340 8168 20349
rect 8576 20340 8628 20392
rect 9588 20340 9640 20392
rect 8300 20204 8352 20256
rect 9588 20204 9640 20256
rect 10692 20408 10744 20460
rect 11612 20272 11664 20324
rect 16488 20408 16540 20460
rect 19248 20544 19300 20596
rect 21456 20544 21508 20596
rect 22192 20544 22244 20596
rect 26332 20544 26384 20596
rect 27620 20544 27672 20596
rect 19800 20476 19852 20528
rect 20628 20476 20680 20528
rect 25504 20476 25556 20528
rect 27436 20519 27488 20528
rect 27436 20485 27445 20519
rect 27445 20485 27479 20519
rect 27479 20485 27488 20519
rect 27436 20476 27488 20485
rect 28080 20519 28132 20528
rect 28080 20485 28089 20519
rect 28089 20485 28123 20519
rect 28123 20485 28132 20519
rect 28080 20476 28132 20485
rect 28172 20519 28224 20528
rect 28172 20485 28181 20519
rect 28181 20485 28215 20519
rect 28215 20485 28224 20519
rect 28172 20476 28224 20485
rect 20536 20408 20588 20460
rect 21456 20451 21508 20460
rect 21456 20417 21465 20451
rect 21465 20417 21499 20451
rect 21499 20417 21508 20451
rect 21456 20408 21508 20417
rect 21640 20408 21692 20460
rect 27988 20451 28040 20460
rect 27988 20417 27997 20451
rect 27997 20417 28031 20451
rect 28031 20417 28040 20451
rect 27988 20408 28040 20417
rect 28356 20451 28408 20460
rect 28356 20417 28365 20451
rect 28365 20417 28399 20451
rect 28399 20417 28408 20451
rect 28356 20408 28408 20417
rect 14188 20383 14240 20392
rect 14188 20349 14197 20383
rect 14197 20349 14231 20383
rect 14231 20349 14240 20383
rect 14188 20340 14240 20349
rect 15936 20340 15988 20392
rect 17040 20340 17092 20392
rect 18880 20340 18932 20392
rect 23480 20383 23532 20392
rect 23480 20349 23489 20383
rect 23489 20349 23523 20383
rect 23523 20349 23532 20383
rect 23480 20340 23532 20349
rect 23756 20383 23808 20392
rect 23756 20349 23765 20383
rect 23765 20349 23799 20383
rect 23799 20349 23808 20383
rect 23756 20340 23808 20349
rect 26700 20340 26752 20392
rect 27252 20340 27304 20392
rect 19432 20272 19484 20324
rect 16212 20204 16264 20256
rect 18236 20204 18288 20256
rect 25504 20272 25556 20324
rect 28448 20272 28500 20324
rect 24400 20204 24452 20256
rect 27988 20204 28040 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 7196 20000 7248 20052
rect 7748 20000 7800 20052
rect 8116 20000 8168 20052
rect 8668 20043 8720 20052
rect 8668 20009 8677 20043
rect 8677 20009 8711 20043
rect 8711 20009 8720 20043
rect 8668 20000 8720 20009
rect 12624 20000 12676 20052
rect 17408 20043 17460 20052
rect 17408 20009 17417 20043
rect 17417 20009 17451 20043
rect 17451 20009 17460 20043
rect 17408 20000 17460 20009
rect 17592 20000 17644 20052
rect 20168 20000 20220 20052
rect 26700 20000 26752 20052
rect 28264 20000 28316 20052
rect 6920 19932 6972 19984
rect 5908 19864 5960 19916
rect 7012 19839 7064 19848
rect 7012 19805 7021 19839
rect 7021 19805 7055 19839
rect 7055 19805 7064 19839
rect 7012 19796 7064 19805
rect 7288 19796 7340 19848
rect 7748 19796 7800 19848
rect 8208 19839 8260 19848
rect 8208 19805 8217 19839
rect 8217 19805 8251 19839
rect 8251 19805 8260 19839
rect 8208 19796 8260 19805
rect 11244 19864 11296 19916
rect 15752 19932 15804 19984
rect 17040 19932 17092 19984
rect 3608 19660 3660 19712
rect 6828 19660 6880 19712
rect 8300 19771 8352 19780
rect 8300 19737 8309 19771
rect 8309 19737 8343 19771
rect 8343 19737 8352 19771
rect 8300 19728 8352 19737
rect 9036 19796 9088 19848
rect 11704 19796 11756 19848
rect 12624 19796 12676 19848
rect 12532 19728 12584 19780
rect 13268 19796 13320 19848
rect 16488 19864 16540 19916
rect 16028 19796 16080 19848
rect 18512 19864 18564 19916
rect 17960 19839 18012 19848
rect 17960 19805 17964 19839
rect 17964 19805 17998 19839
rect 17998 19805 18012 19839
rect 17960 19796 18012 19805
rect 18236 19839 18288 19848
rect 18236 19805 18281 19839
rect 18281 19805 18288 19839
rect 18236 19796 18288 19805
rect 18420 19839 18472 19848
rect 18420 19805 18429 19839
rect 18429 19805 18463 19839
rect 18463 19805 18472 19839
rect 19248 19839 19300 19848
rect 18420 19796 18472 19805
rect 19248 19805 19257 19839
rect 19257 19805 19291 19839
rect 19291 19805 19300 19839
rect 19248 19796 19300 19805
rect 19432 19839 19484 19848
rect 19432 19805 19439 19839
rect 19439 19805 19484 19839
rect 19432 19796 19484 19805
rect 20536 19864 20588 19916
rect 19708 19839 19760 19848
rect 19708 19805 19722 19839
rect 19722 19805 19756 19839
rect 19756 19805 19760 19839
rect 19708 19796 19760 19805
rect 21916 19864 21968 19916
rect 22100 19907 22152 19916
rect 22100 19873 22109 19907
rect 22109 19873 22143 19907
rect 22143 19873 22152 19907
rect 22100 19864 22152 19873
rect 23204 19864 23256 19916
rect 24124 19932 24176 19984
rect 23480 19864 23532 19916
rect 27252 19907 27304 19916
rect 27252 19873 27261 19907
rect 27261 19873 27295 19907
rect 27295 19873 27304 19907
rect 27252 19864 27304 19873
rect 27804 19864 27856 19916
rect 8852 19660 8904 19712
rect 9588 19660 9640 19712
rect 12900 19660 12952 19712
rect 13544 19660 13596 19712
rect 15752 19660 15804 19712
rect 18052 19771 18104 19780
rect 18052 19737 18061 19771
rect 18061 19737 18095 19771
rect 18095 19737 18104 19771
rect 18052 19728 18104 19737
rect 18604 19728 18656 19780
rect 18696 19660 18748 19712
rect 23480 19728 23532 19780
rect 24216 19796 24268 19848
rect 24768 19839 24820 19848
rect 24768 19805 24777 19839
rect 24777 19805 24811 19839
rect 24811 19805 24820 19839
rect 24768 19796 24820 19805
rect 25044 19839 25096 19848
rect 25044 19805 25053 19839
rect 25053 19805 25087 19839
rect 25087 19805 25096 19839
rect 25044 19796 25096 19805
rect 27712 19796 27764 19848
rect 28080 19796 28132 19848
rect 28448 19796 28500 19848
rect 22008 19660 22060 19712
rect 23848 19771 23900 19780
rect 23848 19737 23857 19771
rect 23857 19737 23891 19771
rect 23891 19737 23900 19771
rect 23848 19728 23900 19737
rect 23940 19771 23992 19780
rect 23940 19737 23949 19771
rect 23949 19737 23983 19771
rect 23983 19737 23992 19771
rect 23940 19728 23992 19737
rect 24032 19660 24084 19712
rect 26792 19728 26844 19780
rect 27712 19660 27764 19712
rect 4874 19558 4926 19610
rect 4938 19558 4990 19610
rect 5002 19558 5054 19610
rect 5066 19558 5118 19610
rect 5130 19558 5182 19610
rect 4712 19388 4764 19440
rect 4988 19363 5040 19372
rect 4988 19329 4997 19363
rect 4997 19329 5031 19363
rect 5031 19329 5040 19363
rect 4988 19320 5040 19329
rect 11244 19499 11296 19508
rect 11244 19465 11253 19499
rect 11253 19465 11287 19499
rect 11287 19465 11296 19499
rect 11244 19456 11296 19465
rect 11704 19499 11756 19508
rect 11704 19465 11713 19499
rect 11713 19465 11747 19499
rect 11747 19465 11756 19499
rect 11704 19456 11756 19465
rect 12532 19456 12584 19508
rect 16028 19499 16080 19508
rect 16028 19465 16037 19499
rect 16037 19465 16071 19499
rect 16071 19465 16080 19499
rect 16028 19456 16080 19465
rect 18052 19456 18104 19508
rect 18604 19456 18656 19508
rect 18880 19499 18932 19508
rect 18880 19465 18889 19499
rect 18889 19465 18923 19499
rect 18923 19465 18932 19499
rect 18880 19456 18932 19465
rect 19248 19456 19300 19508
rect 5264 19320 5316 19372
rect 8116 19388 8168 19440
rect 5540 19320 5592 19372
rect 5632 19363 5684 19372
rect 5632 19329 5641 19363
rect 5641 19329 5675 19363
rect 5675 19329 5684 19363
rect 5632 19320 5684 19329
rect 5908 19363 5960 19372
rect 5908 19329 5917 19363
rect 5917 19329 5951 19363
rect 5951 19329 5960 19363
rect 5908 19320 5960 19329
rect 6092 19363 6144 19372
rect 6092 19329 6101 19363
rect 6101 19329 6135 19363
rect 6135 19329 6144 19363
rect 6092 19320 6144 19329
rect 6828 19320 6880 19372
rect 7564 19363 7616 19372
rect 7564 19329 7573 19363
rect 7573 19329 7607 19363
rect 7607 19329 7616 19363
rect 7564 19320 7616 19329
rect 8944 19320 8996 19372
rect 11520 19388 11572 19440
rect 11336 19363 11388 19372
rect 11336 19329 11345 19363
rect 11345 19329 11379 19363
rect 11379 19329 11388 19363
rect 11336 19320 11388 19329
rect 11428 19320 11480 19372
rect 12716 19388 12768 19440
rect 4804 19184 4856 19236
rect 7564 19184 7616 19236
rect 4068 19116 4120 19168
rect 5448 19116 5500 19168
rect 8944 19116 8996 19168
rect 9312 19159 9364 19168
rect 9312 19125 9321 19159
rect 9321 19125 9355 19159
rect 9355 19125 9364 19159
rect 9312 19116 9364 19125
rect 13544 19320 13596 19372
rect 16212 19363 16264 19372
rect 16212 19329 16221 19363
rect 16221 19329 16255 19363
rect 16255 19329 16264 19363
rect 16212 19320 16264 19329
rect 17040 19363 17092 19372
rect 17040 19329 17049 19363
rect 17049 19329 17083 19363
rect 17083 19329 17092 19363
rect 17040 19320 17092 19329
rect 17960 19320 18012 19372
rect 18420 19388 18472 19440
rect 12992 19252 13044 19304
rect 14188 19252 14240 19304
rect 15568 19252 15620 19304
rect 16488 19252 16540 19304
rect 17500 19295 17552 19304
rect 17500 19261 17509 19295
rect 17509 19261 17543 19295
rect 17543 19261 17552 19295
rect 17500 19252 17552 19261
rect 14556 19116 14608 19168
rect 18604 19363 18656 19372
rect 18604 19329 18613 19363
rect 18613 19329 18647 19363
rect 18647 19329 18656 19363
rect 18604 19320 18656 19329
rect 18696 19320 18748 19372
rect 19708 19320 19760 19372
rect 20444 19320 20496 19372
rect 22284 19456 22336 19508
rect 22008 19388 22060 19440
rect 21916 19363 21968 19372
rect 21916 19329 21926 19363
rect 21926 19329 21960 19363
rect 21960 19329 21968 19363
rect 21916 19320 21968 19329
rect 22284 19363 22336 19372
rect 22284 19329 22298 19363
rect 22298 19329 22332 19363
rect 22332 19329 22336 19363
rect 23204 19388 23256 19440
rect 23756 19456 23808 19508
rect 27712 19499 27764 19508
rect 27712 19465 27721 19499
rect 27721 19465 27755 19499
rect 27755 19465 27764 19499
rect 27712 19456 27764 19465
rect 24216 19388 24268 19440
rect 24400 19388 24452 19440
rect 22284 19320 22336 19329
rect 18052 19116 18104 19168
rect 23204 19295 23256 19304
rect 23204 19261 23213 19295
rect 23213 19261 23247 19295
rect 23247 19261 23256 19295
rect 23204 19252 23256 19261
rect 23572 19363 23624 19372
rect 23572 19329 23581 19363
rect 23581 19329 23615 19363
rect 23615 19329 23624 19363
rect 23572 19320 23624 19329
rect 23664 19363 23716 19372
rect 23664 19329 23673 19363
rect 23673 19329 23707 19363
rect 23707 19329 23716 19363
rect 23664 19320 23716 19329
rect 23756 19363 23808 19372
rect 23756 19329 23770 19363
rect 23770 19329 23804 19363
rect 23804 19329 23808 19363
rect 23756 19320 23808 19329
rect 24952 19320 25004 19372
rect 23480 19252 23532 19304
rect 24492 19252 24544 19304
rect 25044 19252 25096 19304
rect 26148 19252 26200 19304
rect 27896 19252 27948 19304
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 5448 18912 5500 18964
rect 6092 18912 6144 18964
rect 8944 18912 8996 18964
rect 11336 18912 11388 18964
rect 5264 18844 5316 18896
rect 4804 18751 4856 18760
rect 4804 18717 4813 18751
rect 4813 18717 4847 18751
rect 4847 18717 4856 18751
rect 4804 18708 4856 18717
rect 4436 18640 4488 18692
rect 5540 18708 5592 18760
rect 5908 18776 5960 18828
rect 5724 18751 5776 18760
rect 5724 18717 5733 18751
rect 5733 18717 5767 18751
rect 5767 18717 5776 18751
rect 5724 18708 5776 18717
rect 6000 18751 6052 18760
rect 6000 18717 6009 18751
rect 6009 18717 6043 18751
rect 6043 18717 6052 18751
rect 6000 18708 6052 18717
rect 11428 18887 11480 18896
rect 11428 18853 11437 18887
rect 11437 18853 11471 18887
rect 11471 18853 11480 18887
rect 11428 18844 11480 18853
rect 10968 18776 11020 18828
rect 11980 18776 12032 18828
rect 12808 18844 12860 18896
rect 15844 18912 15896 18964
rect 18236 18912 18288 18964
rect 18604 18912 18656 18964
rect 23664 18912 23716 18964
rect 27896 18955 27948 18964
rect 27896 18921 27905 18955
rect 27905 18921 27939 18955
rect 27939 18921 27948 18955
rect 27896 18912 27948 18921
rect 8576 18708 8628 18760
rect 9864 18708 9916 18760
rect 11152 18708 11204 18760
rect 4528 18572 4580 18624
rect 7748 18640 7800 18692
rect 11612 18751 11664 18760
rect 11612 18717 11621 18751
rect 11621 18717 11655 18751
rect 11655 18717 11664 18751
rect 11612 18708 11664 18717
rect 11704 18708 11756 18760
rect 12900 18776 12952 18828
rect 19432 18844 19484 18896
rect 23204 18844 23256 18896
rect 14188 18776 14240 18828
rect 17500 18819 17552 18828
rect 17500 18785 17509 18819
rect 17509 18785 17543 18819
rect 17543 18785 17552 18819
rect 17500 18776 17552 18785
rect 18604 18776 18656 18828
rect 20444 18819 20496 18828
rect 20444 18785 20453 18819
rect 20453 18785 20487 18819
rect 20487 18785 20496 18819
rect 20444 18776 20496 18785
rect 22100 18776 22152 18828
rect 23388 18776 23440 18828
rect 23572 18776 23624 18828
rect 23848 18776 23900 18828
rect 12992 18708 13044 18760
rect 5816 18615 5868 18624
rect 5816 18581 5825 18615
rect 5825 18581 5859 18615
rect 5859 18581 5868 18615
rect 5816 18572 5868 18581
rect 8852 18572 8904 18624
rect 13268 18751 13320 18760
rect 13268 18717 13277 18751
rect 13277 18717 13311 18751
rect 13311 18717 13320 18751
rect 13268 18708 13320 18717
rect 14464 18708 14516 18760
rect 14556 18751 14608 18760
rect 14556 18717 14565 18751
rect 14565 18717 14599 18751
rect 14599 18717 14608 18751
rect 14556 18708 14608 18717
rect 16488 18708 16540 18760
rect 17960 18751 18012 18760
rect 17960 18717 17969 18751
rect 17969 18717 18003 18751
rect 18003 18717 18012 18751
rect 17960 18708 18012 18717
rect 23204 18708 23256 18760
rect 11428 18572 11480 18624
rect 12624 18615 12676 18624
rect 12624 18581 12633 18615
rect 12633 18581 12667 18615
rect 12667 18581 12676 18615
rect 12624 18572 12676 18581
rect 12716 18572 12768 18624
rect 13268 18572 13320 18624
rect 14096 18615 14148 18624
rect 14096 18581 14105 18615
rect 14105 18581 14139 18615
rect 14139 18581 14148 18615
rect 14096 18572 14148 18581
rect 15384 18683 15436 18692
rect 15384 18649 15393 18683
rect 15393 18649 15427 18683
rect 15427 18649 15436 18683
rect 15384 18640 15436 18649
rect 19340 18683 19392 18692
rect 14464 18572 14516 18624
rect 15200 18572 15252 18624
rect 16212 18572 16264 18624
rect 16396 18572 16448 18624
rect 19340 18649 19349 18683
rect 19349 18649 19383 18683
rect 19383 18649 19392 18683
rect 19340 18640 19392 18649
rect 20812 18640 20864 18692
rect 21180 18640 21232 18692
rect 22008 18640 22060 18692
rect 24860 18751 24912 18760
rect 24860 18717 24869 18751
rect 24869 18717 24903 18751
rect 24903 18717 24912 18751
rect 24860 18708 24912 18717
rect 26148 18751 26200 18760
rect 26148 18717 26157 18751
rect 26157 18717 26191 18751
rect 26191 18717 26200 18751
rect 26148 18708 26200 18717
rect 25044 18640 25096 18692
rect 25780 18640 25832 18692
rect 26884 18640 26936 18692
rect 16948 18615 17000 18624
rect 16948 18581 16957 18615
rect 16957 18581 16991 18615
rect 16991 18581 17000 18615
rect 16948 18572 17000 18581
rect 18144 18572 18196 18624
rect 22376 18572 22428 18624
rect 4874 18470 4926 18522
rect 4938 18470 4990 18522
rect 5002 18470 5054 18522
rect 5066 18470 5118 18522
rect 5130 18470 5182 18522
rect 4804 18368 4856 18420
rect 5080 18368 5132 18420
rect 5448 18368 5500 18420
rect 3700 18300 3752 18352
rect 4068 18300 4120 18352
rect 5816 18368 5868 18420
rect 7564 18411 7616 18420
rect 7564 18377 7573 18411
rect 7573 18377 7607 18411
rect 7607 18377 7616 18411
rect 7564 18368 7616 18377
rect 4528 18275 4580 18284
rect 4528 18241 4537 18275
rect 4537 18241 4571 18275
rect 4571 18241 4580 18275
rect 4528 18232 4580 18241
rect 4804 18275 4856 18284
rect 4804 18241 4813 18275
rect 4813 18241 4847 18275
rect 4847 18241 4856 18275
rect 4804 18232 4856 18241
rect 5264 18232 5316 18284
rect 5448 18275 5500 18284
rect 5448 18241 5457 18275
rect 5457 18241 5491 18275
rect 5491 18241 5500 18275
rect 5448 18232 5500 18241
rect 5908 18232 5960 18284
rect 7748 18275 7800 18284
rect 7748 18241 7757 18275
rect 7757 18241 7791 18275
rect 7791 18241 7800 18275
rect 7748 18232 7800 18241
rect 14280 18368 14332 18420
rect 15384 18368 15436 18420
rect 16948 18368 17000 18420
rect 1860 18028 1912 18080
rect 4620 18164 4672 18216
rect 4896 18164 4948 18216
rect 4160 18096 4212 18148
rect 4436 18139 4488 18148
rect 4436 18105 4445 18139
rect 4445 18105 4479 18139
rect 4479 18105 4488 18139
rect 4436 18096 4488 18105
rect 4804 18096 4856 18148
rect 3608 18028 3660 18080
rect 5264 18071 5316 18080
rect 5264 18037 5273 18071
rect 5273 18037 5307 18071
rect 5307 18037 5316 18071
rect 5264 18028 5316 18037
rect 5356 18071 5408 18080
rect 5356 18037 5365 18071
rect 5365 18037 5399 18071
rect 5399 18037 5408 18071
rect 5356 18028 5408 18037
rect 5816 18096 5868 18148
rect 5540 18028 5592 18080
rect 5632 18071 5684 18080
rect 5632 18037 5641 18071
rect 5641 18037 5675 18071
rect 5675 18037 5684 18071
rect 5632 18028 5684 18037
rect 6644 18028 6696 18080
rect 8208 18232 8260 18284
rect 8668 18232 8720 18284
rect 11336 18300 11388 18352
rect 12808 18300 12860 18352
rect 15844 18300 15896 18352
rect 17316 18343 17368 18352
rect 17316 18309 17341 18343
rect 17341 18309 17368 18343
rect 19156 18368 19208 18420
rect 20352 18343 20404 18352
rect 17316 18300 17368 18309
rect 20352 18309 20361 18343
rect 20361 18309 20395 18343
rect 20395 18309 20404 18343
rect 20352 18300 20404 18309
rect 10876 18232 10928 18284
rect 10968 18275 11020 18284
rect 10968 18241 10977 18275
rect 10977 18241 11011 18275
rect 11011 18241 11020 18275
rect 10968 18232 11020 18241
rect 11428 18232 11480 18284
rect 8300 18164 8352 18216
rect 8392 18207 8444 18216
rect 8392 18173 8401 18207
rect 8401 18173 8435 18207
rect 8435 18173 8444 18207
rect 8392 18164 8444 18173
rect 8576 18096 8628 18148
rect 8300 18028 8352 18080
rect 8852 18207 8904 18216
rect 8852 18173 8861 18207
rect 8861 18173 8895 18207
rect 8895 18173 8904 18207
rect 8852 18164 8904 18173
rect 9220 18207 9272 18216
rect 9220 18173 9229 18207
rect 9229 18173 9263 18207
rect 9263 18173 9272 18207
rect 9220 18164 9272 18173
rect 10692 18164 10744 18216
rect 12624 18232 12676 18284
rect 15936 18275 15988 18284
rect 15936 18241 15945 18275
rect 15945 18241 15979 18275
rect 15979 18241 15988 18275
rect 15936 18232 15988 18241
rect 16212 18275 16264 18284
rect 16212 18241 16221 18275
rect 16221 18241 16255 18275
rect 16255 18241 16264 18275
rect 16212 18232 16264 18241
rect 18144 18275 18196 18284
rect 18144 18241 18153 18275
rect 18153 18241 18187 18275
rect 18187 18241 18196 18275
rect 18144 18232 18196 18241
rect 19064 18275 19116 18284
rect 19064 18241 19073 18275
rect 19073 18241 19107 18275
rect 19107 18241 19116 18275
rect 19064 18232 19116 18241
rect 20812 18411 20864 18420
rect 20812 18377 20821 18411
rect 20821 18377 20855 18411
rect 20855 18377 20864 18411
rect 20812 18368 20864 18377
rect 22008 18368 22060 18420
rect 24492 18411 24544 18420
rect 24492 18377 24501 18411
rect 24501 18377 24535 18411
rect 24535 18377 24544 18411
rect 24492 18368 24544 18377
rect 24676 18411 24728 18420
rect 24676 18377 24685 18411
rect 24685 18377 24719 18411
rect 24719 18377 24728 18411
rect 24676 18368 24728 18377
rect 25780 18411 25832 18420
rect 25780 18377 25789 18411
rect 25789 18377 25823 18411
rect 25823 18377 25832 18411
rect 25780 18368 25832 18377
rect 24860 18343 24912 18352
rect 24860 18309 24869 18343
rect 24869 18309 24903 18343
rect 24903 18309 24912 18343
rect 24860 18300 24912 18309
rect 9772 18028 9824 18080
rect 10600 18028 10652 18080
rect 14096 18207 14148 18216
rect 14096 18173 14105 18207
rect 14105 18173 14139 18207
rect 14139 18173 14148 18207
rect 14096 18164 14148 18173
rect 15568 18207 15620 18216
rect 15568 18173 15577 18207
rect 15577 18173 15611 18207
rect 15611 18173 15620 18207
rect 15568 18164 15620 18173
rect 14188 18028 14240 18080
rect 14280 18028 14332 18080
rect 22100 18275 22152 18284
rect 22100 18241 22109 18275
rect 22109 18241 22143 18275
rect 22143 18241 22152 18275
rect 22100 18232 22152 18241
rect 22376 18275 22428 18284
rect 22376 18241 22385 18275
rect 22385 18241 22419 18275
rect 22419 18241 22428 18275
rect 22376 18232 22428 18241
rect 24124 18232 24176 18284
rect 25136 18275 25188 18284
rect 25136 18241 25145 18275
rect 25145 18241 25179 18275
rect 25179 18241 25188 18275
rect 25136 18232 25188 18241
rect 25320 18275 25372 18284
rect 25320 18241 25329 18275
rect 25329 18241 25363 18275
rect 25363 18241 25372 18275
rect 25320 18232 25372 18241
rect 22744 18164 22796 18216
rect 23204 18164 23256 18216
rect 24032 18207 24084 18216
rect 24032 18173 24041 18207
rect 24041 18173 24075 18207
rect 24075 18173 24084 18207
rect 24032 18164 24084 18173
rect 25596 18232 25648 18284
rect 25872 18164 25924 18216
rect 17408 18028 17460 18080
rect 17500 18071 17552 18080
rect 17500 18037 17509 18071
rect 17509 18037 17543 18071
rect 17543 18037 17552 18071
rect 17500 18028 17552 18037
rect 19156 18028 19208 18080
rect 19524 18071 19576 18080
rect 19524 18037 19533 18071
rect 19533 18037 19567 18071
rect 19567 18037 19576 18071
rect 19524 18028 19576 18037
rect 20536 18071 20588 18080
rect 20536 18037 20545 18071
rect 20545 18037 20579 18071
rect 20579 18037 20588 18071
rect 20536 18028 20588 18037
rect 21732 18028 21784 18080
rect 25044 18028 25096 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 4068 17824 4120 17876
rect 4620 17824 4672 17876
rect 5356 17824 5408 17876
rect 5448 17824 5500 17876
rect 6000 17867 6052 17876
rect 6000 17833 6009 17867
rect 6009 17833 6043 17867
rect 6043 17833 6052 17867
rect 6000 17824 6052 17833
rect 6920 17824 6972 17876
rect 8392 17824 8444 17876
rect 8668 17824 8720 17876
rect 1860 17731 1912 17740
rect 1860 17697 1869 17731
rect 1869 17697 1903 17731
rect 1903 17697 1912 17731
rect 1860 17688 1912 17697
rect 3700 17620 3752 17672
rect 9864 17824 9916 17876
rect 15568 17824 15620 17876
rect 15936 17824 15988 17876
rect 18604 17867 18656 17876
rect 18604 17833 18613 17867
rect 18613 17833 18647 17867
rect 18647 17833 18656 17867
rect 18604 17824 18656 17833
rect 20536 17824 20588 17876
rect 22100 17824 22152 17876
rect 23388 17824 23440 17876
rect 25136 17824 25188 17876
rect 25320 17824 25372 17876
rect 4988 17688 5040 17740
rect 4620 17620 4672 17672
rect 4712 17663 4764 17672
rect 4712 17629 4721 17663
rect 4721 17629 4755 17663
rect 4755 17629 4764 17663
rect 4712 17620 4764 17629
rect 4896 17620 4948 17672
rect 5080 17663 5132 17672
rect 5080 17629 5084 17663
rect 5084 17629 5118 17663
rect 5118 17629 5132 17663
rect 5080 17620 5132 17629
rect 4712 17484 4764 17536
rect 5080 17484 5132 17536
rect 5264 17595 5316 17604
rect 5264 17561 5273 17595
rect 5273 17561 5307 17595
rect 5307 17561 5316 17595
rect 5264 17552 5316 17561
rect 5540 17663 5592 17672
rect 5540 17629 5549 17663
rect 5549 17629 5583 17663
rect 5583 17629 5592 17663
rect 5540 17620 5592 17629
rect 5724 17620 5776 17672
rect 5816 17663 5868 17672
rect 5816 17629 5825 17663
rect 5825 17629 5859 17663
rect 5859 17629 5868 17663
rect 5816 17620 5868 17629
rect 6184 17552 6236 17604
rect 9680 17756 9732 17808
rect 6552 17663 6604 17672
rect 6552 17629 6561 17663
rect 6561 17629 6595 17663
rect 6595 17629 6604 17663
rect 6552 17620 6604 17629
rect 6644 17663 6696 17672
rect 6644 17629 6653 17663
rect 6653 17629 6687 17663
rect 6687 17629 6696 17663
rect 6644 17620 6696 17629
rect 6828 17663 6880 17672
rect 6828 17629 6837 17663
rect 6837 17629 6871 17663
rect 6871 17629 6880 17663
rect 6828 17620 6880 17629
rect 7012 17620 7064 17672
rect 8392 17552 8444 17604
rect 9312 17688 9364 17740
rect 9128 17620 9180 17672
rect 10600 17731 10652 17740
rect 10600 17697 10609 17731
rect 10609 17697 10643 17731
rect 10643 17697 10652 17731
rect 10600 17688 10652 17697
rect 17868 17688 17920 17740
rect 20536 17688 20588 17740
rect 21732 17731 21784 17740
rect 21732 17697 21741 17731
rect 21741 17697 21775 17731
rect 21775 17697 21784 17731
rect 21732 17688 21784 17697
rect 22100 17688 22152 17740
rect 10876 17620 10928 17672
rect 10140 17552 10192 17604
rect 11244 17663 11296 17672
rect 11244 17629 11253 17663
rect 11253 17629 11287 17663
rect 11287 17629 11296 17663
rect 11244 17620 11296 17629
rect 11428 17663 11480 17672
rect 11428 17629 11437 17663
rect 11437 17629 11471 17663
rect 11471 17629 11480 17663
rect 11428 17620 11480 17629
rect 23388 17620 23440 17672
rect 11060 17552 11112 17604
rect 11980 17552 12032 17604
rect 15844 17552 15896 17604
rect 17408 17552 17460 17604
rect 10048 17527 10100 17536
rect 10048 17493 10057 17527
rect 10057 17493 10091 17527
rect 10091 17493 10100 17527
rect 10048 17484 10100 17493
rect 10232 17484 10284 17536
rect 12348 17484 12400 17536
rect 15568 17484 15620 17536
rect 16488 17484 16540 17536
rect 18512 17552 18564 17604
rect 19156 17552 19208 17604
rect 19432 17552 19484 17604
rect 21180 17552 21232 17604
rect 23940 17663 23992 17672
rect 23940 17629 23949 17663
rect 23949 17629 23983 17663
rect 23983 17629 23992 17663
rect 23940 17620 23992 17629
rect 24124 17663 24176 17672
rect 24124 17629 24133 17663
rect 24133 17629 24167 17663
rect 24167 17629 24176 17663
rect 24124 17620 24176 17629
rect 25320 17688 25372 17740
rect 26148 17688 26200 17740
rect 24676 17663 24728 17672
rect 24676 17629 24685 17663
rect 24685 17629 24719 17663
rect 24719 17629 24728 17663
rect 24676 17620 24728 17629
rect 25136 17663 25188 17672
rect 25136 17629 25145 17663
rect 25145 17629 25179 17663
rect 25179 17629 25188 17663
rect 25136 17620 25188 17629
rect 25596 17663 25648 17672
rect 25596 17629 25605 17663
rect 25605 17629 25639 17663
rect 25639 17629 25648 17663
rect 25596 17620 25648 17629
rect 26792 17595 26844 17604
rect 26792 17561 26801 17595
rect 26801 17561 26835 17595
rect 26835 17561 26844 17595
rect 26792 17552 26844 17561
rect 26884 17552 26936 17604
rect 18788 17484 18840 17536
rect 19248 17484 19300 17536
rect 22376 17484 22428 17536
rect 23204 17527 23256 17536
rect 23204 17493 23213 17527
rect 23213 17493 23247 17527
rect 23247 17493 23256 17527
rect 23204 17484 23256 17493
rect 23296 17484 23348 17536
rect 25044 17527 25096 17536
rect 25044 17493 25053 17527
rect 25053 17493 25087 17527
rect 25087 17493 25096 17527
rect 25044 17484 25096 17493
rect 25136 17484 25188 17536
rect 25780 17527 25832 17536
rect 25780 17493 25789 17527
rect 25789 17493 25823 17527
rect 25823 17493 25832 17527
rect 25780 17484 25832 17493
rect 25872 17484 25924 17536
rect 28264 17527 28316 17536
rect 28264 17493 28273 17527
rect 28273 17493 28307 17527
rect 28307 17493 28316 17527
rect 28264 17484 28316 17493
rect 4874 17382 4926 17434
rect 4938 17382 4990 17434
rect 5002 17382 5054 17434
rect 5066 17382 5118 17434
rect 5130 17382 5182 17434
rect 5264 17323 5316 17332
rect 5264 17289 5273 17323
rect 5273 17289 5307 17323
rect 5307 17289 5316 17323
rect 5264 17280 5316 17289
rect 5540 17280 5592 17332
rect 8760 17280 8812 17332
rect 5264 17144 5316 17196
rect 6000 17212 6052 17264
rect 6552 17212 6604 17264
rect 5448 17144 5500 17196
rect 8392 17212 8444 17264
rect 9220 17280 9272 17332
rect 10140 17323 10192 17332
rect 10140 17289 10149 17323
rect 10149 17289 10183 17323
rect 10183 17289 10192 17323
rect 10140 17280 10192 17289
rect 17408 17323 17460 17332
rect 17408 17289 17417 17323
rect 17417 17289 17451 17323
rect 17451 17289 17460 17323
rect 17408 17280 17460 17289
rect 18512 17280 18564 17332
rect 6920 17187 6972 17196
rect 6920 17153 6929 17187
rect 6929 17153 6963 17187
rect 6963 17153 6972 17187
rect 6920 17144 6972 17153
rect 7012 17187 7064 17196
rect 7012 17153 7021 17187
rect 7021 17153 7055 17187
rect 7055 17153 7064 17187
rect 7012 17144 7064 17153
rect 8484 17187 8536 17196
rect 8484 17153 8493 17187
rect 8493 17153 8527 17187
rect 8527 17153 8536 17187
rect 8484 17144 8536 17153
rect 10048 17212 10100 17264
rect 5724 17119 5776 17128
rect 5724 17085 5733 17119
rect 5733 17085 5767 17119
rect 5767 17085 5776 17119
rect 5724 17076 5776 17085
rect 6460 17008 6512 17060
rect 9312 17187 9364 17196
rect 9312 17153 9321 17187
rect 9321 17153 9355 17187
rect 9355 17153 9364 17187
rect 9312 17144 9364 17153
rect 9496 17187 9548 17196
rect 9496 17153 9505 17187
rect 9505 17153 9539 17187
rect 9539 17153 9548 17187
rect 9496 17144 9548 17153
rect 9772 17187 9824 17196
rect 9772 17153 9781 17187
rect 9781 17153 9815 17187
rect 9815 17153 9824 17187
rect 9772 17144 9824 17153
rect 11060 17212 11112 17264
rect 22284 17280 22336 17332
rect 23296 17280 23348 17332
rect 10232 17187 10284 17196
rect 10232 17153 10241 17187
rect 10241 17153 10275 17187
rect 10275 17153 10284 17187
rect 10232 17144 10284 17153
rect 12348 17187 12400 17196
rect 12348 17153 12357 17187
rect 12357 17153 12391 17187
rect 12391 17153 12400 17187
rect 12348 17144 12400 17153
rect 12440 17144 12492 17196
rect 12808 17144 12860 17196
rect 15844 17144 15896 17196
rect 16028 17144 16080 17196
rect 17500 17144 17552 17196
rect 18144 17144 18196 17196
rect 18512 17144 18564 17196
rect 18604 17144 18656 17196
rect 8760 17008 8812 17060
rect 10600 17008 10652 17060
rect 9588 16983 9640 16992
rect 9588 16949 9597 16983
rect 9597 16949 9631 16983
rect 9631 16949 9640 16983
rect 9588 16940 9640 16949
rect 12164 16983 12216 16992
rect 12164 16949 12173 16983
rect 12173 16949 12207 16983
rect 12207 16949 12216 16983
rect 12164 16940 12216 16949
rect 12808 16940 12860 16992
rect 13912 17119 13964 17128
rect 13912 17085 13921 17119
rect 13921 17085 13955 17119
rect 13955 17085 13964 17119
rect 13912 17076 13964 17085
rect 14188 17119 14240 17128
rect 14188 17085 14197 17119
rect 14197 17085 14231 17119
rect 14231 17085 14240 17119
rect 14188 17076 14240 17085
rect 19248 17187 19300 17196
rect 19248 17153 19257 17187
rect 19257 17153 19291 17187
rect 19291 17153 19300 17187
rect 19248 17144 19300 17153
rect 19432 17187 19484 17196
rect 19432 17153 19441 17187
rect 19441 17153 19475 17187
rect 19475 17153 19484 17187
rect 19432 17144 19484 17153
rect 20628 17144 20680 17196
rect 22652 17212 22704 17264
rect 26884 17212 26936 17264
rect 28080 17255 28132 17264
rect 28080 17221 28089 17255
rect 28089 17221 28123 17255
rect 28123 17221 28132 17255
rect 28080 17212 28132 17221
rect 25596 17187 25648 17196
rect 25596 17153 25605 17187
rect 25605 17153 25639 17187
rect 25639 17153 25648 17187
rect 25596 17144 25648 17153
rect 19524 17076 19576 17128
rect 19984 17076 20036 17128
rect 25412 17076 25464 17128
rect 25872 17076 25924 17128
rect 22468 17008 22520 17060
rect 14740 16940 14792 16992
rect 15476 16983 15528 16992
rect 15476 16949 15485 16983
rect 15485 16949 15519 16983
rect 15519 16949 15528 16983
rect 15476 16940 15528 16949
rect 17316 16940 17368 16992
rect 22284 16940 22336 16992
rect 22376 16983 22428 16992
rect 22376 16949 22385 16983
rect 22385 16949 22419 16983
rect 22419 16949 22428 16983
rect 22376 16940 22428 16949
rect 22560 16983 22612 16992
rect 22560 16949 22569 16983
rect 22569 16949 22603 16983
rect 22603 16949 22612 16983
rect 22560 16940 22612 16949
rect 23940 16940 23992 16992
rect 25044 16940 25096 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 4804 16736 4856 16788
rect 5632 16779 5684 16788
rect 5632 16745 5641 16779
rect 5641 16745 5675 16779
rect 5675 16745 5684 16779
rect 5632 16736 5684 16745
rect 8668 16736 8720 16788
rect 9312 16736 9364 16788
rect 15476 16736 15528 16788
rect 16212 16736 16264 16788
rect 19064 16736 19116 16788
rect 22652 16736 22704 16788
rect 25044 16779 25096 16788
rect 25044 16745 25053 16779
rect 25053 16745 25087 16779
rect 25087 16745 25096 16779
rect 25044 16736 25096 16745
rect 26792 16736 26844 16788
rect 4436 16600 4488 16652
rect 5448 16600 5500 16652
rect 6184 16600 6236 16652
rect 7748 16600 7800 16652
rect 10140 16600 10192 16652
rect 6000 16439 6052 16448
rect 6000 16405 6009 16439
rect 6009 16405 6043 16439
rect 6043 16405 6052 16439
rect 6000 16396 6052 16405
rect 6460 16575 6512 16584
rect 6460 16541 6469 16575
rect 6469 16541 6503 16575
rect 6503 16541 6512 16575
rect 6460 16532 6512 16541
rect 6552 16575 6604 16584
rect 6552 16541 6597 16575
rect 6597 16541 6604 16575
rect 6552 16532 6604 16541
rect 6736 16575 6788 16584
rect 6736 16541 6745 16575
rect 6745 16541 6779 16575
rect 6779 16541 6788 16575
rect 6736 16532 6788 16541
rect 9036 16532 9088 16584
rect 9588 16532 9640 16584
rect 11336 16532 11388 16584
rect 12440 16600 12492 16652
rect 14188 16600 14240 16652
rect 14740 16643 14792 16652
rect 14740 16609 14749 16643
rect 14749 16609 14783 16643
rect 14783 16609 14792 16643
rect 14740 16600 14792 16609
rect 23940 16600 23992 16652
rect 25136 16643 25188 16652
rect 25136 16609 25145 16643
rect 25145 16609 25179 16643
rect 25179 16609 25188 16643
rect 25136 16600 25188 16609
rect 25228 16643 25280 16652
rect 25228 16609 25237 16643
rect 25237 16609 25271 16643
rect 25271 16609 25280 16643
rect 25228 16600 25280 16609
rect 12808 16575 12860 16584
rect 12808 16541 12817 16575
rect 12817 16541 12851 16575
rect 12851 16541 12860 16575
rect 12808 16532 12860 16541
rect 14280 16532 14332 16584
rect 18052 16532 18104 16584
rect 22560 16532 22612 16584
rect 22652 16575 22704 16584
rect 22652 16541 22661 16575
rect 22661 16541 22695 16575
rect 22695 16541 22704 16575
rect 22652 16532 22704 16541
rect 8852 16464 8904 16516
rect 11152 16464 11204 16516
rect 12440 16507 12492 16516
rect 12440 16473 12449 16507
rect 12449 16473 12483 16507
rect 12483 16473 12492 16507
rect 12440 16464 12492 16473
rect 16488 16464 16540 16516
rect 8392 16396 8444 16448
rect 8944 16396 8996 16448
rect 11428 16396 11480 16448
rect 13176 16396 13228 16448
rect 13544 16396 13596 16448
rect 15108 16396 15160 16448
rect 16028 16396 16080 16448
rect 18696 16439 18748 16448
rect 18696 16405 18705 16439
rect 18705 16405 18739 16439
rect 18739 16405 18748 16439
rect 18696 16396 18748 16405
rect 22192 16439 22244 16448
rect 22192 16405 22201 16439
rect 22201 16405 22235 16439
rect 22235 16405 22244 16439
rect 22192 16396 22244 16405
rect 24676 16439 24728 16448
rect 24676 16405 24685 16439
rect 24685 16405 24719 16439
rect 24719 16405 24728 16439
rect 24676 16396 24728 16405
rect 24860 16396 24912 16448
rect 26608 16532 26660 16584
rect 26884 16668 26936 16720
rect 25504 16507 25556 16516
rect 25504 16473 25513 16507
rect 25513 16473 25547 16507
rect 25547 16473 25556 16507
rect 25504 16464 25556 16473
rect 28264 16600 28316 16652
rect 26976 16439 27028 16448
rect 26976 16405 26985 16439
rect 26985 16405 27019 16439
rect 27019 16405 27028 16439
rect 26976 16396 27028 16405
rect 4874 16294 4926 16346
rect 4938 16294 4990 16346
rect 5002 16294 5054 16346
rect 5066 16294 5118 16346
rect 5130 16294 5182 16346
rect 4436 16235 4488 16244
rect 4436 16201 4445 16235
rect 4445 16201 4479 16235
rect 4479 16201 4488 16235
rect 4436 16192 4488 16201
rect 4620 16192 4672 16244
rect 5540 16192 5592 16244
rect 6736 16192 6788 16244
rect 6920 16192 6972 16244
rect 8944 16192 8996 16244
rect 9220 16192 9272 16244
rect 9496 16192 9548 16244
rect 12808 16192 12860 16244
rect 12992 16192 13044 16244
rect 3700 16124 3752 16176
rect 6000 16124 6052 16176
rect 13728 16167 13780 16176
rect 8392 16099 8444 16108
rect 8392 16065 8401 16099
rect 8401 16065 8435 16099
rect 8435 16065 8444 16099
rect 8392 16056 8444 16065
rect 8852 16099 8904 16108
rect 8852 16065 8869 16099
rect 8869 16065 8904 16099
rect 8852 16056 8904 16065
rect 8944 16099 8996 16108
rect 8944 16065 8953 16099
rect 8953 16065 8987 16099
rect 8987 16065 8996 16099
rect 8944 16056 8996 16065
rect 9128 16099 9180 16108
rect 9128 16065 9137 16099
rect 9137 16065 9171 16099
rect 9171 16065 9180 16099
rect 9128 16056 9180 16065
rect 9220 16056 9272 16108
rect 7932 16031 7984 16040
rect 7932 15997 7950 16031
rect 7950 15997 7984 16031
rect 5356 15852 5408 15904
rect 7932 15988 7984 15997
rect 8024 16031 8076 16040
rect 8024 15997 8033 16031
rect 8033 15997 8067 16031
rect 8067 15997 8076 16031
rect 8024 15988 8076 15997
rect 8576 15988 8628 16040
rect 8484 15920 8536 15972
rect 9588 15988 9640 16040
rect 9772 16099 9824 16108
rect 9772 16065 9781 16099
rect 9781 16065 9815 16099
rect 9815 16065 9824 16099
rect 9772 16056 9824 16065
rect 12716 16099 12768 16108
rect 12716 16065 12725 16099
rect 12725 16065 12759 16099
rect 12759 16065 12768 16099
rect 12716 16056 12768 16065
rect 13728 16133 13737 16167
rect 13737 16133 13771 16167
rect 13771 16133 13780 16167
rect 13728 16124 13780 16133
rect 12992 16099 13044 16108
rect 12992 16065 13000 16099
rect 13000 16065 13034 16099
rect 13034 16065 13044 16099
rect 12992 16056 13044 16065
rect 13452 16099 13504 16108
rect 13452 16065 13461 16099
rect 13461 16065 13495 16099
rect 13495 16065 13504 16099
rect 13452 16056 13504 16065
rect 13544 16099 13596 16108
rect 13544 16065 13554 16099
rect 13554 16065 13588 16099
rect 13588 16065 13596 16099
rect 13544 16056 13596 16065
rect 16028 16192 16080 16244
rect 23940 16192 23992 16244
rect 24860 16235 24912 16244
rect 24860 16201 24869 16235
rect 24869 16201 24903 16235
rect 24903 16201 24912 16235
rect 24860 16192 24912 16201
rect 25504 16192 25556 16244
rect 25780 16235 25832 16244
rect 25780 16201 25789 16235
rect 25789 16201 25823 16235
rect 25823 16201 25832 16235
rect 25780 16192 25832 16201
rect 16304 16124 16356 16176
rect 16488 16124 16540 16176
rect 18788 16124 18840 16176
rect 22192 16124 22244 16176
rect 23388 16124 23440 16176
rect 9864 15988 9916 16040
rect 11428 15988 11480 16040
rect 14188 16056 14240 16108
rect 17868 16099 17920 16108
rect 17868 16065 17877 16099
rect 17877 16065 17911 16099
rect 17911 16065 17920 16099
rect 17868 16056 17920 16065
rect 20628 16056 20680 16108
rect 8300 15852 8352 15904
rect 8852 15852 8904 15904
rect 9404 15852 9456 15904
rect 11796 15852 11848 15904
rect 12532 15852 12584 15904
rect 13452 15852 13504 15904
rect 15016 16031 15068 16040
rect 15016 15997 15025 16031
rect 15025 15997 15059 16031
rect 15059 15997 15068 16031
rect 15016 15988 15068 15997
rect 15660 15988 15712 16040
rect 18236 15988 18288 16040
rect 20444 15988 20496 16040
rect 21364 16031 21416 16040
rect 21364 15997 21373 16031
rect 21373 15997 21407 16031
rect 21407 15997 21416 16031
rect 21364 15988 21416 15997
rect 21824 16031 21876 16040
rect 21824 15997 21833 16031
rect 21833 15997 21867 16031
rect 21867 15997 21876 16031
rect 21824 15988 21876 15997
rect 19156 15920 19208 15972
rect 25412 16056 25464 16108
rect 25596 16056 25648 16108
rect 26976 16056 27028 16108
rect 28356 16099 28408 16108
rect 28356 16065 28365 16099
rect 28365 16065 28399 16099
rect 28399 16065 28408 16099
rect 28356 16056 28408 16065
rect 15752 15852 15804 15904
rect 16672 15895 16724 15904
rect 16672 15861 16681 15895
rect 16681 15861 16715 15895
rect 16715 15861 16724 15895
rect 16672 15852 16724 15861
rect 19708 15895 19760 15904
rect 19708 15861 19717 15895
rect 19717 15861 19751 15895
rect 19751 15861 19760 15895
rect 19708 15852 19760 15861
rect 20904 15895 20956 15904
rect 20904 15861 20913 15895
rect 20913 15861 20947 15895
rect 20947 15861 20956 15895
rect 20904 15852 20956 15861
rect 26148 15852 26200 15904
rect 27620 15852 27672 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 9128 15648 9180 15700
rect 12440 15648 12492 15700
rect 13084 15648 13136 15700
rect 13912 15648 13964 15700
rect 15016 15648 15068 15700
rect 16212 15648 16264 15700
rect 18236 15691 18288 15700
rect 18236 15657 18245 15691
rect 18245 15657 18279 15691
rect 18279 15657 18288 15691
rect 18236 15648 18288 15657
rect 20628 15691 20680 15700
rect 20628 15657 20637 15691
rect 20637 15657 20671 15691
rect 20671 15657 20680 15691
rect 20628 15648 20680 15657
rect 20720 15648 20772 15700
rect 21180 15648 21232 15700
rect 21364 15691 21416 15700
rect 21364 15657 21373 15691
rect 21373 15657 21407 15691
rect 21407 15657 21416 15691
rect 21364 15648 21416 15657
rect 14096 15580 14148 15632
rect 15844 15623 15896 15632
rect 15844 15589 15853 15623
rect 15853 15589 15887 15623
rect 15887 15589 15896 15623
rect 15844 15580 15896 15589
rect 18696 15580 18748 15632
rect 22192 15648 22244 15700
rect 23388 15648 23440 15700
rect 8484 15512 8536 15564
rect 10048 15512 10100 15564
rect 11704 15512 11756 15564
rect 11796 15555 11848 15564
rect 11796 15521 11805 15555
rect 11805 15521 11839 15555
rect 11839 15521 11848 15555
rect 11796 15512 11848 15521
rect 9220 15487 9272 15496
rect 9220 15453 9229 15487
rect 9229 15453 9263 15487
rect 9263 15453 9272 15487
rect 9220 15444 9272 15453
rect 9772 15487 9824 15496
rect 9772 15453 9781 15487
rect 9781 15453 9815 15487
rect 9815 15453 9824 15487
rect 9772 15444 9824 15453
rect 9680 15376 9732 15428
rect 10416 15487 10468 15496
rect 10416 15453 10425 15487
rect 10425 15453 10459 15487
rect 10459 15453 10468 15487
rect 10416 15444 10468 15453
rect 11244 15444 11296 15496
rect 12164 15512 12216 15564
rect 12532 15444 12584 15496
rect 13176 15555 13228 15564
rect 13176 15521 13185 15555
rect 13185 15521 13219 15555
rect 13219 15521 13228 15555
rect 13176 15512 13228 15521
rect 16212 15512 16264 15564
rect 16672 15512 16724 15564
rect 13452 15487 13504 15496
rect 13452 15453 13461 15487
rect 13461 15453 13495 15487
rect 13495 15453 13504 15487
rect 13452 15444 13504 15453
rect 15200 15487 15252 15496
rect 15200 15453 15209 15487
rect 15209 15453 15243 15487
rect 15243 15453 15252 15487
rect 15200 15444 15252 15453
rect 15384 15487 15436 15496
rect 15384 15453 15391 15487
rect 15391 15453 15436 15487
rect 15384 15444 15436 15453
rect 15660 15487 15712 15496
rect 15660 15453 15674 15487
rect 15674 15453 15708 15487
rect 15708 15453 15712 15487
rect 15660 15444 15712 15453
rect 15936 15444 15988 15496
rect 19708 15512 19760 15564
rect 19432 15444 19484 15496
rect 19984 15487 20036 15496
rect 19984 15453 19993 15487
rect 19993 15453 20027 15487
rect 20027 15453 20036 15487
rect 19984 15444 20036 15453
rect 21824 15512 21876 15564
rect 25228 15512 25280 15564
rect 13728 15376 13780 15428
rect 15476 15419 15528 15428
rect 15476 15385 15485 15419
rect 15485 15385 15519 15419
rect 15519 15385 15528 15419
rect 15476 15376 15528 15385
rect 15752 15376 15804 15428
rect 18328 15376 18380 15428
rect 6552 15308 6604 15360
rect 7472 15308 7524 15360
rect 12532 15308 12584 15360
rect 18696 15419 18748 15428
rect 18696 15385 18731 15419
rect 18731 15385 18748 15419
rect 18696 15376 18748 15385
rect 18972 15308 19024 15360
rect 19340 15308 19392 15360
rect 20444 15487 20496 15496
rect 20444 15453 20458 15487
rect 20458 15453 20492 15487
rect 20492 15453 20496 15487
rect 20444 15444 20496 15453
rect 20352 15419 20404 15428
rect 20352 15385 20361 15419
rect 20361 15385 20395 15419
rect 20395 15385 20404 15419
rect 20352 15376 20404 15385
rect 21916 15487 21968 15496
rect 21916 15453 21925 15487
rect 21925 15453 21959 15487
rect 21959 15453 21968 15487
rect 21916 15444 21968 15453
rect 24124 15487 24176 15496
rect 24124 15453 24133 15487
rect 24133 15453 24167 15487
rect 24167 15453 24176 15487
rect 24124 15444 24176 15453
rect 26148 15691 26200 15700
rect 26148 15657 26157 15691
rect 26157 15657 26191 15691
rect 26191 15657 26200 15691
rect 26148 15648 26200 15657
rect 26608 15444 26660 15496
rect 27804 15487 27856 15496
rect 27804 15453 27813 15487
rect 27813 15453 27847 15487
rect 27847 15453 27856 15487
rect 27804 15444 27856 15453
rect 22100 15376 22152 15428
rect 22376 15419 22428 15428
rect 22376 15385 22385 15419
rect 22385 15385 22419 15419
rect 22419 15385 22428 15419
rect 22376 15376 22428 15385
rect 23388 15376 23440 15428
rect 24676 15419 24728 15428
rect 24676 15385 24685 15419
rect 24685 15385 24719 15419
rect 24719 15385 24728 15419
rect 24676 15376 24728 15385
rect 27896 15419 27948 15428
rect 21456 15308 21508 15360
rect 27896 15385 27905 15419
rect 27905 15385 27939 15419
rect 27939 15385 27948 15419
rect 27896 15376 27948 15385
rect 28172 15376 28224 15428
rect 27160 15308 27212 15360
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 7472 15104 7524 15156
rect 9036 15104 9088 15156
rect 9588 15147 9640 15156
rect 9588 15113 9597 15147
rect 9597 15113 9631 15147
rect 9631 15113 9640 15147
rect 9588 15104 9640 15113
rect 12624 15104 12676 15156
rect 12992 15104 13044 15156
rect 17868 15104 17920 15156
rect 6276 15036 6328 15088
rect 9496 15036 9548 15088
rect 12900 15036 12952 15088
rect 14096 15079 14148 15088
rect 14096 15045 14105 15079
rect 14105 15045 14139 15079
rect 14139 15045 14148 15079
rect 14096 15036 14148 15045
rect 7012 15011 7064 15020
rect 7012 14977 7021 15011
rect 7021 14977 7055 15011
rect 7055 14977 7064 15011
rect 7012 14968 7064 14977
rect 7748 14968 7800 15020
rect 8024 14968 8076 15020
rect 8392 15011 8444 15020
rect 8392 14977 8401 15011
rect 8401 14977 8435 15011
rect 8435 14977 8444 15011
rect 8392 14968 8444 14977
rect 7656 14900 7708 14952
rect 9128 14968 9180 15020
rect 9220 14943 9272 14952
rect 9220 14909 9229 14943
rect 9229 14909 9263 14943
rect 9263 14909 9272 14943
rect 9220 14900 9272 14909
rect 9588 14968 9640 15020
rect 9680 14968 9732 15020
rect 9772 15011 9824 15020
rect 9772 14977 9781 15011
rect 9781 14977 9815 15011
rect 9815 14977 9824 15011
rect 9772 14968 9824 14977
rect 10048 15011 10100 15020
rect 10048 14977 10057 15011
rect 10057 14977 10091 15011
rect 10091 14977 10100 15011
rect 10048 14968 10100 14977
rect 15844 15011 15896 15020
rect 15844 14977 15853 15011
rect 15853 14977 15887 15011
rect 15887 14977 15896 15011
rect 15844 14968 15896 14977
rect 16212 14968 16264 15020
rect 16488 14968 16540 15020
rect 17868 15011 17920 15020
rect 17868 14977 17877 15011
rect 17877 14977 17911 15011
rect 17911 14977 17920 15011
rect 17868 14968 17920 14977
rect 21916 15104 21968 15156
rect 22376 15104 22428 15156
rect 24124 15104 24176 15156
rect 28080 15104 28132 15156
rect 23388 15036 23440 15088
rect 27896 15079 27948 15088
rect 27896 15045 27905 15079
rect 27905 15045 27939 15079
rect 27939 15045 27948 15079
rect 27896 15036 27948 15045
rect 13360 14943 13412 14952
rect 13360 14909 13369 14943
rect 13369 14909 13403 14943
rect 13403 14909 13412 14943
rect 13360 14900 13412 14909
rect 13820 14900 13872 14952
rect 18236 14900 18288 14952
rect 18788 14900 18840 14952
rect 6552 14764 6604 14816
rect 8116 14832 8168 14884
rect 10324 14832 10376 14884
rect 7932 14764 7984 14816
rect 9864 14764 9916 14816
rect 10048 14764 10100 14816
rect 10416 14764 10468 14816
rect 15660 14807 15712 14816
rect 15660 14773 15669 14807
rect 15669 14773 15703 14807
rect 15703 14773 15712 14807
rect 15660 14764 15712 14773
rect 19432 14764 19484 14816
rect 22468 14968 22520 15020
rect 22652 15011 22704 15020
rect 22652 14977 22661 15011
rect 22661 14977 22695 15011
rect 22695 14977 22704 15011
rect 22652 14968 22704 14977
rect 20904 14900 20956 14952
rect 20628 14764 20680 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 5448 14399 5500 14408
rect 5448 14365 5457 14399
rect 5457 14365 5491 14399
rect 5491 14365 5500 14399
rect 5448 14356 5500 14365
rect 7012 14560 7064 14612
rect 8300 14560 8352 14612
rect 8392 14560 8444 14612
rect 8208 14492 8260 14544
rect 9772 14560 9824 14612
rect 11888 14560 11940 14612
rect 18236 14603 18288 14612
rect 18236 14569 18245 14603
rect 18245 14569 18279 14603
rect 18279 14569 18288 14603
rect 18236 14560 18288 14569
rect 5632 14424 5684 14476
rect 6644 14424 6696 14476
rect 7472 14467 7524 14476
rect 7472 14433 7481 14467
rect 7481 14433 7515 14467
rect 7515 14433 7524 14467
rect 7472 14424 7524 14433
rect 8300 14424 8352 14476
rect 5908 14356 5960 14408
rect 6920 14356 6972 14408
rect 7656 14399 7708 14408
rect 7656 14365 7665 14399
rect 7665 14365 7699 14399
rect 7699 14365 7708 14399
rect 7656 14356 7708 14365
rect 7748 14399 7800 14408
rect 7748 14365 7757 14399
rect 7757 14365 7791 14399
rect 7791 14365 7800 14399
rect 7748 14356 7800 14365
rect 7932 14399 7984 14408
rect 7932 14365 7941 14399
rect 7941 14365 7975 14399
rect 7975 14365 7984 14399
rect 7932 14356 7984 14365
rect 8116 14399 8168 14408
rect 8116 14365 8125 14399
rect 8125 14365 8159 14399
rect 8159 14365 8168 14399
rect 8116 14356 8168 14365
rect 8208 14399 8260 14408
rect 8208 14365 8217 14399
rect 8217 14365 8251 14399
rect 8251 14365 8260 14399
rect 8208 14356 8260 14365
rect 8484 14399 8536 14408
rect 8484 14365 8493 14399
rect 8493 14365 8527 14399
rect 8527 14365 8536 14399
rect 8484 14356 8536 14365
rect 8576 14399 8628 14408
rect 8576 14365 8585 14399
rect 8585 14365 8619 14399
rect 8619 14365 8628 14399
rect 8576 14356 8628 14365
rect 9496 14424 9548 14476
rect 8668 14288 8720 14340
rect 4712 14220 4764 14272
rect 5724 14220 5776 14272
rect 6276 14263 6328 14272
rect 6276 14229 6285 14263
rect 6285 14229 6319 14263
rect 6319 14229 6328 14263
rect 6276 14220 6328 14229
rect 6368 14263 6420 14272
rect 6368 14229 6377 14263
rect 6377 14229 6411 14263
rect 6411 14229 6420 14263
rect 6368 14220 6420 14229
rect 6828 14220 6880 14272
rect 8300 14220 8352 14272
rect 8760 14263 8812 14272
rect 8760 14229 8769 14263
rect 8769 14229 8803 14263
rect 8803 14229 8812 14263
rect 8760 14220 8812 14229
rect 9312 14399 9364 14408
rect 9312 14365 9321 14399
rect 9321 14365 9355 14399
rect 9355 14365 9364 14399
rect 9312 14356 9364 14365
rect 13360 14492 13412 14544
rect 9864 14424 9916 14476
rect 9404 14331 9456 14340
rect 9956 14399 10008 14408
rect 9956 14365 9965 14399
rect 9965 14365 9999 14399
rect 9999 14365 10008 14399
rect 9956 14356 10008 14365
rect 10048 14399 10100 14408
rect 10048 14365 10057 14399
rect 10057 14365 10091 14399
rect 10091 14365 10100 14399
rect 10048 14356 10100 14365
rect 10324 14399 10376 14408
rect 10324 14365 10333 14399
rect 10333 14365 10367 14399
rect 10367 14365 10376 14399
rect 10324 14356 10376 14365
rect 13820 14424 13872 14476
rect 27988 14424 28040 14476
rect 11336 14399 11388 14408
rect 11336 14365 11345 14399
rect 11345 14365 11379 14399
rect 11379 14365 11388 14399
rect 11336 14356 11388 14365
rect 11520 14399 11572 14408
rect 11520 14365 11529 14399
rect 11529 14365 11563 14399
rect 11563 14365 11572 14399
rect 11520 14356 11572 14365
rect 18144 14399 18196 14408
rect 9404 14297 9439 14331
rect 9439 14297 9456 14331
rect 9404 14288 9456 14297
rect 12900 14288 12952 14340
rect 12164 14220 12216 14272
rect 12808 14220 12860 14272
rect 13728 14288 13780 14340
rect 18144 14365 18153 14399
rect 18153 14365 18187 14399
rect 18187 14365 18196 14399
rect 18144 14356 18196 14365
rect 15292 14331 15344 14340
rect 15292 14297 15301 14331
rect 15301 14297 15335 14331
rect 15335 14297 15344 14331
rect 15292 14288 15344 14297
rect 18696 14399 18748 14408
rect 18696 14365 18705 14399
rect 18705 14365 18739 14399
rect 18739 14365 18748 14399
rect 18696 14356 18748 14365
rect 18880 14356 18932 14408
rect 19248 14399 19300 14408
rect 19248 14365 19257 14399
rect 19257 14365 19291 14399
rect 19291 14365 19300 14399
rect 19248 14356 19300 14365
rect 20628 14356 20680 14408
rect 26516 14399 26568 14408
rect 26516 14365 26525 14399
rect 26525 14365 26559 14399
rect 26559 14365 26568 14399
rect 26516 14356 26568 14365
rect 18972 14331 19024 14340
rect 18972 14297 18981 14331
rect 18981 14297 19015 14331
rect 19015 14297 19024 14331
rect 18972 14288 19024 14297
rect 28080 14288 28132 14340
rect 13452 14220 13504 14272
rect 16396 14220 16448 14272
rect 20996 14263 21048 14272
rect 20996 14229 21005 14263
rect 21005 14229 21039 14263
rect 21039 14229 21048 14263
rect 20996 14220 21048 14229
rect 27436 14220 27488 14272
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 5356 14016 5408 14068
rect 4712 13991 4764 14000
rect 4712 13957 4721 13991
rect 4721 13957 4755 13991
rect 4755 13957 4764 13991
rect 4712 13948 4764 13957
rect 6368 14059 6420 14068
rect 6368 14025 6377 14059
rect 6377 14025 6411 14059
rect 6411 14025 6420 14059
rect 6368 14016 6420 14025
rect 11888 14016 11940 14068
rect 5816 13880 5868 13932
rect 6552 13923 6604 13932
rect 6552 13889 6561 13923
rect 6561 13889 6595 13923
rect 6595 13889 6604 13923
rect 6552 13880 6604 13889
rect 6828 13880 6880 13932
rect 7012 13991 7064 14000
rect 7012 13957 7021 13991
rect 7021 13957 7055 13991
rect 7055 13957 7064 13991
rect 7012 13948 7064 13957
rect 6920 13855 6972 13864
rect 6920 13821 6929 13855
rect 6929 13821 6963 13855
rect 6963 13821 6972 13855
rect 6920 13812 6972 13821
rect 7748 13948 7800 14000
rect 8760 13948 8812 14000
rect 8944 13948 8996 14000
rect 10140 13948 10192 14000
rect 16488 14059 16540 14068
rect 16488 14025 16497 14059
rect 16497 14025 16531 14059
rect 16531 14025 16540 14059
rect 16488 14016 16540 14025
rect 18972 14059 19024 14068
rect 18972 14025 18981 14059
rect 18981 14025 19015 14059
rect 19015 14025 19024 14059
rect 18972 14016 19024 14025
rect 19984 14016 20036 14068
rect 20628 14016 20680 14068
rect 6276 13744 6328 13796
rect 6828 13744 6880 13796
rect 8392 13880 8444 13932
rect 11336 13880 11388 13932
rect 12624 13991 12676 14000
rect 12624 13957 12633 13991
rect 12633 13957 12667 13991
rect 12667 13957 12676 13991
rect 12624 13948 12676 13957
rect 12808 13991 12860 14000
rect 12808 13957 12817 13991
rect 12817 13957 12851 13991
rect 12851 13957 12860 13991
rect 12808 13948 12860 13957
rect 12256 13880 12308 13932
rect 8300 13812 8352 13864
rect 11520 13812 11572 13864
rect 16304 13948 16356 14000
rect 18696 13948 18748 14000
rect 22100 13991 22152 14000
rect 22100 13957 22109 13991
rect 22109 13957 22143 13991
rect 22143 13957 22152 13991
rect 22100 13948 22152 13957
rect 12164 13744 12216 13796
rect 12900 13744 12952 13796
rect 13544 13880 13596 13932
rect 13820 13880 13872 13932
rect 17684 13923 17736 13932
rect 17684 13889 17693 13923
rect 17693 13889 17727 13923
rect 17727 13889 17736 13923
rect 17684 13880 17736 13889
rect 19432 13880 19484 13932
rect 21916 13880 21968 13932
rect 22192 13923 22244 13932
rect 22192 13889 22201 13923
rect 22201 13889 22235 13923
rect 22235 13889 22244 13923
rect 22192 13880 22244 13889
rect 26516 14016 26568 14068
rect 27528 14016 27580 14068
rect 28264 14059 28316 14068
rect 28264 14025 28273 14059
rect 28273 14025 28307 14059
rect 28307 14025 28316 14059
rect 28264 14016 28316 14025
rect 27068 13948 27120 14000
rect 13728 13812 13780 13864
rect 15660 13812 15712 13864
rect 16580 13812 16632 13864
rect 18144 13812 18196 13864
rect 19156 13812 19208 13864
rect 20996 13812 21048 13864
rect 25504 13880 25556 13932
rect 27436 13880 27488 13932
rect 27988 13923 28040 13932
rect 27988 13889 27997 13923
rect 27997 13889 28031 13923
rect 28031 13889 28040 13923
rect 27988 13880 28040 13889
rect 18880 13744 18932 13796
rect 13360 13676 13412 13728
rect 17592 13676 17644 13728
rect 19064 13676 19116 13728
rect 25412 13812 25464 13864
rect 27344 13855 27396 13864
rect 27344 13821 27353 13855
rect 27353 13821 27387 13855
rect 27387 13821 27396 13855
rect 27344 13812 27396 13821
rect 22100 13744 22152 13796
rect 27620 13744 27672 13796
rect 22008 13676 22060 13728
rect 24860 13676 24912 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 6828 13515 6880 13524
rect 6828 13481 6837 13515
rect 6837 13481 6871 13515
rect 6871 13481 6880 13515
rect 6828 13472 6880 13481
rect 15936 13515 15988 13524
rect 15936 13481 15945 13515
rect 15945 13481 15979 13515
rect 15979 13481 15988 13515
rect 15936 13472 15988 13481
rect 16580 13472 16632 13524
rect 16488 13404 16540 13456
rect 5356 13336 5408 13388
rect 15200 13268 15252 13320
rect 15660 13336 15712 13388
rect 5632 13200 5684 13252
rect 4620 13132 4672 13184
rect 5816 13200 5868 13252
rect 14464 13200 14516 13252
rect 15476 13268 15528 13320
rect 17592 13379 17644 13388
rect 17592 13345 17601 13379
rect 17601 13345 17635 13379
rect 17635 13345 17644 13379
rect 17592 13336 17644 13345
rect 19248 13336 19300 13388
rect 26516 13379 26568 13388
rect 26516 13345 26525 13379
rect 26525 13345 26559 13379
rect 26559 13345 26568 13379
rect 26516 13336 26568 13345
rect 27804 13336 27856 13388
rect 21548 13311 21600 13320
rect 21548 13277 21557 13311
rect 21557 13277 21591 13311
rect 21591 13277 21600 13311
rect 21548 13268 21600 13277
rect 17132 13200 17184 13252
rect 21824 13243 21876 13252
rect 21824 13209 21833 13243
rect 21833 13209 21867 13243
rect 21867 13209 21876 13243
rect 21824 13200 21876 13209
rect 23204 13200 23256 13252
rect 15752 13132 15804 13184
rect 22192 13132 22244 13184
rect 27804 13200 27856 13252
rect 23388 13175 23440 13184
rect 23388 13141 23397 13175
rect 23397 13141 23431 13175
rect 23431 13141 23440 13175
rect 23388 13132 23440 13141
rect 26976 13132 27028 13184
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 12256 12860 12308 12912
rect 12900 12928 12952 12980
rect 13728 12928 13780 12980
rect 15384 12928 15436 12980
rect 15844 12928 15896 12980
rect 17684 12928 17736 12980
rect 21824 12971 21876 12980
rect 21824 12937 21833 12971
rect 21833 12937 21867 12971
rect 21867 12937 21876 12971
rect 21824 12928 21876 12937
rect 11612 12792 11664 12844
rect 11704 12724 11756 12776
rect 12348 12724 12400 12776
rect 10968 12656 11020 12708
rect 15476 12860 15528 12912
rect 13084 12792 13136 12844
rect 13820 12835 13872 12844
rect 13820 12801 13829 12835
rect 13829 12801 13863 12835
rect 13863 12801 13872 12835
rect 13820 12792 13872 12801
rect 15660 12835 15712 12844
rect 15660 12801 15669 12835
rect 15669 12801 15703 12835
rect 15703 12801 15712 12835
rect 15660 12792 15712 12801
rect 13268 12724 13320 12776
rect 13544 12724 13596 12776
rect 14096 12767 14148 12776
rect 14096 12733 14105 12767
rect 14105 12733 14139 12767
rect 14139 12733 14148 12767
rect 14096 12724 14148 12733
rect 14556 12724 14608 12776
rect 15844 12792 15896 12844
rect 16580 12792 16632 12844
rect 16488 12724 16540 12776
rect 5908 12588 5960 12640
rect 11060 12588 11112 12640
rect 11428 12588 11480 12640
rect 12440 12588 12492 12640
rect 12808 12588 12860 12640
rect 18696 12860 18748 12912
rect 19156 12792 19208 12844
rect 21180 12792 21232 12844
rect 22008 12835 22060 12844
rect 22008 12801 22017 12835
rect 22017 12801 22051 12835
rect 22051 12801 22060 12835
rect 22008 12792 22060 12801
rect 23388 12860 23440 12912
rect 26792 12860 26844 12912
rect 27436 12903 27488 12912
rect 27436 12869 27445 12903
rect 27445 12869 27479 12903
rect 27479 12869 27488 12903
rect 27436 12860 27488 12869
rect 18420 12724 18472 12776
rect 19708 12767 19760 12776
rect 19708 12733 19717 12767
rect 19717 12733 19751 12767
rect 19751 12733 19760 12767
rect 19708 12724 19760 12733
rect 18880 12656 18932 12708
rect 22560 12792 22612 12844
rect 22652 12724 22704 12776
rect 23296 12835 23348 12844
rect 23296 12801 23305 12835
rect 23305 12801 23339 12835
rect 23339 12801 23348 12835
rect 23296 12792 23348 12801
rect 26516 12792 26568 12844
rect 26608 12792 26660 12844
rect 22744 12656 22796 12708
rect 24216 12724 24268 12776
rect 27528 12724 27580 12776
rect 28080 12835 28132 12844
rect 28080 12801 28089 12835
rect 28089 12801 28123 12835
rect 28123 12801 28132 12835
rect 28080 12792 28132 12801
rect 28356 12835 28408 12844
rect 28356 12801 28365 12835
rect 28365 12801 28399 12835
rect 28399 12801 28408 12835
rect 28356 12792 28408 12801
rect 18420 12588 18472 12640
rect 18972 12631 19024 12640
rect 18972 12597 18981 12631
rect 18981 12597 19015 12631
rect 19015 12597 19024 12631
rect 18972 12588 19024 12597
rect 20720 12588 20772 12640
rect 22284 12588 22336 12640
rect 23480 12631 23532 12640
rect 23480 12597 23489 12631
rect 23489 12597 23523 12631
rect 23523 12597 23532 12631
rect 23480 12588 23532 12597
rect 24676 12631 24728 12640
rect 24676 12597 24685 12631
rect 24685 12597 24719 12631
rect 24719 12597 24728 12631
rect 24676 12588 24728 12597
rect 26884 12588 26936 12640
rect 27160 12631 27212 12640
rect 27160 12597 27169 12631
rect 27169 12597 27203 12631
rect 27203 12597 27212 12631
rect 27160 12588 27212 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 5724 12384 5776 12436
rect 12532 12384 12584 12436
rect 12900 12384 12952 12436
rect 13176 12384 13228 12436
rect 10876 12316 10928 12368
rect 4804 12180 4856 12232
rect 5816 12180 5868 12232
rect 6184 12180 6236 12232
rect 5448 12155 5500 12164
rect 5448 12121 5457 12155
rect 5457 12121 5491 12155
rect 5491 12121 5500 12155
rect 5448 12112 5500 12121
rect 5540 12155 5592 12164
rect 5540 12121 5549 12155
rect 5549 12121 5583 12155
rect 5583 12121 5592 12155
rect 5540 12112 5592 12121
rect 5908 12044 5960 12096
rect 6000 12087 6052 12096
rect 6000 12053 6009 12087
rect 6009 12053 6043 12087
rect 6043 12053 6052 12087
rect 6000 12044 6052 12053
rect 9220 12044 9272 12096
rect 10324 12180 10376 12232
rect 10784 12180 10836 12232
rect 11336 12223 11388 12232
rect 11336 12189 11340 12223
rect 11340 12189 11374 12223
rect 11374 12189 11388 12223
rect 11336 12180 11388 12189
rect 11428 12223 11480 12232
rect 11428 12189 11437 12223
rect 11437 12189 11471 12223
rect 11471 12189 11480 12223
rect 11428 12180 11480 12189
rect 11704 12223 11756 12232
rect 11704 12189 11712 12223
rect 11712 12189 11746 12223
rect 11746 12189 11756 12223
rect 11704 12180 11756 12189
rect 12716 12316 12768 12368
rect 13636 12316 13688 12368
rect 14096 12384 14148 12436
rect 18880 12384 18932 12436
rect 19156 12384 19208 12436
rect 18420 12316 18472 12368
rect 20628 12384 20680 12436
rect 23296 12384 23348 12436
rect 12072 12291 12124 12300
rect 12072 12257 12081 12291
rect 12081 12257 12115 12291
rect 12115 12257 12124 12291
rect 12072 12248 12124 12257
rect 12164 12248 12216 12300
rect 15660 12248 15712 12300
rect 18972 12248 19024 12300
rect 11980 12223 12032 12232
rect 11980 12189 11989 12223
rect 11989 12189 12023 12223
rect 12023 12189 12032 12223
rect 11980 12180 12032 12189
rect 12256 12223 12308 12232
rect 12256 12189 12265 12223
rect 12265 12189 12299 12223
rect 12299 12189 12308 12223
rect 12256 12180 12308 12189
rect 12348 12223 12400 12232
rect 12348 12189 12357 12223
rect 12357 12189 12391 12223
rect 12391 12189 12400 12223
rect 12348 12180 12400 12189
rect 11244 12112 11296 12164
rect 11520 12155 11572 12164
rect 11520 12121 11529 12155
rect 11529 12121 11563 12155
rect 11563 12121 11572 12155
rect 11520 12112 11572 12121
rect 12256 12044 12308 12096
rect 12716 12180 12768 12232
rect 12808 12223 12860 12232
rect 12808 12189 12817 12223
rect 12817 12189 12851 12223
rect 12851 12189 12860 12223
rect 12808 12180 12860 12189
rect 13084 12223 13136 12232
rect 13084 12189 13093 12223
rect 13093 12189 13127 12223
rect 13127 12189 13136 12223
rect 13084 12180 13136 12189
rect 13268 12223 13320 12232
rect 13268 12189 13277 12223
rect 13277 12189 13311 12223
rect 13311 12189 13320 12223
rect 13268 12180 13320 12189
rect 13360 12223 13412 12232
rect 13360 12189 13369 12223
rect 13369 12189 13403 12223
rect 13403 12189 13412 12223
rect 13360 12180 13412 12189
rect 14280 12180 14332 12232
rect 14464 12223 14516 12232
rect 14464 12189 14473 12223
rect 14473 12189 14507 12223
rect 14507 12189 14516 12223
rect 14464 12180 14516 12189
rect 14556 12223 14608 12232
rect 14556 12189 14565 12223
rect 14565 12189 14599 12223
rect 14599 12189 14608 12223
rect 14556 12180 14608 12189
rect 15384 12180 15436 12232
rect 18880 12223 18932 12232
rect 18880 12189 18889 12223
rect 18889 12189 18923 12223
rect 18923 12189 18932 12223
rect 18880 12180 18932 12189
rect 20996 12223 21048 12232
rect 20996 12189 21005 12223
rect 21005 12189 21039 12223
rect 21039 12189 21048 12223
rect 20996 12180 21048 12189
rect 21548 12180 21600 12232
rect 13176 12112 13228 12164
rect 14740 12112 14792 12164
rect 20260 12112 20312 12164
rect 20628 12112 20680 12164
rect 21824 12223 21876 12232
rect 21824 12189 21834 12223
rect 21834 12189 21868 12223
rect 21868 12189 21876 12223
rect 21824 12180 21876 12189
rect 22376 12248 22428 12300
rect 24400 12248 24452 12300
rect 26240 12291 26292 12300
rect 26240 12257 26249 12291
rect 26249 12257 26283 12291
rect 26283 12257 26292 12291
rect 26240 12248 26292 12257
rect 26516 12248 26568 12300
rect 22192 12223 22244 12232
rect 22192 12189 22206 12223
rect 22206 12189 22240 12223
rect 22240 12189 22244 12223
rect 22192 12180 22244 12189
rect 12992 12044 13044 12096
rect 13544 12044 13596 12096
rect 15476 12044 15528 12096
rect 18696 12044 18748 12096
rect 22468 12112 22520 12164
rect 22744 12155 22796 12164
rect 22744 12121 22753 12155
rect 22753 12121 22787 12155
rect 22787 12121 22796 12155
rect 22744 12112 22796 12121
rect 22192 12044 22244 12096
rect 23388 12044 23440 12096
rect 25504 12112 25556 12164
rect 24216 12087 24268 12096
rect 24216 12053 24225 12087
rect 24225 12053 24259 12087
rect 24259 12053 24268 12087
rect 24216 12044 24268 12053
rect 27896 12112 27948 12164
rect 27160 12044 27212 12096
rect 28172 12044 28224 12096
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 5356 11840 5408 11892
rect 7748 11840 7800 11892
rect 4620 11772 4672 11824
rect 6920 11772 6972 11824
rect 8208 11772 8260 11824
rect 13636 11840 13688 11892
rect 18512 11840 18564 11892
rect 3608 11679 3660 11688
rect 3608 11645 3617 11679
rect 3617 11645 3651 11679
rect 3651 11645 3660 11679
rect 3608 11636 3660 11645
rect 5816 11679 5868 11688
rect 5816 11645 5825 11679
rect 5825 11645 5859 11679
rect 5859 11645 5868 11679
rect 5816 11636 5868 11645
rect 6092 11747 6144 11756
rect 6092 11713 6101 11747
rect 6101 11713 6135 11747
rect 6135 11713 6144 11747
rect 6092 11704 6144 11713
rect 6368 11704 6420 11756
rect 6276 11636 6328 11688
rect 6552 11704 6604 11756
rect 7012 11636 7064 11688
rect 8024 11704 8076 11756
rect 7840 11636 7892 11688
rect 5172 11543 5224 11552
rect 5172 11509 5181 11543
rect 5181 11509 5215 11543
rect 5215 11509 5224 11543
rect 5172 11500 5224 11509
rect 5724 11500 5776 11552
rect 7104 11500 7156 11552
rect 8300 11543 8352 11552
rect 8300 11509 8309 11543
rect 8309 11509 8343 11543
rect 8343 11509 8352 11543
rect 8300 11500 8352 11509
rect 8944 11500 8996 11552
rect 9864 11679 9916 11688
rect 9864 11645 9873 11679
rect 9873 11645 9907 11679
rect 9907 11645 9916 11679
rect 9864 11636 9916 11645
rect 10416 11636 10468 11688
rect 10968 11704 11020 11756
rect 13820 11772 13872 11824
rect 18696 11815 18748 11824
rect 18696 11781 18705 11815
rect 18705 11781 18739 11815
rect 18739 11781 18748 11815
rect 18696 11772 18748 11781
rect 18880 11840 18932 11892
rect 12992 11747 13044 11756
rect 12992 11713 13001 11747
rect 13001 11713 13035 11747
rect 13035 11713 13044 11747
rect 12992 11704 13044 11713
rect 13176 11747 13228 11756
rect 13176 11713 13185 11747
rect 13185 11713 13219 11747
rect 13219 11713 13228 11747
rect 13176 11704 13228 11713
rect 13268 11747 13320 11756
rect 13268 11713 13277 11747
rect 13277 11713 13311 11747
rect 13311 11713 13320 11747
rect 13268 11704 13320 11713
rect 14372 11704 14424 11756
rect 18420 11747 18472 11756
rect 18420 11713 18429 11747
rect 18429 11713 18463 11747
rect 18463 11713 18472 11747
rect 18420 11704 18472 11713
rect 18604 11747 18656 11756
rect 18604 11713 18611 11747
rect 18611 11713 18656 11747
rect 18604 11704 18656 11713
rect 19708 11840 19760 11892
rect 20260 11840 20312 11892
rect 21456 11840 21508 11892
rect 22652 11883 22704 11892
rect 22652 11849 22661 11883
rect 22661 11849 22695 11883
rect 22695 11849 22704 11883
rect 22652 11840 22704 11849
rect 25504 11840 25556 11892
rect 20720 11772 20772 11824
rect 23388 11772 23440 11824
rect 26240 11772 26292 11824
rect 27344 11883 27396 11892
rect 27344 11849 27353 11883
rect 27353 11849 27387 11883
rect 27387 11849 27396 11883
rect 27344 11840 27396 11849
rect 22284 11704 22336 11756
rect 22376 11747 22428 11756
rect 22376 11713 22385 11747
rect 22385 11713 22419 11747
rect 22419 11713 22428 11747
rect 22376 11704 22428 11713
rect 24400 11747 24452 11756
rect 24400 11713 24409 11747
rect 24409 11713 24443 11747
rect 24443 11713 24452 11747
rect 24400 11704 24452 11713
rect 27896 11772 27948 11824
rect 26884 11704 26936 11756
rect 27160 11747 27212 11756
rect 27160 11713 27169 11747
rect 27169 11713 27203 11747
rect 27203 11713 27212 11747
rect 27160 11704 27212 11713
rect 28356 11747 28408 11756
rect 28356 11713 28365 11747
rect 28365 11713 28399 11747
rect 28399 11713 28408 11747
rect 28356 11704 28408 11713
rect 13084 11636 13136 11688
rect 13728 11636 13780 11688
rect 17868 11636 17920 11688
rect 20260 11636 20312 11688
rect 11060 11568 11112 11620
rect 13268 11568 13320 11620
rect 11704 11500 11756 11552
rect 11980 11500 12032 11552
rect 12532 11500 12584 11552
rect 15200 11568 15252 11620
rect 13544 11500 13596 11552
rect 19248 11500 19300 11552
rect 20996 11636 21048 11688
rect 27436 11636 27488 11688
rect 21548 11568 21600 11620
rect 22652 11568 22704 11620
rect 22560 11500 22612 11552
rect 25044 11543 25096 11552
rect 25044 11509 25053 11543
rect 25053 11509 25087 11543
rect 25087 11509 25096 11543
rect 25044 11500 25096 11509
rect 26516 11500 26568 11552
rect 27068 11500 27120 11552
rect 27344 11500 27396 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 3608 11296 3660 11348
rect 5448 11296 5500 11348
rect 8024 11296 8076 11348
rect 6644 11228 6696 11280
rect 5724 11203 5776 11212
rect 5724 11169 5733 11203
rect 5733 11169 5767 11203
rect 5767 11169 5776 11203
rect 5724 11160 5776 11169
rect 5816 11160 5868 11212
rect 6736 11203 6788 11212
rect 6736 11169 6745 11203
rect 6745 11169 6779 11203
rect 6779 11169 6788 11203
rect 6736 11160 6788 11169
rect 6920 11203 6972 11212
rect 6920 11169 6929 11203
rect 6929 11169 6963 11203
rect 6963 11169 6972 11203
rect 6920 11160 6972 11169
rect 5172 11092 5224 11144
rect 6184 11092 6236 11144
rect 6276 11135 6328 11144
rect 6276 11101 6285 11135
rect 6285 11101 6319 11135
rect 6319 11101 6328 11135
rect 6276 11092 6328 11101
rect 6552 11135 6604 11144
rect 6552 11101 6561 11135
rect 6561 11101 6595 11135
rect 6595 11101 6604 11135
rect 6552 11092 6604 11101
rect 7840 11135 7892 11144
rect 7840 11101 7849 11135
rect 7849 11101 7883 11135
rect 7883 11101 7892 11135
rect 7840 11092 7892 11101
rect 10784 11339 10836 11348
rect 10784 11305 10793 11339
rect 10793 11305 10827 11339
rect 10827 11305 10836 11339
rect 10784 11296 10836 11305
rect 12072 11296 12124 11348
rect 12624 11296 12676 11348
rect 12808 11296 12860 11348
rect 11060 11228 11112 11280
rect 12256 11228 12308 11280
rect 12532 11228 12584 11280
rect 8944 11203 8996 11212
rect 8944 11169 8953 11203
rect 8953 11169 8987 11203
rect 8987 11169 8996 11203
rect 8944 11160 8996 11169
rect 9220 11203 9272 11212
rect 9220 11169 9229 11203
rect 9229 11169 9263 11203
rect 9263 11169 9272 11203
rect 9220 11160 9272 11169
rect 11520 11160 11572 11212
rect 12992 11228 13044 11280
rect 6460 11024 6512 11076
rect 7012 11024 7064 11076
rect 7748 11067 7800 11076
rect 7748 11033 7757 11067
rect 7757 11033 7791 11067
rect 7791 11033 7800 11067
rect 7748 11024 7800 11033
rect 10876 11024 10928 11076
rect 11428 11024 11480 11076
rect 12164 11135 12216 11144
rect 12164 11101 12173 11135
rect 12173 11101 12207 11135
rect 12207 11101 12216 11135
rect 12164 11092 12216 11101
rect 12256 11135 12308 11144
rect 12256 11101 12265 11135
rect 12265 11101 12299 11135
rect 12299 11101 12308 11135
rect 12256 11092 12308 11101
rect 12808 11203 12860 11212
rect 12808 11169 12817 11203
rect 12817 11169 12851 11203
rect 12851 11169 12860 11203
rect 13360 11339 13412 11348
rect 13360 11305 13369 11339
rect 13369 11305 13403 11339
rect 13403 11305 13412 11339
rect 13360 11296 13412 11305
rect 13636 11296 13688 11348
rect 16396 11296 16448 11348
rect 20444 11296 20496 11348
rect 20628 11296 20680 11348
rect 14372 11228 14424 11280
rect 12808 11160 12860 11169
rect 13268 11160 13320 11212
rect 15292 11228 15344 11280
rect 16764 11228 16816 11280
rect 18512 11228 18564 11280
rect 12716 11135 12768 11144
rect 12716 11101 12725 11135
rect 12725 11101 12759 11135
rect 12759 11101 12768 11135
rect 12716 11092 12768 11101
rect 4804 10999 4856 11008
rect 4804 10965 4813 10999
rect 4813 10965 4847 10999
rect 4847 10965 4856 10999
rect 4804 10956 4856 10965
rect 10968 10956 11020 11008
rect 11520 10999 11572 11008
rect 11520 10965 11529 10999
rect 11529 10965 11563 10999
rect 11563 10965 11572 10999
rect 11520 10956 11572 10965
rect 12072 10956 12124 11008
rect 12532 11067 12584 11076
rect 12532 11033 12541 11067
rect 12541 11033 12575 11067
rect 12575 11033 12584 11067
rect 12532 11024 12584 11033
rect 13268 11067 13320 11076
rect 13268 11033 13277 11067
rect 13277 11033 13311 11067
rect 13311 11033 13320 11067
rect 13268 11024 13320 11033
rect 13084 10999 13136 11008
rect 13084 10965 13111 10999
rect 13111 10965 13136 10999
rect 13084 10956 13136 10965
rect 14004 11092 14056 11144
rect 14372 11135 14424 11144
rect 14372 11101 14381 11135
rect 14381 11101 14415 11135
rect 14415 11101 14424 11135
rect 15384 11160 15436 11212
rect 18144 11160 18196 11212
rect 14372 11092 14424 11101
rect 14648 11135 14700 11144
rect 14648 11101 14657 11135
rect 14657 11101 14691 11135
rect 14691 11101 14700 11135
rect 14648 11092 14700 11101
rect 17040 11092 17092 11144
rect 17776 11092 17828 11144
rect 19524 11135 19576 11144
rect 19524 11101 19533 11135
rect 19533 11101 19567 11135
rect 19567 11101 19576 11135
rect 19524 11092 19576 11101
rect 20536 11135 20588 11144
rect 20536 11101 20545 11135
rect 20545 11101 20579 11135
rect 20579 11101 20588 11135
rect 20536 11092 20588 11101
rect 21180 11339 21232 11348
rect 21180 11305 21189 11339
rect 21189 11305 21223 11339
rect 21223 11305 21232 11339
rect 21180 11296 21232 11305
rect 22376 11339 22428 11348
rect 22376 11305 22385 11339
rect 22385 11305 22419 11339
rect 22419 11305 22428 11339
rect 22376 11296 22428 11305
rect 22192 11228 22244 11280
rect 13820 11024 13872 11076
rect 13912 10956 13964 11008
rect 14096 10999 14148 11008
rect 14096 10965 14105 10999
rect 14105 10965 14139 10999
rect 14139 10965 14148 10999
rect 14096 10956 14148 10965
rect 15200 11024 15252 11076
rect 15752 11067 15804 11076
rect 15752 11033 15761 11067
rect 15761 11033 15795 11067
rect 15795 11033 15804 11067
rect 15752 11024 15804 11033
rect 17132 11024 17184 11076
rect 17408 11024 17460 11076
rect 17868 11024 17920 11076
rect 18696 11024 18748 11076
rect 21548 11092 21600 11144
rect 21916 11160 21968 11212
rect 22468 11160 22520 11212
rect 24400 11160 24452 11212
rect 26240 11160 26292 11212
rect 26608 11203 26660 11212
rect 26608 11169 26617 11203
rect 26617 11169 26651 11203
rect 26651 11169 26660 11203
rect 26608 11160 26660 11169
rect 28080 11203 28132 11212
rect 28080 11169 28089 11203
rect 28089 11169 28123 11203
rect 28123 11169 28132 11203
rect 28080 11160 28132 11169
rect 14648 10956 14700 11008
rect 15568 10956 15620 11008
rect 22284 10956 22336 11008
rect 23388 11024 23440 11076
rect 23940 11067 23992 11076
rect 23940 11033 23949 11067
rect 23949 11033 23983 11067
rect 23983 11033 23992 11067
rect 23940 11024 23992 11033
rect 27896 11024 27948 11076
rect 23112 10956 23164 11008
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 4804 10752 4856 10804
rect 6552 10795 6604 10804
rect 6552 10761 6561 10795
rect 6561 10761 6595 10795
rect 6595 10761 6604 10795
rect 6552 10752 6604 10761
rect 13084 10752 13136 10804
rect 15752 10752 15804 10804
rect 16672 10752 16724 10804
rect 7012 10727 7064 10736
rect 7012 10693 7021 10727
rect 7021 10693 7055 10727
rect 7055 10693 7064 10727
rect 7012 10684 7064 10693
rect 5632 10659 5684 10668
rect 5632 10625 5641 10659
rect 5641 10625 5675 10659
rect 5675 10625 5684 10659
rect 5632 10616 5684 10625
rect 5724 10659 5776 10668
rect 5724 10625 5733 10659
rect 5733 10625 5767 10659
rect 5767 10625 5776 10659
rect 5724 10616 5776 10625
rect 5908 10616 5960 10668
rect 6092 10616 6144 10668
rect 6460 10616 6512 10668
rect 8208 10684 8260 10736
rect 8300 10727 8352 10736
rect 8300 10693 8309 10727
rect 8309 10693 8343 10727
rect 8343 10693 8352 10727
rect 8300 10684 8352 10693
rect 8760 10684 8812 10736
rect 11520 10616 11572 10668
rect 12072 10616 12124 10668
rect 13268 10684 13320 10736
rect 16396 10684 16448 10736
rect 18604 10752 18656 10804
rect 22468 10752 22520 10804
rect 17868 10684 17920 10736
rect 18236 10684 18288 10736
rect 12808 10616 12860 10668
rect 14648 10616 14700 10668
rect 15476 10616 15528 10668
rect 21456 10684 21508 10736
rect 22284 10684 22336 10736
rect 23940 10752 23992 10804
rect 26792 10752 26844 10804
rect 19248 10616 19300 10668
rect 19524 10616 19576 10668
rect 22192 10616 22244 10668
rect 22560 10659 22612 10668
rect 22560 10625 22567 10659
rect 22567 10625 22612 10659
rect 22560 10616 22612 10625
rect 24216 10684 24268 10736
rect 26240 10684 26292 10736
rect 26424 10684 26476 10736
rect 26976 10684 27028 10736
rect 23112 10659 23164 10668
rect 23112 10625 23121 10659
rect 23121 10625 23155 10659
rect 23155 10625 23164 10659
rect 23112 10616 23164 10625
rect 23480 10616 23532 10668
rect 6368 10480 6420 10532
rect 6552 10480 6604 10532
rect 7196 10480 7248 10532
rect 10324 10591 10376 10600
rect 10324 10557 10333 10591
rect 10333 10557 10367 10591
rect 10367 10557 10376 10591
rect 10324 10548 10376 10557
rect 10692 10548 10744 10600
rect 11888 10591 11940 10600
rect 11888 10557 11897 10591
rect 11897 10557 11931 10591
rect 11931 10557 11940 10591
rect 11888 10548 11940 10557
rect 13544 10548 13596 10600
rect 14096 10548 14148 10600
rect 12256 10480 12308 10532
rect 12900 10480 12952 10532
rect 14280 10480 14332 10532
rect 8760 10412 8812 10464
rect 9956 10455 10008 10464
rect 9956 10421 9965 10455
rect 9965 10421 9999 10455
rect 9999 10421 10008 10455
rect 9956 10412 10008 10421
rect 15660 10455 15712 10464
rect 15660 10421 15669 10455
rect 15669 10421 15703 10455
rect 15703 10421 15712 10455
rect 15660 10412 15712 10421
rect 16488 10412 16540 10464
rect 17040 10591 17092 10600
rect 17040 10557 17049 10591
rect 17049 10557 17083 10591
rect 17083 10557 17092 10591
rect 17040 10548 17092 10557
rect 18512 10591 18564 10600
rect 18512 10557 18521 10591
rect 18521 10557 18555 10591
rect 18555 10557 18564 10591
rect 18512 10548 18564 10557
rect 20076 10591 20128 10600
rect 20076 10557 20085 10591
rect 20085 10557 20119 10591
rect 20119 10557 20128 10591
rect 20076 10548 20128 10557
rect 24584 10616 24636 10668
rect 27252 10548 27304 10600
rect 27528 10616 27580 10668
rect 18328 10412 18380 10464
rect 21548 10455 21600 10464
rect 21548 10421 21557 10455
rect 21557 10421 21591 10455
rect 21591 10421 21600 10455
rect 21548 10412 21600 10421
rect 21916 10412 21968 10464
rect 27436 10412 27488 10464
rect 27896 10455 27948 10464
rect 27896 10421 27905 10455
rect 27905 10421 27939 10455
rect 27939 10421 27948 10455
rect 27896 10412 27948 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 6092 10208 6144 10260
rect 14004 10208 14056 10260
rect 15660 10251 15712 10260
rect 15660 10217 15669 10251
rect 15669 10217 15703 10251
rect 15703 10217 15712 10251
rect 15660 10208 15712 10217
rect 15936 10208 15988 10260
rect 16396 10251 16448 10260
rect 16396 10217 16405 10251
rect 16405 10217 16439 10251
rect 16439 10217 16448 10251
rect 16396 10208 16448 10217
rect 16672 10208 16724 10260
rect 7656 10183 7708 10192
rect 7656 10149 7665 10183
rect 7665 10149 7699 10183
rect 7699 10149 7708 10183
rect 7656 10140 7708 10149
rect 6276 10072 6328 10124
rect 7288 10072 7340 10124
rect 9956 10072 10008 10124
rect 14188 10072 14240 10124
rect 14556 10072 14608 10124
rect 16856 10072 16908 10124
rect 18144 10115 18196 10124
rect 18144 10081 18153 10115
rect 18153 10081 18187 10115
rect 18187 10081 18196 10115
rect 18144 10072 18196 10081
rect 18328 10072 18380 10124
rect 18512 10208 18564 10260
rect 6000 10004 6052 10056
rect 6644 10047 6696 10056
rect 6644 10013 6653 10047
rect 6653 10013 6687 10047
rect 6687 10013 6696 10047
rect 6644 10004 6696 10013
rect 6736 10047 6788 10056
rect 6736 10013 6745 10047
rect 6745 10013 6779 10047
rect 6779 10013 6788 10047
rect 6736 10004 6788 10013
rect 6920 10047 6972 10056
rect 6920 10013 6929 10047
rect 6929 10013 6963 10047
rect 6963 10013 6972 10047
rect 6920 10004 6972 10013
rect 7196 10047 7248 10056
rect 7196 10013 7205 10047
rect 7205 10013 7239 10047
rect 7239 10013 7248 10047
rect 7196 10004 7248 10013
rect 6828 9936 6880 9988
rect 7840 10047 7892 10056
rect 7840 10013 7849 10047
rect 7849 10013 7883 10047
rect 7883 10013 7892 10047
rect 7840 10004 7892 10013
rect 8760 10004 8812 10056
rect 13636 10004 13688 10056
rect 14280 10047 14332 10056
rect 14280 10013 14289 10047
rect 14289 10013 14323 10047
rect 14323 10013 14332 10047
rect 14280 10004 14332 10013
rect 15936 10047 15988 10056
rect 15936 10013 15945 10047
rect 15945 10013 15979 10047
rect 15979 10013 15988 10047
rect 15936 10004 15988 10013
rect 11888 9936 11940 9988
rect 16488 10004 16540 10056
rect 18512 10047 18564 10056
rect 18512 10013 18521 10047
rect 18521 10013 18555 10047
rect 18555 10013 18564 10047
rect 18512 10004 18564 10013
rect 18604 10047 18656 10056
rect 18604 10013 18613 10047
rect 18613 10013 18647 10047
rect 18647 10013 18656 10047
rect 18604 10004 18656 10013
rect 19524 10072 19576 10124
rect 26240 10072 26292 10124
rect 27344 10072 27396 10124
rect 20444 10047 20496 10056
rect 20444 10013 20453 10047
rect 20453 10013 20487 10047
rect 20487 10013 20496 10047
rect 20444 10004 20496 10013
rect 22744 10004 22796 10056
rect 24584 10047 24636 10056
rect 24584 10013 24593 10047
rect 24593 10013 24627 10047
rect 24627 10013 24636 10047
rect 24584 10004 24636 10013
rect 26424 10047 26476 10056
rect 26424 10013 26433 10047
rect 26433 10013 26467 10047
rect 26467 10013 26476 10047
rect 26424 10004 26476 10013
rect 27896 10004 27948 10056
rect 9956 9868 10008 9920
rect 10692 9911 10744 9920
rect 10692 9877 10701 9911
rect 10701 9877 10735 9911
rect 10735 9877 10744 9911
rect 10692 9868 10744 9877
rect 10876 9868 10928 9920
rect 14464 9868 14516 9920
rect 17408 9936 17460 9988
rect 17868 9979 17920 9988
rect 17868 9945 17877 9979
rect 17877 9945 17911 9979
rect 17911 9945 17920 9979
rect 17868 9936 17920 9945
rect 20352 9936 20404 9988
rect 20720 9979 20772 9988
rect 20720 9945 20729 9979
rect 20729 9945 20763 9979
rect 20763 9945 20772 9979
rect 20720 9936 20772 9945
rect 21824 9936 21876 9988
rect 24768 9936 24820 9988
rect 17040 9868 17092 9920
rect 18236 9911 18288 9920
rect 18236 9877 18245 9911
rect 18245 9877 18279 9911
rect 18279 9877 18288 9911
rect 18236 9868 18288 9877
rect 20904 9911 20956 9920
rect 20904 9877 20913 9911
rect 20913 9877 20947 9911
rect 20947 9877 20956 9911
rect 20904 9868 20956 9877
rect 26332 9911 26384 9920
rect 26332 9877 26341 9911
rect 26341 9877 26375 9911
rect 26375 9877 26384 9911
rect 26332 9868 26384 9877
rect 27528 9868 27580 9920
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 6368 9707 6420 9716
rect 6368 9673 6377 9707
rect 6377 9673 6411 9707
rect 6411 9673 6420 9707
rect 6368 9664 6420 9673
rect 7840 9664 7892 9716
rect 6644 9596 6696 9648
rect 6920 9528 6972 9580
rect 7196 9596 7248 9648
rect 7104 9571 7156 9580
rect 7104 9537 7113 9571
rect 7113 9537 7147 9571
rect 7147 9537 7156 9571
rect 7104 9528 7156 9537
rect 10600 9528 10652 9580
rect 10876 9528 10928 9580
rect 11888 9571 11940 9580
rect 11888 9537 11897 9571
rect 11897 9537 11931 9571
rect 11931 9537 11940 9571
rect 11888 9528 11940 9537
rect 14004 9596 14056 9648
rect 7196 9503 7248 9512
rect 7196 9469 7205 9503
rect 7205 9469 7239 9503
rect 7239 9469 7248 9503
rect 7196 9460 7248 9469
rect 7012 9392 7064 9444
rect 13084 9503 13136 9512
rect 13084 9469 13093 9503
rect 13093 9469 13127 9503
rect 13127 9469 13136 9503
rect 13084 9460 13136 9469
rect 14188 9571 14240 9580
rect 14188 9537 14197 9571
rect 14197 9537 14231 9571
rect 14231 9537 14240 9571
rect 14188 9528 14240 9537
rect 14280 9571 14332 9580
rect 14280 9537 14289 9571
rect 14289 9537 14323 9571
rect 14323 9537 14332 9571
rect 14280 9528 14332 9537
rect 18328 9664 18380 9716
rect 18236 9596 18288 9648
rect 18788 9596 18840 9648
rect 16672 9528 16724 9580
rect 17776 9528 17828 9580
rect 13820 9460 13872 9512
rect 14096 9503 14148 9512
rect 14096 9469 14105 9503
rect 14105 9469 14139 9503
rect 14139 9469 14148 9503
rect 14096 9460 14148 9469
rect 7288 9367 7340 9376
rect 7288 9333 7297 9367
rect 7297 9333 7331 9367
rect 7331 9333 7340 9367
rect 7288 9324 7340 9333
rect 9864 9324 9916 9376
rect 10968 9324 11020 9376
rect 12348 9324 12400 9376
rect 13084 9324 13136 9376
rect 15476 9460 15528 9512
rect 16396 9460 16448 9512
rect 18328 9460 18380 9512
rect 20076 9707 20128 9716
rect 20076 9673 20085 9707
rect 20085 9673 20119 9707
rect 20119 9673 20128 9707
rect 20076 9664 20128 9673
rect 19800 9596 19852 9648
rect 20260 9528 20312 9580
rect 20352 9571 20404 9580
rect 20352 9537 20361 9571
rect 20361 9537 20395 9571
rect 20395 9537 20404 9571
rect 20352 9528 20404 9537
rect 22652 9596 22704 9648
rect 22744 9639 22796 9648
rect 22744 9605 22753 9639
rect 22753 9605 22787 9639
rect 22787 9605 22796 9639
rect 22744 9596 22796 9605
rect 27436 9664 27488 9716
rect 20720 9528 20772 9580
rect 21180 9528 21232 9580
rect 23664 9528 23716 9580
rect 24768 9528 24820 9580
rect 26240 9571 26292 9580
rect 26240 9537 26249 9571
rect 26249 9537 26283 9571
rect 26283 9537 26292 9571
rect 26240 9528 26292 9537
rect 26332 9571 26384 9580
rect 26332 9537 26341 9571
rect 26341 9537 26375 9571
rect 26375 9537 26384 9571
rect 26332 9528 26384 9537
rect 26792 9571 26844 9580
rect 26792 9537 26801 9571
rect 26801 9537 26835 9571
rect 26835 9537 26844 9571
rect 27528 9571 27580 9580
rect 26792 9528 26844 9537
rect 20444 9503 20496 9512
rect 20444 9469 20453 9503
rect 20453 9469 20487 9503
rect 20487 9469 20496 9503
rect 20444 9460 20496 9469
rect 17868 9435 17920 9444
rect 17868 9401 17877 9435
rect 17877 9401 17911 9435
rect 17911 9401 17920 9435
rect 17868 9392 17920 9401
rect 18604 9392 18656 9444
rect 14556 9367 14608 9376
rect 14556 9333 14565 9367
rect 14565 9333 14599 9367
rect 14599 9333 14608 9367
rect 14556 9324 14608 9333
rect 16856 9324 16908 9376
rect 19248 9367 19300 9376
rect 19248 9333 19257 9367
rect 19257 9333 19291 9367
rect 19291 9333 19300 9367
rect 19248 9324 19300 9333
rect 26884 9460 26936 9512
rect 27528 9537 27537 9571
rect 27537 9537 27571 9571
rect 27571 9537 27580 9571
rect 27528 9528 27580 9537
rect 28080 9528 28132 9580
rect 28172 9571 28224 9580
rect 28172 9537 28181 9571
rect 28181 9537 28215 9571
rect 28215 9537 28224 9571
rect 28172 9528 28224 9537
rect 25688 9392 25740 9444
rect 21548 9324 21600 9376
rect 25872 9324 25924 9376
rect 26976 9367 27028 9376
rect 26976 9333 26985 9367
rect 26985 9333 27019 9367
rect 27019 9333 27028 9367
rect 26976 9324 27028 9333
rect 27068 9324 27120 9376
rect 27436 9324 27488 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 6644 9120 6696 9172
rect 7288 9120 7340 9172
rect 6460 9052 6512 9104
rect 5632 8959 5684 8968
rect 5632 8925 5641 8959
rect 5641 8925 5675 8959
rect 5675 8925 5684 8959
rect 5632 8916 5684 8925
rect 7012 8984 7064 9036
rect 14648 9163 14700 9172
rect 14648 9129 14657 9163
rect 14657 9129 14691 9163
rect 14691 9129 14700 9163
rect 14648 9120 14700 9129
rect 16672 9163 16724 9172
rect 16672 9129 16681 9163
rect 16681 9129 16715 9163
rect 16715 9129 16724 9163
rect 16672 9120 16724 9129
rect 17592 9120 17644 9172
rect 19248 9120 19300 9172
rect 19800 9120 19852 9172
rect 6460 8959 6512 8968
rect 6460 8925 6469 8959
rect 6469 8925 6503 8959
rect 6503 8925 6512 8959
rect 6460 8916 6512 8925
rect 9404 8916 9456 8968
rect 10048 8984 10100 9036
rect 5264 8780 5316 8832
rect 6368 8780 6420 8832
rect 7012 8848 7064 8900
rect 8300 8848 8352 8900
rect 9864 8959 9916 8968
rect 9864 8925 9873 8959
rect 9873 8925 9907 8959
rect 9907 8925 9916 8959
rect 9864 8916 9916 8925
rect 9956 8959 10008 8968
rect 9956 8925 9965 8959
rect 9965 8925 9999 8959
rect 9999 8925 10008 8959
rect 9956 8916 10008 8925
rect 15568 9052 15620 9104
rect 20904 9120 20956 9172
rect 26700 9120 26752 9172
rect 26884 9163 26936 9172
rect 26884 9129 26893 9163
rect 26893 9129 26927 9163
rect 26927 9129 26936 9163
rect 26884 9120 26936 9129
rect 25320 9052 25372 9104
rect 26240 9052 26292 9104
rect 27068 9052 27120 9104
rect 28172 9052 28224 9104
rect 10232 8984 10284 9036
rect 12348 9027 12400 9036
rect 12348 8993 12357 9027
rect 12357 8993 12391 9027
rect 12391 8993 12400 9027
rect 12348 8984 12400 8993
rect 15936 8984 15988 9036
rect 17224 8984 17276 9036
rect 17776 8984 17828 9036
rect 18880 8984 18932 9036
rect 20720 8984 20772 9036
rect 21180 8984 21232 9036
rect 22652 9027 22704 9036
rect 22652 8993 22661 9027
rect 22661 8993 22695 9027
rect 22695 8993 22704 9027
rect 22652 8984 22704 8993
rect 24032 8984 24084 9036
rect 25872 9027 25924 9036
rect 25872 8993 25881 9027
rect 25881 8993 25915 9027
rect 25915 8993 25924 9027
rect 25872 8984 25924 8993
rect 10968 8916 11020 8968
rect 11888 8916 11940 8968
rect 14832 8959 14884 8968
rect 14832 8925 14841 8959
rect 14841 8925 14875 8959
rect 14875 8925 14884 8959
rect 14832 8916 14884 8925
rect 15016 8959 15068 8968
rect 15016 8925 15025 8959
rect 15025 8925 15059 8959
rect 15059 8925 15068 8959
rect 15016 8916 15068 8925
rect 9680 8848 9732 8900
rect 10600 8891 10652 8900
rect 10600 8857 10609 8891
rect 10609 8857 10643 8891
rect 10643 8857 10652 8891
rect 10600 8848 10652 8857
rect 12808 8848 12860 8900
rect 15568 8916 15620 8968
rect 16856 8959 16908 8968
rect 16856 8925 16865 8959
rect 16865 8925 16899 8959
rect 16899 8925 16908 8959
rect 16856 8916 16908 8925
rect 20076 8916 20128 8968
rect 20352 8916 20404 8968
rect 20536 8916 20588 8968
rect 22284 8916 22336 8968
rect 24308 8916 24360 8968
rect 24676 8916 24728 8968
rect 25044 8959 25096 8968
rect 25044 8925 25053 8959
rect 25053 8925 25087 8959
rect 25087 8925 25096 8959
rect 25044 8916 25096 8925
rect 15292 8848 15344 8900
rect 16488 8848 16540 8900
rect 21088 8848 21140 8900
rect 24492 8848 24544 8900
rect 25228 8848 25280 8900
rect 26056 8959 26108 8968
rect 26056 8925 26065 8959
rect 26065 8925 26099 8959
rect 26099 8925 26108 8959
rect 26056 8916 26108 8925
rect 26332 8916 26384 8968
rect 26792 8984 26844 9036
rect 26884 8984 26936 9036
rect 26976 8916 27028 8968
rect 27068 8959 27120 8968
rect 27068 8925 27077 8959
rect 27077 8925 27111 8959
rect 27111 8925 27120 8959
rect 27068 8916 27120 8925
rect 27436 8916 27488 8968
rect 28080 8848 28132 8900
rect 7196 8780 7248 8832
rect 9312 8780 9364 8832
rect 14096 8780 14148 8832
rect 15108 8780 15160 8832
rect 15200 8823 15252 8832
rect 15200 8789 15209 8823
rect 15209 8789 15243 8823
rect 15243 8789 15252 8823
rect 15200 8780 15252 8789
rect 15476 8780 15528 8832
rect 19892 8780 19944 8832
rect 20812 8823 20864 8832
rect 20812 8789 20821 8823
rect 20821 8789 20855 8823
rect 20855 8789 20864 8823
rect 20812 8780 20864 8789
rect 22744 8780 22796 8832
rect 24584 8823 24636 8832
rect 24584 8789 24593 8823
rect 24593 8789 24627 8823
rect 24627 8789 24636 8823
rect 24584 8780 24636 8789
rect 24676 8823 24728 8832
rect 24676 8789 24685 8823
rect 24685 8789 24719 8823
rect 24719 8789 24728 8823
rect 24676 8780 24728 8789
rect 26608 8780 26660 8832
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 3240 8508 3292 8560
rect 4620 8508 4672 8560
rect 5264 8619 5316 8628
rect 5264 8585 5273 8619
rect 5273 8585 5307 8619
rect 5307 8585 5316 8619
rect 5264 8576 5316 8585
rect 7012 8576 7064 8628
rect 7380 8576 7432 8628
rect 8392 8619 8444 8628
rect 8392 8585 8401 8619
rect 8401 8585 8435 8619
rect 8435 8585 8444 8619
rect 8392 8576 8444 8585
rect 10692 8576 10744 8628
rect 10968 8576 11020 8628
rect 5632 8508 5684 8560
rect 6460 8508 6512 8560
rect 9312 8551 9364 8560
rect 9312 8517 9321 8551
rect 9321 8517 9355 8551
rect 9355 8517 9364 8551
rect 9312 8508 9364 8517
rect 10324 8508 10376 8560
rect 14556 8576 14608 8628
rect 15016 8576 15068 8628
rect 12808 8508 12860 8560
rect 14188 8508 14240 8560
rect 15568 8576 15620 8628
rect 20536 8619 20588 8628
rect 20536 8585 20545 8619
rect 20545 8585 20579 8619
rect 20579 8585 20588 8619
rect 20536 8576 20588 8585
rect 21088 8619 21140 8628
rect 21088 8585 21103 8619
rect 21103 8585 21137 8619
rect 21137 8585 21140 8619
rect 21088 8576 21140 8585
rect 21824 8576 21876 8628
rect 6552 8483 6604 8492
rect 6552 8449 6561 8483
rect 6561 8449 6595 8483
rect 6595 8449 6604 8483
rect 6552 8440 6604 8449
rect 6828 8483 6880 8492
rect 6828 8449 6837 8483
rect 6837 8449 6871 8483
rect 6871 8449 6880 8483
rect 6828 8440 6880 8449
rect 6920 8483 6972 8492
rect 6920 8449 6929 8483
rect 6929 8449 6963 8483
rect 6963 8449 6972 8483
rect 6920 8440 6972 8449
rect 7012 8483 7064 8492
rect 7012 8449 7021 8483
rect 7021 8449 7055 8483
rect 7055 8449 7064 8483
rect 7012 8440 7064 8449
rect 5356 8415 5408 8424
rect 5356 8381 5365 8415
rect 5365 8381 5399 8415
rect 5399 8381 5408 8415
rect 5356 8372 5408 8381
rect 5448 8415 5500 8424
rect 5448 8381 5457 8415
rect 5457 8381 5491 8415
rect 5491 8381 5500 8415
rect 5448 8372 5500 8381
rect 5908 8372 5960 8424
rect 7288 8483 7340 8492
rect 7288 8449 7297 8483
rect 7297 8449 7331 8483
rect 7331 8449 7340 8483
rect 7288 8440 7340 8449
rect 8300 8483 8352 8492
rect 8300 8449 8309 8483
rect 8309 8449 8343 8483
rect 8343 8449 8352 8483
rect 8300 8440 8352 8449
rect 8760 8372 8812 8424
rect 9404 8372 9456 8424
rect 11888 8372 11940 8424
rect 14924 8483 14976 8492
rect 14924 8449 14933 8483
rect 14933 8449 14967 8483
rect 14967 8449 14976 8483
rect 14924 8440 14976 8449
rect 15292 8483 15344 8492
rect 15292 8449 15301 8483
rect 15301 8449 15335 8483
rect 15335 8449 15344 8483
rect 15292 8440 15344 8449
rect 14188 8415 14240 8424
rect 14188 8381 14197 8415
rect 14197 8381 14231 8415
rect 14231 8381 14240 8415
rect 14188 8372 14240 8381
rect 15568 8483 15620 8492
rect 15568 8449 15577 8483
rect 15577 8449 15611 8483
rect 15611 8449 15620 8483
rect 15568 8440 15620 8449
rect 16396 8508 16448 8560
rect 17408 8508 17460 8560
rect 19708 8551 19760 8560
rect 19708 8517 19717 8551
rect 19717 8517 19751 8551
rect 19751 8517 19760 8551
rect 19708 8508 19760 8517
rect 20168 8551 20220 8560
rect 20168 8517 20177 8551
rect 20177 8517 20211 8551
rect 20211 8517 20220 8551
rect 20168 8508 20220 8517
rect 20352 8551 20404 8560
rect 20352 8517 20377 8551
rect 20377 8517 20404 8551
rect 20352 8508 20404 8517
rect 22744 8576 22796 8628
rect 24124 8576 24176 8628
rect 24584 8576 24636 8628
rect 5724 8236 5776 8288
rect 15752 8415 15804 8424
rect 15752 8381 15761 8415
rect 15761 8381 15795 8415
rect 15795 8381 15804 8415
rect 17224 8483 17276 8492
rect 17224 8449 17233 8483
rect 17233 8449 17267 8483
rect 17267 8449 17276 8483
rect 17224 8440 17276 8449
rect 17500 8483 17552 8492
rect 17500 8449 17509 8483
rect 17509 8449 17543 8483
rect 17543 8449 17552 8483
rect 17500 8440 17552 8449
rect 17592 8483 17644 8492
rect 17592 8449 17601 8483
rect 17601 8449 17635 8483
rect 17635 8449 17644 8483
rect 17592 8440 17644 8449
rect 17684 8483 17736 8492
rect 17684 8449 17693 8483
rect 17693 8449 17727 8483
rect 17727 8449 17736 8483
rect 17684 8440 17736 8449
rect 17868 8483 17920 8492
rect 17868 8449 17877 8483
rect 17877 8449 17911 8483
rect 17911 8449 17920 8483
rect 17868 8440 17920 8449
rect 20076 8483 20128 8492
rect 20076 8449 20085 8483
rect 20085 8449 20119 8483
rect 20119 8449 20128 8483
rect 20076 8440 20128 8449
rect 20536 8440 20588 8492
rect 15752 8372 15804 8381
rect 16764 8372 16816 8424
rect 19432 8372 19484 8424
rect 20168 8372 20220 8424
rect 20260 8372 20312 8424
rect 22284 8440 22336 8492
rect 23940 8440 23992 8492
rect 19800 8304 19852 8356
rect 21088 8372 21140 8424
rect 23664 8415 23716 8424
rect 23664 8381 23673 8415
rect 23673 8381 23707 8415
rect 23707 8381 23716 8415
rect 23664 8372 23716 8381
rect 24216 8372 24268 8424
rect 24676 8508 24728 8560
rect 25044 8508 25096 8560
rect 25228 8483 25280 8492
rect 25228 8449 25237 8483
rect 25237 8449 25271 8483
rect 25271 8449 25280 8483
rect 25228 8440 25280 8449
rect 25320 8483 25372 8492
rect 25320 8449 25329 8483
rect 25329 8449 25363 8483
rect 25363 8449 25372 8483
rect 25320 8440 25372 8449
rect 25688 8483 25740 8492
rect 25688 8449 25697 8483
rect 25697 8449 25731 8483
rect 25731 8449 25740 8483
rect 25688 8440 25740 8449
rect 24768 8372 24820 8424
rect 25044 8415 25096 8424
rect 25044 8381 25053 8415
rect 25053 8381 25087 8415
rect 25087 8381 25096 8415
rect 25044 8372 25096 8381
rect 25412 8372 25464 8424
rect 26056 8483 26108 8492
rect 26056 8449 26065 8483
rect 26065 8449 26099 8483
rect 26099 8449 26108 8483
rect 26056 8440 26108 8449
rect 26332 8372 26384 8424
rect 24676 8304 24728 8356
rect 24952 8304 25004 8356
rect 7288 8279 7340 8288
rect 7288 8245 7297 8279
rect 7297 8245 7331 8279
rect 7331 8245 7340 8279
rect 7288 8236 7340 8245
rect 9496 8236 9548 8288
rect 9864 8236 9916 8288
rect 14924 8236 14976 8288
rect 16120 8279 16172 8288
rect 16120 8245 16129 8279
rect 16129 8245 16163 8279
rect 16163 8245 16172 8279
rect 16120 8236 16172 8245
rect 16672 8279 16724 8288
rect 16672 8245 16681 8279
rect 16681 8245 16715 8279
rect 16715 8245 16724 8279
rect 16672 8236 16724 8245
rect 17316 8279 17368 8288
rect 17316 8245 17325 8279
rect 17325 8245 17359 8279
rect 17359 8245 17368 8279
rect 17316 8236 17368 8245
rect 19524 8279 19576 8288
rect 19524 8245 19533 8279
rect 19533 8245 19567 8279
rect 19567 8245 19576 8279
rect 19524 8236 19576 8245
rect 19892 8236 19944 8288
rect 20260 8236 20312 8288
rect 24308 8279 24360 8288
rect 24308 8245 24317 8279
rect 24317 8245 24351 8279
rect 24351 8245 24360 8279
rect 24308 8236 24360 8245
rect 24400 8236 24452 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 5356 8032 5408 8084
rect 7104 8032 7156 8084
rect 5724 7964 5776 8016
rect 6460 7939 6512 7948
rect 6460 7905 6469 7939
rect 6469 7905 6503 7939
rect 6503 7905 6512 7939
rect 6460 7896 6512 7905
rect 5908 7871 5960 7880
rect 5908 7837 5917 7871
rect 5917 7837 5951 7871
rect 5951 7837 5960 7871
rect 5908 7828 5960 7837
rect 6368 7871 6420 7880
rect 6368 7837 6377 7871
rect 6377 7837 6411 7871
rect 6411 7837 6420 7871
rect 6368 7828 6420 7837
rect 8392 7964 8444 8016
rect 7196 7896 7248 7948
rect 9956 8032 10008 8084
rect 10600 8032 10652 8084
rect 14832 8032 14884 8084
rect 15936 8075 15988 8084
rect 15936 8041 15945 8075
rect 15945 8041 15979 8075
rect 15979 8041 15988 8075
rect 15936 8032 15988 8041
rect 16672 8032 16724 8084
rect 19708 8032 19760 8084
rect 24308 8032 24360 8084
rect 25412 8032 25464 8084
rect 10140 7964 10192 8016
rect 7104 7871 7156 7880
rect 7104 7837 7113 7871
rect 7113 7837 7147 7871
rect 7147 7837 7156 7871
rect 7104 7828 7156 7837
rect 7288 7828 7340 7880
rect 9312 7871 9364 7880
rect 9312 7837 9321 7871
rect 9321 7837 9355 7871
rect 9355 7837 9364 7871
rect 9312 7828 9364 7837
rect 9588 7871 9640 7880
rect 9588 7837 9597 7871
rect 9597 7837 9631 7871
rect 9631 7837 9640 7871
rect 9588 7828 9640 7837
rect 9864 7871 9916 7880
rect 9864 7837 9873 7871
rect 9873 7837 9907 7871
rect 9907 7837 9916 7871
rect 9864 7828 9916 7837
rect 10416 7896 10468 7948
rect 15476 7896 15528 7948
rect 15660 7896 15712 7948
rect 17500 7964 17552 8016
rect 24124 8007 24176 8016
rect 24124 7973 24133 8007
rect 24133 7973 24167 8007
rect 24167 7973 24176 8007
rect 24124 7964 24176 7973
rect 24676 7964 24728 8016
rect 26332 8075 26384 8084
rect 26332 8041 26341 8075
rect 26341 8041 26375 8075
rect 26375 8041 26384 8075
rect 26332 8032 26384 8041
rect 26516 8032 26568 8084
rect 26884 8032 26936 8084
rect 26792 7964 26844 8016
rect 17224 7896 17276 7948
rect 5540 7760 5592 7812
rect 7196 7760 7248 7812
rect 7380 7803 7432 7812
rect 7380 7769 7389 7803
rect 7389 7769 7423 7803
rect 7423 7769 7432 7803
rect 7380 7760 7432 7769
rect 10968 7828 11020 7880
rect 5448 7692 5500 7744
rect 6644 7735 6696 7744
rect 6644 7701 6653 7735
rect 6653 7701 6687 7735
rect 6687 7701 6696 7735
rect 6644 7692 6696 7701
rect 9588 7692 9640 7744
rect 9680 7735 9732 7744
rect 9680 7701 9689 7735
rect 9689 7701 9723 7735
rect 9723 7701 9732 7735
rect 9680 7692 9732 7701
rect 9772 7692 9824 7744
rect 10508 7692 10560 7744
rect 10876 7803 10928 7812
rect 10876 7769 10885 7803
rect 10885 7769 10919 7803
rect 10919 7769 10928 7803
rect 10876 7760 10928 7769
rect 12808 7828 12860 7880
rect 14924 7871 14976 7880
rect 14924 7837 14933 7871
rect 14933 7837 14967 7871
rect 14967 7837 14976 7871
rect 14924 7828 14976 7837
rect 15108 7828 15160 7880
rect 16120 7871 16172 7880
rect 16120 7837 16129 7871
rect 16129 7837 16163 7871
rect 16163 7837 16172 7871
rect 16120 7828 16172 7837
rect 16764 7871 16816 7880
rect 16764 7837 16773 7871
rect 16773 7837 16807 7871
rect 16807 7837 16816 7871
rect 16764 7828 16816 7837
rect 16948 7871 17000 7880
rect 16948 7837 16957 7871
rect 16957 7837 16991 7871
rect 16991 7837 17000 7871
rect 16948 7828 17000 7837
rect 15200 7760 15252 7812
rect 11612 7692 11664 7744
rect 17316 7871 17368 7880
rect 17316 7837 17325 7871
rect 17325 7837 17359 7871
rect 17359 7837 17368 7871
rect 17316 7828 17368 7837
rect 18420 7896 18472 7948
rect 18328 7828 18380 7880
rect 18788 7828 18840 7880
rect 18880 7871 18932 7880
rect 18880 7837 18889 7871
rect 18889 7837 18923 7871
rect 18923 7837 18932 7871
rect 18880 7828 18932 7837
rect 19064 7828 19116 7880
rect 20260 7896 20312 7948
rect 24584 7939 24636 7948
rect 24584 7905 24593 7939
rect 24593 7905 24627 7939
rect 24627 7905 24636 7939
rect 24584 7896 24636 7905
rect 24860 7939 24912 7948
rect 24860 7905 24870 7939
rect 24870 7905 24904 7939
rect 24904 7905 24912 7939
rect 24860 7896 24912 7905
rect 25228 7939 25280 7948
rect 25228 7905 25237 7939
rect 25237 7905 25271 7939
rect 25271 7905 25280 7939
rect 25228 7896 25280 7905
rect 26332 7896 26384 7948
rect 26608 7896 26660 7948
rect 19432 7871 19484 7880
rect 19432 7837 19441 7871
rect 19441 7837 19475 7871
rect 19475 7837 19484 7871
rect 19432 7828 19484 7837
rect 17776 7760 17828 7812
rect 17408 7692 17460 7744
rect 18328 7735 18380 7744
rect 18328 7701 18337 7735
rect 18337 7701 18371 7735
rect 18371 7701 18380 7735
rect 18328 7692 18380 7701
rect 18972 7760 19024 7812
rect 19156 7760 19208 7812
rect 20352 7828 20404 7880
rect 22100 7828 22152 7880
rect 24308 7828 24360 7880
rect 24492 7828 24544 7880
rect 25136 7828 25188 7880
rect 26516 7871 26568 7880
rect 26516 7837 26525 7871
rect 26525 7837 26559 7871
rect 26559 7837 26568 7871
rect 26516 7828 26568 7837
rect 28356 7871 28408 7880
rect 28356 7837 28365 7871
rect 28365 7837 28399 7871
rect 28399 7837 28408 7871
rect 28356 7828 28408 7837
rect 23940 7760 23992 7812
rect 19248 7692 19300 7744
rect 23848 7692 23900 7744
rect 25688 7760 25740 7812
rect 27528 7692 27580 7744
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 5448 7531 5500 7540
rect 5448 7497 5457 7531
rect 5457 7497 5491 7531
rect 5491 7497 5500 7531
rect 5448 7488 5500 7497
rect 6460 7488 6512 7540
rect 9312 7488 9364 7540
rect 11796 7488 11848 7540
rect 5908 7420 5960 7472
rect 4620 7352 4672 7404
rect 5264 7352 5316 7404
rect 6920 7420 6972 7472
rect 6644 7395 6696 7404
rect 6644 7361 6653 7395
rect 6653 7361 6687 7395
rect 6687 7361 6696 7395
rect 6644 7352 6696 7361
rect 10416 7420 10468 7472
rect 11612 7420 11664 7472
rect 12072 7420 12124 7472
rect 17868 7488 17920 7540
rect 18328 7488 18380 7540
rect 15016 7420 15068 7472
rect 17132 7420 17184 7472
rect 7380 7352 7432 7404
rect 10968 7395 11020 7404
rect 3240 7327 3292 7336
rect 3240 7293 3249 7327
rect 3249 7293 3283 7327
rect 3283 7293 3292 7327
rect 3240 7284 3292 7293
rect 5356 7284 5408 7336
rect 6460 7284 6512 7336
rect 7196 7284 7248 7336
rect 8300 7284 8352 7336
rect 8760 7327 8812 7336
rect 8760 7293 8769 7327
rect 8769 7293 8803 7327
rect 8803 7293 8812 7327
rect 8760 7284 8812 7293
rect 9036 7327 9088 7336
rect 9036 7293 9045 7327
rect 9045 7293 9079 7327
rect 9079 7293 9088 7327
rect 9036 7284 9088 7293
rect 10968 7361 10977 7395
rect 10977 7361 11011 7395
rect 11011 7361 11020 7395
rect 10968 7352 11020 7361
rect 11152 7284 11204 7336
rect 12440 7395 12492 7404
rect 12440 7361 12449 7395
rect 12449 7361 12483 7395
rect 12483 7361 12492 7395
rect 12440 7352 12492 7361
rect 13636 7352 13688 7404
rect 18420 7463 18472 7472
rect 18420 7429 18429 7463
rect 18429 7429 18463 7463
rect 18463 7429 18472 7463
rect 18420 7420 18472 7429
rect 17960 7395 18012 7404
rect 17960 7361 17969 7395
rect 17969 7361 18003 7395
rect 18003 7361 18012 7395
rect 17960 7352 18012 7361
rect 18052 7395 18104 7404
rect 18052 7361 18061 7395
rect 18061 7361 18095 7395
rect 18095 7361 18104 7395
rect 18052 7352 18104 7361
rect 12348 7284 12400 7336
rect 12716 7284 12768 7336
rect 12992 7327 13044 7336
rect 12992 7293 13001 7327
rect 13001 7293 13035 7327
rect 13035 7293 13044 7327
rect 12992 7284 13044 7293
rect 18512 7395 18564 7404
rect 18512 7361 18521 7395
rect 18521 7361 18555 7395
rect 18555 7361 18564 7395
rect 18512 7352 18564 7361
rect 18696 7395 18748 7404
rect 18696 7361 18704 7395
rect 18704 7361 18738 7395
rect 18738 7361 18748 7395
rect 18696 7352 18748 7361
rect 19432 7488 19484 7540
rect 22100 7488 22152 7540
rect 24308 7488 24360 7540
rect 25228 7488 25280 7540
rect 19156 7463 19208 7472
rect 19156 7429 19165 7463
rect 19165 7429 19199 7463
rect 19199 7429 19208 7463
rect 19156 7420 19208 7429
rect 19248 7463 19300 7472
rect 19248 7429 19257 7463
rect 19257 7429 19291 7463
rect 19291 7429 19300 7463
rect 19248 7420 19300 7429
rect 19524 7420 19576 7472
rect 21456 7420 21508 7472
rect 24676 7420 24728 7472
rect 18604 7284 18656 7336
rect 17776 7216 17828 7268
rect 17960 7216 18012 7268
rect 9496 7148 9548 7200
rect 9588 7148 9640 7200
rect 10692 7148 10744 7200
rect 12532 7148 12584 7200
rect 24400 7395 24452 7404
rect 24400 7361 24409 7395
rect 24409 7361 24443 7395
rect 24443 7361 24452 7395
rect 24400 7352 24452 7361
rect 26056 7488 26108 7540
rect 25688 7463 25740 7472
rect 25688 7429 25697 7463
rect 25697 7429 25731 7463
rect 25731 7429 25740 7463
rect 25688 7420 25740 7429
rect 26332 7395 26384 7404
rect 26332 7361 26341 7395
rect 26341 7361 26375 7395
rect 26375 7361 26384 7395
rect 26332 7352 26384 7361
rect 26424 7395 26476 7404
rect 26424 7361 26433 7395
rect 26433 7361 26467 7395
rect 26467 7361 26476 7395
rect 26424 7352 26476 7361
rect 26240 7284 26292 7336
rect 28356 7395 28408 7404
rect 28356 7361 28365 7395
rect 28365 7361 28399 7395
rect 28399 7361 28408 7395
rect 28356 7352 28408 7361
rect 26332 7216 26384 7268
rect 21180 7148 21232 7200
rect 24400 7191 24452 7200
rect 24400 7157 24409 7191
rect 24409 7157 24443 7191
rect 24443 7157 24452 7191
rect 24400 7148 24452 7157
rect 25504 7148 25556 7200
rect 27896 7148 27948 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 9036 6944 9088 6996
rect 10508 6987 10560 6996
rect 10508 6953 10517 6987
rect 10517 6953 10551 6987
rect 10551 6953 10560 6987
rect 10508 6944 10560 6953
rect 11980 6944 12032 6996
rect 12164 6987 12216 6996
rect 12164 6953 12194 6987
rect 12194 6953 12216 6987
rect 12164 6944 12216 6953
rect 12348 6944 12400 6996
rect 18052 6944 18104 6996
rect 11520 6876 11572 6928
rect 18328 6876 18380 6928
rect 19064 6944 19116 6996
rect 27528 6944 27580 6996
rect 10968 6851 11020 6860
rect 10968 6817 10977 6851
rect 10977 6817 11011 6851
rect 11011 6817 11020 6851
rect 10968 6808 11020 6817
rect 10048 6740 10100 6792
rect 10232 6783 10284 6792
rect 10232 6749 10241 6783
rect 10241 6749 10275 6783
rect 10275 6749 10284 6783
rect 10232 6740 10284 6749
rect 10692 6783 10744 6792
rect 10692 6749 10701 6783
rect 10701 6749 10735 6783
rect 10735 6749 10744 6783
rect 10692 6740 10744 6749
rect 11152 6783 11204 6792
rect 11152 6749 11161 6783
rect 11161 6749 11195 6783
rect 11195 6749 11204 6783
rect 11152 6740 11204 6749
rect 12532 6808 12584 6860
rect 17684 6808 17736 6860
rect 11520 6783 11572 6792
rect 11520 6749 11529 6783
rect 11529 6749 11563 6783
rect 11563 6749 11572 6783
rect 11520 6740 11572 6749
rect 11888 6783 11940 6792
rect 11888 6749 11897 6783
rect 11897 6749 11931 6783
rect 11931 6749 11940 6783
rect 11888 6740 11940 6749
rect 18788 6808 18840 6860
rect 18604 6783 18656 6792
rect 10784 6672 10836 6724
rect 11244 6604 11296 6656
rect 12440 6604 12492 6656
rect 12624 6672 12676 6724
rect 17224 6672 17276 6724
rect 18604 6749 18613 6783
rect 18613 6749 18647 6783
rect 18647 6749 18656 6783
rect 18604 6740 18656 6749
rect 18236 6715 18288 6724
rect 18236 6681 18245 6715
rect 18245 6681 18279 6715
rect 18279 6681 18288 6715
rect 18236 6672 18288 6681
rect 18880 6740 18932 6792
rect 28264 6783 28316 6792
rect 28264 6749 28273 6783
rect 28273 6749 28307 6783
rect 28307 6749 28316 6783
rect 28264 6740 28316 6749
rect 19156 6672 19208 6724
rect 23572 6672 23624 6724
rect 24216 6672 24268 6724
rect 26700 6672 26752 6724
rect 27252 6672 27304 6724
rect 13636 6647 13688 6656
rect 13636 6613 13645 6647
rect 13645 6613 13679 6647
rect 13679 6613 13688 6647
rect 13636 6604 13688 6613
rect 19800 6604 19852 6656
rect 24124 6604 24176 6656
rect 26608 6604 26660 6656
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 12164 6400 12216 6452
rect 12716 6443 12768 6452
rect 12716 6409 12725 6443
rect 12725 6409 12759 6443
rect 12759 6409 12768 6443
rect 12716 6400 12768 6409
rect 12808 6400 12860 6452
rect 22284 6400 22336 6452
rect 23572 6443 23624 6452
rect 23572 6409 23581 6443
rect 23581 6409 23615 6443
rect 23615 6409 23624 6443
rect 23572 6400 23624 6409
rect 24860 6443 24912 6452
rect 24860 6409 24869 6443
rect 24869 6409 24903 6443
rect 24903 6409 24912 6443
rect 24860 6400 24912 6409
rect 27160 6443 27212 6452
rect 27160 6409 27169 6443
rect 27169 6409 27203 6443
rect 27203 6409 27212 6443
rect 27160 6400 27212 6409
rect 13452 6375 13504 6384
rect 13452 6341 13461 6375
rect 13461 6341 13495 6375
rect 13495 6341 13504 6375
rect 13452 6332 13504 6341
rect 14924 6332 14976 6384
rect 16580 6332 16632 6384
rect 20444 6332 20496 6384
rect 22560 6332 22612 6384
rect 11520 6264 11572 6316
rect 11980 6307 12032 6316
rect 11980 6273 11989 6307
rect 11989 6273 12023 6307
rect 12023 6273 12032 6307
rect 11980 6264 12032 6273
rect 12716 6264 12768 6316
rect 13636 6264 13688 6316
rect 13912 6264 13964 6316
rect 14740 6264 14792 6316
rect 15936 6264 15988 6316
rect 12532 6196 12584 6248
rect 11796 6128 11848 6180
rect 15384 6196 15436 6248
rect 15200 6128 15252 6180
rect 16212 6307 16264 6316
rect 16212 6273 16221 6307
rect 16221 6273 16255 6307
rect 16255 6273 16264 6307
rect 16212 6264 16264 6273
rect 16396 6307 16448 6316
rect 16396 6273 16405 6307
rect 16405 6273 16439 6307
rect 16439 6273 16448 6307
rect 16396 6264 16448 6273
rect 16856 6196 16908 6248
rect 18512 6264 18564 6316
rect 23848 6307 23900 6316
rect 23848 6273 23857 6307
rect 23857 6273 23891 6307
rect 23891 6273 23900 6307
rect 23848 6264 23900 6273
rect 24032 6307 24084 6316
rect 24032 6273 24041 6307
rect 24041 6273 24075 6307
rect 24075 6273 24084 6307
rect 24032 6264 24084 6273
rect 24124 6307 24176 6316
rect 24124 6273 24133 6307
rect 24133 6273 24167 6307
rect 24167 6273 24176 6307
rect 24124 6264 24176 6273
rect 24584 6307 24636 6316
rect 24584 6273 24593 6307
rect 24593 6273 24627 6307
rect 24627 6273 24636 6307
rect 24584 6264 24636 6273
rect 25044 6264 25096 6316
rect 18696 6196 18748 6248
rect 19064 6196 19116 6248
rect 21180 6196 21232 6248
rect 16028 6128 16080 6180
rect 16672 6171 16724 6180
rect 16672 6137 16681 6171
rect 16681 6137 16715 6171
rect 16715 6137 16724 6171
rect 16672 6128 16724 6137
rect 17316 6128 17368 6180
rect 23480 6128 23532 6180
rect 24768 6128 24820 6180
rect 26240 6307 26292 6316
rect 26240 6273 26249 6307
rect 26249 6273 26283 6307
rect 26283 6273 26292 6307
rect 26240 6264 26292 6273
rect 26792 6264 26844 6316
rect 26240 6128 26292 6180
rect 27620 6307 27672 6316
rect 27620 6273 27629 6307
rect 27629 6273 27663 6307
rect 27663 6273 27672 6307
rect 27620 6264 27672 6273
rect 28356 6307 28408 6316
rect 28356 6273 28365 6307
rect 28365 6273 28399 6307
rect 28399 6273 28408 6307
rect 28356 6264 28408 6273
rect 27988 6196 28040 6248
rect 27896 6128 27948 6180
rect 13084 6060 13136 6112
rect 13728 6060 13780 6112
rect 15476 6060 15528 6112
rect 15752 6103 15804 6112
rect 15752 6069 15761 6103
rect 15761 6069 15795 6103
rect 15795 6069 15804 6103
rect 15752 6060 15804 6069
rect 23756 6060 23808 6112
rect 26148 6103 26200 6112
rect 26148 6069 26157 6103
rect 26157 6069 26191 6103
rect 26191 6069 26200 6103
rect 26148 6060 26200 6069
rect 27528 6103 27580 6112
rect 27528 6069 27537 6103
rect 27537 6069 27571 6103
rect 27571 6069 27580 6103
rect 27528 6060 27580 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 16948 5856 17000 5908
rect 17224 5856 17276 5908
rect 24584 5856 24636 5908
rect 6920 5788 6972 5840
rect 14740 5831 14792 5840
rect 14740 5797 14749 5831
rect 14749 5797 14783 5831
rect 14783 5797 14792 5831
rect 14740 5788 14792 5797
rect 15476 5831 15528 5840
rect 15476 5797 15485 5831
rect 15485 5797 15519 5831
rect 15519 5797 15528 5831
rect 15476 5788 15528 5797
rect 24216 5788 24268 5840
rect 25044 5856 25096 5908
rect 26148 5856 26200 5908
rect 26516 5856 26568 5908
rect 26700 5856 26752 5908
rect 6460 5695 6512 5704
rect 6460 5661 6469 5695
rect 6469 5661 6503 5695
rect 6503 5661 6512 5695
rect 6460 5652 6512 5661
rect 16672 5763 16724 5772
rect 14924 5695 14976 5704
rect 14924 5661 14933 5695
rect 14933 5661 14967 5695
rect 14967 5661 14976 5695
rect 14924 5652 14976 5661
rect 15936 5652 15988 5704
rect 11152 5584 11204 5636
rect 16672 5729 16681 5763
rect 16681 5729 16715 5763
rect 16715 5729 16724 5763
rect 16672 5720 16724 5729
rect 17500 5763 17552 5772
rect 17500 5729 17509 5763
rect 17509 5729 17543 5763
rect 17543 5729 17552 5763
rect 17500 5720 17552 5729
rect 16212 5652 16264 5704
rect 16948 5652 17000 5704
rect 6644 5559 6696 5568
rect 6644 5525 6653 5559
rect 6653 5525 6687 5559
rect 6687 5525 6696 5559
rect 6644 5516 6696 5525
rect 7472 5516 7524 5568
rect 10232 5516 10284 5568
rect 13084 5516 13136 5568
rect 15292 5516 15344 5568
rect 16304 5584 16356 5636
rect 17316 5695 17368 5704
rect 17316 5661 17325 5695
rect 17325 5661 17359 5695
rect 17359 5661 17368 5695
rect 17316 5652 17368 5661
rect 17684 5695 17736 5704
rect 17684 5661 17693 5695
rect 17693 5661 17727 5695
rect 17727 5661 17736 5695
rect 17684 5652 17736 5661
rect 21180 5695 21232 5704
rect 21180 5661 21189 5695
rect 21189 5661 21223 5695
rect 21223 5661 21232 5695
rect 21180 5652 21232 5661
rect 22560 5652 22612 5704
rect 23480 5695 23532 5704
rect 23480 5661 23489 5695
rect 23489 5661 23523 5695
rect 23523 5661 23532 5695
rect 23480 5652 23532 5661
rect 23756 5695 23808 5704
rect 23756 5661 23765 5695
rect 23765 5661 23799 5695
rect 23799 5661 23808 5695
rect 23756 5652 23808 5661
rect 24860 5788 24912 5840
rect 24400 5720 24452 5772
rect 24676 5695 24728 5704
rect 24676 5661 24685 5695
rect 24685 5661 24719 5695
rect 24719 5661 24728 5695
rect 24676 5652 24728 5661
rect 24860 5695 24912 5704
rect 24860 5661 24869 5695
rect 24869 5661 24903 5695
rect 24903 5661 24912 5695
rect 24860 5652 24912 5661
rect 25044 5695 25096 5704
rect 25044 5661 25053 5695
rect 25053 5661 25087 5695
rect 25087 5661 25096 5695
rect 25044 5652 25096 5661
rect 27988 5763 28040 5772
rect 27988 5729 27997 5763
rect 27997 5729 28031 5763
rect 28031 5729 28040 5763
rect 27988 5720 28040 5729
rect 25412 5652 25464 5704
rect 17776 5516 17828 5568
rect 24400 5559 24452 5568
rect 24400 5525 24409 5559
rect 24409 5525 24443 5559
rect 24443 5525 24452 5559
rect 24400 5516 24452 5525
rect 25504 5627 25556 5636
rect 25504 5593 25513 5627
rect 25513 5593 25547 5627
rect 25547 5593 25556 5627
rect 25504 5584 25556 5593
rect 26240 5627 26292 5636
rect 26240 5593 26249 5627
rect 26249 5593 26283 5627
rect 26283 5593 26292 5627
rect 26240 5584 26292 5593
rect 28264 5695 28316 5704
rect 28264 5661 28273 5695
rect 28273 5661 28307 5695
rect 28307 5661 28316 5695
rect 28264 5652 28316 5661
rect 27252 5584 27304 5636
rect 26516 5559 26568 5568
rect 26516 5525 26525 5559
rect 26525 5525 26559 5559
rect 26559 5525 26568 5559
rect 26516 5516 26568 5525
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 6644 5312 6696 5364
rect 6736 5312 6788 5364
rect 5264 5244 5316 5296
rect 5724 5176 5776 5228
rect 6552 5244 6604 5296
rect 6184 5176 6236 5228
rect 7472 5244 7524 5296
rect 6920 5219 6972 5228
rect 6920 5185 6937 5219
rect 6937 5185 6972 5219
rect 6920 5176 6972 5185
rect 3332 5151 3384 5160
rect 3332 5117 3341 5151
rect 3341 5117 3375 5151
rect 3375 5117 3384 5151
rect 3332 5108 3384 5117
rect 3608 5151 3660 5160
rect 3608 5117 3617 5151
rect 3617 5117 3651 5151
rect 3651 5117 3660 5151
rect 3608 5108 3660 5117
rect 4988 5040 5040 5092
rect 5908 5151 5960 5160
rect 5908 5117 5917 5151
rect 5917 5117 5951 5151
rect 5951 5117 5960 5151
rect 5908 5108 5960 5117
rect 6276 5108 6328 5160
rect 6460 5108 6512 5160
rect 7104 5219 7156 5228
rect 7104 5185 7113 5219
rect 7113 5185 7147 5219
rect 7147 5185 7156 5219
rect 7104 5176 7156 5185
rect 7564 5176 7616 5228
rect 7472 5108 7524 5160
rect 6552 5040 6604 5092
rect 8024 5219 8076 5228
rect 8024 5185 8033 5219
rect 8033 5185 8067 5219
rect 8067 5185 8076 5219
rect 8024 5176 8076 5185
rect 9220 5244 9272 5296
rect 12348 5312 12400 5364
rect 15200 5312 15252 5364
rect 15568 5312 15620 5364
rect 15936 5312 15988 5364
rect 9588 5287 9640 5296
rect 9588 5253 9623 5287
rect 9623 5253 9640 5287
rect 9588 5244 9640 5253
rect 11796 5244 11848 5296
rect 12440 5244 12492 5296
rect 13176 5244 13228 5296
rect 16488 5244 16540 5296
rect 16856 5287 16908 5296
rect 16856 5253 16865 5287
rect 16865 5253 16899 5287
rect 16899 5253 16908 5287
rect 16856 5244 16908 5253
rect 17224 5355 17276 5364
rect 17224 5321 17233 5355
rect 17233 5321 17267 5355
rect 17267 5321 17276 5355
rect 17224 5312 17276 5321
rect 18512 5312 18564 5364
rect 19064 5355 19116 5364
rect 19064 5321 19073 5355
rect 19073 5321 19107 5355
rect 19107 5321 19116 5355
rect 19064 5312 19116 5321
rect 19432 5312 19484 5364
rect 20444 5312 20496 5364
rect 17960 5244 18012 5296
rect 8484 5176 8536 5228
rect 7932 5151 7984 5160
rect 7932 5117 7941 5151
rect 7941 5117 7975 5151
rect 7975 5117 7984 5151
rect 7932 5108 7984 5117
rect 8852 5219 8904 5228
rect 8852 5185 8861 5219
rect 8861 5185 8895 5219
rect 8895 5185 8904 5219
rect 8852 5176 8904 5185
rect 9312 5219 9364 5228
rect 9312 5185 9321 5219
rect 9321 5185 9355 5219
rect 9355 5185 9364 5219
rect 9312 5176 9364 5185
rect 9404 5219 9456 5228
rect 9404 5185 9413 5219
rect 9413 5185 9447 5219
rect 9447 5185 9456 5219
rect 9404 5176 9456 5185
rect 7748 5040 7800 5092
rect 9588 5108 9640 5160
rect 12716 5176 12768 5228
rect 12992 5176 13044 5228
rect 15292 5219 15344 5228
rect 15292 5185 15301 5219
rect 15301 5185 15335 5219
rect 15335 5185 15344 5219
rect 15292 5176 15344 5185
rect 15568 5219 15620 5228
rect 15568 5185 15577 5219
rect 15577 5185 15611 5219
rect 15611 5185 15620 5219
rect 15568 5176 15620 5185
rect 15844 5176 15896 5228
rect 12256 5108 12308 5160
rect 9220 5040 9272 5092
rect 10140 5040 10192 5092
rect 10692 5040 10744 5092
rect 15384 5040 15436 5092
rect 5540 4972 5592 5024
rect 6460 4972 6512 5024
rect 7656 4972 7708 5024
rect 9128 5015 9180 5024
rect 9128 4981 9137 5015
rect 9137 4981 9171 5015
rect 9171 4981 9180 5015
rect 9128 4972 9180 4981
rect 12992 5015 13044 5024
rect 12992 4981 13001 5015
rect 13001 4981 13035 5015
rect 13035 4981 13044 5015
rect 12992 4972 13044 4981
rect 16580 5176 16632 5228
rect 16948 5219 17000 5228
rect 16948 5185 16957 5219
rect 16957 5185 16991 5219
rect 16991 5185 17000 5219
rect 16948 5176 17000 5185
rect 17316 5176 17368 5228
rect 18052 5219 18104 5228
rect 18052 5185 18061 5219
rect 18061 5185 18095 5219
rect 18095 5185 18104 5219
rect 18052 5176 18104 5185
rect 19524 5244 19576 5296
rect 19800 5287 19852 5296
rect 19800 5253 19809 5287
rect 19809 5253 19843 5287
rect 19843 5253 19852 5287
rect 19800 5244 19852 5253
rect 18788 5219 18840 5228
rect 17592 5108 17644 5160
rect 17684 5040 17736 5092
rect 18788 5185 18797 5219
rect 18797 5185 18831 5219
rect 18831 5185 18840 5219
rect 18788 5176 18840 5185
rect 18880 5219 18932 5228
rect 18880 5185 18889 5219
rect 18889 5185 18923 5219
rect 18923 5185 18932 5219
rect 18880 5176 18932 5185
rect 19432 5151 19484 5160
rect 19432 5117 19441 5151
rect 19441 5117 19475 5151
rect 19475 5117 19484 5151
rect 19432 5108 19484 5117
rect 22284 5312 22336 5364
rect 23756 5312 23808 5364
rect 24860 5312 24912 5364
rect 22560 5244 22612 5296
rect 24400 5244 24452 5296
rect 24676 5244 24728 5296
rect 25964 5312 26016 5364
rect 27620 5312 27672 5364
rect 27988 5312 28040 5364
rect 26240 5244 26292 5296
rect 23848 5176 23900 5228
rect 24952 5176 25004 5228
rect 25044 5219 25096 5228
rect 25044 5185 25053 5219
rect 25053 5185 25087 5219
rect 25087 5185 25096 5219
rect 25044 5176 25096 5185
rect 25504 5176 25556 5228
rect 26516 5219 26568 5228
rect 26516 5185 26525 5219
rect 26525 5185 26559 5219
rect 26559 5185 26568 5219
rect 26516 5176 26568 5185
rect 28356 5219 28408 5228
rect 28356 5185 28365 5219
rect 28365 5185 28399 5219
rect 28399 5185 28408 5219
rect 28356 5176 28408 5185
rect 19616 5040 19668 5092
rect 16672 4972 16724 5024
rect 18880 4972 18932 5024
rect 18972 4972 19024 5024
rect 20168 5040 20220 5092
rect 22192 5040 22244 5092
rect 23572 5151 23624 5160
rect 23572 5117 23581 5151
rect 23581 5117 23615 5151
rect 23615 5117 23624 5151
rect 23572 5108 23624 5117
rect 24860 5151 24912 5160
rect 24860 5117 24869 5151
rect 24869 5117 24903 5151
rect 24903 5117 24912 5151
rect 24860 5108 24912 5117
rect 26792 5108 26844 5160
rect 24400 5015 24452 5024
rect 24400 4981 24409 5015
rect 24409 4981 24443 5015
rect 24443 4981 24452 5015
rect 24400 4972 24452 4981
rect 25504 5015 25556 5024
rect 25504 4981 25513 5015
rect 25513 4981 25547 5015
rect 25547 4981 25556 5015
rect 25504 4972 25556 4981
rect 26332 4972 26384 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 3608 4768 3660 4820
rect 5356 4768 5408 4820
rect 5908 4768 5960 4820
rect 6184 4768 6236 4820
rect 6092 4632 6144 4684
rect 6552 4768 6604 4820
rect 7012 4768 7064 4820
rect 8024 4768 8076 4820
rect 9312 4768 9364 4820
rect 9404 4768 9456 4820
rect 6460 4700 6512 4752
rect 4988 4607 5040 4616
rect 4988 4573 4997 4607
rect 4997 4573 5031 4607
rect 5031 4573 5040 4607
rect 4988 4564 5040 4573
rect 5448 4564 5500 4616
rect 5816 4496 5868 4548
rect 6460 4607 6512 4616
rect 6460 4573 6469 4607
rect 6469 4573 6503 4607
rect 6503 4573 6512 4607
rect 6460 4564 6512 4573
rect 7472 4700 7524 4752
rect 7564 4700 7616 4752
rect 7012 4607 7064 4616
rect 7012 4573 7021 4607
rect 7021 4573 7055 4607
rect 7055 4573 7064 4607
rect 7012 4564 7064 4573
rect 8484 4675 8536 4684
rect 8484 4641 8493 4675
rect 8493 4641 8527 4675
rect 8527 4641 8536 4675
rect 8484 4632 8536 4641
rect 9588 4700 9640 4752
rect 9864 4632 9916 4684
rect 7748 4496 7800 4548
rect 8300 4564 8352 4616
rect 8392 4607 8444 4616
rect 8392 4573 8401 4607
rect 8401 4573 8435 4607
rect 8435 4573 8444 4607
rect 8392 4564 8444 4573
rect 8668 4607 8720 4616
rect 8668 4573 8677 4607
rect 8677 4573 8711 4607
rect 8711 4573 8720 4607
rect 8668 4564 8720 4573
rect 8760 4564 8812 4616
rect 9220 4607 9272 4616
rect 9220 4573 9229 4607
rect 9229 4573 9263 4607
rect 9263 4573 9272 4607
rect 9220 4564 9272 4573
rect 9496 4607 9548 4616
rect 9496 4573 9505 4607
rect 9505 4573 9539 4607
rect 9539 4573 9548 4607
rect 9496 4564 9548 4573
rect 9588 4607 9640 4616
rect 9588 4573 9597 4607
rect 9597 4573 9631 4607
rect 9631 4573 9640 4607
rect 9588 4564 9640 4573
rect 10140 4564 10192 4616
rect 10692 4607 10744 4616
rect 10692 4573 10701 4607
rect 10701 4573 10735 4607
rect 10735 4573 10744 4607
rect 10692 4564 10744 4573
rect 13912 4768 13964 4820
rect 16120 4811 16172 4820
rect 16120 4777 16129 4811
rect 16129 4777 16163 4811
rect 16163 4777 16172 4811
rect 16120 4768 16172 4777
rect 16396 4811 16448 4820
rect 16396 4777 16405 4811
rect 16405 4777 16439 4811
rect 16439 4777 16448 4811
rect 16396 4768 16448 4777
rect 18052 4768 18104 4820
rect 18512 4811 18564 4820
rect 18512 4777 18521 4811
rect 18521 4777 18555 4811
rect 18555 4777 18564 4811
rect 18512 4768 18564 4777
rect 24860 4768 24912 4820
rect 25504 4768 25556 4820
rect 25872 4768 25924 4820
rect 26240 4768 26292 4820
rect 12624 4700 12676 4752
rect 12440 4632 12492 4684
rect 12992 4675 13044 4684
rect 10508 4496 10560 4548
rect 12164 4607 12216 4616
rect 12164 4573 12173 4607
rect 12173 4573 12207 4607
rect 12207 4573 12216 4607
rect 12164 4564 12216 4573
rect 12992 4641 13001 4675
rect 13001 4641 13035 4675
rect 13035 4641 13044 4675
rect 12992 4632 13044 4641
rect 15568 4700 15620 4752
rect 16948 4700 17000 4752
rect 18696 4700 18748 4752
rect 15752 4675 15804 4684
rect 15752 4641 15761 4675
rect 15761 4641 15795 4675
rect 15795 4641 15804 4675
rect 15752 4632 15804 4641
rect 16488 4675 16540 4684
rect 16488 4641 16497 4675
rect 16497 4641 16531 4675
rect 16531 4641 16540 4675
rect 16488 4632 16540 4641
rect 12624 4607 12676 4616
rect 12624 4573 12633 4607
rect 12633 4573 12667 4607
rect 12667 4573 12676 4607
rect 12624 4564 12676 4573
rect 12808 4607 12860 4616
rect 12808 4573 12817 4607
rect 12817 4573 12851 4607
rect 12851 4573 12860 4607
rect 12808 4564 12860 4573
rect 12900 4607 12952 4616
rect 12900 4573 12909 4607
rect 12909 4573 12943 4607
rect 12943 4573 12952 4607
rect 12900 4564 12952 4573
rect 13176 4607 13228 4616
rect 13176 4573 13185 4607
rect 13185 4573 13219 4607
rect 13219 4573 13228 4607
rect 13176 4564 13228 4573
rect 13452 4607 13504 4616
rect 13452 4573 13461 4607
rect 13461 4573 13495 4607
rect 13495 4573 13504 4607
rect 13452 4564 13504 4573
rect 13636 4607 13688 4616
rect 13636 4573 13645 4607
rect 13645 4573 13679 4607
rect 13679 4573 13688 4607
rect 13636 4564 13688 4573
rect 13728 4607 13780 4616
rect 13728 4573 13737 4607
rect 13737 4573 13771 4607
rect 13771 4573 13780 4607
rect 13728 4564 13780 4573
rect 14556 4564 14608 4616
rect 15844 4607 15896 4616
rect 15844 4573 15853 4607
rect 15853 4573 15887 4607
rect 15887 4573 15896 4607
rect 15844 4564 15896 4573
rect 16212 4607 16264 4616
rect 16212 4573 16221 4607
rect 16221 4573 16255 4607
rect 16255 4573 16264 4607
rect 16212 4564 16264 4573
rect 16580 4564 16632 4616
rect 7564 4471 7616 4480
rect 7564 4437 7573 4471
rect 7573 4437 7607 4471
rect 7607 4437 7616 4471
rect 7564 4428 7616 4437
rect 7932 4428 7984 4480
rect 11980 4428 12032 4480
rect 12992 4428 13044 4480
rect 13360 4539 13412 4548
rect 13360 4505 13369 4539
rect 13369 4505 13403 4539
rect 13403 4505 13412 4539
rect 13360 4496 13412 4505
rect 15200 4496 15252 4548
rect 17316 4632 17368 4684
rect 19432 4700 19484 4752
rect 16856 4564 16908 4616
rect 17040 4607 17092 4616
rect 17040 4573 17049 4607
rect 17049 4573 17083 4607
rect 17083 4573 17092 4607
rect 17040 4564 17092 4573
rect 17224 4607 17276 4616
rect 17224 4573 17233 4607
rect 17233 4573 17267 4607
rect 17267 4573 17276 4607
rect 17224 4564 17276 4573
rect 19800 4632 19852 4684
rect 24400 4700 24452 4752
rect 23572 4632 23624 4684
rect 19064 4564 19116 4616
rect 13820 4471 13872 4480
rect 13820 4437 13829 4471
rect 13829 4437 13863 4471
rect 13863 4437 13872 4471
rect 13820 4428 13872 4437
rect 17132 4428 17184 4480
rect 19248 4539 19300 4548
rect 19248 4505 19257 4539
rect 19257 4505 19291 4539
rect 19291 4505 19300 4539
rect 19248 4496 19300 4505
rect 19616 4607 19668 4616
rect 19616 4573 19625 4607
rect 19625 4573 19659 4607
rect 19659 4573 19668 4607
rect 19616 4564 19668 4573
rect 20168 4607 20220 4616
rect 20168 4573 20177 4607
rect 20177 4573 20211 4607
rect 20211 4573 20220 4607
rect 20168 4564 20220 4573
rect 20444 4607 20496 4616
rect 20444 4573 20453 4607
rect 20453 4573 20487 4607
rect 20487 4573 20496 4607
rect 20444 4564 20496 4573
rect 22560 4496 22612 4548
rect 18788 4428 18840 4480
rect 19524 4471 19576 4480
rect 19524 4437 19533 4471
rect 19533 4437 19567 4471
rect 19567 4437 19576 4471
rect 19524 4428 19576 4437
rect 19984 4471 20036 4480
rect 19984 4437 19993 4471
rect 19993 4437 20027 4471
rect 20027 4437 20036 4471
rect 19984 4428 20036 4437
rect 20260 4471 20312 4480
rect 20260 4437 20269 4471
rect 20269 4437 20303 4471
rect 20303 4437 20312 4471
rect 20260 4428 20312 4437
rect 20996 4428 21048 4480
rect 25964 4607 26016 4616
rect 25964 4573 25973 4607
rect 25973 4573 26007 4607
rect 26007 4573 26016 4607
rect 25964 4564 26016 4573
rect 26700 4632 26752 4684
rect 27988 4675 28040 4684
rect 27988 4641 27997 4675
rect 27997 4641 28031 4675
rect 28031 4641 28040 4675
rect 27988 4632 28040 4641
rect 26608 4564 26660 4616
rect 28264 4607 28316 4616
rect 28264 4573 28273 4607
rect 28273 4573 28307 4607
rect 28307 4573 28316 4607
rect 28264 4564 28316 4573
rect 27252 4496 27304 4548
rect 26240 4428 26292 4480
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 6184 4267 6236 4276
rect 6184 4233 6193 4267
rect 6193 4233 6227 4267
rect 6227 4233 6236 4267
rect 6184 4224 6236 4233
rect 6276 4224 6328 4276
rect 5356 4156 5408 4208
rect 6000 4131 6052 4140
rect 6000 4097 6009 4131
rect 6009 4097 6043 4131
rect 6043 4097 6052 4131
rect 6000 4088 6052 4097
rect 6460 4088 6512 4140
rect 6736 4199 6788 4208
rect 6736 4165 6745 4199
rect 6745 4165 6779 4199
rect 6779 4165 6788 4199
rect 6736 4156 6788 4165
rect 7196 4156 7248 4208
rect 8300 4224 8352 4276
rect 9128 4224 9180 4276
rect 12072 4224 12124 4276
rect 12348 4224 12400 4276
rect 8392 4156 8444 4208
rect 5816 4063 5868 4072
rect 5816 4029 5825 4063
rect 5825 4029 5859 4063
rect 5859 4029 5868 4063
rect 5816 4020 5868 4029
rect 6644 4020 6696 4072
rect 7104 4131 7156 4140
rect 7104 4097 7113 4131
rect 7113 4097 7147 4131
rect 7147 4097 7156 4131
rect 7104 4088 7156 4097
rect 7288 4131 7340 4140
rect 7288 4097 7297 4131
rect 7297 4097 7331 4131
rect 7331 4097 7340 4131
rect 7288 4088 7340 4097
rect 8852 4156 8904 4208
rect 10600 4156 10652 4208
rect 11980 4199 12032 4208
rect 11980 4165 11989 4199
rect 11989 4165 12023 4199
rect 12023 4165 12032 4199
rect 11980 4156 12032 4165
rect 13728 4224 13780 4276
rect 8760 4088 8812 4140
rect 8576 4020 8628 4072
rect 9864 4088 9916 4140
rect 10508 4088 10560 4140
rect 11428 4088 11480 4140
rect 12992 4199 13044 4208
rect 12992 4165 13001 4199
rect 13001 4165 13035 4199
rect 13035 4165 13044 4199
rect 12992 4156 13044 4165
rect 13360 4156 13412 4208
rect 7564 3952 7616 4004
rect 7840 3952 7892 4004
rect 10232 4020 10284 4072
rect 11980 4020 12032 4072
rect 12348 4063 12400 4072
rect 12348 4029 12357 4063
rect 12357 4029 12391 4063
rect 12391 4029 12400 4063
rect 12348 4020 12400 4029
rect 6920 3927 6972 3936
rect 6920 3893 6929 3927
rect 6929 3893 6963 3927
rect 6963 3893 6972 3927
rect 6920 3884 6972 3893
rect 7656 3884 7708 3936
rect 8760 3927 8812 3936
rect 8760 3893 8769 3927
rect 8769 3893 8803 3927
rect 8803 3893 8812 3927
rect 8760 3884 8812 3893
rect 10876 3884 10928 3936
rect 13360 3995 13412 4004
rect 13360 3961 13369 3995
rect 13369 3961 13403 3995
rect 13403 3961 13412 3995
rect 13360 3952 13412 3961
rect 13544 4063 13596 4072
rect 13544 4029 13553 4063
rect 13553 4029 13587 4063
rect 13587 4029 13596 4063
rect 13544 4020 13596 4029
rect 13820 4131 13872 4140
rect 13820 4097 13829 4131
rect 13829 4097 13863 4131
rect 13863 4097 13872 4131
rect 13820 4088 13872 4097
rect 13912 4131 13964 4140
rect 13912 4097 13921 4131
rect 13921 4097 13955 4131
rect 13955 4097 13964 4131
rect 13912 4088 13964 4097
rect 17040 4224 17092 4276
rect 17224 4224 17276 4276
rect 15844 4156 15896 4208
rect 16396 4156 16448 4208
rect 19524 4224 19576 4276
rect 22560 4224 22612 4276
rect 14556 4131 14608 4140
rect 14556 4097 14565 4131
rect 14565 4097 14599 4131
rect 14599 4097 14608 4131
rect 14556 4088 14608 4097
rect 16580 4088 16632 4140
rect 16672 4131 16724 4140
rect 16672 4097 16681 4131
rect 16681 4097 16715 4131
rect 16715 4097 16724 4131
rect 16672 4088 16724 4097
rect 18880 4156 18932 4208
rect 17500 4088 17552 4140
rect 17960 4131 18012 4140
rect 17960 4097 17969 4131
rect 17969 4097 18003 4131
rect 18003 4097 18012 4131
rect 17960 4088 18012 4097
rect 15752 4020 15804 4072
rect 15936 4020 15988 4072
rect 16764 4020 16816 4072
rect 19708 4156 19760 4208
rect 19892 4088 19944 4140
rect 20168 4088 20220 4140
rect 20260 4131 20312 4140
rect 20260 4097 20269 4131
rect 20269 4097 20303 4131
rect 20303 4097 20312 4131
rect 20260 4088 20312 4097
rect 20628 4131 20680 4140
rect 20628 4097 20637 4131
rect 20637 4097 20671 4131
rect 20671 4097 20680 4131
rect 20628 4088 20680 4097
rect 20996 4131 21048 4140
rect 20996 4097 21005 4131
rect 21005 4097 21039 4131
rect 21039 4097 21048 4131
rect 20996 4088 21048 4097
rect 23572 4156 23624 4208
rect 25964 4224 26016 4276
rect 26240 4224 26292 4276
rect 26792 4224 26844 4276
rect 26608 4156 26660 4208
rect 25872 4131 25924 4140
rect 25872 4097 25881 4131
rect 25881 4097 25915 4131
rect 25915 4097 25924 4131
rect 25872 4088 25924 4097
rect 25964 4088 26016 4140
rect 27620 4088 27672 4140
rect 27712 4088 27764 4140
rect 13636 3952 13688 4004
rect 12716 3884 12768 3936
rect 12900 3884 12952 3936
rect 15200 3884 15252 3936
rect 16304 3927 16356 3936
rect 16304 3893 16313 3927
rect 16313 3893 16347 3927
rect 16347 3893 16356 3927
rect 16304 3884 16356 3893
rect 16580 3884 16632 3936
rect 18512 4020 18564 4072
rect 17592 3952 17644 4004
rect 19432 4020 19484 4072
rect 23296 4063 23348 4072
rect 23296 4029 23305 4063
rect 23305 4029 23339 4063
rect 23339 4029 23348 4063
rect 23296 4020 23348 4029
rect 25412 4063 25464 4072
rect 25412 4029 25421 4063
rect 25421 4029 25455 4063
rect 25455 4029 25464 4063
rect 25412 4020 25464 4029
rect 18328 3884 18380 3936
rect 25596 3952 25648 4004
rect 19984 3884 20036 3936
rect 20536 3884 20588 3936
rect 25688 3884 25740 3936
rect 26516 4020 26568 4072
rect 27252 3952 27304 4004
rect 27436 3952 27488 4004
rect 28172 3952 28224 4004
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 5816 3680 5868 3732
rect 9588 3680 9640 3732
rect 11428 3680 11480 3732
rect 11612 3680 11664 3732
rect 7196 3612 7248 3664
rect 7840 3655 7892 3664
rect 7840 3621 7849 3655
rect 7849 3621 7883 3655
rect 7883 3621 7892 3655
rect 7840 3612 7892 3621
rect 3332 3544 3384 3596
rect 6644 3587 6696 3596
rect 6644 3553 6653 3587
rect 6653 3553 6687 3587
rect 6687 3553 6696 3587
rect 6644 3544 6696 3553
rect 6920 3476 6972 3528
rect 7656 3519 7708 3528
rect 7656 3485 7665 3519
rect 7665 3485 7699 3519
rect 7699 3485 7708 3519
rect 7656 3476 7708 3485
rect 10876 3587 10928 3596
rect 10876 3553 10885 3587
rect 10885 3553 10919 3587
rect 10919 3553 10928 3587
rect 10876 3544 10928 3553
rect 11796 3612 11848 3664
rect 13728 3723 13780 3732
rect 13728 3689 13737 3723
rect 13737 3689 13771 3723
rect 13771 3689 13780 3723
rect 13728 3680 13780 3689
rect 11520 3587 11572 3596
rect 11520 3553 11529 3587
rect 11529 3553 11563 3587
rect 11563 3553 11572 3587
rect 11520 3544 11572 3553
rect 11428 3519 11480 3528
rect 11428 3485 11437 3519
rect 11437 3485 11471 3519
rect 11471 3485 11480 3519
rect 11428 3476 11480 3485
rect 5264 3340 5316 3392
rect 8208 3408 8260 3460
rect 10416 3408 10468 3460
rect 11980 3587 12032 3596
rect 11980 3553 11989 3587
rect 11989 3553 12023 3587
rect 12023 3553 12032 3587
rect 11980 3544 12032 3553
rect 12624 3544 12676 3596
rect 13360 3476 13412 3528
rect 15476 3680 15528 3732
rect 17592 3680 17644 3732
rect 17960 3680 18012 3732
rect 19248 3723 19300 3732
rect 19248 3689 19257 3723
rect 19257 3689 19291 3723
rect 19291 3689 19300 3723
rect 19248 3680 19300 3689
rect 19800 3680 19852 3732
rect 20628 3680 20680 3732
rect 16212 3655 16264 3664
rect 16212 3621 16221 3655
rect 16221 3621 16255 3655
rect 16255 3621 16264 3655
rect 16212 3612 16264 3621
rect 17040 3612 17092 3664
rect 15200 3519 15252 3528
rect 15200 3485 15209 3519
rect 15209 3485 15243 3519
rect 15243 3485 15252 3519
rect 15200 3476 15252 3485
rect 15476 3519 15528 3528
rect 15476 3485 15485 3519
rect 15485 3485 15519 3519
rect 15519 3485 15528 3519
rect 15476 3476 15528 3485
rect 12256 3451 12308 3460
rect 12256 3417 12265 3451
rect 12265 3417 12299 3451
rect 12299 3417 12308 3451
rect 12256 3408 12308 3417
rect 16028 3476 16080 3528
rect 16580 3519 16632 3528
rect 16580 3485 16586 3519
rect 16586 3485 16620 3519
rect 16620 3485 16632 3519
rect 16580 3476 16632 3485
rect 16948 3476 17000 3528
rect 10508 3340 10560 3392
rect 12992 3340 13044 3392
rect 13544 3340 13596 3392
rect 14096 3383 14148 3392
rect 14096 3349 14105 3383
rect 14105 3349 14139 3383
rect 14139 3349 14148 3383
rect 14096 3340 14148 3349
rect 15752 3383 15804 3392
rect 15752 3349 15761 3383
rect 15761 3349 15795 3383
rect 15795 3349 15804 3383
rect 15752 3340 15804 3349
rect 16028 3340 16080 3392
rect 16120 3340 16172 3392
rect 16856 3408 16908 3460
rect 17132 3408 17184 3460
rect 17408 3476 17460 3528
rect 20996 3612 21048 3664
rect 19708 3587 19760 3596
rect 19708 3553 19717 3587
rect 19717 3553 19751 3587
rect 19751 3553 19760 3587
rect 19708 3544 19760 3553
rect 19800 3587 19852 3596
rect 19800 3553 19809 3587
rect 19809 3553 19843 3587
rect 19843 3553 19852 3587
rect 19800 3544 19852 3553
rect 21548 3544 21600 3596
rect 25320 3612 25372 3664
rect 25964 3612 26016 3664
rect 26332 3680 26384 3732
rect 26516 3723 26568 3732
rect 26516 3689 26525 3723
rect 26525 3689 26559 3723
rect 26559 3689 26568 3723
rect 26516 3680 26568 3689
rect 26884 3612 26936 3664
rect 23572 3544 23624 3596
rect 28264 3587 28316 3596
rect 28264 3553 28273 3587
rect 28273 3553 28307 3587
rect 28307 3553 28316 3587
rect 28264 3544 28316 3553
rect 20168 3519 20220 3528
rect 16948 3340 17000 3392
rect 20168 3485 20177 3519
rect 20177 3485 20211 3519
rect 20211 3485 20220 3519
rect 20168 3476 20220 3485
rect 20536 3519 20588 3528
rect 20536 3485 20545 3519
rect 20545 3485 20579 3519
rect 20579 3485 20588 3519
rect 20536 3476 20588 3485
rect 21272 3519 21324 3528
rect 21272 3485 21281 3519
rect 21281 3485 21315 3519
rect 21315 3485 21324 3519
rect 21272 3476 21324 3485
rect 22836 3476 22888 3528
rect 23296 3519 23348 3528
rect 23296 3485 23305 3519
rect 23305 3485 23339 3519
rect 23339 3485 23348 3519
rect 23296 3476 23348 3485
rect 23388 3519 23440 3528
rect 23388 3485 23397 3519
rect 23397 3485 23431 3519
rect 23431 3485 23440 3519
rect 23388 3476 23440 3485
rect 25320 3519 25372 3528
rect 25320 3485 25329 3519
rect 25329 3485 25363 3519
rect 25363 3485 25372 3519
rect 25320 3476 25372 3485
rect 19340 3408 19392 3460
rect 19892 3408 19944 3460
rect 21548 3451 21600 3460
rect 21548 3417 21557 3451
rect 21557 3417 21591 3451
rect 21591 3417 21600 3451
rect 21548 3408 21600 3417
rect 22560 3408 22612 3460
rect 23940 3408 23992 3460
rect 19432 3340 19484 3392
rect 24308 3340 24360 3392
rect 24400 3340 24452 3392
rect 25596 3408 25648 3460
rect 25688 3451 25740 3460
rect 25688 3417 25697 3451
rect 25697 3417 25731 3451
rect 25731 3417 25740 3451
rect 25688 3408 25740 3417
rect 26240 3519 26292 3528
rect 26240 3485 26249 3519
rect 26249 3485 26283 3519
rect 26283 3485 26292 3519
rect 26240 3476 26292 3485
rect 26516 3408 26568 3460
rect 27436 3408 27488 3460
rect 27896 3408 27948 3460
rect 27160 3340 27212 3392
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 6000 3136 6052 3188
rect 6644 3068 6696 3120
rect 11612 3136 11664 3188
rect 12256 3136 12308 3188
rect 12900 3179 12952 3188
rect 12900 3145 12909 3179
rect 12909 3145 12943 3179
rect 12943 3145 12952 3179
rect 12900 3136 12952 3145
rect 13360 3179 13412 3188
rect 13360 3145 13369 3179
rect 13369 3145 13403 3179
rect 13403 3145 13412 3179
rect 13360 3136 13412 3145
rect 16396 3179 16448 3188
rect 16396 3145 16405 3179
rect 16405 3145 16439 3179
rect 16439 3145 16448 3179
rect 16396 3136 16448 3145
rect 16764 3179 16816 3188
rect 16764 3145 16773 3179
rect 16773 3145 16807 3179
rect 16807 3145 16816 3179
rect 16764 3136 16816 3145
rect 18972 3136 19024 3188
rect 19524 3179 19576 3188
rect 19524 3145 19533 3179
rect 19533 3145 19567 3179
rect 19567 3145 19576 3179
rect 19524 3136 19576 3145
rect 8760 3068 8812 3120
rect 10416 3068 10468 3120
rect 10508 3068 10560 3120
rect 8208 3043 8260 3052
rect 8208 3009 8217 3043
rect 8217 3009 8251 3043
rect 8251 3009 8260 3043
rect 8208 3000 8260 3009
rect 14096 3068 14148 3120
rect 14464 3111 14516 3120
rect 14464 3077 14473 3111
rect 14473 3077 14507 3111
rect 14507 3077 14516 3111
rect 14464 3068 14516 3077
rect 16304 3068 16356 3120
rect 7012 2932 7064 2984
rect 9864 2932 9916 2984
rect 12808 2932 12860 2984
rect 13084 2975 13136 2984
rect 13084 2941 13093 2975
rect 13093 2941 13127 2975
rect 13127 2941 13136 2975
rect 13084 2932 13136 2941
rect 16764 3000 16816 3052
rect 16948 3043 17000 3052
rect 16948 3009 16957 3043
rect 16957 3009 16991 3043
rect 16991 3009 17000 3043
rect 16948 3000 17000 3009
rect 17132 3043 17184 3052
rect 17132 3009 17141 3043
rect 17141 3009 17175 3043
rect 17175 3009 17184 3043
rect 17132 3000 17184 3009
rect 19340 3000 19392 3052
rect 19616 3000 19668 3052
rect 20536 3068 20588 3120
rect 22560 3068 22612 3120
rect 23848 3136 23900 3188
rect 25320 3136 25372 3188
rect 26240 3136 26292 3188
rect 26424 3179 26476 3188
rect 26424 3145 26433 3179
rect 26433 3145 26467 3179
rect 26467 3145 26476 3179
rect 26424 3136 26476 3145
rect 27712 3179 27764 3188
rect 27712 3145 27721 3179
rect 27721 3145 27755 3179
rect 27755 3145 27764 3179
rect 27712 3136 27764 3145
rect 24400 3068 24452 3120
rect 19984 3000 20036 3052
rect 21272 3000 21324 3052
rect 23572 3000 23624 3052
rect 28172 3111 28224 3120
rect 28172 3077 28181 3111
rect 28181 3077 28215 3111
rect 28215 3077 28224 3111
rect 28172 3068 28224 3077
rect 25964 3000 26016 3052
rect 17040 2932 17092 2984
rect 13452 2864 13504 2916
rect 22192 2932 22244 2984
rect 23388 2932 23440 2984
rect 14556 2796 14608 2848
rect 18328 2796 18380 2848
rect 21456 2796 21508 2848
rect 25688 2932 25740 2984
rect 27528 3043 27580 3052
rect 27528 3009 27537 3043
rect 27537 3009 27571 3043
rect 27571 3009 27580 3043
rect 27528 3000 27580 3009
rect 27620 2864 27672 2916
rect 23940 2839 23992 2848
rect 23940 2805 23970 2839
rect 23970 2805 23992 2839
rect 23940 2796 23992 2805
rect 26516 2796 26568 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 21548 2635 21600 2644
rect 21548 2601 21557 2635
rect 21557 2601 21591 2635
rect 21591 2601 21600 2635
rect 21548 2592 21600 2601
rect 22192 2635 22244 2644
rect 22192 2601 22201 2635
rect 22201 2601 22235 2635
rect 22235 2601 22244 2635
rect 22192 2592 22244 2601
rect 22836 2635 22888 2644
rect 22836 2601 22845 2635
rect 22845 2601 22879 2635
rect 22879 2601 22888 2635
rect 22836 2592 22888 2601
rect 23940 2592 23992 2644
rect 21272 2388 21324 2440
rect 21916 2388 21968 2440
rect 22560 2388 22612 2440
rect 23204 2388 23256 2440
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
<< metal2 >>
rect 4874 29404 5182 29413
rect 4874 29402 4880 29404
rect 4936 29402 4960 29404
rect 5016 29402 5040 29404
rect 5096 29402 5120 29404
rect 5176 29402 5182 29404
rect 4936 29350 4938 29402
rect 5118 29350 5120 29402
rect 4874 29348 4880 29350
rect 4936 29348 4960 29350
rect 5016 29348 5040 29350
rect 5096 29348 5120 29350
rect 5176 29348 5182 29350
rect 4874 29339 5182 29348
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4874 28316 5182 28325
rect 4874 28314 4880 28316
rect 4936 28314 4960 28316
rect 5016 28314 5040 28316
rect 5096 28314 5120 28316
rect 5176 28314 5182 28316
rect 4936 28262 4938 28314
rect 5118 28262 5120 28314
rect 4874 28260 4880 28262
rect 4936 28260 4960 28262
rect 5016 28260 5040 28262
rect 5096 28260 5120 28262
rect 5176 28260 5182 28262
rect 4874 28251 5182 28260
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4874 27228 5182 27237
rect 4874 27226 4880 27228
rect 4936 27226 4960 27228
rect 5016 27226 5040 27228
rect 5096 27226 5120 27228
rect 5176 27226 5182 27228
rect 4936 27174 4938 27226
rect 5118 27174 5120 27226
rect 4874 27172 4880 27174
rect 4936 27172 4960 27174
rect 5016 27172 5040 27174
rect 5096 27172 5120 27174
rect 5176 27172 5182 27174
rect 4874 27163 5182 27172
rect 110 27024 166 27033
rect 110 26959 166 26968
rect 124 14385 152 26959
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4874 26140 5182 26149
rect 4874 26138 4880 26140
rect 4936 26138 4960 26140
rect 5016 26138 5040 26140
rect 5096 26138 5120 26140
rect 5176 26138 5182 26140
rect 4936 26086 4938 26138
rect 5118 26086 5120 26138
rect 4874 26084 4880 26086
rect 4936 26084 4960 26086
rect 5016 26084 5040 26086
rect 5096 26084 5120 26086
rect 5176 26084 5182 26086
rect 4874 26075 5182 26084
rect 17776 25968 17828 25974
rect 17776 25910 17828 25916
rect 22836 25968 22888 25974
rect 22836 25910 22888 25916
rect 7840 25900 7892 25906
rect 7840 25842 7892 25848
rect 8576 25900 8628 25906
rect 8576 25842 8628 25848
rect 9588 25900 9640 25906
rect 9588 25842 9640 25848
rect 10324 25900 10376 25906
rect 10324 25842 10376 25848
rect 15292 25900 15344 25906
rect 15292 25842 15344 25848
rect 17684 25900 17736 25906
rect 17684 25842 17736 25848
rect 5540 25696 5592 25702
rect 5540 25638 5592 25644
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 5448 25356 5500 25362
rect 5448 25298 5500 25304
rect 4712 25288 4764 25294
rect 4712 25230 4764 25236
rect 4724 24886 4752 25230
rect 4874 25052 5182 25061
rect 4874 25050 4880 25052
rect 4936 25050 4960 25052
rect 5016 25050 5040 25052
rect 5096 25050 5120 25052
rect 5176 25050 5182 25052
rect 4936 24998 4938 25050
rect 5118 24998 5120 25050
rect 4874 24996 4880 24998
rect 4936 24996 4960 24998
rect 5016 24996 5040 24998
rect 5096 24996 5120 24998
rect 5176 24996 5182 24998
rect 4874 24987 5182 24996
rect 4712 24880 4764 24886
rect 4712 24822 4764 24828
rect 4804 24744 4856 24750
rect 4804 24686 4856 24692
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4816 21962 4844 24686
rect 5460 24614 5488 25298
rect 5552 25226 5580 25638
rect 7852 25294 7880 25842
rect 8392 25696 8444 25702
rect 8392 25638 8444 25644
rect 8404 25362 8432 25638
rect 8588 25498 8616 25842
rect 8944 25832 8996 25838
rect 8944 25774 8996 25780
rect 8956 25498 8984 25774
rect 8576 25492 8628 25498
rect 8576 25434 8628 25440
rect 8944 25492 8996 25498
rect 8944 25434 8996 25440
rect 8392 25356 8444 25362
rect 8392 25298 8444 25304
rect 9600 25294 9628 25842
rect 9772 25696 9824 25702
rect 9772 25638 9824 25644
rect 7840 25288 7892 25294
rect 7840 25230 7892 25236
rect 8760 25288 8812 25294
rect 8760 25230 8812 25236
rect 9588 25288 9640 25294
rect 9588 25230 9640 25236
rect 5540 25220 5592 25226
rect 5540 25162 5592 25168
rect 5908 25220 5960 25226
rect 5908 25162 5960 25168
rect 5920 24750 5948 25162
rect 6920 25152 6972 25158
rect 6920 25094 6972 25100
rect 7196 25152 7248 25158
rect 7196 25094 7248 25100
rect 6932 24886 6960 25094
rect 6920 24880 6972 24886
rect 6920 24822 6972 24828
rect 5908 24744 5960 24750
rect 5908 24686 5960 24692
rect 5448 24608 5500 24614
rect 5448 24550 5500 24556
rect 5460 24274 5488 24550
rect 5448 24268 5500 24274
rect 5448 24210 5500 24216
rect 5920 24070 5948 24686
rect 6920 24268 6972 24274
rect 6920 24210 6972 24216
rect 5908 24064 5960 24070
rect 5908 24006 5960 24012
rect 4874 23964 5182 23973
rect 4874 23962 4880 23964
rect 4936 23962 4960 23964
rect 5016 23962 5040 23964
rect 5096 23962 5120 23964
rect 5176 23962 5182 23964
rect 4936 23910 4938 23962
rect 5118 23910 5120 23962
rect 4874 23908 4880 23910
rect 4936 23908 4960 23910
rect 5016 23908 5040 23910
rect 5096 23908 5120 23910
rect 5176 23908 5182 23910
rect 4874 23899 5182 23908
rect 4874 22876 5182 22885
rect 4874 22874 4880 22876
rect 4936 22874 4960 22876
rect 5016 22874 5040 22876
rect 5096 22874 5120 22876
rect 5176 22874 5182 22876
rect 4936 22822 4938 22874
rect 5118 22822 5120 22874
rect 4874 22820 4880 22822
rect 4936 22820 4960 22822
rect 5016 22820 5040 22822
rect 5096 22820 5120 22822
rect 5176 22820 5182 22822
rect 4874 22811 5182 22820
rect 6932 22098 6960 24210
rect 7208 24138 7236 25094
rect 7852 24954 7880 25230
rect 7840 24948 7892 24954
rect 7840 24890 7892 24896
rect 8772 24410 8800 25230
rect 9680 25152 9732 25158
rect 9680 25094 9732 25100
rect 9588 24744 9640 24750
rect 9588 24686 9640 24692
rect 9128 24608 9180 24614
rect 9128 24550 9180 24556
rect 8760 24404 8812 24410
rect 8760 24346 8812 24352
rect 7196 24132 7248 24138
rect 7196 24074 7248 24080
rect 9140 23730 9168 24550
rect 9600 24274 9628 24686
rect 9692 24682 9720 25094
rect 9680 24676 9732 24682
rect 9680 24618 9732 24624
rect 9588 24268 9640 24274
rect 9588 24210 9640 24216
rect 9220 24132 9272 24138
rect 9220 24074 9272 24080
rect 9232 23866 9260 24074
rect 9220 23860 9272 23866
rect 9220 23802 9272 23808
rect 9784 23730 9812 25638
rect 9956 25424 10008 25430
rect 9956 25366 10008 25372
rect 9864 25152 9916 25158
rect 9864 25094 9916 25100
rect 9876 24614 9904 25094
rect 9968 24682 9996 25366
rect 10336 24886 10364 25842
rect 11980 25832 12032 25838
rect 11980 25774 12032 25780
rect 11060 25696 11112 25702
rect 11060 25638 11112 25644
rect 10692 25288 10744 25294
rect 10692 25230 10744 25236
rect 10416 25152 10468 25158
rect 10416 25094 10468 25100
rect 10324 24880 10376 24886
rect 10324 24822 10376 24828
rect 10428 24818 10456 25094
rect 10048 24812 10100 24818
rect 10048 24754 10100 24760
rect 10416 24812 10468 24818
rect 10416 24754 10468 24760
rect 9956 24676 10008 24682
rect 9956 24618 10008 24624
rect 9864 24608 9916 24614
rect 9864 24550 9916 24556
rect 9876 23798 9904 24550
rect 10060 23866 10088 24754
rect 10428 24410 10456 24754
rect 10416 24404 10468 24410
rect 10416 24346 10468 24352
rect 10704 24274 10732 25230
rect 10968 25220 11020 25226
rect 10968 25162 11020 25168
rect 10980 24954 11008 25162
rect 10968 24948 11020 24954
rect 10968 24890 11020 24896
rect 11072 24750 11100 25638
rect 11992 25498 12020 25774
rect 11980 25492 12032 25498
rect 11980 25434 12032 25440
rect 11520 24812 11572 24818
rect 11520 24754 11572 24760
rect 11060 24744 11112 24750
rect 11060 24686 11112 24692
rect 10968 24608 11020 24614
rect 10968 24550 11020 24556
rect 10692 24268 10744 24274
rect 10692 24210 10744 24216
rect 10048 23860 10100 23866
rect 10048 23802 10100 23808
rect 9864 23792 9916 23798
rect 9864 23734 9916 23740
rect 9128 23724 9180 23730
rect 9128 23666 9180 23672
rect 9772 23724 9824 23730
rect 9772 23666 9824 23672
rect 10980 23186 11008 24550
rect 11060 24404 11112 24410
rect 11060 24346 11112 24352
rect 11072 23730 11100 24346
rect 11244 24132 11296 24138
rect 11244 24074 11296 24080
rect 11060 23724 11112 23730
rect 11060 23666 11112 23672
rect 11152 23520 11204 23526
rect 11152 23462 11204 23468
rect 10968 23180 11020 23186
rect 10968 23122 11020 23128
rect 11164 23118 11192 23462
rect 11256 23322 11284 24074
rect 11532 23594 11560 24754
rect 11796 24744 11848 24750
rect 11796 24686 11848 24692
rect 11808 24274 11836 24686
rect 11796 24268 11848 24274
rect 11796 24210 11848 24216
rect 11702 24168 11758 24177
rect 11702 24103 11704 24112
rect 11756 24103 11758 24112
rect 11704 24074 11756 24080
rect 11612 24064 11664 24070
rect 11612 24006 11664 24012
rect 11624 23730 11652 24006
rect 11612 23724 11664 23730
rect 11612 23666 11664 23672
rect 11520 23588 11572 23594
rect 11520 23530 11572 23536
rect 11244 23316 11296 23322
rect 11244 23258 11296 23264
rect 11152 23112 11204 23118
rect 11152 23054 11204 23060
rect 8116 22704 8168 22710
rect 8116 22646 8168 22652
rect 7748 22636 7800 22642
rect 7748 22578 7800 22584
rect 6920 22092 6972 22098
rect 6920 22034 6972 22040
rect 5814 21992 5870 22001
rect 4804 21956 4856 21962
rect 4804 21898 4856 21904
rect 5540 21956 5592 21962
rect 5814 21927 5870 21936
rect 6276 21956 6328 21962
rect 5540 21898 5592 21904
rect 4068 21888 4120 21894
rect 4068 21830 4120 21836
rect 4080 21554 4108 21830
rect 4068 21548 4120 21554
rect 4068 21490 4120 21496
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4712 20868 4764 20874
rect 4712 20810 4764 20816
rect 3608 20392 3660 20398
rect 3608 20334 3660 20340
rect 3620 19718 3648 20334
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 3608 19712 3660 19718
rect 3608 19654 3660 19660
rect 3620 18086 3648 19654
rect 4724 19446 4752 20810
rect 4816 20602 4844 21898
rect 4874 21788 5182 21797
rect 4874 21786 4880 21788
rect 4936 21786 4960 21788
rect 5016 21786 5040 21788
rect 5096 21786 5120 21788
rect 5176 21786 5182 21788
rect 4936 21734 4938 21786
rect 5118 21734 5120 21786
rect 4874 21732 4880 21734
rect 4936 21732 4960 21734
rect 5016 21732 5040 21734
rect 5096 21732 5120 21734
rect 5176 21732 5182 21734
rect 4874 21723 5182 21732
rect 5552 21690 5580 21898
rect 5540 21684 5592 21690
rect 5540 21626 5592 21632
rect 4988 21616 5040 21622
rect 4988 21558 5040 21564
rect 5000 20874 5028 21558
rect 5368 21554 5672 21570
rect 5828 21554 5856 21927
rect 6276 21898 6328 21904
rect 5080 21548 5132 21554
rect 5080 21490 5132 21496
rect 5356 21548 5672 21554
rect 5408 21542 5672 21548
rect 5356 21490 5408 21496
rect 5092 21010 5120 21490
rect 5356 21412 5408 21418
rect 5356 21354 5408 21360
rect 5080 21004 5132 21010
rect 5080 20946 5132 20952
rect 5368 20942 5396 21354
rect 5172 20936 5224 20942
rect 5356 20936 5408 20942
rect 5224 20896 5304 20924
rect 5172 20878 5224 20884
rect 4988 20868 5040 20874
rect 4988 20810 5040 20816
rect 4874 20700 5182 20709
rect 4874 20698 4880 20700
rect 4936 20698 4960 20700
rect 5016 20698 5040 20700
rect 5096 20698 5120 20700
rect 5176 20698 5182 20700
rect 4936 20646 4938 20698
rect 5118 20646 5120 20698
rect 4874 20644 4880 20646
rect 4936 20644 4960 20646
rect 5016 20644 5040 20646
rect 5096 20644 5120 20646
rect 5176 20644 5182 20646
rect 4874 20635 5182 20644
rect 4804 20596 4856 20602
rect 4804 20538 4856 20544
rect 5276 20262 5304 20896
rect 5356 20878 5408 20884
rect 5540 20936 5592 20942
rect 5540 20878 5592 20884
rect 5552 20618 5580 20878
rect 5644 20788 5672 21542
rect 5816 21548 5868 21554
rect 5816 21490 5868 21496
rect 6092 21548 6144 21554
rect 6092 21490 6144 21496
rect 5724 21480 5776 21486
rect 5724 21422 5776 21428
rect 5736 21146 5764 21422
rect 5724 21140 5776 21146
rect 5724 21082 5776 21088
rect 5828 20942 5856 21490
rect 6104 21350 6132 21490
rect 6092 21344 6144 21350
rect 6092 21286 6144 21292
rect 6184 21344 6236 21350
rect 6184 21286 6236 21292
rect 6196 20942 6224 21286
rect 6288 21146 6316 21898
rect 7012 21888 7064 21894
rect 7012 21830 7064 21836
rect 6920 21548 6972 21554
rect 6920 21490 6972 21496
rect 6932 21350 6960 21490
rect 6920 21344 6972 21350
rect 6920 21286 6972 21292
rect 6276 21140 6328 21146
rect 6276 21082 6328 21088
rect 5816 20936 5868 20942
rect 5816 20878 5868 20884
rect 6184 20936 6236 20942
rect 6184 20878 6236 20884
rect 5908 20868 5960 20874
rect 5908 20810 5960 20816
rect 6368 20868 6420 20874
rect 6368 20810 6420 20816
rect 5644 20760 5856 20788
rect 5368 20590 5580 20618
rect 5264 20256 5316 20262
rect 5264 20198 5316 20204
rect 4874 19612 5182 19621
rect 4874 19610 4880 19612
rect 4936 19610 4960 19612
rect 5016 19610 5040 19612
rect 5096 19610 5120 19612
rect 5176 19610 5182 19612
rect 4936 19558 4938 19610
rect 5118 19558 5120 19610
rect 4874 19556 4880 19558
rect 4936 19556 4960 19558
rect 5016 19556 5040 19558
rect 5096 19556 5120 19558
rect 5176 19556 5182 19558
rect 4874 19547 5182 19556
rect 4712 19440 4764 19446
rect 4712 19382 4764 19388
rect 5262 19408 5318 19417
rect 4068 19168 4120 19174
rect 4068 19110 4120 19116
rect 4080 18358 4108 19110
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4436 18692 4488 18698
rect 4436 18634 4488 18640
rect 3700 18352 3752 18358
rect 3700 18294 3752 18300
rect 4068 18352 4120 18358
rect 4068 18294 4120 18300
rect 1860 18080 1912 18086
rect 1860 18022 1912 18028
rect 3608 18080 3660 18086
rect 3608 18022 3660 18028
rect 1872 17746 1900 18022
rect 1860 17740 1912 17746
rect 1860 17682 1912 17688
rect 3712 17678 3740 18294
rect 4080 18154 4200 18170
rect 4448 18154 4476 18634
rect 4528 18624 4580 18630
rect 4528 18566 4580 18572
rect 4540 18290 4568 18566
rect 4528 18284 4580 18290
rect 4528 18226 4580 18232
rect 4620 18216 4672 18222
rect 4620 18158 4672 18164
rect 4080 18148 4212 18154
rect 4080 18142 4160 18148
rect 4080 17882 4108 18142
rect 4160 18090 4212 18096
rect 4436 18148 4488 18154
rect 4436 18090 4488 18096
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4632 17882 4660 18158
rect 4068 17876 4120 17882
rect 4068 17818 4120 17824
rect 4620 17876 4672 17882
rect 4620 17818 4672 17824
rect 4724 17678 4752 19382
rect 4988 19372 5040 19378
rect 5262 19343 5264 19352
rect 4988 19314 5040 19320
rect 5316 19343 5318 19352
rect 5264 19314 5316 19320
rect 5000 19258 5028 19314
rect 5368 19258 5396 20590
rect 5828 20534 5856 20760
rect 5920 20602 5948 20810
rect 5908 20596 5960 20602
rect 5908 20538 5960 20544
rect 5448 20528 5500 20534
rect 5448 20470 5500 20476
rect 5816 20528 5868 20534
rect 5816 20470 5868 20476
rect 4804 19236 4856 19242
rect 5000 19230 5396 19258
rect 4804 19178 4856 19184
rect 4816 18766 4844 19178
rect 5264 18896 5316 18902
rect 5264 18838 5316 18844
rect 4804 18760 4856 18766
rect 4804 18702 4856 18708
rect 4816 18426 4844 18702
rect 4874 18524 5182 18533
rect 4874 18522 4880 18524
rect 4936 18522 4960 18524
rect 5016 18522 5040 18524
rect 5096 18522 5120 18524
rect 5176 18522 5182 18524
rect 4936 18470 4938 18522
rect 5118 18470 5120 18522
rect 4874 18468 4880 18470
rect 4936 18468 4960 18470
rect 5016 18468 5040 18470
rect 5096 18468 5120 18470
rect 5176 18468 5182 18470
rect 4874 18459 5182 18468
rect 4804 18420 4856 18426
rect 4804 18362 4856 18368
rect 5080 18420 5132 18426
rect 5080 18362 5132 18368
rect 4816 18290 5028 18306
rect 4804 18284 5028 18290
rect 4856 18278 5028 18284
rect 4804 18226 4856 18232
rect 4896 18216 4948 18222
rect 4896 18158 4948 18164
rect 4804 18148 4856 18154
rect 4804 18090 4856 18096
rect 3700 17672 3752 17678
rect 3700 17614 3752 17620
rect 4620 17672 4672 17678
rect 4620 17614 4672 17620
rect 4712 17672 4764 17678
rect 4712 17614 4764 17620
rect 3712 16182 3740 17614
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4436 16652 4488 16658
rect 4436 16594 4488 16600
rect 4448 16250 4476 16594
rect 4632 16250 4660 17614
rect 4712 17536 4764 17542
rect 4712 17478 4764 17484
rect 4436 16244 4488 16250
rect 4436 16186 4488 16192
rect 4620 16244 4672 16250
rect 4620 16186 4672 16192
rect 3700 16176 3752 16182
rect 3700 16118 3752 16124
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 110 14376 166 14385
rect 4724 14362 4752 17478
rect 4816 16794 4844 18090
rect 4908 17678 4936 18158
rect 5000 17746 5028 18278
rect 4988 17740 5040 17746
rect 4988 17682 5040 17688
rect 5092 17678 5120 18362
rect 5276 18290 5304 18838
rect 5264 18284 5316 18290
rect 5264 18226 5316 18232
rect 5368 18170 5396 19230
rect 5460 19174 5488 20470
rect 5724 20460 5776 20466
rect 5724 20402 5776 20408
rect 5540 20392 5592 20398
rect 5736 20346 5764 20402
rect 5540 20334 5592 20340
rect 5552 19378 5580 20334
rect 5644 20318 5764 20346
rect 5644 20262 5672 20318
rect 5632 20256 5684 20262
rect 5632 20198 5684 20204
rect 5644 19394 5672 20198
rect 5920 19922 5948 20538
rect 6380 20534 6408 20810
rect 6932 20534 6960 21286
rect 7024 20874 7052 21830
rect 7564 21548 7616 21554
rect 7564 21490 7616 21496
rect 7196 21412 7248 21418
rect 7196 21354 7248 21360
rect 7012 20868 7064 20874
rect 7012 20810 7064 20816
rect 6368 20528 6420 20534
rect 6368 20470 6420 20476
rect 6920 20528 6972 20534
rect 6920 20470 6972 20476
rect 6932 19990 6960 20470
rect 7024 20262 7052 20810
rect 7208 20466 7236 21354
rect 7576 20874 7604 21490
rect 7564 20868 7616 20874
rect 7564 20810 7616 20816
rect 7196 20460 7248 20466
rect 7196 20402 7248 20408
rect 7288 20460 7340 20466
rect 7288 20402 7340 20408
rect 7012 20256 7064 20262
rect 7012 20198 7064 20204
rect 6920 19984 6972 19990
rect 6920 19926 6972 19932
rect 5908 19916 5960 19922
rect 5908 19858 5960 19864
rect 6828 19712 6880 19718
rect 6828 19654 6880 19660
rect 5644 19378 5948 19394
rect 6840 19378 6868 19654
rect 5540 19372 5592 19378
rect 5540 19314 5592 19320
rect 5632 19372 5960 19378
rect 5684 19366 5908 19372
rect 5632 19314 5684 19320
rect 5908 19314 5960 19320
rect 6092 19372 6144 19378
rect 6092 19314 6144 19320
rect 6828 19372 6880 19378
rect 6828 19314 6880 19320
rect 5448 19168 5500 19174
rect 5448 19110 5500 19116
rect 5448 18964 5500 18970
rect 5448 18906 5500 18912
rect 5460 18426 5488 18906
rect 5540 18760 5592 18766
rect 5540 18702 5592 18708
rect 5448 18420 5500 18426
rect 5448 18362 5500 18368
rect 5460 18290 5488 18362
rect 5448 18284 5500 18290
rect 5448 18226 5500 18232
rect 5184 18142 5396 18170
rect 4896 17672 4948 17678
rect 4896 17614 4948 17620
rect 5080 17672 5132 17678
rect 5080 17614 5132 17620
rect 5080 17536 5132 17542
rect 5184 17524 5212 18142
rect 5264 18080 5316 18086
rect 5264 18022 5316 18028
rect 5356 18080 5408 18086
rect 5356 18022 5408 18028
rect 5276 17762 5304 18022
rect 5368 17882 5396 18022
rect 5460 17882 5488 18226
rect 5552 18086 5580 18702
rect 5644 18086 5672 19314
rect 6104 18970 6132 19314
rect 6092 18964 6144 18970
rect 6092 18906 6144 18912
rect 5908 18828 5960 18834
rect 5908 18770 5960 18776
rect 5724 18760 5776 18766
rect 5724 18702 5776 18708
rect 5540 18080 5592 18086
rect 5540 18022 5592 18028
rect 5632 18080 5684 18086
rect 5632 18022 5684 18028
rect 5356 17876 5408 17882
rect 5356 17818 5408 17824
rect 5448 17876 5500 17882
rect 5448 17818 5500 17824
rect 5276 17734 5396 17762
rect 5264 17604 5316 17610
rect 5264 17546 5316 17552
rect 5132 17496 5212 17524
rect 5080 17478 5132 17484
rect 4874 17436 5182 17445
rect 4874 17434 4880 17436
rect 4936 17434 4960 17436
rect 5016 17434 5040 17436
rect 5096 17434 5120 17436
rect 5176 17434 5182 17436
rect 4936 17382 4938 17434
rect 5118 17382 5120 17434
rect 4874 17380 4880 17382
rect 4936 17380 4960 17382
rect 5016 17380 5040 17382
rect 5096 17380 5120 17382
rect 5176 17380 5182 17382
rect 4874 17371 5182 17380
rect 5276 17338 5304 17546
rect 5264 17332 5316 17338
rect 5264 17274 5316 17280
rect 5264 17196 5316 17202
rect 5368 17184 5396 17734
rect 5460 17202 5488 17818
rect 5736 17678 5764 18702
rect 5816 18624 5868 18630
rect 5816 18566 5868 18572
rect 5828 18426 5856 18566
rect 5816 18420 5868 18426
rect 5816 18362 5868 18368
rect 5920 18290 5948 18770
rect 6000 18760 6052 18766
rect 6000 18702 6052 18708
rect 5908 18284 5960 18290
rect 5908 18226 5960 18232
rect 5816 18148 5868 18154
rect 5816 18090 5868 18096
rect 5828 17678 5856 18090
rect 6012 17882 6040 18702
rect 6644 18080 6696 18086
rect 6644 18022 6696 18028
rect 6000 17876 6052 17882
rect 6000 17818 6052 17824
rect 5540 17672 5592 17678
rect 5540 17614 5592 17620
rect 5724 17672 5776 17678
rect 5724 17614 5776 17620
rect 5816 17672 5868 17678
rect 5816 17614 5868 17620
rect 5552 17338 5580 17614
rect 5540 17332 5592 17338
rect 5540 17274 5592 17280
rect 5316 17156 5396 17184
rect 5448 17196 5500 17202
rect 5264 17138 5316 17144
rect 5448 17138 5500 17144
rect 4804 16788 4856 16794
rect 4804 16730 4856 16736
rect 5460 16658 5488 17138
rect 5736 17134 5764 17614
rect 6012 17270 6040 17818
rect 6656 17678 6684 18022
rect 6932 17882 6960 19926
rect 7024 19854 7052 20198
rect 7208 20058 7236 20402
rect 7196 20052 7248 20058
rect 7196 19994 7248 20000
rect 7300 19854 7328 20402
rect 7576 20398 7604 20810
rect 7564 20392 7616 20398
rect 7564 20334 7616 20340
rect 7012 19848 7064 19854
rect 7012 19790 7064 19796
rect 7288 19848 7340 19854
rect 7288 19790 7340 19796
rect 7576 19378 7604 20334
rect 7760 20058 7788 22578
rect 7840 22500 7892 22506
rect 7840 22442 7892 22448
rect 7852 22094 7880 22442
rect 8128 22098 8156 22646
rect 9680 22636 9732 22642
rect 9680 22578 9732 22584
rect 9036 22432 9088 22438
rect 9036 22374 9088 22380
rect 7932 22094 7984 22098
rect 7852 22092 7984 22094
rect 7852 22066 7932 22092
rect 7932 22034 7984 22040
rect 8116 22092 8168 22098
rect 8116 22034 8168 22040
rect 7944 21962 7972 22034
rect 7840 21956 7892 21962
rect 7840 21898 7892 21904
rect 7932 21956 7984 21962
rect 7932 21898 7984 21904
rect 7852 21690 7880 21898
rect 7840 21684 7892 21690
rect 7840 21626 7892 21632
rect 7852 20942 7880 21626
rect 7840 20936 7892 20942
rect 7840 20878 7892 20884
rect 8128 20602 8156 22034
rect 8576 22024 8628 22030
rect 8576 21966 8628 21972
rect 8392 20936 8444 20942
rect 8392 20878 8444 20884
rect 8208 20800 8260 20806
rect 8208 20742 8260 20748
rect 8116 20596 8168 20602
rect 8116 20538 8168 20544
rect 8116 20392 8168 20398
rect 8116 20334 8168 20340
rect 8128 20058 8156 20334
rect 7748 20052 7800 20058
rect 7748 19994 7800 20000
rect 8116 20052 8168 20058
rect 8116 19994 8168 20000
rect 8220 19854 8248 20742
rect 8404 20534 8432 20878
rect 8588 20534 8616 21966
rect 8668 21480 8720 21486
rect 8668 21422 8720 21428
rect 8392 20528 8444 20534
rect 8392 20470 8444 20476
rect 8576 20528 8628 20534
rect 8576 20470 8628 20476
rect 8588 20398 8616 20470
rect 8576 20392 8628 20398
rect 8576 20334 8628 20340
rect 8300 20256 8352 20262
rect 8300 20198 8352 20204
rect 7748 19848 7800 19854
rect 7748 19790 7800 19796
rect 8208 19848 8260 19854
rect 8208 19790 8260 19796
rect 7564 19372 7616 19378
rect 7564 19314 7616 19320
rect 7564 19236 7616 19242
rect 7564 19178 7616 19184
rect 7576 18426 7604 19178
rect 7760 18698 7788 19790
rect 8312 19786 8340 20198
rect 8300 19780 8352 19786
rect 8300 19722 8352 19728
rect 8116 19440 8168 19446
rect 8116 19382 8168 19388
rect 7748 18692 7800 18698
rect 7748 18634 7800 18640
rect 7564 18420 7616 18426
rect 7564 18362 7616 18368
rect 7760 18290 7788 18634
rect 7748 18284 7800 18290
rect 8128 18272 8156 19382
rect 8208 18284 8260 18290
rect 8128 18244 8208 18272
rect 7748 18226 7800 18232
rect 8208 18226 8260 18232
rect 6920 17876 6972 17882
rect 6920 17818 6972 17824
rect 6552 17672 6604 17678
rect 6552 17614 6604 17620
rect 6644 17672 6696 17678
rect 6644 17614 6696 17620
rect 6828 17672 6880 17678
rect 7012 17672 7064 17678
rect 6880 17620 6960 17626
rect 6828 17614 6960 17620
rect 7012 17614 7064 17620
rect 6184 17604 6236 17610
rect 6184 17546 6236 17552
rect 6000 17264 6052 17270
rect 6000 17206 6052 17212
rect 5724 17128 5776 17134
rect 5724 17070 5776 17076
rect 5632 16788 5684 16794
rect 5632 16730 5684 16736
rect 5448 16652 5500 16658
rect 5448 16594 5500 16600
rect 4874 16348 5182 16357
rect 4874 16346 4880 16348
rect 4936 16346 4960 16348
rect 5016 16346 5040 16348
rect 5096 16346 5120 16348
rect 5176 16346 5182 16348
rect 4936 16294 4938 16346
rect 5118 16294 5120 16346
rect 4874 16292 4880 16294
rect 4936 16292 4960 16294
rect 5016 16292 5040 16294
rect 5096 16292 5120 16294
rect 5176 16292 5182 16294
rect 4874 16283 5182 16292
rect 5540 16244 5592 16250
rect 5460 16204 5540 16232
rect 5356 15904 5408 15910
rect 5356 15846 5408 15852
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 4724 14334 4844 14362
rect 110 14311 166 14320
rect 4712 14272 4764 14278
rect 4712 14214 4764 14220
rect 4724 14006 4752 14214
rect 4712 14000 4764 14006
rect 4712 13942 4764 13948
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4620 13184 4672 13190
rect 4620 13126 4672 13132
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4632 11830 4660 13126
rect 4816 12238 4844 14334
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 5368 14074 5396 15846
rect 5460 14521 5488 16204
rect 5540 16186 5592 16192
rect 5446 14512 5502 14521
rect 5644 14482 5672 16730
rect 6196 16658 6224 17546
rect 6564 17270 6592 17614
rect 6840 17598 6960 17614
rect 6552 17264 6604 17270
rect 6552 17206 6604 17212
rect 6932 17202 6960 17598
rect 7024 17202 7052 17614
rect 6920 17196 6972 17202
rect 6920 17138 6972 17144
rect 7012 17196 7064 17202
rect 7012 17138 7064 17144
rect 6460 17060 6512 17066
rect 6460 17002 6512 17008
rect 6184 16652 6236 16658
rect 6184 16594 6236 16600
rect 6472 16590 6500 17002
rect 6460 16584 6512 16590
rect 6460 16526 6512 16532
rect 6552 16584 6604 16590
rect 6552 16526 6604 16532
rect 6736 16584 6788 16590
rect 6736 16526 6788 16532
rect 6000 16448 6052 16454
rect 6000 16390 6052 16396
rect 6012 16182 6040 16390
rect 6000 16176 6052 16182
rect 6000 16118 6052 16124
rect 6564 15366 6592 16526
rect 6748 16250 6776 16526
rect 6932 16250 6960 17138
rect 6736 16244 6788 16250
rect 6736 16186 6788 16192
rect 6920 16244 6972 16250
rect 6920 16186 6972 16192
rect 6552 15360 6604 15366
rect 6552 15302 6604 15308
rect 6276 15088 6328 15094
rect 6276 15030 6328 15036
rect 5446 14447 5502 14456
rect 5632 14476 5684 14482
rect 5460 14414 5488 14447
rect 5632 14418 5684 14424
rect 5448 14408 5500 14414
rect 5448 14350 5500 14356
rect 5908 14408 5960 14414
rect 5908 14350 5960 14356
rect 5724 14272 5776 14278
rect 5724 14214 5776 14220
rect 5356 14068 5408 14074
rect 5356 14010 5408 14016
rect 5368 13394 5396 14010
rect 5356 13388 5408 13394
rect 5356 13330 5408 13336
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 4804 12232 4856 12238
rect 4804 12174 4856 12180
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 5368 11898 5396 13330
rect 5736 13274 5764 14214
rect 5816 13932 5868 13938
rect 5816 13874 5868 13880
rect 5644 13258 5764 13274
rect 5828 13258 5856 13874
rect 5632 13252 5764 13258
rect 5684 13246 5764 13252
rect 5816 13252 5868 13258
rect 5632 13194 5684 13200
rect 5816 13194 5868 13200
rect 5920 13138 5948 14350
rect 6288 14278 6316 15030
rect 7024 15026 7052 17138
rect 7760 16658 7788 18226
rect 8312 18222 8340 19722
rect 8588 18766 8616 20334
rect 8680 20058 8708 21422
rect 8668 20052 8720 20058
rect 8668 19994 8720 20000
rect 9048 19854 9076 22374
rect 9588 21956 9640 21962
rect 9588 21898 9640 21904
rect 9128 21888 9180 21894
rect 9128 21830 9180 21836
rect 9140 20942 9168 21830
rect 9600 21554 9628 21898
rect 9220 21548 9272 21554
rect 9220 21490 9272 21496
rect 9588 21548 9640 21554
rect 9588 21490 9640 21496
rect 9232 21010 9260 21490
rect 9220 21004 9272 21010
rect 9220 20946 9272 20952
rect 9128 20936 9180 20942
rect 9128 20878 9180 20884
rect 9312 20936 9364 20942
rect 9312 20878 9364 20884
rect 9324 20806 9352 20878
rect 9312 20800 9364 20806
rect 9364 20760 9444 20788
rect 9312 20742 9364 20748
rect 9416 20602 9444 20760
rect 9404 20596 9456 20602
rect 9404 20538 9456 20544
rect 9586 20496 9642 20505
rect 9586 20431 9642 20440
rect 9600 20398 9628 20431
rect 9588 20392 9640 20398
rect 9588 20334 9640 20340
rect 9588 20256 9640 20262
rect 9588 20198 9640 20204
rect 9036 19848 9088 19854
rect 9036 19790 9088 19796
rect 9600 19718 9628 20198
rect 8852 19712 8904 19718
rect 8852 19654 8904 19660
rect 9588 19712 9640 19718
rect 9588 19654 9640 19660
rect 8864 19417 8892 19654
rect 8850 19408 8906 19417
rect 8850 19343 8906 19352
rect 8944 19372 8996 19378
rect 8576 18760 8628 18766
rect 8576 18702 8628 18708
rect 8864 18630 8892 19343
rect 8944 19314 8996 19320
rect 8956 19174 8984 19314
rect 8944 19168 8996 19174
rect 8944 19110 8996 19116
rect 9312 19168 9364 19174
rect 9312 19110 9364 19116
rect 8956 18970 8984 19110
rect 8944 18964 8996 18970
rect 8944 18906 8996 18912
rect 8852 18624 8904 18630
rect 8852 18566 8904 18572
rect 8668 18284 8720 18290
rect 8668 18226 8720 18232
rect 8300 18216 8352 18222
rect 8300 18158 8352 18164
rect 8392 18216 8444 18222
rect 8392 18158 8444 18164
rect 8300 18080 8352 18086
rect 8300 18022 8352 18028
rect 8312 17762 8340 18022
rect 8404 17882 8432 18158
rect 8576 18148 8628 18154
rect 8576 18090 8628 18096
rect 8392 17876 8444 17882
rect 8392 17818 8444 17824
rect 8588 17762 8616 18090
rect 8680 17882 8708 18226
rect 8864 18222 8892 18566
rect 8852 18216 8904 18222
rect 8852 18158 8904 18164
rect 9220 18216 9272 18222
rect 9220 18158 9272 18164
rect 8668 17876 8720 17882
rect 8668 17818 8720 17824
rect 8312 17734 8432 17762
rect 8588 17734 8708 17762
rect 8404 17610 8432 17734
rect 8392 17604 8444 17610
rect 8392 17546 8444 17552
rect 8404 17270 8432 17546
rect 8392 17264 8444 17270
rect 8392 17206 8444 17212
rect 7748 16652 7800 16658
rect 7748 16594 7800 16600
rect 8404 16454 8432 17206
rect 8484 17196 8536 17202
rect 8484 17138 8536 17144
rect 8392 16448 8444 16454
rect 8392 16390 8444 16396
rect 8404 16114 8432 16390
rect 8392 16108 8444 16114
rect 8392 16050 8444 16056
rect 7932 16040 7984 16046
rect 7932 15982 7984 15988
rect 8024 16040 8076 16046
rect 8024 15982 8076 15988
rect 7472 15360 7524 15366
rect 7472 15302 7524 15308
rect 7484 15162 7512 15302
rect 7472 15156 7524 15162
rect 7472 15098 7524 15104
rect 7012 15020 7064 15026
rect 7012 14962 7064 14968
rect 6552 14816 6604 14822
rect 6552 14758 6604 14764
rect 6276 14272 6328 14278
rect 6276 14214 6328 14220
rect 6368 14272 6420 14278
rect 6368 14214 6420 14220
rect 6288 13802 6316 14214
rect 6380 14074 6408 14214
rect 6368 14068 6420 14074
rect 6368 14010 6420 14016
rect 6564 13938 6592 14758
rect 7012 14612 7064 14618
rect 7012 14554 7064 14560
rect 6644 14476 6696 14482
rect 6644 14418 6696 14424
rect 6552 13932 6604 13938
rect 6552 13874 6604 13880
rect 6276 13796 6328 13802
rect 6276 13738 6328 13744
rect 5736 13110 5948 13138
rect 5736 12442 5764 13110
rect 5908 12640 5960 12646
rect 5908 12582 5960 12588
rect 5724 12436 5776 12442
rect 5724 12378 5776 12384
rect 5816 12232 5868 12238
rect 5816 12174 5868 12180
rect 5448 12164 5500 12170
rect 5448 12106 5500 12112
rect 5540 12164 5592 12170
rect 5540 12106 5592 12112
rect 5356 11892 5408 11898
rect 5356 11834 5408 11840
rect 4620 11824 4672 11830
rect 4620 11766 4672 11772
rect 3608 11688 3660 11694
rect 3608 11630 3660 11636
rect 3620 11354 3648 11630
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 3608 11348 3660 11354
rect 3608 11290 3660 11296
rect 4632 10713 4660 11766
rect 5172 11552 5224 11558
rect 5172 11494 5224 11500
rect 5184 11150 5212 11494
rect 5460 11354 5488 12106
rect 5448 11348 5500 11354
rect 5448 11290 5500 11296
rect 5172 11144 5224 11150
rect 5172 11086 5224 11092
rect 4804 11008 4856 11014
rect 4804 10950 4856 10956
rect 4816 10810 4844 10950
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 5552 10826 5580 12106
rect 5828 11694 5856 12174
rect 5920 12102 5948 12582
rect 6184 12232 6236 12238
rect 6184 12174 6236 12180
rect 5908 12096 5960 12102
rect 5908 12038 5960 12044
rect 6000 12096 6052 12102
rect 6000 12038 6052 12044
rect 5816 11688 5868 11694
rect 5816 11630 5868 11636
rect 5724 11552 5776 11558
rect 5724 11494 5776 11500
rect 5736 11218 5764 11494
rect 5828 11218 5856 11630
rect 5724 11212 5776 11218
rect 5724 11154 5776 11160
rect 5816 11212 5868 11218
rect 5816 11154 5868 11160
rect 4804 10804 4856 10810
rect 4804 10746 4856 10752
rect 5552 10798 5764 10826
rect 4618 10704 4674 10713
rect 4618 10639 4674 10648
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4632 8566 4660 10639
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 5264 8832 5316 8838
rect 5264 8774 5316 8780
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 5276 8634 5304 8774
rect 5264 8628 5316 8634
rect 5264 8570 5316 8576
rect 3240 8560 3292 8566
rect 3240 8502 3292 8508
rect 4620 8560 4672 8566
rect 4620 8502 4672 8508
rect 3252 7342 3280 8502
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4632 7410 4660 8502
rect 5356 8424 5408 8430
rect 5356 8366 5408 8372
rect 5448 8424 5500 8430
rect 5448 8366 5500 8372
rect 5368 8090 5396 8366
rect 5356 8084 5408 8090
rect 5356 8026 5408 8032
rect 5460 7834 5488 8366
rect 5368 7806 5488 7834
rect 5552 7818 5580 10798
rect 5736 10674 5764 10798
rect 5920 10674 5948 12038
rect 5632 10668 5684 10674
rect 5632 10610 5684 10616
rect 5724 10668 5776 10674
rect 5724 10610 5776 10616
rect 5908 10668 5960 10674
rect 5908 10610 5960 10616
rect 5644 8974 5672 10610
rect 6012 10062 6040 12038
rect 6092 11756 6144 11762
rect 6092 11698 6144 11704
rect 6104 10674 6132 11698
rect 6196 11150 6224 12174
rect 6368 11756 6420 11762
rect 6368 11698 6420 11704
rect 6552 11756 6604 11762
rect 6552 11698 6604 11704
rect 6276 11688 6328 11694
rect 6276 11630 6328 11636
rect 6288 11150 6316 11630
rect 6184 11144 6236 11150
rect 6184 11086 6236 11092
rect 6276 11144 6328 11150
rect 6276 11086 6328 11092
rect 6092 10668 6144 10674
rect 6092 10610 6144 10616
rect 6104 10266 6132 10610
rect 6092 10260 6144 10266
rect 6092 10202 6144 10208
rect 6288 10130 6316 11086
rect 6380 10538 6408 11698
rect 6564 11150 6592 11698
rect 6656 11286 6684 14418
rect 6920 14408 6972 14414
rect 6920 14350 6972 14356
rect 6828 14272 6880 14278
rect 6828 14214 6880 14220
rect 6840 13938 6868 14214
rect 6828 13932 6880 13938
rect 6828 13874 6880 13880
rect 6932 13870 6960 14350
rect 7024 14006 7052 14554
rect 7484 14482 7512 15098
rect 7748 15020 7800 15026
rect 7748 14962 7800 14968
rect 7656 14952 7708 14958
rect 7656 14894 7708 14900
rect 7472 14476 7524 14482
rect 7472 14418 7524 14424
rect 7668 14414 7696 14894
rect 7760 14414 7788 14962
rect 7944 14822 7972 15982
rect 8036 15026 8064 15982
rect 8496 15978 8524 17138
rect 8680 16794 8708 17734
rect 8760 17332 8812 17338
rect 8760 17274 8812 17280
rect 8772 17066 8800 17274
rect 8760 17060 8812 17066
rect 8760 17002 8812 17008
rect 8668 16788 8720 16794
rect 8668 16730 8720 16736
rect 8576 16040 8628 16046
rect 8576 15982 8628 15988
rect 8484 15972 8536 15978
rect 8484 15914 8536 15920
rect 8300 15904 8352 15910
rect 8588 15858 8616 15982
rect 8300 15846 8352 15852
rect 8024 15020 8076 15026
rect 8024 14962 8076 14968
rect 8116 14884 8168 14890
rect 8116 14826 8168 14832
rect 7932 14816 7984 14822
rect 7932 14758 7984 14764
rect 7944 14414 7972 14758
rect 8128 14414 8156 14826
rect 8312 14618 8340 15846
rect 8496 15830 8616 15858
rect 8496 15570 8524 15830
rect 8484 15564 8536 15570
rect 8484 15506 8536 15512
rect 8392 15020 8444 15026
rect 8392 14962 8444 14968
rect 8404 14618 8432 14962
rect 8300 14612 8352 14618
rect 8300 14554 8352 14560
rect 8392 14612 8444 14618
rect 8392 14554 8444 14560
rect 8208 14544 8260 14550
rect 8208 14486 8260 14492
rect 8220 14414 8248 14486
rect 8300 14476 8352 14482
rect 8300 14418 8352 14424
rect 7656 14408 7708 14414
rect 7656 14350 7708 14356
rect 7748 14408 7800 14414
rect 7748 14350 7800 14356
rect 7932 14408 7984 14414
rect 7932 14350 7984 14356
rect 8116 14408 8168 14414
rect 8116 14350 8168 14356
rect 8208 14408 8260 14414
rect 8208 14350 8260 14356
rect 7012 14000 7064 14006
rect 7012 13942 7064 13948
rect 6920 13864 6972 13870
rect 6920 13806 6972 13812
rect 6828 13796 6880 13802
rect 6828 13738 6880 13744
rect 6840 13530 6868 13738
rect 6828 13524 6880 13530
rect 6828 13466 6880 13472
rect 6932 12434 6960 13806
rect 6932 12406 7052 12434
rect 6920 11824 6972 11830
rect 6920 11766 6972 11772
rect 6644 11280 6696 11286
rect 6644 11222 6696 11228
rect 6932 11218 6960 11766
rect 7024 11694 7052 12406
rect 7012 11688 7064 11694
rect 7012 11630 7064 11636
rect 7104 11552 7156 11558
rect 7104 11494 7156 11500
rect 6736 11212 6788 11218
rect 6736 11154 6788 11160
rect 6920 11212 6972 11218
rect 6920 11154 6972 11160
rect 6552 11144 6604 11150
rect 6552 11086 6604 11092
rect 6460 11076 6512 11082
rect 6460 11018 6512 11024
rect 6472 10674 6500 11018
rect 6552 10804 6604 10810
rect 6552 10746 6604 10752
rect 6460 10668 6512 10674
rect 6460 10610 6512 10616
rect 6564 10538 6592 10746
rect 6368 10532 6420 10538
rect 6368 10474 6420 10480
rect 6552 10532 6604 10538
rect 6552 10474 6604 10480
rect 6276 10124 6328 10130
rect 6276 10066 6328 10072
rect 6000 10056 6052 10062
rect 6000 9998 6052 10004
rect 6380 9722 6408 10474
rect 6748 10062 6776 11154
rect 7012 11076 7064 11082
rect 7012 11018 7064 11024
rect 7024 10742 7052 11018
rect 7012 10736 7064 10742
rect 7012 10678 7064 10684
rect 7116 10554 7144 11494
rect 6932 10526 7144 10554
rect 7196 10532 7248 10538
rect 6932 10062 6960 10526
rect 7196 10474 7248 10480
rect 7208 10062 7236 10474
rect 7668 10198 7696 14350
rect 7760 14006 7788 14350
rect 8312 14278 8340 14418
rect 8300 14272 8352 14278
rect 8300 14214 8352 14220
rect 7748 14000 7800 14006
rect 7748 13942 7800 13948
rect 8404 13938 8432 14554
rect 8496 14414 8524 15506
rect 8574 14512 8630 14521
rect 8574 14447 8630 14456
rect 8588 14414 8616 14447
rect 8484 14408 8536 14414
rect 8484 14350 8536 14356
rect 8576 14408 8628 14414
rect 8576 14350 8628 14356
rect 8680 14346 8708 16730
rect 8864 16522 8892 18158
rect 9128 17672 9180 17678
rect 9128 17614 9180 17620
rect 9036 16584 9088 16590
rect 9036 16526 9088 16532
rect 8852 16516 8904 16522
rect 8852 16458 8904 16464
rect 8864 16114 8892 16458
rect 8944 16448 8996 16454
rect 8944 16390 8996 16396
rect 8956 16250 8984 16390
rect 8944 16244 8996 16250
rect 8944 16186 8996 16192
rect 8852 16108 8904 16114
rect 8852 16050 8904 16056
rect 8944 16108 8996 16114
rect 9048 16096 9076 16526
rect 9140 16114 9168 17614
rect 9232 17338 9260 18158
rect 9324 17746 9352 19110
rect 9692 17814 9720 22578
rect 10968 22024 11020 22030
rect 10968 21966 11020 21972
rect 11428 22024 11480 22030
rect 11428 21966 11480 21972
rect 9864 21480 9916 21486
rect 9864 21422 9916 21428
rect 9772 20800 9824 20806
rect 9772 20742 9824 20748
rect 9784 20466 9812 20742
rect 9876 20602 9904 21422
rect 10980 21418 11008 21966
rect 10968 21412 11020 21418
rect 10968 21354 11020 21360
rect 9956 20868 10008 20874
rect 9956 20810 10008 20816
rect 9864 20596 9916 20602
rect 9864 20538 9916 20544
rect 9772 20460 9824 20466
rect 9772 20402 9824 20408
rect 9864 18760 9916 18766
rect 9968 18748 9996 20810
rect 10980 20534 11008 21354
rect 11440 21146 11468 21966
rect 11428 21140 11480 21146
rect 11428 21082 11480 21088
rect 11152 20936 11204 20942
rect 11152 20878 11204 20884
rect 10968 20528 11020 20534
rect 10968 20470 11020 20476
rect 10692 20460 10744 20466
rect 10692 20402 10744 20408
rect 9916 18720 9996 18748
rect 9864 18702 9916 18708
rect 9772 18080 9824 18086
rect 9772 18022 9824 18028
rect 9680 17808 9732 17814
rect 9680 17750 9732 17756
rect 9312 17740 9364 17746
rect 9312 17682 9364 17688
rect 9220 17332 9272 17338
rect 9220 17274 9272 17280
rect 9784 17202 9812 18022
rect 9876 17882 9904 18702
rect 10704 18222 10732 20402
rect 10968 18828 11020 18834
rect 10968 18770 11020 18776
rect 10980 18290 11008 18770
rect 11164 18766 11192 20878
rect 11244 19916 11296 19922
rect 11244 19858 11296 19864
rect 11256 19514 11284 19858
rect 11244 19508 11296 19514
rect 11244 19450 11296 19456
rect 11532 19446 11560 23530
rect 11716 21622 11744 24074
rect 11992 23662 12020 25434
rect 12992 25424 13044 25430
rect 12992 25366 13044 25372
rect 12624 25220 12676 25226
rect 12624 25162 12676 25168
rect 12532 25152 12584 25158
rect 12532 25094 12584 25100
rect 12544 24750 12572 25094
rect 12532 24744 12584 24750
rect 12532 24686 12584 24692
rect 12636 24177 12664 25162
rect 13004 24732 13032 25366
rect 13820 25288 13872 25294
rect 13820 25230 13872 25236
rect 14372 25288 14424 25294
rect 14372 25230 14424 25236
rect 15200 25288 15252 25294
rect 15200 25230 15252 25236
rect 13636 25220 13688 25226
rect 13636 25162 13688 25168
rect 13360 24880 13412 24886
rect 13360 24822 13412 24828
rect 13084 24744 13136 24750
rect 13004 24704 13084 24732
rect 12808 24608 12860 24614
rect 12808 24550 12860 24556
rect 12820 24342 12848 24550
rect 12808 24336 12860 24342
rect 12808 24278 12860 24284
rect 12622 24168 12678 24177
rect 12622 24103 12678 24112
rect 12164 23724 12216 23730
rect 12164 23666 12216 23672
rect 11980 23656 12032 23662
rect 11980 23598 12032 23604
rect 12176 23594 12204 23666
rect 12164 23588 12216 23594
rect 12164 23530 12216 23536
rect 12072 22432 12124 22438
rect 12072 22374 12124 22380
rect 12084 22030 12112 22374
rect 12072 22024 12124 22030
rect 12070 21992 12072 22001
rect 12124 21992 12126 22001
rect 12070 21927 12126 21936
rect 12440 21956 12492 21962
rect 12440 21898 12492 21904
rect 11796 21888 11848 21894
rect 11796 21830 11848 21836
rect 11888 21888 11940 21894
rect 11888 21830 11940 21836
rect 11808 21622 11836 21830
rect 11704 21616 11756 21622
rect 11704 21558 11756 21564
rect 11796 21616 11848 21622
rect 11796 21558 11848 21564
rect 11900 20942 11928 21830
rect 12452 21146 12480 21898
rect 12716 21888 12768 21894
rect 12716 21830 12768 21836
rect 12440 21140 12492 21146
rect 12440 21082 12492 21088
rect 12728 20942 12756 21830
rect 11888 20936 11940 20942
rect 11888 20878 11940 20884
rect 12716 20936 12768 20942
rect 12716 20878 12768 20884
rect 12716 20800 12768 20806
rect 12716 20742 12768 20748
rect 11612 20324 11664 20330
rect 11612 20266 11664 20272
rect 11520 19440 11572 19446
rect 11520 19382 11572 19388
rect 11336 19372 11388 19378
rect 11336 19314 11388 19320
rect 11428 19372 11480 19378
rect 11428 19314 11480 19320
rect 11348 18970 11376 19314
rect 11336 18964 11388 18970
rect 11336 18906 11388 18912
rect 11440 18902 11468 19314
rect 11428 18896 11480 18902
rect 11428 18838 11480 18844
rect 11624 18766 11652 20266
rect 12624 20052 12676 20058
rect 12624 19994 12676 20000
rect 12636 19854 12664 19994
rect 11704 19848 11756 19854
rect 11704 19790 11756 19796
rect 12624 19848 12676 19854
rect 12624 19790 12676 19796
rect 11716 19514 11744 19790
rect 12532 19780 12584 19786
rect 12532 19722 12584 19728
rect 12544 19514 12572 19722
rect 11704 19508 11756 19514
rect 11704 19450 11756 19456
rect 12532 19508 12584 19514
rect 12532 19450 12584 19456
rect 12728 19446 12756 20742
rect 12716 19440 12768 19446
rect 12716 19382 12768 19388
rect 11980 18828 12032 18834
rect 11980 18770 12032 18776
rect 11152 18760 11204 18766
rect 11612 18760 11664 18766
rect 11204 18720 11284 18748
rect 11152 18702 11204 18708
rect 10876 18284 10928 18290
rect 10876 18226 10928 18232
rect 10968 18284 11020 18290
rect 10968 18226 11020 18232
rect 10692 18216 10744 18222
rect 10692 18158 10744 18164
rect 10600 18080 10652 18086
rect 10600 18022 10652 18028
rect 9864 17876 9916 17882
rect 9864 17818 9916 17824
rect 10612 17746 10640 18022
rect 10600 17740 10652 17746
rect 10600 17682 10652 17688
rect 10704 17626 10732 18158
rect 10888 17678 10916 18226
rect 11256 17678 11284 18720
rect 11612 18702 11664 18708
rect 11704 18760 11756 18766
rect 11704 18702 11756 18708
rect 11428 18624 11480 18630
rect 11428 18566 11480 18572
rect 11336 18352 11388 18358
rect 11336 18294 11388 18300
rect 10140 17604 10192 17610
rect 10140 17546 10192 17552
rect 10612 17598 10732 17626
rect 10876 17672 10928 17678
rect 10876 17614 10928 17620
rect 11244 17672 11296 17678
rect 11244 17614 11296 17620
rect 10048 17536 10100 17542
rect 10048 17478 10100 17484
rect 10060 17270 10088 17478
rect 10152 17338 10180 17546
rect 10232 17536 10284 17542
rect 10232 17478 10284 17484
rect 10140 17332 10192 17338
rect 10140 17274 10192 17280
rect 10048 17264 10100 17270
rect 10048 17206 10100 17212
rect 9312 17196 9364 17202
rect 9312 17138 9364 17144
rect 9496 17196 9548 17202
rect 9496 17138 9548 17144
rect 9772 17196 9824 17202
rect 9772 17138 9824 17144
rect 9324 16794 9352 17138
rect 9312 16788 9364 16794
rect 9312 16730 9364 16736
rect 9508 16250 9536 17138
rect 9588 16992 9640 16998
rect 9588 16934 9640 16940
rect 9600 16590 9628 16934
rect 10152 16658 10180 17274
rect 10244 17202 10272 17478
rect 10232 17196 10284 17202
rect 10232 17138 10284 17144
rect 10612 17066 10640 17598
rect 10600 17060 10652 17066
rect 10600 17002 10652 17008
rect 10140 16652 10192 16658
rect 10140 16594 10192 16600
rect 9588 16584 9640 16590
rect 9588 16526 9640 16532
rect 9220 16244 9272 16250
rect 9220 16186 9272 16192
rect 9496 16244 9548 16250
rect 9496 16186 9548 16192
rect 9232 16114 9260 16186
rect 8996 16068 9076 16096
rect 8944 16050 8996 16056
rect 8864 15910 8892 16050
rect 8852 15904 8904 15910
rect 8852 15846 8904 15852
rect 9048 15348 9076 16068
rect 9128 16108 9180 16114
rect 9128 16050 9180 16056
rect 9220 16108 9272 16114
rect 9772 16108 9824 16114
rect 9220 16050 9272 16056
rect 9692 16068 9772 16096
rect 9140 15706 9168 16050
rect 9128 15700 9180 15706
rect 9128 15642 9180 15648
rect 9232 15502 9260 16050
rect 9588 16040 9640 16046
rect 9588 15982 9640 15988
rect 9404 15904 9456 15910
rect 9404 15846 9456 15852
rect 9220 15496 9272 15502
rect 9220 15438 9272 15444
rect 9048 15320 9352 15348
rect 9048 15162 9076 15320
rect 9036 15156 9088 15162
rect 9036 15098 9088 15104
rect 9126 15056 9182 15065
rect 9126 14991 9128 15000
rect 9180 14991 9182 15000
rect 9128 14962 9180 14968
rect 9220 14952 9272 14958
rect 9218 14920 9220 14929
rect 9272 14920 9274 14929
rect 9218 14855 9274 14864
rect 9324 14414 9352 15320
rect 9312 14408 9364 14414
rect 9312 14350 9364 14356
rect 9416 14346 9444 15846
rect 9600 15162 9628 15982
rect 9692 15434 9720 16068
rect 9772 16050 9824 16056
rect 9864 16040 9916 16046
rect 9864 15982 9916 15988
rect 9772 15496 9824 15502
rect 9772 15438 9824 15444
rect 9680 15428 9732 15434
rect 9680 15370 9732 15376
rect 9588 15156 9640 15162
rect 9588 15098 9640 15104
rect 9496 15088 9548 15094
rect 9496 15030 9548 15036
rect 9586 15056 9642 15065
rect 9508 14482 9536 15030
rect 9692 15026 9720 15370
rect 9784 15026 9812 15438
rect 9586 14991 9588 15000
rect 9640 14991 9642 15000
rect 9680 15020 9732 15026
rect 9588 14962 9640 14968
rect 9680 14962 9732 14968
rect 9772 15020 9824 15026
rect 9772 14962 9824 14968
rect 9784 14618 9812 14962
rect 9876 14822 9904 15982
rect 10048 15564 10100 15570
rect 10048 15506 10100 15512
rect 10060 15042 10088 15506
rect 10416 15496 10468 15502
rect 10416 15438 10468 15444
rect 9968 15026 10088 15042
rect 9968 15020 10100 15026
rect 9968 15014 10048 15020
rect 9864 14816 9916 14822
rect 9864 14758 9916 14764
rect 9772 14612 9824 14618
rect 9772 14554 9824 14560
rect 9876 14482 9904 14758
rect 9496 14476 9548 14482
rect 9496 14418 9548 14424
rect 9864 14476 9916 14482
rect 9864 14418 9916 14424
rect 9968 14414 9996 15014
rect 10048 14962 10100 14968
rect 10046 14920 10102 14929
rect 10046 14855 10102 14864
rect 10324 14884 10376 14890
rect 10060 14822 10088 14855
rect 10324 14826 10376 14832
rect 10048 14816 10100 14822
rect 10048 14758 10100 14764
rect 10060 14414 10088 14758
rect 10336 14414 10364 14826
rect 10428 14822 10456 15438
rect 10416 14816 10468 14822
rect 10416 14758 10468 14764
rect 9956 14408 10008 14414
rect 9956 14350 10008 14356
rect 10048 14408 10100 14414
rect 10048 14350 10100 14356
rect 10324 14408 10376 14414
rect 10324 14350 10376 14356
rect 8668 14340 8720 14346
rect 8668 14282 8720 14288
rect 9404 14340 9456 14346
rect 9404 14282 9456 14288
rect 8760 14272 8812 14278
rect 8760 14214 8812 14220
rect 8772 14006 8800 14214
rect 8760 14000 8812 14006
rect 8944 14000 8996 14006
rect 8760 13942 8812 13948
rect 8864 13960 8944 13988
rect 8392 13932 8444 13938
rect 8392 13874 8444 13880
rect 8300 13864 8352 13870
rect 8300 13806 8352 13812
rect 8312 12434 8340 13806
rect 8220 12406 8340 12434
rect 7748 11892 7800 11898
rect 7748 11834 7800 11840
rect 7760 11082 7788 11834
rect 8220 11830 8248 12406
rect 8208 11824 8260 11830
rect 8208 11766 8260 11772
rect 8024 11756 8076 11762
rect 8024 11698 8076 11704
rect 7840 11688 7892 11694
rect 7840 11630 7892 11636
rect 7852 11150 7880 11630
rect 8036 11354 8064 11698
rect 8024 11348 8076 11354
rect 8024 11290 8076 11296
rect 7840 11144 7892 11150
rect 7840 11086 7892 11092
rect 7748 11076 7800 11082
rect 7748 11018 7800 11024
rect 8220 10742 8248 11766
rect 8300 11552 8352 11558
rect 8300 11494 8352 11500
rect 8312 10742 8340 11494
rect 8208 10736 8260 10742
rect 8208 10678 8260 10684
rect 8300 10736 8352 10742
rect 8760 10736 8812 10742
rect 8300 10678 8352 10684
rect 8758 10704 8760 10713
rect 8864 10724 8892 13960
rect 9968 13988 9996 14350
rect 10140 14000 10192 14006
rect 9968 13960 10140 13988
rect 8944 13942 8996 13948
rect 10140 13942 10192 13948
rect 10324 12232 10376 12238
rect 10324 12174 10376 12180
rect 9220 12096 9272 12102
rect 9220 12038 9272 12044
rect 8944 11552 8996 11558
rect 8944 11494 8996 11500
rect 8956 11218 8984 11494
rect 9232 11218 9260 12038
rect 9864 11688 9916 11694
rect 9864 11630 9916 11636
rect 9876 11393 9904 11630
rect 9862 11384 9918 11393
rect 9862 11319 9918 11328
rect 8944 11212 8996 11218
rect 8944 11154 8996 11160
rect 9220 11212 9272 11218
rect 9220 11154 9272 11160
rect 8812 10704 8892 10724
rect 8814 10696 8892 10704
rect 8758 10639 8814 10648
rect 10336 10606 10364 12174
rect 10416 11688 10468 11694
rect 10416 11630 10468 11636
rect 10324 10600 10376 10606
rect 10324 10542 10376 10548
rect 8760 10464 8812 10470
rect 8760 10406 8812 10412
rect 9956 10464 10008 10470
rect 9956 10406 10008 10412
rect 7656 10192 7708 10198
rect 7656 10134 7708 10140
rect 7288 10124 7340 10130
rect 7288 10066 7340 10072
rect 6644 10056 6696 10062
rect 6644 9998 6696 10004
rect 6736 10056 6788 10062
rect 6736 9998 6788 10004
rect 6920 10056 6972 10062
rect 6920 9998 6972 10004
rect 7196 10056 7248 10062
rect 7196 9998 7248 10004
rect 6368 9716 6420 9722
rect 6368 9658 6420 9664
rect 6656 9654 6684 9998
rect 6828 9988 6880 9994
rect 6828 9930 6880 9936
rect 6644 9648 6696 9654
rect 6644 9590 6696 9596
rect 6656 9178 6684 9590
rect 6644 9172 6696 9178
rect 6644 9114 6696 9120
rect 6460 9104 6512 9110
rect 6460 9046 6512 9052
rect 6472 8974 6500 9046
rect 5632 8968 5684 8974
rect 5632 8910 5684 8916
rect 6460 8968 6512 8974
rect 6460 8910 6512 8916
rect 5644 8566 5672 8910
rect 6368 8832 6420 8838
rect 6368 8774 6420 8780
rect 5632 8560 5684 8566
rect 5632 8502 5684 8508
rect 5908 8424 5960 8430
rect 5908 8366 5960 8372
rect 5724 8288 5776 8294
rect 5724 8230 5776 8236
rect 5736 8022 5764 8230
rect 5724 8016 5776 8022
rect 5724 7958 5776 7964
rect 5540 7812 5592 7818
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 4620 7404 4672 7410
rect 4620 7346 4672 7352
rect 5264 7404 5316 7410
rect 5264 7346 5316 7352
rect 3240 7336 3292 7342
rect 3292 7296 3372 7324
rect 3240 7278 3292 7284
rect 3344 5166 3372 7296
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 5276 5302 5304 7346
rect 5368 7342 5396 7806
rect 5540 7754 5592 7760
rect 5448 7744 5500 7750
rect 5448 7686 5500 7692
rect 5460 7546 5488 7686
rect 5448 7540 5500 7546
rect 5448 7482 5500 7488
rect 5356 7336 5408 7342
rect 5356 7278 5408 7284
rect 5264 5296 5316 5302
rect 5264 5238 5316 5244
rect 3332 5160 3384 5166
rect 3332 5102 3384 5108
rect 3608 5160 3660 5166
rect 3608 5102 3660 5108
rect 3344 3602 3372 5102
rect 3620 4826 3648 5102
rect 4988 5092 5040 5098
rect 4988 5034 5040 5040
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 3608 4820 3660 4826
rect 3608 4762 3660 4768
rect 5000 4622 5028 5034
rect 4988 4616 5040 4622
rect 4988 4558 5040 4564
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 3332 3596 3384 3602
rect 3332 3538 3384 3544
rect 5276 3398 5304 5238
rect 5368 4826 5396 7278
rect 5736 5234 5764 7958
rect 5920 7886 5948 8366
rect 6380 7886 6408 8774
rect 6472 8566 6500 8910
rect 6460 8560 6512 8566
rect 6460 8502 6512 8508
rect 6550 8528 6606 8537
rect 6840 8498 6868 9930
rect 7208 9654 7236 9998
rect 7196 9648 7248 9654
rect 7196 9590 7248 9596
rect 6920 9580 6972 9586
rect 6920 9522 6972 9528
rect 7104 9580 7156 9586
rect 7104 9522 7156 9528
rect 6932 8498 6960 9522
rect 7012 9444 7064 9450
rect 7012 9386 7064 9392
rect 7024 9042 7052 9386
rect 7012 9036 7064 9042
rect 7012 8978 7064 8984
rect 7012 8900 7064 8906
rect 7012 8842 7064 8848
rect 7024 8634 7052 8842
rect 7012 8628 7064 8634
rect 7012 8570 7064 8576
rect 6550 8463 6552 8472
rect 6604 8463 6606 8472
rect 6828 8492 6880 8498
rect 6552 8434 6604 8440
rect 6828 8434 6880 8440
rect 6920 8492 6972 8498
rect 6920 8434 6972 8440
rect 7012 8492 7064 8498
rect 7116 8480 7144 9522
rect 7196 9512 7248 9518
rect 7196 9454 7248 9460
rect 7208 8838 7236 9454
rect 7300 9382 7328 10066
rect 8772 10062 8800 10406
rect 9968 10130 9996 10406
rect 9956 10124 10008 10130
rect 9956 10066 10008 10072
rect 7840 10056 7892 10062
rect 7840 9998 7892 10004
rect 8760 10056 8812 10062
rect 8760 9998 8812 10004
rect 7852 9722 7880 9998
rect 7840 9716 7892 9722
rect 7840 9658 7892 9664
rect 7288 9376 7340 9382
rect 7288 9318 7340 9324
rect 7288 9172 7340 9178
rect 7288 9114 7340 9120
rect 7196 8832 7248 8838
rect 7196 8774 7248 8780
rect 7300 8537 7328 9114
rect 8300 8900 8352 8906
rect 8300 8842 8352 8848
rect 7380 8628 7432 8634
rect 7380 8570 7432 8576
rect 7064 8452 7144 8480
rect 7286 8528 7342 8537
rect 7286 8463 7288 8472
rect 7012 8434 7064 8440
rect 6840 8401 6868 8434
rect 6826 8392 6882 8401
rect 6826 8327 6882 8336
rect 6460 7948 6512 7954
rect 6460 7890 6512 7896
rect 5908 7880 5960 7886
rect 5908 7822 5960 7828
rect 6368 7880 6420 7886
rect 6368 7822 6420 7828
rect 5920 7478 5948 7822
rect 6472 7546 6500 7890
rect 6644 7744 6696 7750
rect 6644 7686 6696 7692
rect 6460 7540 6512 7546
rect 6460 7482 6512 7488
rect 5908 7472 5960 7478
rect 5908 7414 5960 7420
rect 6656 7410 6684 7686
rect 6932 7478 6960 8434
rect 7116 8090 7144 8452
rect 7340 8463 7342 8472
rect 7288 8434 7340 8440
rect 7194 8392 7250 8401
rect 7194 8327 7250 8336
rect 7104 8084 7156 8090
rect 7104 8026 7156 8032
rect 7116 7886 7144 8026
rect 7208 7954 7236 8327
rect 7288 8288 7340 8294
rect 7288 8230 7340 8236
rect 7196 7948 7248 7954
rect 7196 7890 7248 7896
rect 7300 7886 7328 8230
rect 7104 7880 7156 7886
rect 7104 7822 7156 7828
rect 7288 7880 7340 7886
rect 7288 7822 7340 7828
rect 7392 7818 7420 8570
rect 8312 8498 8340 8842
rect 8392 8628 8444 8634
rect 8392 8570 8444 8576
rect 8300 8492 8352 8498
rect 8300 8434 8352 8440
rect 7654 8392 7710 8401
rect 7654 8327 7710 8336
rect 7196 7812 7248 7818
rect 7196 7754 7248 7760
rect 7380 7812 7432 7818
rect 7380 7754 7432 7760
rect 6920 7472 6972 7478
rect 6920 7414 6972 7420
rect 6644 7404 6696 7410
rect 6644 7346 6696 7352
rect 7208 7342 7236 7754
rect 7392 7410 7420 7754
rect 7380 7404 7432 7410
rect 7380 7346 7432 7352
rect 6460 7336 6512 7342
rect 6460 7278 6512 7284
rect 7196 7336 7248 7342
rect 7196 7278 7248 7284
rect 6472 5710 6500 7278
rect 6920 5840 6972 5846
rect 6920 5782 6972 5788
rect 6460 5704 6512 5710
rect 6460 5646 6512 5652
rect 5724 5228 5776 5234
rect 5724 5170 5776 5176
rect 6184 5228 6236 5234
rect 6184 5170 6236 5176
rect 5908 5160 5960 5166
rect 5908 5102 5960 5108
rect 5540 5024 5592 5030
rect 5540 4966 5592 4972
rect 5356 4820 5408 4826
rect 5356 4762 5408 4768
rect 5368 4214 5396 4762
rect 5448 4616 5500 4622
rect 5552 4604 5580 4966
rect 5920 4826 5948 5102
rect 6196 4826 6224 5170
rect 6472 5166 6500 5646
rect 6644 5568 6696 5574
rect 6932 5545 6960 5782
rect 6644 5510 6696 5516
rect 6918 5536 6974 5545
rect 6656 5370 6684 5510
rect 6918 5471 6974 5480
rect 6644 5364 6696 5370
rect 6644 5306 6696 5312
rect 6736 5364 6788 5370
rect 6736 5306 6788 5312
rect 6552 5296 6604 5302
rect 6748 5250 6776 5306
rect 6604 5244 6776 5250
rect 6552 5238 6776 5244
rect 6564 5222 6776 5238
rect 6932 5234 6960 5471
rect 6276 5160 6328 5166
rect 6276 5102 6328 5108
rect 6460 5160 6512 5166
rect 6460 5102 6512 5108
rect 5908 4820 5960 4826
rect 5908 4762 5960 4768
rect 6184 4820 6236 4826
rect 6184 4762 6236 4768
rect 6090 4720 6146 4729
rect 6090 4655 6092 4664
rect 6144 4655 6146 4664
rect 6092 4626 6144 4632
rect 5500 4576 5580 4604
rect 5448 4558 5500 4564
rect 5816 4548 5868 4554
rect 5816 4490 5868 4496
rect 5356 4208 5408 4214
rect 5356 4150 5408 4156
rect 5828 4078 5856 4490
rect 6196 4282 6224 4762
rect 6288 4282 6316 5102
rect 6472 5030 6500 5102
rect 6552 5092 6604 5098
rect 6552 5034 6604 5040
rect 6460 5024 6512 5030
rect 6460 4966 6512 4972
rect 6564 4826 6592 5034
rect 6552 4820 6604 4826
rect 6552 4762 6604 4768
rect 6460 4752 6512 4758
rect 6460 4694 6512 4700
rect 6472 4622 6500 4694
rect 6460 4616 6512 4622
rect 6460 4558 6512 4564
rect 6184 4276 6236 4282
rect 6184 4218 6236 4224
rect 6276 4276 6328 4282
rect 6276 4218 6328 4224
rect 6472 4146 6500 4558
rect 6748 4214 6776 5222
rect 6920 5228 6972 5234
rect 7104 5228 7156 5234
rect 6920 5170 6972 5176
rect 7024 5188 7104 5216
rect 7024 4826 7052 5188
rect 7104 5170 7156 5176
rect 7208 5114 7236 7278
rect 7472 5568 7524 5574
rect 7472 5510 7524 5516
rect 7484 5302 7512 5510
rect 7472 5296 7524 5302
rect 7472 5238 7524 5244
rect 7484 5166 7512 5238
rect 7564 5228 7616 5234
rect 7564 5170 7616 5176
rect 7116 5086 7236 5114
rect 7472 5160 7524 5166
rect 7472 5102 7524 5108
rect 7012 4820 7064 4826
rect 7012 4762 7064 4768
rect 7024 4622 7052 4762
rect 7116 4729 7144 5086
rect 7484 4758 7512 5102
rect 7576 4758 7604 5170
rect 7668 5030 7696 8327
rect 8404 8022 8432 8570
rect 8772 8430 8800 9998
rect 9956 9920 10008 9926
rect 9956 9862 10008 9868
rect 9864 9376 9916 9382
rect 9864 9318 9916 9324
rect 9876 8974 9904 9318
rect 9968 8974 9996 9862
rect 10428 9674 10456 11630
rect 10336 9646 10456 9674
rect 10060 9042 10180 9058
rect 10048 9036 10180 9042
rect 10100 9030 10180 9036
rect 10048 8978 10100 8984
rect 9404 8968 9456 8974
rect 9404 8910 9456 8916
rect 9864 8968 9916 8974
rect 9864 8910 9916 8916
rect 9956 8968 10008 8974
rect 9956 8910 10008 8916
rect 9312 8832 9364 8838
rect 9312 8774 9364 8780
rect 9324 8566 9352 8774
rect 9312 8560 9364 8566
rect 9312 8502 9364 8508
rect 9416 8430 9444 8910
rect 9680 8900 9732 8906
rect 9680 8842 9732 8848
rect 8760 8424 8812 8430
rect 8760 8366 8812 8372
rect 9404 8424 9456 8430
rect 9404 8366 9456 8372
rect 8392 8016 8444 8022
rect 8392 7958 8444 7964
rect 8772 7342 8800 8366
rect 9496 8288 9548 8294
rect 9496 8230 9548 8236
rect 9312 7880 9364 7886
rect 9312 7822 9364 7828
rect 9324 7546 9352 7822
rect 9312 7540 9364 7546
rect 9312 7482 9364 7488
rect 8300 7336 8352 7342
rect 8300 7278 8352 7284
rect 8760 7336 8812 7342
rect 8760 7278 8812 7284
rect 9036 7336 9088 7342
rect 9036 7278 9088 7284
rect 8312 6882 8340 7278
rect 9048 7002 9076 7278
rect 9508 7206 9536 8230
rect 9692 7993 9720 8842
rect 9876 8294 9904 8910
rect 10152 8378 10180 9030
rect 10232 9036 10284 9042
rect 10232 8978 10284 8984
rect 9968 8350 10180 8378
rect 9864 8288 9916 8294
rect 9864 8230 9916 8236
rect 9968 8090 9996 8350
rect 9956 8084 10008 8090
rect 9956 8026 10008 8032
rect 9968 7993 9996 8026
rect 10140 8016 10192 8022
rect 9678 7984 9734 7993
rect 9678 7919 9734 7928
rect 9954 7984 10010 7993
rect 10140 7958 10192 7964
rect 9954 7919 10010 7928
rect 9588 7880 9640 7886
rect 9864 7880 9916 7886
rect 9640 7840 9812 7868
rect 9588 7822 9640 7828
rect 9784 7750 9812 7840
rect 9916 7857 9996 7868
rect 9916 7848 10010 7857
rect 9916 7840 9954 7848
rect 9864 7822 9916 7828
rect 9954 7783 10010 7792
rect 9588 7744 9640 7750
rect 9680 7744 9732 7750
rect 9588 7686 9640 7692
rect 9678 7712 9680 7721
rect 9772 7744 9824 7750
rect 9732 7712 9734 7721
rect 9600 7206 9628 7686
rect 9772 7686 9824 7692
rect 9678 7647 9734 7656
rect 9496 7200 9548 7206
rect 9496 7142 9548 7148
rect 9588 7200 9640 7206
rect 9588 7142 9640 7148
rect 9036 6996 9088 7002
rect 9036 6938 9088 6944
rect 8220 6854 8340 6882
rect 8024 5228 8076 5234
rect 8024 5170 8076 5176
rect 7932 5160 7984 5166
rect 7932 5102 7984 5108
rect 7748 5092 7800 5098
rect 7748 5034 7800 5040
rect 7656 5024 7708 5030
rect 7656 4966 7708 4972
rect 7472 4752 7524 4758
rect 7102 4720 7158 4729
rect 7472 4694 7524 4700
rect 7564 4752 7616 4758
rect 7564 4694 7616 4700
rect 7102 4655 7158 4664
rect 7012 4616 7064 4622
rect 7012 4558 7064 4564
rect 6736 4208 6788 4214
rect 6736 4150 6788 4156
rect 6000 4140 6052 4146
rect 6000 4082 6052 4088
rect 6460 4140 6512 4146
rect 6460 4082 6512 4088
rect 5816 4072 5868 4078
rect 5816 4014 5868 4020
rect 5828 3738 5856 4014
rect 5816 3732 5868 3738
rect 5816 3674 5868 3680
rect 5264 3392 5316 3398
rect 5264 3334 5316 3340
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 6012 3194 6040 4082
rect 6644 4072 6696 4078
rect 6644 4014 6696 4020
rect 6656 3602 6684 4014
rect 6920 3936 6972 3942
rect 6920 3878 6972 3884
rect 6644 3596 6696 3602
rect 6644 3538 6696 3544
rect 6000 3188 6052 3194
rect 6000 3130 6052 3136
rect 6656 3126 6684 3538
rect 6932 3534 6960 3878
rect 6920 3528 6972 3534
rect 6920 3470 6972 3476
rect 6644 3120 6696 3126
rect 6644 3062 6696 3068
rect 7024 2990 7052 4558
rect 7116 4146 7144 4655
rect 7760 4554 7788 5034
rect 7748 4548 7800 4554
rect 7748 4490 7800 4496
rect 7944 4486 7972 5102
rect 8036 4826 8064 5170
rect 8024 4820 8076 4826
rect 8024 4762 8076 4768
rect 7564 4480 7616 4486
rect 7564 4422 7616 4428
rect 7932 4480 7984 4486
rect 7932 4422 7984 4428
rect 7196 4208 7248 4214
rect 7196 4150 7248 4156
rect 7286 4176 7342 4185
rect 7104 4140 7156 4146
rect 7104 4082 7156 4088
rect 7208 3670 7236 4150
rect 7286 4111 7288 4120
rect 7340 4111 7342 4120
rect 7288 4082 7340 4088
rect 7576 4010 7604 4422
rect 7564 4004 7616 4010
rect 7564 3946 7616 3952
rect 7840 4004 7892 4010
rect 7840 3946 7892 3952
rect 7656 3936 7708 3942
rect 7656 3878 7708 3884
rect 7196 3664 7248 3670
rect 7196 3606 7248 3612
rect 7668 3534 7696 3878
rect 7852 3670 7880 3946
rect 7840 3664 7892 3670
rect 7840 3606 7892 3612
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 8220 3466 8248 6854
rect 9508 5386 9536 7142
rect 9508 5358 9628 5386
rect 9600 5302 9628 5358
rect 9220 5296 9272 5302
rect 9220 5238 9272 5244
rect 9588 5296 9640 5302
rect 9588 5238 9640 5244
rect 8484 5228 8536 5234
rect 8852 5228 8904 5234
rect 8536 5188 8616 5216
rect 8484 5170 8536 5176
rect 8482 4720 8538 4729
rect 8482 4655 8484 4664
rect 8536 4655 8538 4664
rect 8484 4626 8536 4632
rect 8300 4616 8352 4622
rect 8300 4558 8352 4564
rect 8392 4616 8444 4622
rect 8392 4558 8444 4564
rect 8312 4282 8340 4558
rect 8300 4276 8352 4282
rect 8300 4218 8352 4224
rect 8404 4214 8432 4558
rect 8392 4208 8444 4214
rect 8392 4150 8444 4156
rect 8588 4078 8616 5188
rect 8852 5170 8904 5176
rect 8668 4616 8720 4622
rect 8666 4584 8668 4593
rect 8760 4616 8812 4622
rect 8720 4584 8722 4593
rect 8760 4558 8812 4564
rect 8666 4519 8722 4528
rect 8772 4146 8800 4558
rect 8864 4214 8892 5170
rect 9232 5098 9260 5238
rect 9312 5228 9364 5234
rect 9312 5170 9364 5176
rect 9404 5228 9456 5234
rect 9404 5170 9456 5176
rect 9220 5092 9272 5098
rect 9220 5034 9272 5040
rect 9128 5024 9180 5030
rect 9128 4966 9180 4972
rect 9140 4282 9168 4966
rect 9232 4622 9260 5034
rect 9324 4826 9352 5170
rect 9416 4826 9444 5170
rect 9588 5160 9640 5166
rect 9588 5102 9640 5108
rect 9312 4820 9364 4826
rect 9312 4762 9364 4768
rect 9404 4820 9456 4826
rect 9404 4762 9456 4768
rect 9600 4758 9628 5102
rect 9588 4752 9640 4758
rect 9494 4720 9550 4729
rect 9588 4694 9640 4700
rect 9494 4655 9550 4664
rect 9508 4622 9536 4655
rect 9600 4622 9628 4694
rect 9864 4684 9916 4690
rect 9864 4626 9916 4632
rect 9220 4616 9272 4622
rect 9220 4558 9272 4564
rect 9496 4616 9548 4622
rect 9496 4558 9548 4564
rect 9588 4616 9640 4622
rect 9876 4593 9904 4626
rect 9588 4558 9640 4564
rect 9862 4584 9918 4593
rect 9128 4276 9180 4282
rect 9128 4218 9180 4224
rect 8852 4208 8904 4214
rect 8852 4150 8904 4156
rect 8760 4140 8812 4146
rect 8760 4082 8812 4088
rect 8576 4072 8628 4078
rect 8576 4014 8628 4020
rect 8760 3936 8812 3942
rect 8760 3878 8812 3884
rect 8208 3460 8260 3466
rect 8208 3402 8260 3408
rect 8220 3058 8248 3402
rect 8772 3126 8800 3878
rect 9600 3738 9628 4558
rect 9862 4519 9918 4528
rect 9968 4185 9996 7783
rect 10048 6792 10100 6798
rect 10152 6780 10180 7958
rect 10244 6798 10272 8978
rect 10336 8566 10364 9646
rect 10612 9586 10640 17002
rect 10888 12434 10916 17614
rect 11060 17604 11112 17610
rect 11060 17546 11112 17552
rect 11072 17270 11100 17546
rect 11060 17264 11112 17270
rect 11060 17206 11112 17212
rect 11152 16516 11204 16522
rect 11256 16504 11284 17614
rect 11348 16590 11376 18294
rect 11440 18290 11468 18566
rect 11428 18284 11480 18290
rect 11428 18226 11480 18232
rect 11440 17678 11468 18226
rect 11428 17672 11480 17678
rect 11428 17614 11480 17620
rect 11336 16584 11388 16590
rect 11336 16526 11388 16532
rect 11204 16476 11284 16504
rect 11152 16458 11204 16464
rect 11428 16448 11480 16454
rect 11428 16390 11480 16396
rect 11440 16046 11468 16390
rect 11428 16040 11480 16046
rect 11428 15982 11480 15988
rect 11244 15496 11296 15502
rect 11244 15438 11296 15444
rect 10968 12708 11020 12714
rect 10968 12650 11020 12656
rect 10704 12406 10916 12434
rect 10704 10690 10732 12406
rect 10876 12368 10928 12374
rect 10876 12310 10928 12316
rect 10784 12232 10836 12238
rect 10784 12174 10836 12180
rect 10796 11354 10824 12174
rect 10784 11348 10836 11354
rect 10784 11290 10836 11296
rect 10888 11082 10916 12310
rect 10980 11762 11008 12650
rect 11060 12640 11112 12646
rect 11060 12582 11112 12588
rect 10968 11756 11020 11762
rect 11072 11744 11100 12582
rect 11256 12170 11284 15438
rect 11336 14408 11388 14414
rect 11336 14350 11388 14356
rect 11348 13938 11376 14350
rect 11336 13932 11388 13938
rect 11336 13874 11388 13880
rect 11440 13818 11468 15982
rect 11520 14408 11572 14414
rect 11520 14350 11572 14356
rect 11532 13870 11560 14350
rect 11348 13790 11468 13818
rect 11520 13864 11572 13870
rect 11520 13806 11572 13812
rect 11348 12238 11376 13790
rect 11624 12850 11652 18702
rect 11716 15570 11744 18702
rect 11992 17610 12020 18770
rect 12728 18748 12756 19382
rect 12820 18902 12848 24278
rect 13004 24138 13032 24704
rect 13084 24686 13136 24692
rect 13096 24274 13308 24290
rect 13084 24268 13320 24274
rect 13136 24262 13268 24268
rect 13084 24210 13136 24216
rect 13268 24210 13320 24216
rect 12992 24132 13044 24138
rect 12992 24074 13044 24080
rect 13004 23730 13032 24074
rect 12992 23724 13044 23730
rect 12992 23666 13044 23672
rect 13280 22710 13308 24210
rect 13372 24177 13400 24822
rect 13452 24812 13504 24818
rect 13452 24754 13504 24760
rect 13358 24168 13414 24177
rect 13358 24103 13414 24112
rect 13372 24070 13400 24103
rect 13360 24064 13412 24070
rect 13360 24006 13412 24012
rect 13464 23798 13492 24754
rect 13648 24682 13676 25162
rect 13832 24818 13860 25230
rect 13820 24812 13872 24818
rect 13820 24754 13872 24760
rect 14096 24812 14148 24818
rect 14096 24754 14148 24760
rect 14188 24812 14240 24818
rect 14188 24754 14240 24760
rect 13636 24676 13688 24682
rect 13636 24618 13688 24624
rect 13832 24614 13860 24754
rect 13820 24608 13872 24614
rect 13820 24550 13872 24556
rect 13832 24410 13860 24550
rect 14108 24410 14136 24754
rect 13820 24404 13872 24410
rect 13820 24346 13872 24352
rect 14096 24404 14148 24410
rect 14096 24346 14148 24352
rect 14200 23866 14228 24754
rect 14384 24682 14412 25230
rect 14556 25152 14608 25158
rect 14556 25094 14608 25100
rect 14372 24676 14424 24682
rect 14372 24618 14424 24624
rect 14568 24138 14596 25094
rect 15212 24614 15240 25230
rect 15200 24608 15252 24614
rect 15200 24550 15252 24556
rect 15212 24274 15240 24550
rect 15304 24410 15332 25842
rect 16948 25832 17000 25838
rect 16948 25774 17000 25780
rect 15476 25696 15528 25702
rect 15476 25638 15528 25644
rect 15488 25362 15516 25638
rect 15476 25356 15528 25362
rect 15476 25298 15528 25304
rect 16028 25220 16080 25226
rect 16028 25162 16080 25168
rect 15384 24948 15436 24954
rect 15384 24890 15436 24896
rect 15396 24614 15424 24890
rect 16040 24886 16068 25162
rect 16960 25158 16988 25774
rect 17592 25288 17644 25294
rect 17592 25230 17644 25236
rect 16948 25152 17000 25158
rect 16948 25094 17000 25100
rect 16028 24880 16080 24886
rect 16028 24822 16080 24828
rect 16212 24812 16264 24818
rect 16212 24754 16264 24760
rect 16764 24812 16816 24818
rect 16764 24754 16816 24760
rect 15384 24608 15436 24614
rect 15384 24550 15436 24556
rect 16224 24410 16252 24754
rect 16304 24676 16356 24682
rect 16304 24618 16356 24624
rect 15292 24404 15344 24410
rect 15292 24346 15344 24352
rect 16212 24404 16264 24410
rect 16212 24346 16264 24352
rect 15844 24336 15896 24342
rect 15844 24278 15896 24284
rect 15200 24268 15252 24274
rect 15200 24210 15252 24216
rect 15660 24200 15712 24206
rect 15660 24142 15712 24148
rect 14556 24132 14608 24138
rect 14556 24074 14608 24080
rect 14188 23860 14240 23866
rect 14188 23802 14240 23808
rect 13452 23792 13504 23798
rect 13452 23734 13504 23740
rect 15672 23508 15700 24142
rect 15488 23480 15700 23508
rect 15384 23248 15436 23254
rect 15384 23190 15436 23196
rect 15108 23112 15160 23118
rect 15108 23054 15160 23060
rect 13268 22704 13320 22710
rect 13268 22646 13320 22652
rect 13084 22636 13136 22642
rect 13084 22578 13136 22584
rect 12900 21956 12952 21962
rect 12900 21898 12952 21904
rect 12912 21554 12940 21898
rect 12900 21548 12952 21554
rect 12952 21508 13032 21536
rect 12900 21490 12952 21496
rect 12900 21344 12952 21350
rect 12900 21286 12952 21292
rect 12912 20942 12940 21286
rect 12900 20936 12952 20942
rect 12900 20878 12952 20884
rect 13004 20806 13032 21508
rect 13096 21418 13124 22578
rect 13176 22094 13228 22098
rect 13280 22094 13308 22646
rect 14096 22636 14148 22642
rect 14096 22578 14148 22584
rect 13176 22092 13308 22094
rect 13228 22066 13308 22092
rect 13176 22034 13228 22040
rect 13188 22003 13216 22034
rect 13280 21554 13308 22066
rect 14108 21690 14136 22578
rect 15016 22568 15068 22574
rect 15120 22556 15148 23054
rect 15292 23044 15344 23050
rect 15292 22986 15344 22992
rect 15304 22778 15332 22986
rect 15292 22772 15344 22778
rect 15292 22714 15344 22720
rect 15396 22642 15424 23190
rect 15292 22636 15344 22642
rect 15292 22578 15344 22584
rect 15384 22636 15436 22642
rect 15384 22578 15436 22584
rect 15068 22528 15148 22556
rect 15016 22510 15068 22516
rect 14372 22432 14424 22438
rect 14372 22374 14424 22380
rect 14096 21684 14148 21690
rect 14096 21626 14148 21632
rect 13268 21548 13320 21554
rect 13268 21490 13320 21496
rect 13084 21412 13136 21418
rect 13084 21354 13136 21360
rect 12992 20800 13044 20806
rect 12992 20742 13044 20748
rect 14108 20602 14136 21626
rect 14384 21486 14412 22374
rect 15120 21894 15148 22528
rect 15200 22432 15252 22438
rect 15200 22374 15252 22380
rect 15108 21888 15160 21894
rect 15108 21830 15160 21836
rect 14372 21480 14424 21486
rect 14372 21422 14424 21428
rect 14384 20874 14412 21422
rect 14832 21344 14884 21350
rect 14832 21286 14884 21292
rect 14844 21010 14872 21286
rect 14832 21004 14884 21010
rect 14832 20946 14884 20952
rect 15212 20942 15240 22374
rect 15200 20936 15252 20942
rect 15200 20878 15252 20884
rect 14372 20868 14424 20874
rect 14372 20810 14424 20816
rect 14096 20596 14148 20602
rect 14096 20538 14148 20544
rect 15304 20505 15332 22578
rect 15488 22438 15516 23480
rect 15752 23180 15804 23186
rect 15752 23122 15804 23128
rect 15568 22976 15620 22982
rect 15568 22918 15620 22924
rect 15580 22506 15608 22918
rect 15568 22500 15620 22506
rect 15568 22442 15620 22448
rect 15476 22432 15528 22438
rect 15476 22374 15528 22380
rect 15488 21962 15516 22374
rect 15476 21956 15528 21962
rect 15476 21898 15528 21904
rect 15476 21480 15528 21486
rect 15476 21422 15528 21428
rect 15488 21146 15516 21422
rect 15476 21140 15528 21146
rect 15476 21082 15528 21088
rect 13082 20496 13138 20505
rect 13082 20431 13138 20440
rect 15290 20496 15346 20505
rect 15290 20431 15346 20440
rect 12900 19712 12952 19718
rect 12900 19654 12952 19660
rect 12808 18896 12860 18902
rect 12808 18838 12860 18844
rect 12912 18834 12940 19654
rect 12992 19304 13044 19310
rect 12992 19246 13044 19252
rect 12900 18828 12952 18834
rect 12900 18770 12952 18776
rect 13004 18766 13032 19246
rect 12992 18760 13044 18766
rect 12728 18720 12848 18748
rect 12624 18624 12676 18630
rect 12624 18566 12676 18572
rect 12716 18624 12768 18630
rect 12716 18566 12768 18572
rect 12636 18290 12664 18566
rect 12624 18284 12676 18290
rect 12624 18226 12676 18232
rect 11980 17604 12032 17610
rect 11980 17546 12032 17552
rect 11796 15904 11848 15910
rect 11796 15846 11848 15852
rect 11808 15570 11836 15846
rect 11704 15564 11756 15570
rect 11704 15506 11756 15512
rect 11796 15564 11848 15570
rect 11796 15506 11848 15512
rect 11612 12844 11664 12850
rect 11612 12786 11664 12792
rect 11428 12640 11480 12646
rect 11428 12582 11480 12588
rect 11440 12238 11468 12582
rect 11336 12232 11388 12238
rect 11336 12174 11388 12180
rect 11428 12232 11480 12238
rect 11428 12174 11480 12180
rect 11244 12164 11296 12170
rect 11244 12106 11296 12112
rect 11072 11716 11284 11744
rect 10968 11698 11020 11704
rect 11060 11620 11112 11626
rect 11060 11562 11112 11568
rect 11072 11286 11100 11562
rect 11060 11280 11112 11286
rect 11060 11222 11112 11228
rect 10876 11076 10928 11082
rect 10876 11018 10928 11024
rect 10704 10662 10824 10690
rect 10692 10600 10744 10606
rect 10692 10542 10744 10548
rect 10704 9926 10732 10542
rect 10692 9920 10744 9926
rect 10692 9862 10744 9868
rect 10600 9580 10652 9586
rect 10600 9522 10652 9528
rect 10600 8900 10652 8906
rect 10600 8842 10652 8848
rect 10324 8560 10376 8566
rect 10324 8502 10376 8508
rect 10336 7460 10364 8502
rect 10612 8090 10640 8842
rect 10796 8650 10824 10662
rect 10888 9926 10916 11018
rect 10968 11008 11020 11014
rect 10968 10950 11020 10956
rect 10876 9920 10928 9926
rect 10876 9862 10928 9868
rect 10876 9580 10928 9586
rect 10876 9522 10928 9528
rect 10704 8634 10824 8650
rect 10692 8628 10824 8634
rect 10744 8622 10824 8628
rect 10692 8570 10744 8576
rect 10600 8084 10652 8090
rect 10600 8026 10652 8032
rect 10414 7984 10470 7993
rect 10414 7919 10416 7928
rect 10468 7919 10470 7928
rect 10416 7890 10468 7896
rect 10508 7744 10560 7750
rect 10508 7686 10560 7692
rect 10416 7472 10468 7478
rect 10336 7432 10416 7460
rect 10416 7414 10468 7420
rect 10100 6752 10180 6780
rect 10232 6792 10284 6798
rect 10048 6734 10100 6740
rect 10232 6734 10284 6740
rect 10244 5574 10272 6734
rect 10232 5568 10284 5574
rect 10232 5510 10284 5516
rect 10140 5092 10192 5098
rect 10140 5034 10192 5040
rect 10152 4622 10180 5034
rect 10140 4616 10192 4622
rect 10140 4558 10192 4564
rect 9954 4176 10010 4185
rect 9864 4140 9916 4146
rect 9954 4111 10010 4120
rect 9864 4082 9916 4088
rect 9588 3732 9640 3738
rect 9588 3674 9640 3680
rect 8760 3120 8812 3126
rect 8760 3062 8812 3068
rect 8208 3052 8260 3058
rect 8208 2994 8260 3000
rect 9876 2990 9904 4082
rect 10244 4078 10272 5510
rect 10232 4072 10284 4078
rect 10232 4014 10284 4020
rect 10428 3466 10456 7414
rect 10520 7002 10548 7686
rect 10692 7200 10744 7206
rect 10692 7142 10744 7148
rect 10508 6996 10560 7002
rect 10508 6938 10560 6944
rect 10704 6798 10732 7142
rect 10692 6792 10744 6798
rect 10692 6734 10744 6740
rect 10796 6730 10824 8622
rect 10888 7857 10916 9522
rect 10980 9382 11008 10950
rect 10968 9376 11020 9382
rect 10968 9318 11020 9324
rect 10968 8968 11020 8974
rect 10968 8910 11020 8916
rect 10980 8634 11008 8910
rect 10968 8628 11020 8634
rect 10968 8570 11020 8576
rect 10980 7886 11008 8570
rect 10968 7880 11020 7886
rect 10874 7848 10930 7857
rect 10968 7822 11020 7828
rect 10874 7783 10876 7792
rect 10928 7783 10930 7792
rect 10876 7754 10928 7760
rect 10968 7404 11020 7410
rect 10968 7346 11020 7352
rect 10980 6866 11008 7346
rect 11152 7336 11204 7342
rect 11152 7278 11204 7284
rect 10968 6860 11020 6866
rect 10968 6802 11020 6808
rect 11164 6798 11192 7278
rect 11152 6792 11204 6798
rect 11152 6734 11204 6740
rect 10784 6724 10836 6730
rect 10784 6666 10836 6672
rect 11164 5642 11192 6734
rect 11256 6662 11284 11716
rect 11440 11082 11468 12174
rect 11520 12164 11572 12170
rect 11520 12106 11572 12112
rect 11532 11218 11560 12106
rect 11520 11212 11572 11218
rect 11520 11154 11572 11160
rect 11428 11076 11480 11082
rect 11428 11018 11480 11024
rect 11520 11008 11572 11014
rect 11520 10950 11572 10956
rect 11532 10674 11560 10950
rect 11520 10668 11572 10674
rect 11520 10610 11572 10616
rect 11624 7750 11652 12786
rect 11716 12782 11744 15506
rect 11888 14612 11940 14618
rect 11888 14554 11940 14560
rect 11900 14074 11928 14554
rect 11888 14068 11940 14074
rect 11888 14010 11940 14016
rect 11704 12776 11756 12782
rect 11704 12718 11756 12724
rect 11704 12232 11756 12238
rect 11704 12174 11756 12180
rect 11716 11558 11744 12174
rect 11704 11552 11756 11558
rect 11704 11494 11756 11500
rect 11900 10606 11928 14010
rect 11992 12434 12020 17546
rect 12348 17536 12400 17542
rect 12348 17478 12400 17484
rect 12360 17202 12388 17478
rect 12348 17196 12400 17202
rect 12348 17138 12400 17144
rect 12440 17196 12492 17202
rect 12440 17138 12492 17144
rect 12164 16992 12216 16998
rect 12164 16934 12216 16940
rect 12176 15570 12204 16934
rect 12452 16658 12480 17138
rect 12440 16652 12492 16658
rect 12440 16594 12492 16600
rect 12440 16516 12492 16522
rect 12440 16458 12492 16464
rect 12452 15706 12480 16458
rect 12728 16114 12756 18566
rect 12820 18358 12848 18720
rect 12992 18702 13044 18708
rect 12808 18352 12860 18358
rect 12808 18294 12860 18300
rect 12820 17202 12848 18294
rect 12808 17196 12860 17202
rect 12808 17138 12860 17144
rect 12820 17082 12848 17138
rect 12820 17054 12940 17082
rect 12808 16992 12860 16998
rect 12808 16934 12860 16940
rect 12820 16590 12848 16934
rect 12808 16584 12860 16590
rect 12808 16526 12860 16532
rect 12820 16250 12848 16526
rect 12808 16244 12860 16250
rect 12808 16186 12860 16192
rect 12716 16108 12768 16114
rect 12716 16050 12768 16056
rect 12532 15904 12584 15910
rect 12532 15846 12584 15852
rect 12440 15700 12492 15706
rect 12440 15642 12492 15648
rect 12164 15564 12216 15570
rect 12164 15506 12216 15512
rect 12544 15502 12572 15846
rect 12532 15496 12584 15502
rect 12532 15438 12584 15444
rect 12532 15360 12584 15366
rect 12532 15302 12584 15308
rect 12164 14272 12216 14278
rect 12164 14214 12216 14220
rect 12176 13802 12204 14214
rect 12256 13932 12308 13938
rect 12256 13874 12308 13880
rect 12164 13796 12216 13802
rect 12164 13738 12216 13744
rect 12268 12918 12296 13874
rect 12256 12912 12308 12918
rect 12256 12854 12308 12860
rect 11992 12406 12112 12434
rect 12084 12306 12112 12406
rect 12072 12300 12124 12306
rect 12072 12242 12124 12248
rect 12164 12300 12216 12306
rect 12164 12242 12216 12248
rect 11980 12232 12032 12238
rect 11980 12174 12032 12180
rect 11992 11558 12020 12174
rect 11980 11552 12032 11558
rect 11980 11494 12032 11500
rect 11992 11234 12020 11494
rect 12084 11354 12112 12242
rect 12072 11348 12124 11354
rect 12072 11290 12124 11296
rect 11992 11206 12112 11234
rect 12084 11014 12112 11206
rect 12176 11150 12204 12242
rect 12268 12238 12296 12854
rect 12348 12776 12400 12782
rect 12348 12718 12400 12724
rect 12360 12238 12388 12718
rect 12440 12640 12492 12646
rect 12440 12582 12492 12588
rect 12256 12232 12308 12238
rect 12256 12174 12308 12180
rect 12348 12232 12400 12238
rect 12348 12174 12400 12180
rect 12256 12096 12308 12102
rect 12256 12038 12308 12044
rect 12268 11286 12296 12038
rect 12256 11280 12308 11286
rect 12256 11222 12308 11228
rect 12164 11144 12216 11150
rect 12164 11086 12216 11092
rect 12256 11144 12308 11150
rect 12256 11086 12308 11092
rect 12072 11008 12124 11014
rect 12072 10950 12124 10956
rect 12084 10674 12112 10950
rect 12072 10668 12124 10674
rect 12072 10610 12124 10616
rect 11888 10600 11940 10606
rect 11888 10542 11940 10548
rect 12268 10538 12296 11086
rect 12256 10532 12308 10538
rect 12256 10474 12308 10480
rect 11888 9988 11940 9994
rect 11888 9930 11940 9936
rect 11900 9586 11928 9930
rect 12360 9874 12388 12174
rect 12452 11098 12480 12582
rect 12544 12442 12572 15302
rect 12624 15156 12676 15162
rect 12624 15098 12676 15104
rect 12636 14006 12664 15098
rect 12912 15094 12940 17054
rect 13004 16250 13032 18702
rect 12992 16244 13044 16250
rect 12992 16186 13044 16192
rect 12992 16108 13044 16114
rect 12992 16050 13044 16056
rect 13004 15162 13032 16050
rect 13096 15706 13124 20431
rect 14188 20392 14240 20398
rect 14188 20334 14240 20340
rect 13268 19848 13320 19854
rect 13268 19790 13320 19796
rect 13280 18766 13308 19790
rect 13544 19712 13596 19718
rect 13544 19654 13596 19660
rect 13556 19378 13584 19654
rect 13544 19372 13596 19378
rect 13544 19314 13596 19320
rect 14200 19310 14228 20334
rect 15764 19990 15792 23122
rect 15856 23118 15884 24278
rect 16028 24268 16080 24274
rect 16028 24210 16080 24216
rect 16040 23730 16068 24210
rect 16224 24206 16252 24346
rect 16212 24200 16264 24206
rect 16212 24142 16264 24148
rect 16224 23866 16252 24142
rect 16316 24138 16344 24618
rect 16304 24132 16356 24138
rect 16304 24074 16356 24080
rect 16212 23860 16264 23866
rect 16212 23802 16264 23808
rect 16316 23730 16344 24074
rect 16776 23866 16804 24754
rect 16856 24608 16908 24614
rect 16856 24550 16908 24556
rect 16764 23860 16816 23866
rect 16764 23802 16816 23808
rect 16868 23730 16896 24550
rect 16960 24410 16988 25094
rect 17040 24812 17092 24818
rect 17040 24754 17092 24760
rect 16948 24404 17000 24410
rect 16948 24346 17000 24352
rect 17052 24342 17080 24754
rect 17132 24744 17184 24750
rect 17132 24686 17184 24692
rect 17040 24336 17092 24342
rect 17040 24278 17092 24284
rect 16028 23724 16080 23730
rect 16028 23666 16080 23672
rect 16120 23724 16172 23730
rect 16120 23666 16172 23672
rect 16304 23724 16356 23730
rect 16304 23666 16356 23672
rect 16856 23724 16908 23730
rect 16856 23666 16908 23672
rect 16132 23118 16160 23666
rect 17144 23594 17172 24686
rect 17408 24608 17460 24614
rect 17408 24550 17460 24556
rect 17420 24410 17448 24550
rect 17408 24404 17460 24410
rect 17408 24346 17460 24352
rect 17604 24274 17632 25230
rect 17696 24682 17724 25842
rect 17788 24886 17816 25910
rect 21180 25832 21232 25838
rect 21180 25774 21232 25780
rect 19524 25696 19576 25702
rect 19524 25638 19576 25644
rect 19536 25362 19564 25638
rect 21192 25498 21220 25774
rect 21456 25764 21508 25770
rect 21456 25706 21508 25712
rect 21180 25492 21232 25498
rect 21180 25434 21232 25440
rect 19524 25356 19576 25362
rect 19524 25298 19576 25304
rect 19248 25288 19300 25294
rect 19248 25230 19300 25236
rect 21272 25288 21324 25294
rect 21272 25230 21324 25236
rect 17868 24948 17920 24954
rect 17868 24890 17920 24896
rect 17776 24880 17828 24886
rect 17776 24822 17828 24828
rect 17880 24698 17908 24890
rect 19260 24818 19288 25230
rect 20536 25220 20588 25226
rect 20536 25162 20588 25168
rect 19248 24812 19300 24818
rect 19248 24754 19300 24760
rect 19156 24744 19208 24750
rect 17684 24676 17736 24682
rect 17880 24670 18000 24698
rect 19156 24686 19208 24692
rect 17684 24618 17736 24624
rect 17868 24608 17920 24614
rect 17868 24550 17920 24556
rect 17592 24268 17644 24274
rect 17592 24210 17644 24216
rect 17604 23662 17632 24210
rect 17880 23798 17908 24550
rect 17972 24154 18000 24670
rect 19168 24410 19196 24686
rect 19156 24404 19208 24410
rect 19156 24346 19208 24352
rect 19524 24268 19576 24274
rect 19524 24210 19576 24216
rect 17972 24138 18092 24154
rect 17972 24132 18104 24138
rect 17972 24126 18052 24132
rect 17972 23798 18000 24126
rect 18052 24074 18104 24080
rect 19432 24064 19484 24070
rect 19432 24006 19484 24012
rect 17868 23792 17920 23798
rect 17868 23734 17920 23740
rect 17960 23792 18012 23798
rect 17960 23734 18012 23740
rect 17592 23656 17644 23662
rect 17592 23598 17644 23604
rect 17132 23588 17184 23594
rect 17132 23530 17184 23536
rect 17144 23186 17172 23530
rect 17604 23186 17632 23598
rect 17132 23180 17184 23186
rect 17132 23122 17184 23128
rect 17592 23180 17644 23186
rect 17592 23122 17644 23128
rect 15844 23112 15896 23118
rect 15844 23054 15896 23060
rect 16120 23112 16172 23118
rect 16120 23054 16172 23060
rect 15856 22710 15884 23054
rect 15844 22704 15896 22710
rect 15844 22646 15896 22652
rect 15936 22568 15988 22574
rect 15936 22510 15988 22516
rect 15948 22234 15976 22510
rect 15936 22228 15988 22234
rect 15936 22170 15988 22176
rect 15948 21962 15976 22170
rect 16132 22166 16160 23054
rect 17500 23044 17552 23050
rect 17500 22986 17552 22992
rect 16488 22500 16540 22506
rect 16488 22442 16540 22448
rect 16500 22234 16528 22442
rect 16672 22432 16724 22438
rect 16672 22374 16724 22380
rect 16488 22228 16540 22234
rect 16488 22170 16540 22176
rect 16120 22160 16172 22166
rect 16120 22102 16172 22108
rect 16132 22030 16160 22102
rect 16120 22024 16172 22030
rect 16120 21966 16172 21972
rect 15936 21956 15988 21962
rect 15936 21898 15988 21904
rect 16500 21690 16528 22170
rect 16684 22030 16712 22374
rect 16672 22024 16724 22030
rect 16672 21966 16724 21972
rect 16488 21684 16540 21690
rect 16488 21626 16540 21632
rect 16304 21616 16356 21622
rect 16304 21558 16356 21564
rect 15844 20936 15896 20942
rect 15844 20878 15896 20884
rect 15752 19984 15804 19990
rect 15752 19926 15804 19932
rect 15752 19712 15804 19718
rect 15752 19654 15804 19660
rect 14188 19304 14240 19310
rect 14188 19246 14240 19252
rect 15568 19304 15620 19310
rect 15568 19246 15620 19252
rect 14200 18834 14228 19246
rect 14556 19168 14608 19174
rect 14556 19110 14608 19116
rect 14188 18828 14240 18834
rect 14188 18770 14240 18776
rect 13268 18760 13320 18766
rect 13268 18702 13320 18708
rect 13268 18624 13320 18630
rect 13268 18566 13320 18572
rect 14096 18624 14148 18630
rect 14096 18566 14148 18572
rect 13176 16448 13228 16454
rect 13176 16390 13228 16396
rect 13084 15700 13136 15706
rect 13084 15642 13136 15648
rect 13188 15570 13216 16390
rect 13176 15564 13228 15570
rect 13176 15506 13228 15512
rect 12992 15156 13044 15162
rect 12992 15098 13044 15104
rect 12900 15088 12952 15094
rect 12900 15030 12952 15036
rect 12912 14346 12940 15030
rect 12900 14340 12952 14346
rect 12900 14282 12952 14288
rect 12808 14272 12860 14278
rect 12808 14214 12860 14220
rect 12820 14006 12848 14214
rect 13280 14090 13308 18566
rect 14108 18222 14136 18566
rect 14096 18216 14148 18222
rect 14096 18158 14148 18164
rect 14200 18086 14228 18770
rect 14568 18766 14596 19110
rect 14464 18760 14516 18766
rect 14464 18702 14516 18708
rect 14556 18760 14608 18766
rect 14556 18702 14608 18708
rect 14476 18630 14504 18702
rect 15384 18692 15436 18698
rect 15384 18634 15436 18640
rect 14464 18624 14516 18630
rect 14464 18566 14516 18572
rect 15200 18624 15252 18630
rect 15200 18566 15252 18572
rect 14280 18420 14332 18426
rect 14280 18362 14332 18368
rect 14292 18086 14320 18362
rect 14188 18080 14240 18086
rect 14188 18022 14240 18028
rect 14280 18080 14332 18086
rect 14280 18022 14332 18028
rect 14200 17134 14228 18022
rect 13912 17128 13964 17134
rect 13912 17070 13964 17076
rect 14188 17128 14240 17134
rect 14188 17070 14240 17076
rect 13544 16448 13596 16454
rect 13464 16408 13544 16436
rect 13464 16114 13492 16408
rect 13544 16390 13596 16396
rect 13728 16176 13780 16182
rect 13728 16118 13780 16124
rect 13452 16108 13504 16114
rect 13452 16050 13504 16056
rect 13544 16108 13596 16114
rect 13544 16050 13596 16056
rect 13452 15904 13504 15910
rect 13452 15846 13504 15852
rect 13464 15502 13492 15846
rect 13452 15496 13504 15502
rect 13452 15438 13504 15444
rect 13360 14952 13412 14958
rect 13360 14894 13412 14900
rect 13372 14550 13400 14894
rect 13360 14544 13412 14550
rect 13360 14486 13412 14492
rect 13452 14272 13504 14278
rect 13556 14260 13584 16050
rect 13740 15434 13768 16118
rect 13924 15706 13952 17070
rect 14200 16658 14228 17070
rect 14188 16652 14240 16658
rect 14188 16594 14240 16600
rect 14200 16114 14228 16594
rect 14292 16590 14320 18022
rect 14740 16992 14792 16998
rect 14740 16934 14792 16940
rect 14752 16658 14780 16934
rect 14740 16652 14792 16658
rect 14740 16594 14792 16600
rect 14280 16584 14332 16590
rect 14280 16526 14332 16532
rect 15108 16448 15160 16454
rect 15212 16436 15240 18566
rect 15396 18426 15424 18634
rect 15384 18420 15436 18426
rect 15384 18362 15436 18368
rect 15580 18222 15608 19246
rect 15764 18850 15792 19654
rect 15856 18970 15884 20878
rect 15936 20800 15988 20806
rect 15936 20742 15988 20748
rect 15948 20398 15976 20742
rect 16316 20534 16344 21558
rect 17512 21146 17540 22986
rect 17604 22098 17632 23122
rect 17972 23050 18000 23734
rect 19444 23730 19472 24006
rect 19432 23724 19484 23730
rect 19432 23666 19484 23672
rect 19536 23610 19564 24210
rect 20168 24200 20220 24206
rect 20168 24142 20220 24148
rect 19616 24064 19668 24070
rect 19616 24006 19668 24012
rect 19708 24064 19760 24070
rect 19708 24006 19760 24012
rect 19628 23798 19656 24006
rect 19720 23866 19748 24006
rect 20180 23866 20208 24142
rect 19708 23860 19760 23866
rect 19708 23802 19760 23808
rect 20168 23860 20220 23866
rect 20168 23802 20220 23808
rect 19616 23792 19668 23798
rect 19616 23734 19668 23740
rect 19800 23724 19852 23730
rect 19800 23666 19852 23672
rect 19616 23656 19668 23662
rect 19536 23604 19616 23610
rect 19536 23598 19668 23604
rect 19536 23582 19656 23598
rect 19340 23112 19392 23118
rect 19340 23054 19392 23060
rect 17960 23044 18012 23050
rect 17960 22986 18012 22992
rect 17972 22778 18000 22986
rect 17960 22772 18012 22778
rect 17960 22714 18012 22720
rect 18880 22772 18932 22778
rect 18880 22714 18932 22720
rect 17592 22092 17644 22098
rect 17592 22034 17644 22040
rect 18892 21962 18920 22714
rect 19248 22092 19300 22098
rect 19248 22034 19300 22040
rect 17592 21956 17644 21962
rect 17592 21898 17644 21904
rect 18880 21956 18932 21962
rect 18880 21898 18932 21904
rect 17500 21140 17552 21146
rect 17500 21082 17552 21088
rect 17408 20800 17460 20806
rect 17408 20742 17460 20748
rect 16396 20596 16448 20602
rect 16396 20538 16448 20544
rect 16304 20528 16356 20534
rect 16304 20470 16356 20476
rect 15936 20392 15988 20398
rect 15936 20334 15988 20340
rect 16212 20256 16264 20262
rect 16212 20198 16264 20204
rect 16028 19848 16080 19854
rect 16028 19790 16080 19796
rect 16040 19514 16068 19790
rect 16028 19508 16080 19514
rect 16028 19450 16080 19456
rect 16224 19378 16252 20198
rect 16212 19372 16264 19378
rect 16212 19314 16264 19320
rect 15844 18964 15896 18970
rect 15844 18906 15896 18912
rect 15764 18822 15884 18850
rect 15856 18358 15884 18822
rect 16408 18630 16436 20538
rect 16488 20460 16540 20466
rect 16488 20402 16540 20408
rect 16500 19922 16528 20402
rect 17040 20392 17092 20398
rect 17040 20334 17092 20340
rect 17052 19990 17080 20334
rect 17420 20058 17448 20742
rect 17604 20058 17632 21898
rect 18892 21622 18920 21898
rect 19260 21622 19288 22034
rect 19352 21894 19380 23054
rect 19524 22432 19576 22438
rect 19524 22374 19576 22380
rect 19536 22234 19564 22374
rect 19524 22228 19576 22234
rect 19524 22170 19576 22176
rect 19340 21888 19392 21894
rect 19340 21830 19392 21836
rect 18880 21616 18932 21622
rect 18880 21558 18932 21564
rect 19248 21616 19300 21622
rect 19248 21558 19300 21564
rect 19260 21010 19288 21558
rect 19340 21548 19392 21554
rect 19340 21490 19392 21496
rect 19248 21004 19300 21010
rect 19248 20946 19300 20952
rect 17960 20936 18012 20942
rect 17960 20878 18012 20884
rect 17408 20052 17460 20058
rect 17408 19994 17460 20000
rect 17592 20052 17644 20058
rect 17592 19994 17644 20000
rect 17040 19984 17092 19990
rect 17040 19926 17092 19932
rect 16488 19916 16540 19922
rect 16488 19858 16540 19864
rect 16500 19310 16528 19858
rect 17052 19378 17080 19926
rect 17972 19854 18000 20878
rect 18420 20868 18472 20874
rect 18420 20810 18472 20816
rect 18236 20256 18288 20262
rect 18236 20198 18288 20204
rect 18248 19854 18276 20198
rect 18432 19854 18460 20810
rect 19260 20602 19288 20946
rect 19248 20596 19300 20602
rect 19248 20538 19300 20544
rect 18880 20392 18932 20398
rect 18880 20334 18932 20340
rect 19352 20346 19380 21490
rect 19628 21486 19656 23582
rect 19812 23322 19840 23666
rect 19800 23316 19852 23322
rect 19800 23258 19852 23264
rect 20352 22568 20404 22574
rect 20352 22510 20404 22516
rect 19800 21956 19852 21962
rect 19800 21898 19852 21904
rect 19616 21480 19668 21486
rect 19616 21422 19668 21428
rect 19812 20534 19840 21898
rect 20364 21690 20392 22510
rect 20548 21962 20576 25162
rect 21284 24410 21312 25230
rect 21364 25152 21416 25158
rect 21364 25094 21416 25100
rect 21376 24750 21404 25094
rect 21364 24744 21416 24750
rect 21364 24686 21416 24692
rect 21272 24404 21324 24410
rect 21272 24346 21324 24352
rect 21468 24342 21496 25706
rect 21548 25492 21600 25498
rect 21548 25434 21600 25440
rect 21560 24682 21588 25434
rect 22100 25288 22152 25294
rect 22100 25230 22152 25236
rect 22112 24954 22140 25230
rect 22100 24948 22152 24954
rect 22100 24890 22152 24896
rect 22468 24812 22520 24818
rect 22848 24800 22876 25910
rect 23296 25832 23348 25838
rect 23296 25774 23348 25780
rect 24032 25832 24084 25838
rect 24032 25774 24084 25780
rect 24308 25832 24360 25838
rect 24308 25774 24360 25780
rect 22928 25696 22980 25702
rect 22928 25638 22980 25644
rect 22940 25294 22968 25638
rect 22928 25288 22980 25294
rect 22928 25230 22980 25236
rect 22520 24772 22876 24800
rect 22468 24754 22520 24760
rect 22284 24744 22336 24750
rect 22284 24686 22336 24692
rect 21548 24676 21600 24682
rect 21548 24618 21600 24624
rect 22008 24676 22060 24682
rect 22008 24618 22060 24624
rect 21456 24336 21508 24342
rect 21456 24278 21508 24284
rect 21180 24268 21232 24274
rect 21180 24210 21232 24216
rect 21088 24200 21140 24206
rect 21088 24142 21140 24148
rect 20996 24064 21048 24070
rect 20996 24006 21048 24012
rect 21008 23730 21036 24006
rect 21100 23866 21128 24142
rect 21088 23860 21140 23866
rect 21088 23802 21140 23808
rect 21192 23730 21220 24210
rect 21468 24206 21496 24278
rect 21560 24206 21588 24618
rect 21732 24608 21784 24614
rect 21732 24550 21784 24556
rect 21744 24206 21772 24550
rect 22020 24342 22048 24618
rect 22008 24336 22060 24342
rect 22008 24278 22060 24284
rect 21456 24200 21508 24206
rect 21456 24142 21508 24148
rect 21548 24200 21600 24206
rect 21548 24142 21600 24148
rect 21732 24200 21784 24206
rect 21732 24142 21784 24148
rect 21272 24132 21324 24138
rect 21272 24074 21324 24080
rect 21284 23798 21312 24074
rect 21640 24064 21692 24070
rect 21640 24006 21692 24012
rect 21272 23792 21324 23798
rect 21272 23734 21324 23740
rect 21652 23730 21680 24006
rect 20996 23724 21048 23730
rect 20996 23666 21048 23672
rect 21180 23724 21232 23730
rect 21180 23666 21232 23672
rect 21364 23724 21416 23730
rect 21364 23666 21416 23672
rect 21640 23724 21692 23730
rect 21692 23684 21772 23712
rect 21640 23666 21692 23672
rect 20812 23656 20864 23662
rect 20812 23598 20864 23604
rect 20824 23254 20852 23598
rect 20812 23248 20864 23254
rect 20812 23190 20864 23196
rect 21376 23050 21404 23666
rect 21640 23520 21692 23526
rect 21640 23462 21692 23468
rect 21652 23118 21680 23462
rect 21744 23186 21772 23684
rect 22020 23662 22048 24278
rect 22296 24206 22324 24686
rect 22284 24200 22336 24206
rect 22284 24142 22336 24148
rect 22848 24138 22876 24772
rect 22836 24132 22888 24138
rect 22756 24092 22836 24120
rect 22008 23656 22060 23662
rect 22008 23598 22060 23604
rect 22100 23520 22152 23526
rect 22100 23462 22152 23468
rect 21732 23180 21784 23186
rect 21732 23122 21784 23128
rect 22112 23118 22140 23462
rect 21640 23112 21692 23118
rect 21640 23054 21692 23060
rect 22100 23112 22152 23118
rect 22100 23054 22152 23060
rect 20996 23044 21048 23050
rect 20996 22986 21048 22992
rect 21364 23044 21416 23050
rect 21364 22986 21416 22992
rect 20536 21956 20588 21962
rect 20536 21898 20588 21904
rect 20352 21684 20404 21690
rect 20352 21626 20404 21632
rect 20168 20868 20220 20874
rect 20168 20810 20220 20816
rect 19800 20528 19852 20534
rect 19800 20470 19852 20476
rect 18512 19916 18564 19922
rect 18512 19858 18564 19864
rect 17960 19848 18012 19854
rect 17960 19790 18012 19796
rect 18236 19848 18288 19854
rect 18236 19790 18288 19796
rect 18420 19848 18472 19854
rect 18420 19790 18472 19796
rect 18052 19780 18104 19786
rect 18052 19722 18104 19728
rect 18064 19514 18092 19722
rect 18052 19508 18104 19514
rect 18052 19450 18104 19456
rect 18432 19446 18460 19790
rect 18420 19440 18472 19446
rect 18420 19382 18472 19388
rect 17040 19372 17092 19378
rect 17040 19314 17092 19320
rect 17960 19372 18012 19378
rect 17960 19314 18012 19320
rect 16488 19304 16540 19310
rect 16488 19246 16540 19252
rect 17500 19304 17552 19310
rect 17500 19246 17552 19252
rect 17512 18834 17540 19246
rect 17500 18828 17552 18834
rect 17500 18770 17552 18776
rect 16488 18760 16540 18766
rect 16488 18702 16540 18708
rect 16212 18624 16264 18630
rect 16212 18566 16264 18572
rect 16396 18624 16448 18630
rect 16396 18566 16448 18572
rect 15844 18352 15896 18358
rect 15844 18294 15896 18300
rect 15568 18216 15620 18222
rect 15568 18158 15620 18164
rect 15580 17882 15608 18158
rect 15568 17876 15620 17882
rect 15568 17818 15620 17824
rect 15856 17610 15884 18294
rect 16224 18290 16252 18566
rect 15936 18284 15988 18290
rect 15936 18226 15988 18232
rect 16212 18284 16264 18290
rect 16212 18226 16264 18232
rect 15948 17882 15976 18226
rect 15936 17876 15988 17882
rect 15936 17818 15988 17824
rect 15844 17604 15896 17610
rect 15764 17564 15844 17592
rect 15568 17536 15620 17542
rect 15488 17496 15568 17524
rect 15488 16998 15516 17496
rect 15568 17478 15620 17484
rect 15476 16992 15528 16998
rect 15476 16934 15528 16940
rect 15488 16794 15516 16934
rect 15476 16788 15528 16794
rect 15476 16730 15528 16736
rect 15160 16408 15240 16436
rect 15108 16390 15160 16396
rect 14188 16108 14240 16114
rect 14188 16050 14240 16056
rect 15016 16040 15068 16046
rect 15016 15982 15068 15988
rect 15028 15706 15056 15982
rect 13912 15700 13964 15706
rect 13912 15642 13964 15648
rect 15016 15700 15068 15706
rect 15016 15642 15068 15648
rect 14096 15632 14148 15638
rect 14096 15574 14148 15580
rect 13728 15428 13780 15434
rect 13728 15370 13780 15376
rect 14108 15094 14136 15574
rect 15212 15502 15240 16408
rect 15660 16040 15712 16046
rect 15660 15982 15712 15988
rect 15672 15502 15700 15982
rect 15764 15910 15792 17564
rect 15844 17546 15896 17552
rect 15844 17196 15896 17202
rect 15844 17138 15896 17144
rect 16028 17196 16080 17202
rect 16028 17138 16080 17144
rect 15752 15904 15804 15910
rect 15752 15846 15804 15852
rect 15200 15496 15252 15502
rect 15200 15438 15252 15444
rect 15384 15496 15436 15502
rect 15384 15438 15436 15444
rect 15660 15496 15712 15502
rect 15660 15438 15712 15444
rect 14096 15088 14148 15094
rect 14096 15030 14148 15036
rect 13820 14952 13872 14958
rect 13820 14894 13872 14900
rect 13832 14482 13860 14894
rect 13820 14476 13872 14482
rect 13820 14418 13872 14424
rect 13728 14340 13780 14346
rect 13728 14282 13780 14288
rect 13504 14232 13584 14260
rect 13452 14214 13504 14220
rect 13280 14062 13492 14090
rect 12624 14000 12676 14006
rect 12624 13942 12676 13948
rect 12808 14000 12860 14006
rect 12808 13942 12860 13948
rect 12900 13796 12952 13802
rect 12900 13738 12952 13744
rect 12912 12986 12940 13738
rect 13360 13728 13412 13734
rect 13360 13670 13412 13676
rect 12900 12980 12952 12986
rect 12900 12922 12952 12928
rect 12808 12640 12860 12646
rect 12808 12582 12860 12588
rect 12532 12436 12584 12442
rect 12532 12378 12584 12384
rect 12716 12368 12768 12374
rect 12716 12310 12768 12316
rect 12728 12238 12756 12310
rect 12820 12238 12848 12582
rect 12912 12442 12940 12922
rect 13084 12844 13136 12850
rect 13084 12786 13136 12792
rect 12900 12436 12952 12442
rect 13096 12434 13124 12786
rect 13268 12776 13320 12782
rect 13268 12718 13320 12724
rect 12900 12378 12952 12384
rect 13004 12406 13124 12434
rect 13176 12436 13228 12442
rect 13004 12288 13032 12406
rect 13176 12378 13228 12384
rect 13188 12322 13216 12378
rect 12912 12260 13032 12288
rect 13096 12294 13216 12322
rect 12716 12232 12768 12238
rect 12716 12174 12768 12180
rect 12808 12232 12860 12238
rect 12808 12174 12860 12180
rect 12532 11552 12584 11558
rect 12532 11494 12584 11500
rect 12544 11286 12572 11494
rect 12806 11384 12862 11393
rect 12624 11348 12676 11354
rect 12806 11319 12808 11328
rect 12624 11290 12676 11296
rect 12860 11319 12862 11328
rect 12808 11290 12860 11296
rect 12532 11280 12584 11286
rect 12532 11222 12584 11228
rect 12636 11234 12664 11290
rect 12636 11206 12756 11234
rect 12728 11150 12756 11206
rect 12808 11212 12860 11218
rect 12808 11154 12860 11160
rect 12716 11144 12768 11150
rect 12452 11082 12572 11098
rect 12716 11086 12768 11092
rect 12452 11076 12584 11082
rect 12452 11070 12532 11076
rect 12532 11018 12584 11024
rect 12820 10674 12848 11154
rect 12808 10668 12860 10674
rect 12808 10610 12860 10616
rect 12912 10538 12940 12260
rect 13096 12238 13124 12294
rect 13280 12238 13308 12718
rect 13372 12238 13400 13670
rect 13084 12232 13136 12238
rect 13084 12174 13136 12180
rect 13268 12232 13320 12238
rect 13268 12174 13320 12180
rect 13360 12232 13412 12238
rect 13360 12174 13412 12180
rect 12992 12096 13044 12102
rect 12992 12038 13044 12044
rect 13004 11762 13032 12038
rect 12992 11756 13044 11762
rect 12992 11698 13044 11704
rect 13096 11694 13124 12174
rect 13176 12164 13228 12170
rect 13176 12106 13228 12112
rect 13188 11762 13216 12106
rect 13176 11756 13228 11762
rect 13176 11698 13228 11704
rect 13268 11756 13320 11762
rect 13268 11698 13320 11704
rect 13084 11688 13136 11694
rect 13084 11630 13136 11636
rect 12992 11280 13044 11286
rect 13188 11268 13216 11698
rect 13280 11626 13308 11698
rect 13268 11620 13320 11626
rect 13268 11562 13320 11568
rect 13044 11240 13216 11268
rect 12992 11222 13044 11228
rect 13280 11218 13308 11562
rect 13372 11354 13400 12174
rect 13360 11348 13412 11354
rect 13360 11290 13412 11296
rect 13268 11212 13320 11218
rect 13268 11154 13320 11160
rect 13268 11076 13320 11082
rect 13268 11018 13320 11024
rect 13084 11008 13136 11014
rect 13084 10950 13136 10956
rect 13096 10810 13124 10950
rect 13084 10804 13136 10810
rect 13084 10746 13136 10752
rect 13280 10742 13308 11018
rect 13268 10736 13320 10742
rect 13268 10678 13320 10684
rect 12900 10532 12952 10538
rect 12900 10474 12952 10480
rect 12268 9846 12388 9874
rect 11888 9580 11940 9586
rect 11888 9522 11940 9528
rect 11900 8974 11928 9522
rect 11888 8968 11940 8974
rect 11888 8910 11940 8916
rect 11900 8430 11928 8910
rect 11888 8424 11940 8430
rect 11888 8366 11940 8372
rect 11612 7744 11664 7750
rect 11612 7686 11664 7692
rect 11624 7478 11652 7686
rect 11796 7540 11848 7546
rect 11796 7482 11848 7488
rect 11612 7472 11664 7478
rect 11612 7414 11664 7420
rect 11520 6928 11572 6934
rect 11520 6870 11572 6876
rect 11532 6798 11560 6870
rect 11520 6792 11572 6798
rect 11520 6734 11572 6740
rect 11244 6656 11296 6662
rect 11244 6598 11296 6604
rect 11532 6322 11560 6734
rect 11520 6316 11572 6322
rect 11520 6258 11572 6264
rect 11808 6186 11836 7482
rect 11900 6798 11928 8366
rect 12072 7472 12124 7478
rect 12072 7414 12124 7420
rect 11980 6996 12032 7002
rect 11980 6938 12032 6944
rect 11888 6792 11940 6798
rect 11888 6734 11940 6740
rect 11796 6180 11848 6186
rect 11796 6122 11848 6128
rect 11152 5636 11204 5642
rect 11152 5578 11204 5584
rect 11808 5302 11836 6122
rect 11796 5296 11848 5302
rect 11796 5238 11848 5244
rect 10692 5092 10744 5098
rect 10692 5034 10744 5040
rect 10704 4622 10732 5034
rect 11518 4720 11574 4729
rect 11518 4655 11574 4664
rect 10692 4616 10744 4622
rect 10692 4558 10744 4564
rect 10508 4548 10560 4554
rect 10508 4490 10560 4496
rect 10520 4146 10548 4490
rect 10704 4298 10732 4558
rect 10612 4270 10732 4298
rect 10612 4214 10640 4270
rect 10600 4208 10652 4214
rect 10600 4150 10652 4156
rect 10508 4140 10560 4146
rect 10508 4082 10560 4088
rect 11428 4140 11480 4146
rect 11428 4082 11480 4088
rect 10876 3936 10928 3942
rect 10876 3878 10928 3884
rect 10888 3602 10916 3878
rect 11440 3738 11468 4082
rect 11428 3732 11480 3738
rect 11428 3674 11480 3680
rect 10876 3596 10928 3602
rect 10876 3538 10928 3544
rect 11440 3534 11468 3674
rect 11532 3602 11560 4655
rect 11612 3732 11664 3738
rect 11612 3674 11664 3680
rect 11520 3596 11572 3602
rect 11520 3538 11572 3544
rect 11428 3528 11480 3534
rect 11428 3470 11480 3476
rect 10416 3460 10468 3466
rect 10416 3402 10468 3408
rect 10428 3126 10456 3402
rect 10508 3392 10560 3398
rect 10508 3334 10560 3340
rect 10520 3126 10548 3334
rect 11624 3194 11652 3674
rect 11796 3664 11848 3670
rect 11900 3618 11928 6734
rect 11992 6322 12020 6938
rect 11980 6316 12032 6322
rect 11980 6258 12032 6264
rect 11980 4480 12032 4486
rect 11980 4422 12032 4428
rect 11992 4214 12020 4422
rect 12084 4282 12112 7414
rect 12164 6996 12216 7002
rect 12164 6938 12216 6944
rect 12176 6458 12204 6938
rect 12164 6452 12216 6458
rect 12164 6394 12216 6400
rect 12268 5166 12296 9846
rect 13084 9512 13136 9518
rect 13084 9454 13136 9460
rect 13096 9382 13124 9454
rect 12348 9376 12400 9382
rect 12348 9318 12400 9324
rect 13084 9376 13136 9382
rect 13084 9318 13136 9324
rect 12360 9042 12388 9318
rect 12348 9036 12400 9042
rect 12348 8978 12400 8984
rect 12808 8900 12860 8906
rect 12808 8842 12860 8848
rect 12820 8566 12848 8842
rect 12808 8560 12860 8566
rect 12636 8520 12808 8548
rect 12440 7404 12492 7410
rect 12440 7346 12492 7352
rect 12348 7336 12400 7342
rect 12348 7278 12400 7284
rect 12360 7002 12388 7278
rect 12348 6996 12400 7002
rect 12348 6938 12400 6944
rect 12360 5370 12388 6938
rect 12452 6662 12480 7346
rect 12532 7200 12584 7206
rect 12532 7142 12584 7148
rect 12544 6866 12572 7142
rect 12532 6860 12584 6866
rect 12532 6802 12584 6808
rect 12440 6656 12492 6662
rect 12440 6598 12492 6604
rect 12544 6254 12572 6802
rect 12636 6730 12664 8520
rect 12808 8502 12860 8508
rect 12808 7880 12860 7886
rect 12808 7822 12860 7828
rect 12716 7336 12768 7342
rect 12716 7278 12768 7284
rect 12624 6724 12676 6730
rect 12624 6666 12676 6672
rect 12532 6248 12584 6254
rect 12532 6190 12584 6196
rect 12636 6100 12664 6666
rect 12728 6458 12756 7278
rect 12820 6458 12848 7822
rect 12992 7336 13044 7342
rect 12992 7278 13044 7284
rect 12716 6452 12768 6458
rect 12716 6394 12768 6400
rect 12808 6452 12860 6458
rect 12808 6394 12860 6400
rect 12716 6316 12768 6322
rect 12716 6258 12768 6264
rect 12544 6072 12664 6100
rect 12348 5364 12400 5370
rect 12348 5306 12400 5312
rect 12256 5160 12308 5166
rect 12256 5102 12308 5108
rect 12164 4616 12216 4622
rect 12162 4584 12164 4593
rect 12216 4584 12218 4593
rect 12162 4519 12218 4528
rect 12360 4282 12388 5306
rect 12440 5296 12492 5302
rect 12440 5238 12492 5244
rect 12452 4690 12480 5238
rect 12440 4684 12492 4690
rect 12440 4626 12492 4632
rect 12072 4276 12124 4282
rect 12072 4218 12124 4224
rect 12348 4276 12400 4282
rect 12348 4218 12400 4224
rect 11980 4208 12032 4214
rect 11980 4150 12032 4156
rect 11980 4072 12032 4078
rect 11978 4040 11980 4049
rect 12348 4072 12400 4078
rect 12032 4040 12034 4049
rect 12348 4014 12400 4020
rect 11978 3975 12034 3984
rect 12360 3777 12388 4014
rect 12346 3768 12402 3777
rect 12346 3703 12402 3712
rect 11848 3612 12020 3618
rect 11796 3606 12020 3612
rect 11808 3602 12020 3606
rect 11808 3596 12032 3602
rect 11808 3590 11980 3596
rect 12544 3584 12572 6072
rect 12728 5234 12756 6258
rect 13004 5953 13032 7278
rect 13464 6390 13492 14062
rect 13556 13938 13584 14232
rect 13544 13932 13596 13938
rect 13544 13874 13596 13880
rect 13556 12782 13584 13874
rect 13740 13870 13768 14282
rect 13832 13938 13860 14418
rect 13820 13932 13872 13938
rect 13820 13874 13872 13880
rect 13728 13864 13780 13870
rect 13728 13806 13780 13812
rect 13740 12986 13768 13806
rect 13728 12980 13780 12986
rect 13728 12922 13780 12928
rect 13544 12776 13596 12782
rect 13544 12718 13596 12724
rect 13740 12628 13768 12922
rect 13832 12850 13860 13874
rect 15212 13326 15240 15438
rect 15290 14376 15346 14385
rect 15290 14311 15292 14320
rect 15344 14311 15346 14320
rect 15292 14282 15344 14288
rect 15200 13320 15252 13326
rect 15200 13262 15252 13268
rect 14464 13252 14516 13258
rect 14464 13194 14516 13200
rect 13820 12844 13872 12850
rect 13820 12786 13872 12792
rect 13648 12600 13768 12628
rect 13648 12434 13676 12600
rect 13556 12406 13676 12434
rect 13726 12472 13782 12481
rect 13726 12407 13782 12416
rect 13556 12102 13584 12406
rect 13636 12368 13688 12374
rect 13740 12322 13768 12407
rect 13688 12316 13768 12322
rect 13636 12310 13768 12316
rect 13648 12294 13768 12310
rect 13544 12096 13596 12102
rect 13544 12038 13596 12044
rect 13636 11892 13688 11898
rect 13636 11834 13688 11840
rect 13544 11552 13596 11558
rect 13544 11494 13596 11500
rect 13556 10606 13584 11494
rect 13648 11354 13676 11834
rect 13832 11830 13860 12786
rect 14096 12776 14148 12782
rect 14096 12718 14148 12724
rect 14108 12442 14136 12718
rect 14096 12436 14148 12442
rect 14096 12378 14148 12384
rect 14476 12238 14504 13194
rect 15396 12986 15424 15438
rect 15764 15434 15792 15846
rect 15856 15638 15884 17138
rect 16040 16454 16068 17138
rect 16212 16788 16264 16794
rect 16212 16730 16264 16736
rect 16028 16448 16080 16454
rect 16028 16390 16080 16396
rect 16040 16250 16068 16390
rect 16028 16244 16080 16250
rect 16028 16186 16080 16192
rect 16224 15706 16252 16730
rect 16304 16176 16356 16182
rect 16304 16118 16356 16124
rect 16212 15700 16264 15706
rect 16212 15642 16264 15648
rect 15844 15632 15896 15638
rect 15844 15574 15896 15580
rect 16224 15570 16252 15642
rect 16212 15564 16264 15570
rect 16212 15506 16264 15512
rect 15936 15496 15988 15502
rect 15936 15438 15988 15444
rect 15476 15428 15528 15434
rect 15476 15370 15528 15376
rect 15752 15428 15804 15434
rect 15752 15370 15804 15376
rect 15488 13326 15516 15370
rect 15660 14816 15712 14822
rect 15660 14758 15712 14764
rect 15672 13870 15700 14758
rect 15660 13864 15712 13870
rect 15660 13806 15712 13812
rect 15660 13388 15712 13394
rect 15660 13330 15712 13336
rect 15476 13320 15528 13326
rect 15476 13262 15528 13268
rect 15384 12980 15436 12986
rect 15384 12922 15436 12928
rect 14556 12776 14608 12782
rect 14556 12718 14608 12724
rect 14568 12238 14596 12718
rect 15396 12238 15424 12922
rect 15488 12918 15516 13262
rect 15476 12912 15528 12918
rect 15476 12854 15528 12860
rect 15488 12481 15516 12854
rect 15672 12850 15700 13330
rect 15764 13190 15792 15370
rect 15844 15020 15896 15026
rect 15844 14962 15896 14968
rect 15752 13184 15804 13190
rect 15752 13126 15804 13132
rect 15764 12866 15792 13126
rect 15856 12986 15884 14962
rect 15948 13530 15976 15438
rect 16224 15026 16252 15506
rect 16212 15020 16264 15026
rect 16212 14962 16264 14968
rect 16316 14006 16344 16118
rect 16408 14278 16436 18566
rect 16500 17542 16528 18702
rect 16948 18624 17000 18630
rect 16948 18566 17000 18572
rect 16960 18426 16988 18566
rect 16948 18420 17000 18426
rect 16948 18362 17000 18368
rect 17316 18352 17368 18358
rect 17316 18294 17368 18300
rect 16488 17536 16540 17542
rect 16488 17478 16540 17484
rect 16500 16522 16528 17478
rect 17328 16998 17356 18294
rect 17512 18170 17540 18770
rect 17972 18766 18000 19314
rect 18052 19168 18104 19174
rect 18052 19110 18104 19116
rect 17960 18760 18012 18766
rect 17960 18702 18012 18708
rect 17420 18142 17540 18170
rect 17420 18086 17448 18142
rect 17408 18080 17460 18086
rect 17408 18022 17460 18028
rect 17500 18080 17552 18086
rect 17500 18022 17552 18028
rect 17408 17604 17460 17610
rect 17408 17546 17460 17552
rect 17420 17338 17448 17546
rect 17408 17332 17460 17338
rect 17408 17274 17460 17280
rect 17512 17202 17540 18022
rect 17868 17740 17920 17746
rect 17868 17682 17920 17688
rect 17500 17196 17552 17202
rect 17500 17138 17552 17144
rect 17316 16992 17368 16998
rect 17316 16934 17368 16940
rect 16488 16516 16540 16522
rect 16488 16458 16540 16464
rect 16500 16182 16528 16458
rect 16488 16176 16540 16182
rect 16488 16118 16540 16124
rect 17880 16114 17908 17682
rect 18064 16590 18092 19110
rect 18236 18964 18288 18970
rect 18288 18924 18368 18952
rect 18236 18906 18288 18912
rect 18144 18624 18196 18630
rect 18144 18566 18196 18572
rect 18156 18290 18184 18566
rect 18144 18284 18196 18290
rect 18144 18226 18196 18232
rect 18156 17202 18184 18226
rect 18144 17196 18196 17202
rect 18144 17138 18196 17144
rect 18052 16584 18104 16590
rect 18052 16526 18104 16532
rect 17868 16108 17920 16114
rect 17868 16050 17920 16056
rect 16672 15904 16724 15910
rect 16672 15846 16724 15852
rect 16684 15570 16712 15846
rect 16672 15564 16724 15570
rect 16672 15506 16724 15512
rect 17880 15162 17908 16050
rect 18236 16040 18288 16046
rect 18236 15982 18288 15988
rect 18248 15706 18276 15982
rect 18236 15700 18288 15706
rect 18236 15642 18288 15648
rect 18340 15434 18368 18924
rect 18524 17610 18552 19858
rect 18604 19780 18656 19786
rect 18604 19722 18656 19728
rect 18616 19514 18644 19722
rect 18696 19712 18748 19718
rect 18696 19654 18748 19660
rect 18604 19508 18656 19514
rect 18604 19450 18656 19456
rect 18708 19378 18736 19654
rect 18892 19514 18920 20334
rect 19352 20330 19472 20346
rect 19352 20324 19484 20330
rect 19352 20318 19432 20324
rect 19248 19848 19300 19854
rect 19248 19790 19300 19796
rect 19260 19514 19288 19790
rect 18880 19508 18932 19514
rect 18880 19450 18932 19456
rect 19248 19508 19300 19514
rect 19248 19450 19300 19456
rect 18604 19372 18656 19378
rect 18604 19314 18656 19320
rect 18696 19372 18748 19378
rect 18696 19314 18748 19320
rect 18616 18970 18644 19314
rect 18604 18964 18656 18970
rect 18604 18906 18656 18912
rect 18604 18828 18656 18834
rect 18604 18770 18656 18776
rect 18616 17882 18644 18770
rect 19352 18698 19380 20318
rect 19432 20266 19484 20272
rect 20180 20058 20208 20810
rect 20548 20466 20576 21898
rect 21008 21894 21036 22986
rect 22112 22710 22140 23054
rect 22100 22704 22152 22710
rect 22100 22646 22152 22652
rect 22376 22568 22428 22574
rect 22376 22510 22428 22516
rect 21824 22432 21876 22438
rect 21824 22374 21876 22380
rect 21836 22234 21864 22374
rect 21824 22228 21876 22234
rect 21824 22170 21876 22176
rect 20996 21888 21048 21894
rect 20996 21830 21048 21836
rect 21008 21690 21036 21830
rect 22388 21690 22416 22510
rect 22756 21894 22784 24092
rect 22836 24074 22888 24080
rect 22940 23798 22968 25230
rect 23020 25152 23072 25158
rect 23020 25094 23072 25100
rect 23032 24818 23060 25094
rect 23308 24954 23336 25774
rect 23756 25356 23808 25362
rect 23756 25298 23808 25304
rect 23768 24954 23796 25298
rect 23296 24948 23348 24954
rect 23296 24890 23348 24896
rect 23756 24948 23808 24954
rect 23756 24890 23808 24896
rect 23020 24812 23072 24818
rect 23020 24754 23072 24760
rect 24044 24274 24072 25774
rect 24320 25498 24348 25774
rect 25780 25696 25832 25702
rect 25780 25638 25832 25644
rect 24308 25492 24360 25498
rect 24308 25434 24360 25440
rect 24860 25356 24912 25362
rect 24860 25298 24912 25304
rect 24872 24818 24900 25298
rect 25136 25152 25188 25158
rect 25136 25094 25188 25100
rect 25148 24818 25176 25094
rect 25688 24880 25740 24886
rect 25688 24822 25740 24828
rect 24860 24812 24912 24818
rect 24860 24754 24912 24760
rect 25136 24812 25188 24818
rect 25136 24754 25188 24760
rect 24032 24268 24084 24274
rect 24032 24210 24084 24216
rect 22928 23792 22980 23798
rect 22928 23734 22980 23740
rect 22836 23112 22888 23118
rect 22836 23054 22888 23060
rect 22848 22506 22876 23054
rect 23940 22976 23992 22982
rect 23940 22918 23992 22924
rect 23952 22642 23980 22918
rect 23940 22636 23992 22642
rect 23940 22578 23992 22584
rect 23480 22568 23532 22574
rect 23480 22510 23532 22516
rect 22836 22500 22888 22506
rect 22836 22442 22888 22448
rect 22848 22234 22876 22442
rect 23020 22432 23072 22438
rect 23020 22374 23072 22380
rect 22836 22228 22888 22234
rect 22836 22170 22888 22176
rect 22744 21888 22796 21894
rect 22744 21830 22796 21836
rect 22848 21706 22876 22170
rect 20996 21684 21048 21690
rect 20996 21626 21048 21632
rect 22376 21684 22428 21690
rect 22376 21626 22428 21632
rect 22664 21678 22876 21706
rect 22664 21622 22692 21678
rect 23032 21622 23060 22374
rect 23492 21894 23520 22510
rect 24044 22098 24072 24210
rect 24584 22704 24636 22710
rect 24584 22646 24636 22652
rect 24032 22092 24084 22098
rect 24032 22034 24084 22040
rect 23112 21888 23164 21894
rect 23112 21830 23164 21836
rect 23480 21888 23532 21894
rect 23480 21830 23532 21836
rect 23664 21888 23716 21894
rect 23664 21830 23716 21836
rect 22652 21616 22704 21622
rect 22652 21558 22704 21564
rect 23020 21616 23072 21622
rect 23020 21558 23072 21564
rect 22192 21548 22244 21554
rect 22192 21490 22244 21496
rect 21456 21480 21508 21486
rect 21456 21422 21508 21428
rect 20628 20868 20680 20874
rect 20628 20810 20680 20816
rect 20640 20534 20668 20810
rect 21468 20602 21496 21422
rect 21640 20800 21692 20806
rect 21640 20742 21692 20748
rect 21456 20596 21508 20602
rect 21456 20538 21508 20544
rect 20628 20528 20680 20534
rect 20628 20470 20680 20476
rect 21652 20466 21680 20742
rect 22204 20602 22232 21490
rect 22744 21480 22796 21486
rect 22744 21422 22796 21428
rect 22756 21010 22784 21422
rect 22744 21004 22796 21010
rect 22744 20946 22796 20952
rect 23124 20942 23152 21830
rect 23676 21146 23704 21830
rect 24044 21690 24072 22034
rect 24216 22024 24268 22030
rect 24216 21966 24268 21972
rect 24032 21684 24084 21690
rect 24032 21626 24084 21632
rect 23664 21140 23716 21146
rect 23664 21082 23716 21088
rect 24044 21010 24072 21626
rect 24228 21486 24256 21966
rect 24596 21962 24624 22646
rect 24872 22624 24900 24754
rect 25596 24268 25648 24274
rect 25596 24210 25648 24216
rect 25608 23866 25636 24210
rect 25596 23860 25648 23866
rect 25596 23802 25648 23808
rect 25700 23730 25728 24822
rect 25792 24614 25820 25638
rect 26148 25288 26200 25294
rect 26148 25230 26200 25236
rect 26332 25288 26384 25294
rect 26332 25230 26384 25236
rect 27160 25288 27212 25294
rect 27160 25230 27212 25236
rect 26160 24834 26188 25230
rect 26160 24806 26280 24834
rect 25780 24608 25832 24614
rect 25780 24550 25832 24556
rect 26252 24342 26280 24806
rect 26344 24682 26372 25230
rect 27172 24954 27200 25230
rect 27804 25152 27856 25158
rect 27804 25094 27856 25100
rect 26424 24948 26476 24954
rect 26424 24890 26476 24896
rect 27160 24948 27212 24954
rect 27160 24890 27212 24896
rect 26332 24676 26384 24682
rect 26332 24618 26384 24624
rect 26240 24336 26292 24342
rect 26240 24278 26292 24284
rect 26436 24206 26464 24890
rect 26976 24812 27028 24818
rect 26976 24754 27028 24760
rect 27160 24812 27212 24818
rect 27160 24754 27212 24760
rect 26792 24608 26844 24614
rect 26792 24550 26844 24556
rect 26804 24274 26832 24550
rect 26988 24410 27016 24754
rect 26976 24404 27028 24410
rect 26976 24346 27028 24352
rect 26516 24268 26568 24274
rect 26516 24210 26568 24216
rect 26792 24268 26844 24274
rect 26792 24210 26844 24216
rect 25872 24200 25924 24206
rect 26424 24200 26476 24206
rect 25872 24142 25924 24148
rect 26344 24160 26424 24188
rect 25884 23866 25912 24142
rect 26148 24064 26200 24070
rect 26344 24018 26372 24160
rect 26424 24142 26476 24148
rect 26200 24012 26372 24018
rect 26148 24006 26372 24012
rect 26424 24064 26476 24070
rect 26424 24006 26476 24012
rect 26160 23990 26372 24006
rect 25872 23860 25924 23866
rect 25872 23802 25924 23808
rect 26344 23798 26372 23990
rect 26332 23792 26384 23798
rect 26332 23734 26384 23740
rect 26436 23730 26464 24006
rect 25688 23724 25740 23730
rect 25688 23666 25740 23672
rect 26424 23724 26476 23730
rect 26424 23666 26476 23672
rect 25044 23520 25096 23526
rect 25044 23462 25096 23468
rect 24952 22636 25004 22642
rect 24872 22596 24952 22624
rect 24872 22438 24900 22596
rect 24952 22578 25004 22584
rect 25056 22574 25084 23462
rect 26436 23118 26464 23666
rect 26528 23186 26556 24210
rect 27172 23730 27200 24754
rect 27816 24138 27844 25094
rect 27896 24812 27948 24818
rect 27896 24754 27948 24760
rect 27804 24132 27856 24138
rect 27804 24074 27856 24080
rect 27160 23724 27212 23730
rect 27160 23666 27212 23672
rect 26884 23588 26936 23594
rect 26884 23530 26936 23536
rect 26896 23186 26924 23530
rect 26516 23180 26568 23186
rect 26516 23122 26568 23128
rect 26884 23180 26936 23186
rect 26884 23122 26936 23128
rect 26424 23112 26476 23118
rect 26424 23054 26476 23060
rect 26332 22976 26384 22982
rect 26332 22918 26384 22924
rect 25228 22636 25280 22642
rect 25228 22578 25280 22584
rect 25044 22568 25096 22574
rect 25044 22510 25096 22516
rect 24860 22432 24912 22438
rect 24860 22374 24912 22380
rect 24584 21956 24636 21962
rect 24584 21898 24636 21904
rect 24596 21690 24624 21898
rect 24584 21684 24636 21690
rect 24584 21626 24636 21632
rect 25056 21622 25084 22510
rect 25240 21894 25268 22578
rect 26344 22574 26372 22918
rect 26424 22636 26476 22642
rect 26424 22578 26476 22584
rect 25596 22568 25648 22574
rect 25596 22510 25648 22516
rect 26332 22568 26384 22574
rect 26332 22510 26384 22516
rect 25504 21956 25556 21962
rect 25504 21898 25556 21904
rect 25228 21888 25280 21894
rect 25228 21830 25280 21836
rect 25044 21616 25096 21622
rect 25044 21558 25096 21564
rect 25240 21486 25268 21830
rect 25516 21690 25544 21898
rect 25608 21690 25636 22510
rect 26148 22432 26200 22438
rect 26148 22374 26200 22380
rect 26160 22234 26188 22374
rect 26148 22228 26200 22234
rect 26148 22170 26200 22176
rect 26436 21690 26464 22578
rect 26528 21962 26556 23122
rect 27816 23050 27844 24074
rect 27908 23662 27936 24754
rect 27988 24608 28040 24614
rect 27988 24550 28040 24556
rect 28000 23798 28028 24550
rect 27988 23792 28040 23798
rect 27988 23734 28040 23740
rect 27896 23656 27948 23662
rect 27896 23598 27948 23604
rect 27908 23322 27936 23598
rect 27896 23316 27948 23322
rect 27896 23258 27948 23264
rect 27804 23044 27856 23050
rect 27804 22986 27856 22992
rect 27436 22568 27488 22574
rect 27436 22510 27488 22516
rect 27620 22568 27672 22574
rect 27620 22510 27672 22516
rect 26608 22500 26660 22506
rect 26608 22442 26660 22448
rect 26516 21956 26568 21962
rect 26516 21898 26568 21904
rect 25504 21684 25556 21690
rect 25504 21626 25556 21632
rect 25596 21684 25648 21690
rect 25596 21626 25648 21632
rect 26424 21684 26476 21690
rect 26424 21626 26476 21632
rect 24216 21480 24268 21486
rect 24216 21422 24268 21428
rect 25228 21480 25280 21486
rect 25228 21422 25280 21428
rect 24032 21004 24084 21010
rect 24032 20946 24084 20952
rect 24768 21004 24820 21010
rect 24768 20946 24820 20952
rect 23112 20936 23164 20942
rect 23112 20878 23164 20884
rect 22284 20868 22336 20874
rect 22284 20810 22336 20816
rect 24400 20868 24452 20874
rect 24400 20810 24452 20816
rect 22192 20596 22244 20602
rect 22192 20538 22244 20544
rect 20536 20460 20588 20466
rect 20536 20402 20588 20408
rect 21456 20460 21508 20466
rect 21456 20402 21508 20408
rect 21640 20460 21692 20466
rect 21640 20402 21692 20408
rect 20168 20052 20220 20058
rect 20168 19994 20220 20000
rect 20536 19916 20588 19922
rect 20536 19858 20588 19864
rect 19432 19848 19484 19854
rect 19432 19790 19484 19796
rect 19708 19848 19760 19854
rect 19708 19790 19760 19796
rect 19444 18902 19472 19790
rect 19720 19417 19748 19790
rect 19706 19408 19762 19417
rect 19706 19343 19708 19352
rect 19760 19343 19762 19352
rect 20444 19372 20496 19378
rect 19708 19314 19760 19320
rect 20444 19314 20496 19320
rect 19432 18896 19484 18902
rect 19432 18838 19484 18844
rect 20456 18834 20484 19314
rect 20444 18828 20496 18834
rect 20444 18770 20496 18776
rect 19340 18692 19392 18698
rect 19340 18634 19392 18640
rect 19156 18420 19208 18426
rect 19156 18362 19208 18368
rect 19064 18284 19116 18290
rect 19064 18226 19116 18232
rect 18604 17876 18656 17882
rect 18604 17818 18656 17824
rect 18512 17604 18564 17610
rect 18512 17546 18564 17552
rect 18524 17354 18552 17546
rect 18432 17338 18552 17354
rect 18432 17332 18564 17338
rect 18432 17326 18512 17332
rect 18328 15428 18380 15434
rect 18328 15370 18380 15376
rect 17868 15156 17920 15162
rect 17868 15098 17920 15104
rect 17880 15026 17908 15098
rect 16488 15020 16540 15026
rect 16488 14962 16540 14968
rect 17868 15020 17920 15026
rect 17868 14962 17920 14968
rect 16396 14272 16448 14278
rect 16396 14214 16448 14220
rect 16304 14000 16356 14006
rect 16304 13942 16356 13948
rect 15936 13524 15988 13530
rect 15936 13466 15988 13472
rect 15844 12980 15896 12986
rect 15844 12922 15896 12928
rect 15764 12850 15884 12866
rect 15660 12844 15712 12850
rect 15764 12844 15896 12850
rect 15764 12838 15844 12844
rect 15660 12786 15712 12792
rect 15844 12786 15896 12792
rect 15474 12472 15530 12481
rect 15474 12407 15530 12416
rect 15672 12306 15700 12786
rect 15660 12300 15712 12306
rect 15660 12242 15712 12248
rect 14280 12232 14332 12238
rect 14280 12174 14332 12180
rect 14464 12232 14516 12238
rect 14464 12174 14516 12180
rect 14556 12232 14608 12238
rect 14556 12174 14608 12180
rect 15384 12232 15436 12238
rect 15384 12174 15436 12180
rect 13820 11824 13872 11830
rect 13820 11766 13872 11772
rect 13728 11688 13780 11694
rect 13728 11630 13780 11636
rect 13636 11348 13688 11354
rect 13636 11290 13688 11296
rect 13544 10600 13596 10606
rect 13544 10542 13596 10548
rect 13648 10062 13676 11290
rect 13636 10056 13688 10062
rect 13636 9998 13688 10004
rect 13636 7404 13688 7410
rect 13636 7346 13688 7352
rect 13648 6662 13676 7346
rect 13636 6656 13688 6662
rect 13636 6598 13688 6604
rect 13452 6384 13504 6390
rect 13452 6326 13504 6332
rect 13648 6322 13676 6598
rect 13636 6316 13688 6322
rect 13636 6258 13688 6264
rect 13740 6118 13768 11630
rect 14004 11144 14056 11150
rect 14004 11086 14056 11092
rect 13820 11076 13872 11082
rect 13820 11018 13872 11024
rect 13832 9518 13860 11018
rect 13912 11008 13964 11014
rect 13912 10950 13964 10956
rect 13820 9512 13872 9518
rect 13820 9454 13872 9460
rect 13924 6322 13952 10950
rect 14016 10266 14044 11086
rect 14096 11008 14148 11014
rect 14096 10950 14148 10956
rect 14108 10606 14136 10950
rect 14096 10600 14148 10606
rect 14096 10542 14148 10548
rect 14292 10538 14320 12174
rect 14372 11756 14424 11762
rect 14372 11698 14424 11704
rect 14384 11286 14412 11698
rect 14372 11280 14424 11286
rect 14372 11222 14424 11228
rect 14384 11150 14412 11222
rect 14372 11144 14424 11150
rect 14372 11086 14424 11092
rect 14280 10532 14332 10538
rect 14280 10474 14332 10480
rect 14004 10260 14056 10266
rect 14004 10202 14056 10208
rect 14016 9654 14044 10202
rect 14188 10124 14240 10130
rect 14188 10066 14240 10072
rect 14004 9648 14056 9654
rect 14004 9590 14056 9596
rect 14200 9586 14228 10066
rect 14292 10062 14320 10474
rect 14568 10130 14596 12174
rect 14740 12164 14792 12170
rect 14740 12106 14792 12112
rect 14648 11144 14700 11150
rect 14752 11132 14780 12106
rect 15200 11620 15252 11626
rect 15200 11562 15252 11568
rect 14700 11104 14780 11132
rect 14648 11086 14700 11092
rect 14660 11014 14688 11086
rect 15212 11082 15240 11562
rect 15292 11280 15344 11286
rect 15292 11222 15344 11228
rect 15304 11098 15332 11222
rect 15396 11218 15424 12174
rect 15476 12096 15528 12102
rect 15476 12038 15528 12044
rect 15384 11212 15436 11218
rect 15384 11154 15436 11160
rect 15200 11076 15252 11082
rect 15304 11070 15424 11098
rect 15200 11018 15252 11024
rect 14648 11008 14700 11014
rect 14648 10950 14700 10956
rect 14648 10668 14700 10674
rect 14648 10610 14700 10616
rect 14556 10124 14608 10130
rect 14556 10066 14608 10072
rect 14280 10056 14332 10062
rect 14280 9998 14332 10004
rect 14292 9586 14320 9998
rect 14464 9920 14516 9926
rect 14464 9862 14516 9868
rect 14188 9580 14240 9586
rect 14188 9522 14240 9528
rect 14280 9580 14332 9586
rect 14280 9522 14332 9528
rect 14096 9512 14148 9518
rect 14096 9454 14148 9460
rect 14108 8838 14136 9454
rect 14096 8832 14148 8838
rect 14096 8774 14148 8780
rect 14200 8566 14228 9522
rect 14188 8560 14240 8566
rect 14188 8502 14240 8508
rect 14200 8430 14228 8502
rect 14188 8424 14240 8430
rect 14188 8366 14240 8372
rect 13912 6316 13964 6322
rect 13912 6258 13964 6264
rect 13084 6112 13136 6118
rect 13084 6054 13136 6060
rect 13728 6112 13780 6118
rect 13728 6054 13780 6060
rect 12990 5944 13046 5953
rect 12990 5879 13046 5888
rect 13004 5234 13032 5879
rect 13096 5574 13124 6054
rect 13084 5568 13136 5574
rect 13084 5510 13136 5516
rect 12716 5228 12768 5234
rect 12716 5170 12768 5176
rect 12992 5228 13044 5234
rect 12992 5170 13044 5176
rect 12624 4752 12676 4758
rect 12624 4694 12676 4700
rect 12636 4622 12664 4694
rect 12624 4616 12676 4622
rect 12624 4558 12676 4564
rect 12728 3942 12756 5170
rect 12992 5024 13044 5030
rect 12992 4966 13044 4972
rect 13004 4690 13032 4966
rect 12992 4684 13044 4690
rect 12992 4626 13044 4632
rect 12808 4616 12860 4622
rect 12808 4558 12860 4564
rect 12900 4616 12952 4622
rect 12900 4558 12952 4564
rect 12716 3936 12768 3942
rect 12716 3878 12768 3884
rect 12624 3596 12676 3602
rect 12544 3556 12624 3584
rect 11980 3538 12032 3544
rect 12624 3538 12676 3544
rect 12256 3460 12308 3466
rect 12256 3402 12308 3408
rect 12268 3194 12296 3402
rect 11612 3188 11664 3194
rect 11612 3130 11664 3136
rect 12256 3188 12308 3194
rect 12256 3130 12308 3136
rect 10416 3120 10468 3126
rect 10416 3062 10468 3068
rect 10508 3120 10560 3126
rect 10508 3062 10560 3068
rect 12820 2990 12848 4558
rect 12912 4026 12940 4558
rect 12992 4480 13044 4486
rect 12992 4422 13044 4428
rect 13004 4214 13032 4422
rect 12992 4208 13044 4214
rect 12992 4150 13044 4156
rect 12912 3998 13032 4026
rect 12900 3936 12952 3942
rect 12900 3878 12952 3884
rect 12912 3194 12940 3878
rect 13004 3398 13032 3998
rect 12992 3392 13044 3398
rect 12992 3334 13044 3340
rect 12900 3188 12952 3194
rect 12900 3130 12952 3136
rect 13096 2990 13124 5510
rect 13176 5296 13228 5302
rect 13176 5238 13228 5244
rect 13188 4622 13216 5238
rect 13912 4820 13964 4826
rect 13912 4762 13964 4768
rect 13176 4616 13228 4622
rect 13452 4616 13504 4622
rect 13176 4558 13228 4564
rect 13358 4584 13414 4593
rect 13452 4558 13504 4564
rect 13636 4616 13688 4622
rect 13636 4558 13688 4564
rect 13728 4616 13780 4622
rect 13728 4558 13780 4564
rect 13358 4519 13360 4528
rect 13412 4519 13414 4528
rect 13360 4490 13412 4496
rect 13372 4214 13400 4490
rect 13360 4208 13412 4214
rect 13360 4150 13412 4156
rect 13358 4040 13414 4049
rect 13358 3975 13360 3984
rect 13412 3975 13414 3984
rect 13360 3946 13412 3952
rect 13360 3528 13412 3534
rect 13360 3470 13412 3476
rect 13372 3194 13400 3470
rect 13360 3188 13412 3194
rect 13360 3130 13412 3136
rect 7012 2984 7064 2990
rect 7012 2926 7064 2932
rect 9864 2984 9916 2990
rect 9864 2926 9916 2932
rect 12808 2984 12860 2990
rect 12808 2926 12860 2932
rect 13084 2984 13136 2990
rect 13084 2926 13136 2932
rect 13464 2922 13492 4558
rect 13544 4072 13596 4078
rect 13544 4014 13596 4020
rect 13556 3398 13584 4014
rect 13648 4010 13676 4558
rect 13740 4282 13768 4558
rect 13820 4480 13872 4486
rect 13820 4422 13872 4428
rect 13728 4276 13780 4282
rect 13728 4218 13780 4224
rect 13636 4004 13688 4010
rect 13636 3946 13688 3952
rect 13740 3777 13768 4218
rect 13832 4146 13860 4422
rect 13924 4146 13952 4762
rect 13820 4140 13872 4146
rect 13820 4082 13872 4088
rect 13912 4140 13964 4146
rect 13912 4082 13964 4088
rect 13726 3768 13782 3777
rect 13726 3703 13728 3712
rect 13780 3703 13782 3712
rect 13728 3674 13780 3680
rect 13544 3392 13596 3398
rect 13544 3334 13596 3340
rect 14096 3392 14148 3398
rect 14096 3334 14148 3340
rect 14108 3126 14136 3334
rect 14476 3233 14504 9862
rect 14556 9376 14608 9382
rect 14556 9318 14608 9324
rect 14568 8634 14596 9318
rect 14660 9178 14688 10610
rect 14648 9172 14700 9178
rect 14648 9114 14700 9120
rect 14832 8968 14884 8974
rect 14832 8910 14884 8916
rect 15016 8968 15068 8974
rect 15016 8910 15068 8916
rect 14556 8628 14608 8634
rect 14556 8570 14608 8576
rect 14844 8090 14872 8910
rect 15028 8634 15056 8910
rect 15292 8900 15344 8906
rect 15292 8842 15344 8848
rect 15108 8832 15160 8838
rect 15108 8774 15160 8780
rect 15200 8832 15252 8838
rect 15200 8774 15252 8780
rect 15016 8628 15068 8634
rect 15016 8570 15068 8576
rect 14924 8492 14976 8498
rect 14976 8452 15056 8480
rect 14924 8434 14976 8440
rect 14924 8288 14976 8294
rect 14924 8230 14976 8236
rect 14832 8084 14884 8090
rect 14832 8026 14884 8032
rect 14936 7886 14964 8230
rect 14924 7880 14976 7886
rect 14924 7822 14976 7828
rect 15028 7478 15056 8452
rect 15120 7886 15148 8774
rect 15108 7880 15160 7886
rect 15108 7822 15160 7828
rect 15212 7818 15240 8774
rect 15304 8498 15332 8842
rect 15292 8492 15344 8498
rect 15292 8434 15344 8440
rect 15200 7812 15252 7818
rect 15200 7754 15252 7760
rect 15016 7472 15068 7478
rect 15016 7414 15068 7420
rect 14924 6384 14976 6390
rect 14924 6326 14976 6332
rect 14740 6316 14792 6322
rect 14740 6258 14792 6264
rect 14752 5846 14780 6258
rect 14740 5840 14792 5846
rect 14740 5782 14792 5788
rect 14936 5710 14964 6326
rect 15396 6254 15424 11070
rect 15488 10674 15516 12038
rect 16408 11354 16436 14214
rect 16500 14074 16528 14962
rect 18236 14952 18288 14958
rect 18236 14894 18288 14900
rect 18248 14618 18276 14894
rect 18236 14612 18288 14618
rect 18236 14554 18288 14560
rect 18144 14408 18196 14414
rect 18144 14350 18196 14356
rect 16488 14068 16540 14074
rect 16488 14010 16540 14016
rect 16500 13462 16528 14010
rect 17684 13932 17736 13938
rect 17684 13874 17736 13880
rect 16580 13864 16632 13870
rect 16580 13806 16632 13812
rect 16592 13530 16620 13806
rect 17592 13728 17644 13734
rect 17592 13670 17644 13676
rect 16580 13524 16632 13530
rect 16580 13466 16632 13472
rect 16488 13456 16540 13462
rect 16488 13398 16540 13404
rect 16592 12850 16620 13466
rect 17604 13394 17632 13670
rect 17592 13388 17644 13394
rect 17592 13330 17644 13336
rect 17132 13252 17184 13258
rect 17132 13194 17184 13200
rect 16580 12844 16632 12850
rect 16580 12786 16632 12792
rect 16488 12776 16540 12782
rect 16488 12718 16540 12724
rect 16396 11348 16448 11354
rect 16396 11290 16448 11296
rect 16500 11268 16528 12718
rect 16764 11280 16816 11286
rect 16500 11240 16764 11268
rect 15752 11076 15804 11082
rect 15752 11018 15804 11024
rect 15568 11008 15620 11014
rect 15568 10950 15620 10956
rect 15476 10668 15528 10674
rect 15476 10610 15528 10616
rect 15488 9518 15516 10610
rect 15580 10146 15608 10950
rect 15764 10810 15792 11018
rect 15752 10804 15804 10810
rect 15752 10746 15804 10752
rect 16396 10736 16448 10742
rect 16396 10678 16448 10684
rect 15660 10464 15712 10470
rect 15660 10406 15712 10412
rect 15672 10266 15700 10406
rect 16408 10266 16436 10678
rect 16500 10470 16528 11240
rect 16764 11222 16816 11228
rect 17040 11144 17092 11150
rect 17040 11086 17092 11092
rect 16672 10804 16724 10810
rect 16672 10746 16724 10752
rect 16488 10464 16540 10470
rect 16488 10406 16540 10412
rect 15660 10260 15712 10266
rect 15660 10202 15712 10208
rect 15936 10260 15988 10266
rect 15936 10202 15988 10208
rect 16396 10260 16448 10266
rect 16396 10202 16448 10208
rect 15580 10118 15700 10146
rect 15476 9512 15528 9518
rect 15476 9454 15528 9460
rect 15488 8838 15516 9454
rect 15568 9104 15620 9110
rect 15568 9046 15620 9052
rect 15580 8974 15608 9046
rect 15568 8968 15620 8974
rect 15568 8910 15620 8916
rect 15476 8832 15528 8838
rect 15476 8774 15528 8780
rect 15580 8634 15608 8910
rect 15568 8628 15620 8634
rect 15568 8570 15620 8576
rect 15580 8498 15608 8570
rect 15568 8492 15620 8498
rect 15568 8434 15620 8440
rect 15476 7948 15528 7954
rect 15476 7890 15528 7896
rect 15488 7857 15516 7890
rect 15474 7848 15530 7857
rect 15474 7783 15530 7792
rect 15384 6248 15436 6254
rect 15384 6190 15436 6196
rect 15200 6180 15252 6186
rect 15200 6122 15252 6128
rect 14924 5704 14976 5710
rect 14924 5646 14976 5652
rect 15212 5370 15240 6122
rect 15476 6112 15528 6118
rect 15476 6054 15528 6060
rect 15488 5846 15516 6054
rect 15476 5840 15528 5846
rect 15476 5782 15528 5788
rect 15292 5568 15344 5574
rect 15292 5510 15344 5516
rect 15200 5364 15252 5370
rect 15200 5306 15252 5312
rect 14556 4616 14608 4622
rect 14556 4558 14608 4564
rect 14568 4146 14596 4558
rect 15212 4554 15240 5306
rect 15304 5234 15332 5510
rect 15580 5370 15608 8434
rect 15672 7954 15700 10118
rect 15948 10062 15976 10202
rect 15936 10056 15988 10062
rect 15936 9998 15988 10004
rect 16408 9518 16436 10202
rect 16500 10062 16528 10406
rect 16684 10266 16712 10746
rect 17052 10606 17080 11086
rect 17144 11082 17172 13194
rect 17696 12986 17724 13874
rect 18156 13870 18184 14350
rect 18144 13864 18196 13870
rect 18144 13806 18196 13812
rect 17684 12980 17736 12986
rect 17684 12922 17736 12928
rect 18432 12782 18460 17326
rect 18512 17274 18564 17280
rect 18616 17202 18644 17818
rect 18788 17536 18840 17542
rect 18788 17478 18840 17484
rect 18512 17196 18564 17202
rect 18512 17138 18564 17144
rect 18604 17196 18656 17202
rect 18604 17138 18656 17144
rect 18524 15416 18552 17138
rect 18696 16448 18748 16454
rect 18696 16390 18748 16396
rect 18708 15638 18736 16390
rect 18800 16182 18828 17478
rect 19076 16794 19104 18226
rect 19168 18086 19196 18362
rect 20352 18352 20404 18358
rect 20352 18294 20404 18300
rect 19156 18080 19208 18086
rect 19156 18022 19208 18028
rect 19524 18080 19576 18086
rect 19524 18022 19576 18028
rect 19168 17610 19196 18022
rect 19156 17604 19208 17610
rect 19156 17546 19208 17552
rect 19432 17604 19484 17610
rect 19432 17546 19484 17552
rect 19064 16788 19116 16794
rect 19064 16730 19116 16736
rect 18788 16176 18840 16182
rect 18788 16118 18840 16124
rect 18696 15632 18748 15638
rect 18696 15574 18748 15580
rect 18696 15428 18748 15434
rect 18524 15388 18696 15416
rect 18696 15370 18748 15376
rect 18800 14958 18828 16118
rect 19168 15978 19196 17546
rect 19248 17536 19300 17542
rect 19248 17478 19300 17484
rect 19260 17202 19288 17478
rect 19444 17202 19472 17546
rect 19248 17196 19300 17202
rect 19248 17138 19300 17144
rect 19432 17196 19484 17202
rect 19432 17138 19484 17144
rect 19536 17134 19564 18022
rect 19524 17128 19576 17134
rect 19524 17070 19576 17076
rect 19984 17128 20036 17134
rect 19984 17070 20036 17076
rect 19156 15972 19208 15978
rect 19156 15914 19208 15920
rect 19168 15858 19196 15914
rect 19076 15830 19196 15858
rect 19708 15904 19760 15910
rect 19708 15846 19760 15852
rect 18972 15360 19024 15366
rect 18972 15302 19024 15308
rect 18788 14952 18840 14958
rect 18788 14894 18840 14900
rect 18984 14498 19012 15302
rect 18892 14470 19012 14498
rect 18892 14414 18920 14470
rect 18696 14408 18748 14414
rect 18696 14350 18748 14356
rect 18880 14408 18932 14414
rect 18880 14350 18932 14356
rect 18708 14006 18736 14350
rect 18972 14340 19024 14346
rect 18972 14282 19024 14288
rect 18984 14074 19012 14282
rect 18972 14068 19024 14074
rect 18972 14010 19024 14016
rect 18696 14000 18748 14006
rect 19076 13954 19104 15830
rect 19720 15570 19748 15846
rect 19708 15564 19760 15570
rect 19708 15506 19760 15512
rect 19996 15502 20024 17070
rect 19432 15496 19484 15502
rect 19432 15438 19484 15444
rect 19984 15496 20036 15502
rect 19984 15438 20036 15444
rect 19340 15360 19392 15366
rect 18696 13942 18748 13948
rect 18892 13926 19104 13954
rect 19168 15308 19340 15314
rect 19168 15302 19392 15308
rect 19168 15286 19380 15302
rect 18892 13802 18920 13926
rect 19168 13870 19196 15286
rect 19444 14822 19472 15438
rect 19432 14816 19484 14822
rect 19432 14758 19484 14764
rect 19248 14408 19300 14414
rect 19248 14350 19300 14356
rect 19156 13864 19208 13870
rect 19156 13806 19208 13812
rect 18880 13796 18932 13802
rect 18880 13738 18932 13744
rect 18696 12912 18748 12918
rect 18696 12854 18748 12860
rect 18420 12776 18472 12782
rect 18472 12736 18552 12764
rect 18420 12718 18472 12724
rect 18420 12640 18472 12646
rect 18420 12582 18472 12588
rect 18432 12374 18460 12582
rect 18420 12368 18472 12374
rect 18420 12310 18472 12316
rect 18432 11762 18460 12310
rect 18524 11898 18552 12736
rect 18708 12102 18736 12854
rect 18892 12714 18920 13738
rect 19064 13728 19116 13734
rect 19064 13670 19116 13676
rect 18880 12708 18932 12714
rect 18880 12650 18932 12656
rect 18892 12442 18920 12650
rect 18972 12640 19024 12646
rect 18972 12582 19024 12588
rect 18880 12436 18932 12442
rect 18880 12378 18932 12384
rect 18984 12306 19012 12582
rect 18972 12300 19024 12306
rect 18972 12242 19024 12248
rect 18880 12232 18932 12238
rect 18880 12174 18932 12180
rect 18696 12096 18748 12102
rect 18696 12038 18748 12044
rect 18512 11892 18564 11898
rect 18512 11834 18564 11840
rect 18420 11756 18472 11762
rect 18420 11698 18472 11704
rect 17868 11688 17920 11694
rect 17868 11630 17920 11636
rect 17776 11144 17828 11150
rect 17776 11086 17828 11092
rect 17132 11076 17184 11082
rect 17132 11018 17184 11024
rect 17408 11076 17460 11082
rect 17408 11018 17460 11024
rect 17040 10600 17092 10606
rect 17040 10542 17092 10548
rect 16672 10260 16724 10266
rect 16672 10202 16724 10208
rect 16488 10056 16540 10062
rect 16488 9998 16540 10004
rect 16396 9512 16448 9518
rect 16396 9454 16448 9460
rect 15936 9036 15988 9042
rect 15936 8978 15988 8984
rect 15752 8424 15804 8430
rect 15750 8392 15752 8401
rect 15804 8392 15806 8401
rect 15750 8327 15806 8336
rect 15948 8090 15976 8978
rect 16408 8566 16436 9454
rect 16500 8906 16528 9998
rect 16684 9586 16712 10202
rect 16856 10124 16908 10130
rect 16856 10066 16908 10072
rect 16672 9580 16724 9586
rect 16672 9522 16724 9528
rect 16684 9178 16712 9522
rect 16868 9382 16896 10066
rect 17052 9926 17080 10542
rect 17420 9994 17448 11018
rect 17408 9988 17460 9994
rect 17408 9930 17460 9936
rect 17040 9920 17092 9926
rect 17040 9862 17092 9868
rect 17788 9586 17816 11086
rect 17880 11082 17908 11630
rect 18524 11286 18552 11834
rect 18708 11830 18736 12038
rect 18892 11898 18920 12174
rect 18880 11892 18932 11898
rect 18880 11834 18932 11840
rect 18696 11824 18748 11830
rect 18696 11766 18748 11772
rect 18604 11756 18656 11762
rect 18604 11698 18656 11704
rect 18512 11280 18564 11286
rect 18512 11222 18564 11228
rect 18144 11212 18196 11218
rect 18144 11154 18196 11160
rect 17868 11076 17920 11082
rect 17868 11018 17920 11024
rect 17880 10742 17908 11018
rect 17868 10736 17920 10742
rect 17868 10678 17920 10684
rect 18156 10724 18184 11154
rect 18616 10810 18644 11698
rect 18708 11082 18736 11766
rect 18696 11076 18748 11082
rect 18696 11018 18748 11024
rect 18604 10804 18656 10810
rect 18604 10746 18656 10752
rect 18236 10736 18288 10742
rect 18156 10696 18236 10724
rect 18156 10130 18184 10696
rect 18236 10678 18288 10684
rect 18512 10600 18564 10606
rect 18512 10542 18564 10548
rect 18328 10464 18380 10470
rect 18328 10406 18380 10412
rect 18340 10130 18368 10406
rect 18524 10266 18552 10542
rect 18512 10260 18564 10266
rect 18512 10202 18564 10208
rect 18616 10146 18644 10746
rect 18144 10124 18196 10130
rect 18144 10066 18196 10072
rect 18328 10124 18380 10130
rect 18328 10066 18380 10072
rect 18524 10118 18644 10146
rect 17868 9988 17920 9994
rect 17868 9930 17920 9936
rect 17776 9580 17828 9586
rect 17776 9522 17828 9528
rect 16856 9376 16908 9382
rect 16856 9318 16908 9324
rect 16672 9172 16724 9178
rect 16672 9114 16724 9120
rect 16868 8974 16896 9318
rect 17592 9172 17644 9178
rect 17592 9114 17644 9120
rect 17224 9036 17276 9042
rect 17224 8978 17276 8984
rect 16856 8968 16908 8974
rect 16856 8910 16908 8916
rect 16488 8900 16540 8906
rect 16488 8842 16540 8848
rect 16396 8560 16448 8566
rect 16396 8502 16448 8508
rect 17236 8498 17264 8978
rect 17408 8560 17460 8566
rect 17408 8502 17460 8508
rect 17224 8492 17276 8498
rect 17224 8434 17276 8440
rect 16764 8424 16816 8430
rect 16764 8366 16816 8372
rect 16120 8288 16172 8294
rect 16120 8230 16172 8236
rect 16672 8288 16724 8294
rect 16672 8230 16724 8236
rect 15936 8084 15988 8090
rect 15936 8026 15988 8032
rect 15660 7948 15712 7954
rect 15660 7890 15712 7896
rect 16132 7886 16160 8230
rect 16684 8090 16712 8230
rect 16672 8084 16724 8090
rect 16672 8026 16724 8032
rect 16776 7886 16804 8366
rect 17236 7954 17264 8434
rect 17316 8288 17368 8294
rect 17316 8230 17368 8236
rect 17224 7948 17276 7954
rect 17224 7890 17276 7896
rect 17328 7886 17356 8230
rect 16120 7880 16172 7886
rect 16120 7822 16172 7828
rect 16764 7880 16816 7886
rect 16764 7822 16816 7828
rect 16948 7880 17000 7886
rect 16948 7822 17000 7828
rect 17316 7880 17368 7886
rect 17316 7822 17368 7828
rect 16580 6384 16632 6390
rect 16580 6326 16632 6332
rect 16960 6338 16988 7822
rect 17420 7750 17448 8502
rect 17604 8498 17632 9114
rect 17788 9042 17816 9522
rect 17880 9450 17908 9930
rect 18236 9920 18288 9926
rect 18236 9862 18288 9868
rect 18248 9654 18276 9862
rect 18340 9722 18368 10066
rect 18524 10062 18552 10118
rect 18512 10056 18564 10062
rect 18512 9998 18564 10004
rect 18604 10056 18656 10062
rect 18604 9998 18656 10004
rect 18328 9716 18380 9722
rect 18328 9658 18380 9664
rect 18236 9648 18288 9654
rect 18236 9590 18288 9596
rect 18340 9518 18368 9658
rect 18328 9512 18380 9518
rect 18328 9454 18380 9460
rect 18616 9450 18644 9998
rect 18788 9648 18840 9654
rect 18788 9590 18840 9596
rect 17868 9444 17920 9450
rect 17868 9386 17920 9392
rect 18604 9444 18656 9450
rect 18604 9386 18656 9392
rect 17776 9036 17828 9042
rect 17776 8978 17828 8984
rect 17500 8492 17552 8498
rect 17500 8434 17552 8440
rect 17592 8492 17644 8498
rect 17592 8434 17644 8440
rect 17684 8492 17736 8498
rect 17684 8434 17736 8440
rect 17868 8492 17920 8498
rect 17868 8434 17920 8440
rect 17512 8022 17540 8434
rect 17500 8016 17552 8022
rect 17500 7958 17552 7964
rect 17408 7744 17460 7750
rect 17408 7686 17460 7692
rect 17132 7472 17184 7478
rect 17132 7414 17184 7420
rect 15936 6316 15988 6322
rect 16212 6316 16264 6322
rect 15988 6276 16212 6304
rect 15936 6258 15988 6264
rect 16212 6258 16264 6264
rect 16396 6316 16448 6322
rect 16396 6258 16448 6264
rect 16028 6180 16080 6186
rect 16028 6122 16080 6128
rect 15752 6112 15804 6118
rect 15750 6080 15752 6089
rect 15804 6080 15806 6089
rect 15750 6015 15806 6024
rect 15568 5364 15620 5370
rect 15568 5306 15620 5312
rect 15292 5228 15344 5234
rect 15292 5170 15344 5176
rect 15568 5228 15620 5234
rect 15568 5170 15620 5176
rect 15384 5092 15436 5098
rect 15384 5034 15436 5040
rect 15396 5001 15424 5034
rect 15382 4992 15438 5001
rect 15382 4927 15438 4936
rect 15580 4758 15608 5170
rect 15568 4752 15620 4758
rect 15568 4694 15620 4700
rect 15764 4690 15792 6015
rect 15936 5704 15988 5710
rect 15936 5646 15988 5652
rect 15948 5370 15976 5646
rect 15936 5364 15988 5370
rect 15936 5306 15988 5312
rect 15842 5264 15898 5273
rect 15842 5199 15844 5208
rect 15896 5199 15898 5208
rect 15844 5170 15896 5176
rect 15752 4684 15804 4690
rect 15752 4626 15804 4632
rect 15844 4616 15896 4622
rect 15844 4558 15896 4564
rect 15200 4548 15252 4554
rect 15200 4490 15252 4496
rect 15856 4214 15884 4558
rect 15844 4208 15896 4214
rect 15844 4150 15896 4156
rect 14556 4140 14608 4146
rect 14556 4082 14608 4088
rect 14462 3224 14518 3233
rect 14462 3159 14518 3168
rect 14476 3126 14504 3159
rect 14096 3120 14148 3126
rect 14096 3062 14148 3068
rect 14464 3120 14516 3126
rect 14464 3062 14516 3068
rect 13452 2916 13504 2922
rect 13452 2858 13504 2864
rect 14568 2854 14596 4082
rect 15948 4078 15976 5306
rect 16040 4865 16068 6122
rect 16212 5704 16264 5710
rect 16212 5646 16264 5652
rect 16118 5536 16174 5545
rect 16118 5471 16174 5480
rect 16026 4856 16082 4865
rect 16132 4826 16160 5471
rect 16026 4791 16082 4800
rect 16120 4820 16172 4826
rect 16120 4762 16172 4768
rect 16224 4622 16252 5646
rect 16304 5636 16356 5642
rect 16304 5578 16356 5584
rect 16212 4616 16264 4622
rect 16212 4558 16264 4564
rect 15752 4072 15804 4078
rect 15752 4014 15804 4020
rect 15936 4072 15988 4078
rect 15936 4014 15988 4020
rect 16210 4040 16266 4049
rect 15200 3936 15252 3942
rect 15200 3878 15252 3884
rect 15212 3534 15240 3878
rect 15476 3732 15528 3738
rect 15476 3674 15528 3680
rect 15488 3534 15516 3674
rect 15200 3528 15252 3534
rect 15200 3470 15252 3476
rect 15476 3528 15528 3534
rect 15476 3470 15528 3476
rect 15764 3398 15792 4014
rect 16210 3975 16266 3984
rect 16118 3904 16174 3913
rect 16118 3839 16174 3848
rect 16028 3528 16080 3534
rect 16028 3470 16080 3476
rect 16040 3398 16068 3470
rect 16132 3398 16160 3839
rect 16224 3670 16252 3975
rect 16316 3942 16344 5578
rect 16408 4826 16436 6258
rect 16488 5296 16540 5302
rect 16592 5273 16620 6326
rect 16960 6310 17080 6338
rect 16856 6248 16908 6254
rect 16856 6190 16908 6196
rect 16672 6180 16724 6186
rect 16672 6122 16724 6128
rect 16684 5778 16712 6122
rect 16672 5772 16724 5778
rect 16672 5714 16724 5720
rect 16868 5302 16896 6190
rect 16948 5908 17000 5914
rect 16948 5850 17000 5856
rect 16960 5817 16988 5850
rect 16946 5808 17002 5817
rect 16946 5743 17002 5752
rect 16948 5704 17000 5710
rect 16948 5646 17000 5652
rect 16856 5296 16908 5302
rect 16488 5238 16540 5244
rect 16578 5264 16634 5273
rect 16396 4820 16448 4826
rect 16396 4762 16448 4768
rect 16500 4690 16528 5238
rect 16856 5238 16908 5244
rect 16960 5234 16988 5646
rect 16578 5199 16580 5208
rect 16632 5199 16634 5208
rect 16948 5228 17000 5234
rect 16580 5170 16632 5176
rect 16948 5170 17000 5176
rect 16488 4684 16540 4690
rect 16488 4626 16540 4632
rect 16592 4622 16620 5170
rect 16672 5024 16724 5030
rect 16672 4966 16724 4972
rect 16580 4616 16632 4622
rect 16580 4558 16632 4564
rect 16396 4208 16448 4214
rect 16396 4150 16448 4156
rect 16304 3936 16356 3942
rect 16304 3878 16356 3884
rect 16212 3664 16264 3670
rect 16212 3606 16264 3612
rect 15752 3392 15804 3398
rect 15752 3334 15804 3340
rect 16028 3392 16080 3398
rect 16028 3334 16080 3340
rect 16120 3392 16172 3398
rect 16120 3334 16172 3340
rect 16316 3126 16344 3878
rect 16408 3194 16436 4150
rect 16592 4146 16620 4558
rect 16684 4146 16712 4966
rect 16960 4842 16988 5170
rect 17052 5001 17080 6310
rect 17038 4992 17094 5001
rect 17038 4927 17094 4936
rect 16868 4814 16988 4842
rect 16868 4622 16896 4814
rect 16948 4752 17000 4758
rect 16948 4694 17000 4700
rect 16856 4616 16908 4622
rect 16856 4558 16908 4564
rect 16580 4140 16632 4146
rect 16580 4082 16632 4088
rect 16672 4140 16724 4146
rect 16672 4082 16724 4088
rect 16592 3942 16620 4082
rect 16764 4072 16816 4078
rect 16764 4014 16816 4020
rect 16580 3936 16632 3942
rect 16580 3878 16632 3884
rect 16592 3534 16620 3878
rect 16580 3528 16632 3534
rect 16580 3470 16632 3476
rect 16776 3194 16804 4014
rect 16868 3466 16896 4558
rect 16960 3534 16988 4694
rect 17040 4616 17092 4622
rect 17040 4558 17092 4564
rect 17052 4282 17080 4558
rect 17144 4486 17172 7414
rect 17224 6724 17276 6730
rect 17224 6666 17276 6672
rect 17236 5953 17264 6666
rect 17316 6180 17368 6186
rect 17316 6122 17368 6128
rect 17222 5944 17278 5953
rect 17222 5879 17224 5888
rect 17276 5879 17278 5888
rect 17224 5850 17276 5856
rect 17222 5808 17278 5817
rect 17222 5743 17278 5752
rect 17236 5370 17264 5743
rect 17328 5710 17356 6122
rect 17316 5704 17368 5710
rect 17316 5646 17368 5652
rect 17224 5364 17276 5370
rect 17224 5306 17276 5312
rect 17316 5228 17368 5234
rect 17316 5170 17368 5176
rect 17328 4690 17356 5170
rect 17316 4684 17368 4690
rect 17316 4626 17368 4632
rect 17224 4616 17276 4622
rect 17224 4558 17276 4564
rect 17132 4480 17184 4486
rect 17132 4422 17184 4428
rect 17236 4282 17264 4558
rect 17040 4276 17092 4282
rect 17040 4218 17092 4224
rect 17224 4276 17276 4282
rect 17224 4218 17276 4224
rect 17040 3664 17092 3670
rect 17040 3606 17092 3612
rect 16948 3528 17000 3534
rect 16948 3470 17000 3476
rect 16856 3460 16908 3466
rect 16856 3402 16908 3408
rect 16948 3392 17000 3398
rect 16948 3334 17000 3340
rect 16396 3188 16448 3194
rect 16396 3130 16448 3136
rect 16764 3188 16816 3194
rect 16764 3130 16816 3136
rect 16304 3120 16356 3126
rect 16960 3074 16988 3334
rect 16304 3062 16356 3068
rect 16776 3058 16988 3074
rect 16764 3052 17000 3058
rect 16816 3046 16948 3052
rect 16764 2994 16816 3000
rect 16948 2994 17000 3000
rect 17052 2990 17080 3606
rect 17328 3516 17356 4626
rect 17420 4049 17448 7686
rect 17696 6866 17724 8434
rect 17776 7812 17828 7818
rect 17776 7754 17828 7760
rect 17788 7274 17816 7754
rect 17880 7546 17908 8434
rect 18420 7948 18472 7954
rect 18420 7890 18472 7896
rect 18328 7880 18380 7886
rect 18248 7828 18328 7834
rect 18248 7822 18380 7828
rect 18248 7806 18368 7822
rect 17868 7540 17920 7546
rect 17868 7482 17920 7488
rect 17960 7404 18012 7410
rect 17960 7346 18012 7352
rect 18052 7404 18104 7410
rect 18052 7346 18104 7352
rect 17972 7274 18000 7346
rect 17776 7268 17828 7274
rect 17776 7210 17828 7216
rect 17960 7268 18012 7274
rect 17960 7210 18012 7216
rect 17684 6860 17736 6866
rect 17684 6802 17736 6808
rect 17498 6080 17554 6089
rect 17498 6015 17554 6024
rect 17512 5778 17540 6015
rect 17500 5772 17552 5778
rect 17500 5714 17552 5720
rect 17684 5704 17736 5710
rect 17684 5646 17736 5652
rect 17592 5160 17644 5166
rect 17592 5102 17644 5108
rect 17498 4992 17554 5001
rect 17498 4927 17554 4936
rect 17512 4146 17540 4927
rect 17500 4140 17552 4146
rect 17500 4082 17552 4088
rect 17406 4040 17462 4049
rect 17604 4010 17632 5102
rect 17696 5098 17724 5646
rect 17788 5574 17816 7210
rect 18064 7002 18092 7346
rect 18052 6996 18104 7002
rect 18052 6938 18104 6944
rect 18248 6730 18276 7806
rect 18328 7744 18380 7750
rect 18328 7686 18380 7692
rect 18340 7546 18368 7686
rect 18328 7540 18380 7546
rect 18328 7482 18380 7488
rect 18432 7478 18460 7890
rect 18800 7886 18828 9590
rect 18880 9036 18932 9042
rect 18880 8978 18932 8984
rect 18892 7886 18920 8978
rect 19076 7886 19104 13670
rect 19260 13394 19288 14350
rect 19444 13938 19472 14758
rect 19996 14074 20024 15438
rect 20364 15434 20392 18294
rect 20456 17728 20484 18770
rect 20548 18086 20576 19858
rect 20812 18692 20864 18698
rect 20812 18634 20864 18640
rect 21180 18692 21232 18698
rect 21180 18634 21232 18640
rect 20824 18426 20852 18634
rect 20812 18420 20864 18426
rect 20812 18362 20864 18368
rect 20536 18080 20588 18086
rect 20536 18022 20588 18028
rect 20548 17882 20576 18022
rect 20536 17876 20588 17882
rect 20588 17836 20668 17864
rect 20536 17818 20588 17824
rect 20536 17740 20588 17746
rect 20456 17700 20536 17728
rect 20536 17682 20588 17688
rect 20640 17202 20668 17836
rect 21192 17610 21220 18634
rect 21180 17604 21232 17610
rect 21180 17546 21232 17552
rect 20628 17196 20680 17202
rect 20628 17138 20680 17144
rect 20628 16108 20680 16114
rect 20628 16050 20680 16056
rect 20444 16040 20496 16046
rect 20444 15982 20496 15988
rect 20456 15502 20484 15982
rect 20640 15706 20668 16050
rect 20904 15904 20956 15910
rect 20904 15846 20956 15852
rect 20628 15700 20680 15706
rect 20628 15642 20680 15648
rect 20720 15700 20772 15706
rect 20720 15642 20772 15648
rect 20444 15496 20496 15502
rect 20444 15438 20496 15444
rect 20352 15428 20404 15434
rect 20352 15370 20404 15376
rect 20628 14816 20680 14822
rect 20732 14770 20760 15642
rect 20916 14958 20944 15846
rect 21192 15706 21220 17546
rect 21364 16040 21416 16046
rect 21364 15982 21416 15988
rect 21376 15706 21404 15982
rect 21180 15700 21232 15706
rect 21180 15642 21232 15648
rect 21364 15700 21416 15706
rect 21364 15642 21416 15648
rect 21468 15366 21496 20402
rect 21916 19916 21968 19922
rect 21916 19858 21968 19864
rect 22100 19916 22152 19922
rect 22100 19858 22152 19864
rect 21928 19378 21956 19858
rect 22008 19712 22060 19718
rect 22008 19654 22060 19660
rect 22020 19446 22048 19654
rect 22008 19440 22060 19446
rect 22008 19382 22060 19388
rect 21916 19372 21968 19378
rect 21916 19314 21968 19320
rect 22112 18834 22140 19858
rect 22296 19514 22324 20810
rect 23480 20392 23532 20398
rect 23480 20334 23532 20340
rect 23756 20392 23808 20398
rect 23756 20334 23808 20340
rect 23492 19922 23520 20334
rect 23204 19916 23256 19922
rect 23204 19858 23256 19864
rect 23480 19916 23532 19922
rect 23480 19858 23532 19864
rect 22284 19508 22336 19514
rect 22284 19450 22336 19456
rect 23216 19446 23244 19858
rect 23480 19780 23532 19786
rect 23480 19722 23532 19728
rect 23204 19440 23256 19446
rect 22282 19408 22338 19417
rect 23204 19382 23256 19388
rect 22282 19343 22284 19352
rect 22336 19343 22338 19352
rect 22284 19314 22336 19320
rect 23492 19310 23520 19722
rect 23768 19514 23796 20334
rect 24412 20262 24440 20810
rect 24400 20256 24452 20262
rect 24400 20198 24452 20204
rect 24124 19984 24176 19990
rect 24124 19926 24176 19932
rect 23848 19780 23900 19786
rect 23848 19722 23900 19728
rect 23940 19780 23992 19786
rect 23940 19722 23992 19728
rect 23756 19508 23808 19514
rect 23756 19450 23808 19456
rect 23754 19408 23810 19417
rect 23572 19372 23624 19378
rect 23572 19314 23624 19320
rect 23664 19372 23716 19378
rect 23754 19343 23756 19352
rect 23664 19314 23716 19320
rect 23808 19343 23810 19352
rect 23756 19314 23808 19320
rect 23204 19304 23256 19310
rect 23204 19246 23256 19252
rect 23480 19304 23532 19310
rect 23480 19246 23532 19252
rect 23216 18902 23244 19246
rect 23204 18896 23256 18902
rect 23204 18838 23256 18844
rect 23584 18834 23612 19314
rect 23676 18970 23704 19314
rect 23664 18964 23716 18970
rect 23664 18906 23716 18912
rect 23860 18834 23888 19722
rect 22100 18828 22152 18834
rect 22100 18770 22152 18776
rect 23388 18828 23440 18834
rect 23388 18770 23440 18776
rect 23572 18828 23624 18834
rect 23572 18770 23624 18776
rect 23848 18828 23900 18834
rect 23848 18770 23900 18776
rect 23204 18760 23256 18766
rect 23204 18702 23256 18708
rect 22008 18692 22060 18698
rect 22008 18634 22060 18640
rect 22020 18426 22048 18634
rect 22376 18624 22428 18630
rect 22376 18566 22428 18572
rect 22008 18420 22060 18426
rect 22008 18362 22060 18368
rect 22388 18290 22416 18566
rect 22100 18284 22152 18290
rect 22100 18226 22152 18232
rect 22376 18284 22428 18290
rect 22376 18226 22428 18232
rect 21732 18080 21784 18086
rect 21732 18022 21784 18028
rect 21744 17746 21772 18022
rect 22112 17882 22140 18226
rect 23216 18222 23244 18702
rect 22744 18216 22796 18222
rect 22744 18158 22796 18164
rect 23204 18216 23256 18222
rect 23204 18158 23256 18164
rect 22100 17876 22152 17882
rect 22100 17818 22152 17824
rect 21732 17740 21784 17746
rect 21732 17682 21784 17688
rect 22100 17740 22152 17746
rect 22100 17682 22152 17688
rect 21824 16040 21876 16046
rect 21824 15982 21876 15988
rect 21836 15570 21864 15982
rect 21824 15564 21876 15570
rect 21824 15506 21876 15512
rect 21916 15496 21968 15502
rect 21916 15438 21968 15444
rect 21456 15360 21508 15366
rect 21456 15302 21508 15308
rect 21928 15162 21956 15438
rect 22112 15434 22140 17682
rect 22376 17536 22428 17542
rect 22376 17478 22428 17484
rect 22284 17332 22336 17338
rect 22284 17274 22336 17280
rect 22296 16998 22324 17274
rect 22388 16998 22416 17478
rect 22652 17264 22704 17270
rect 22652 17206 22704 17212
rect 22468 17060 22520 17066
rect 22468 17002 22520 17008
rect 22284 16992 22336 16998
rect 22284 16934 22336 16940
rect 22376 16992 22428 16998
rect 22376 16934 22428 16940
rect 22192 16448 22244 16454
rect 22192 16390 22244 16396
rect 22204 16182 22232 16390
rect 22192 16176 22244 16182
rect 22192 16118 22244 16124
rect 22192 15700 22244 15706
rect 22192 15642 22244 15648
rect 22100 15428 22152 15434
rect 22100 15370 22152 15376
rect 21916 15156 21968 15162
rect 21916 15098 21968 15104
rect 20904 14952 20956 14958
rect 20904 14894 20956 14900
rect 20680 14764 20760 14770
rect 20628 14758 20760 14764
rect 20640 14742 20760 14758
rect 20732 14498 20760 14742
rect 20640 14470 20760 14498
rect 20640 14414 20668 14470
rect 20628 14408 20680 14414
rect 20628 14350 20680 14356
rect 20996 14272 21048 14278
rect 20996 14214 21048 14220
rect 19984 14068 20036 14074
rect 19984 14010 20036 14016
rect 20628 14068 20680 14074
rect 20628 14010 20680 14016
rect 19432 13932 19484 13938
rect 19432 13874 19484 13880
rect 19248 13388 19300 13394
rect 19248 13330 19300 13336
rect 19156 12844 19208 12850
rect 19156 12786 19208 12792
rect 19168 12442 19196 12786
rect 19156 12436 19208 12442
rect 19156 12378 19208 12384
rect 19260 11558 19288 13330
rect 19248 11552 19300 11558
rect 19248 11494 19300 11500
rect 19260 10674 19288 11494
rect 19248 10668 19300 10674
rect 19248 10610 19300 10616
rect 19248 9376 19300 9382
rect 19248 9318 19300 9324
rect 19260 9178 19288 9318
rect 19248 9172 19300 9178
rect 19248 9114 19300 9120
rect 19444 8430 19472 13874
rect 19708 12776 19760 12782
rect 19708 12718 19760 12724
rect 19720 11898 19748 12718
rect 20640 12442 20668 14010
rect 21008 13870 21036 14214
rect 21928 13938 21956 15098
rect 22112 14006 22140 15370
rect 22100 14000 22152 14006
rect 22100 13942 22152 13948
rect 22204 13938 22232 15642
rect 22376 15428 22428 15434
rect 22376 15370 22428 15376
rect 22388 15162 22416 15370
rect 22376 15156 22428 15162
rect 22376 15098 22428 15104
rect 22480 15026 22508 17002
rect 22560 16992 22612 16998
rect 22560 16934 22612 16940
rect 22572 16590 22600 16934
rect 22664 16794 22692 17206
rect 22652 16788 22704 16794
rect 22652 16730 22704 16736
rect 22756 16674 22784 18158
rect 23216 17542 23244 18158
rect 23400 17882 23428 18770
rect 23388 17876 23440 17882
rect 23388 17818 23440 17824
rect 23952 17678 23980 19722
rect 24032 19712 24084 19718
rect 24032 19654 24084 19660
rect 24044 18222 24072 19654
rect 24136 18290 24164 19926
rect 24216 19848 24268 19854
rect 24216 19790 24268 19796
rect 24228 19446 24256 19790
rect 24412 19446 24440 20198
rect 24780 19854 24808 20946
rect 25516 20942 25544 21626
rect 26620 21554 26648 22442
rect 26976 22432 27028 22438
rect 26976 22374 27028 22380
rect 26988 22234 27016 22374
rect 26976 22228 27028 22234
rect 26976 22170 27028 22176
rect 27344 21888 27396 21894
rect 27344 21830 27396 21836
rect 27356 21622 27384 21830
rect 27344 21616 27396 21622
rect 27344 21558 27396 21564
rect 26608 21548 26660 21554
rect 26608 21490 26660 21496
rect 26332 21480 26384 21486
rect 26332 21422 26384 21428
rect 25504 20936 25556 20942
rect 25504 20878 25556 20884
rect 25516 20534 25544 20878
rect 26344 20602 26372 21422
rect 26792 21412 26844 21418
rect 26792 21354 26844 21360
rect 26804 21010 26832 21354
rect 27160 21344 27212 21350
rect 27160 21286 27212 21292
rect 26792 21004 26844 21010
rect 26792 20946 26844 20952
rect 26792 20868 26844 20874
rect 26792 20810 26844 20816
rect 26332 20596 26384 20602
rect 26332 20538 26384 20544
rect 25504 20528 25556 20534
rect 25504 20470 25556 20476
rect 25516 20330 25544 20470
rect 26700 20392 26752 20398
rect 26700 20334 26752 20340
rect 25504 20324 25556 20330
rect 25504 20266 25556 20272
rect 26712 20058 26740 20334
rect 26700 20052 26752 20058
rect 26700 19994 26752 20000
rect 24768 19848 24820 19854
rect 24768 19790 24820 19796
rect 25044 19848 25096 19854
rect 25044 19790 25096 19796
rect 24216 19440 24268 19446
rect 24216 19382 24268 19388
rect 24400 19440 24452 19446
rect 24400 19382 24452 19388
rect 24952 19372 25004 19378
rect 24952 19314 25004 19320
rect 24492 19304 24544 19310
rect 24492 19246 24544 19252
rect 24504 18426 24532 19246
rect 24860 18760 24912 18766
rect 24860 18702 24912 18708
rect 24492 18420 24544 18426
rect 24492 18362 24544 18368
rect 24676 18420 24728 18426
rect 24676 18362 24728 18368
rect 24124 18284 24176 18290
rect 24124 18226 24176 18232
rect 24032 18216 24084 18222
rect 24032 18158 24084 18164
rect 24136 17678 24164 18226
rect 24688 17678 24716 18362
rect 24872 18358 24900 18702
rect 24860 18352 24912 18358
rect 24860 18294 24912 18300
rect 23388 17672 23440 17678
rect 23388 17614 23440 17620
rect 23940 17672 23992 17678
rect 23940 17614 23992 17620
rect 24124 17672 24176 17678
rect 24124 17614 24176 17620
rect 24676 17672 24728 17678
rect 24676 17614 24728 17620
rect 24964 17626 24992 19314
rect 25056 19310 25084 19790
rect 26804 19786 26832 20810
rect 27172 20754 27200 21286
rect 27172 20726 27292 20754
rect 27264 20398 27292 20726
rect 27356 20516 27384 21558
rect 27448 21554 27476 22510
rect 27436 21548 27488 21554
rect 27436 21490 27488 21496
rect 27632 20602 27660 22510
rect 27816 22094 27844 22986
rect 27896 22636 27948 22642
rect 27896 22578 27948 22584
rect 27724 22066 27844 22094
rect 27620 20596 27672 20602
rect 27620 20538 27672 20544
rect 27436 20528 27488 20534
rect 27356 20488 27436 20516
rect 27436 20470 27488 20476
rect 27252 20392 27304 20398
rect 27252 20334 27304 20340
rect 27264 19922 27292 20334
rect 27252 19916 27304 19922
rect 27252 19858 27304 19864
rect 27724 19854 27752 22066
rect 27804 20800 27856 20806
rect 27908 20788 27936 22578
rect 28000 22506 28028 23734
rect 28356 22704 28408 22710
rect 28356 22646 28408 22652
rect 27988 22500 28040 22506
rect 27988 22442 28040 22448
rect 27856 20760 27936 20788
rect 27804 20742 27856 20748
rect 27816 19922 27844 20742
rect 28000 20466 28028 22442
rect 28080 22432 28132 22438
rect 28080 22374 28132 22380
rect 28092 20534 28120 22374
rect 28264 21480 28316 21486
rect 28264 21422 28316 21428
rect 28172 21344 28224 21350
rect 28172 21286 28224 21292
rect 28184 20534 28212 21286
rect 28080 20528 28132 20534
rect 28080 20470 28132 20476
rect 28172 20528 28224 20534
rect 28172 20470 28224 20476
rect 27988 20460 28040 20466
rect 27988 20402 28040 20408
rect 27988 20256 28040 20262
rect 27988 20198 28040 20204
rect 27804 19916 27856 19922
rect 27804 19858 27856 19864
rect 27712 19848 27764 19854
rect 27712 19790 27764 19796
rect 26792 19780 26844 19786
rect 26792 19722 26844 19728
rect 25044 19304 25096 19310
rect 25044 19246 25096 19252
rect 26148 19304 26200 19310
rect 26148 19246 26200 19252
rect 26160 18766 26188 19246
rect 26148 18760 26200 18766
rect 26148 18702 26200 18708
rect 25044 18692 25096 18698
rect 25044 18634 25096 18640
rect 25780 18692 25832 18698
rect 25780 18634 25832 18640
rect 25056 18086 25084 18634
rect 25792 18426 25820 18634
rect 25780 18420 25832 18426
rect 25780 18362 25832 18368
rect 25136 18284 25188 18290
rect 25136 18226 25188 18232
rect 25320 18284 25372 18290
rect 25320 18226 25372 18232
rect 25596 18284 25648 18290
rect 25596 18226 25648 18232
rect 25044 18080 25096 18086
rect 25044 18022 25096 18028
rect 25056 17762 25084 18022
rect 25148 17882 25176 18226
rect 25332 17882 25360 18226
rect 25136 17876 25188 17882
rect 25136 17818 25188 17824
rect 25320 17876 25372 17882
rect 25320 17818 25372 17824
rect 25056 17734 25176 17762
rect 25148 17678 25176 17734
rect 25320 17740 25372 17746
rect 25240 17700 25320 17728
rect 25136 17672 25188 17678
rect 23204 17536 23256 17542
rect 23204 17478 23256 17484
rect 23296 17536 23348 17542
rect 23296 17478 23348 17484
rect 23308 17338 23336 17478
rect 23296 17332 23348 17338
rect 23296 17274 23348 17280
rect 22664 16646 22784 16674
rect 22664 16590 22692 16646
rect 22560 16584 22612 16590
rect 22560 16526 22612 16532
rect 22652 16584 22704 16590
rect 22652 16526 22704 16532
rect 22664 15026 22692 16526
rect 23400 16182 23428 17614
rect 23952 16998 23980 17614
rect 23940 16992 23992 16998
rect 23940 16934 23992 16940
rect 23952 16658 23980 16934
rect 23940 16652 23992 16658
rect 23940 16594 23992 16600
rect 23952 16250 23980 16594
rect 23940 16244 23992 16250
rect 23940 16186 23992 16192
rect 23388 16176 23440 16182
rect 23388 16118 23440 16124
rect 23400 15706 23428 16118
rect 23388 15700 23440 15706
rect 23388 15642 23440 15648
rect 23400 15434 23428 15642
rect 24136 15502 24164 17614
rect 24964 17598 25084 17626
rect 25136 17614 25188 17620
rect 25056 17542 25084 17598
rect 25148 17542 25176 17614
rect 25044 17536 25096 17542
rect 25044 17478 25096 17484
rect 25136 17536 25188 17542
rect 25136 17478 25188 17484
rect 25056 17354 25084 17478
rect 25056 17326 25176 17354
rect 25044 16992 25096 16998
rect 25044 16934 25096 16940
rect 25056 16794 25084 16934
rect 25044 16788 25096 16794
rect 25044 16730 25096 16736
rect 25148 16658 25176 17326
rect 25240 16658 25268 17700
rect 25320 17682 25372 17688
rect 25608 17678 25636 18226
rect 25872 18216 25924 18222
rect 25872 18158 25924 18164
rect 25596 17672 25648 17678
rect 25596 17614 25648 17620
rect 25608 17202 25636 17614
rect 25884 17542 25912 18158
rect 26160 17746 26188 18702
rect 26804 18680 26832 19722
rect 27712 19712 27764 19718
rect 27712 19654 27764 19660
rect 27724 19514 27752 19654
rect 27712 19508 27764 19514
rect 27712 19450 27764 19456
rect 27896 19304 27948 19310
rect 27896 19246 27948 19252
rect 27908 18970 27936 19246
rect 27896 18964 27948 18970
rect 27896 18906 27948 18912
rect 26884 18692 26936 18698
rect 26804 18652 26884 18680
rect 26884 18634 26936 18640
rect 26148 17740 26200 17746
rect 26148 17682 26200 17688
rect 26896 17610 26924 18634
rect 26792 17604 26844 17610
rect 26792 17546 26844 17552
rect 26884 17604 26936 17610
rect 26884 17546 26936 17552
rect 25780 17536 25832 17542
rect 25780 17478 25832 17484
rect 25872 17536 25924 17542
rect 25872 17478 25924 17484
rect 25596 17196 25648 17202
rect 25596 17138 25648 17144
rect 25412 17128 25464 17134
rect 25412 17070 25464 17076
rect 25136 16652 25188 16658
rect 25136 16594 25188 16600
rect 25228 16652 25280 16658
rect 25228 16594 25280 16600
rect 24676 16448 24728 16454
rect 24676 16390 24728 16396
rect 24860 16448 24912 16454
rect 24860 16390 24912 16396
rect 24124 15496 24176 15502
rect 24124 15438 24176 15444
rect 23388 15428 23440 15434
rect 23388 15370 23440 15376
rect 23400 15094 23428 15370
rect 24136 15162 24164 15438
rect 24688 15434 24716 16390
rect 24872 16250 24900 16390
rect 24860 16244 24912 16250
rect 24860 16186 24912 16192
rect 25240 15570 25268 16594
rect 25424 16114 25452 17070
rect 25504 16516 25556 16522
rect 25504 16458 25556 16464
rect 25516 16250 25544 16458
rect 25504 16244 25556 16250
rect 25504 16186 25556 16192
rect 25608 16114 25636 17138
rect 25792 16250 25820 17478
rect 25884 17134 25912 17478
rect 25872 17128 25924 17134
rect 25872 17070 25924 17076
rect 26804 16794 26832 17546
rect 26896 17270 26924 17546
rect 26884 17264 26936 17270
rect 26884 17206 26936 17212
rect 26792 16788 26844 16794
rect 26792 16730 26844 16736
rect 26896 16726 26924 17206
rect 26884 16720 26936 16726
rect 26884 16662 26936 16668
rect 26608 16584 26660 16590
rect 26608 16526 26660 16532
rect 25780 16244 25832 16250
rect 25780 16186 25832 16192
rect 25412 16108 25464 16114
rect 25412 16050 25464 16056
rect 25596 16108 25648 16114
rect 25596 16050 25648 16056
rect 25228 15564 25280 15570
rect 25228 15506 25280 15512
rect 24676 15428 24728 15434
rect 24676 15370 24728 15376
rect 24124 15156 24176 15162
rect 24124 15098 24176 15104
rect 23388 15088 23440 15094
rect 23388 15030 23440 15036
rect 22468 15020 22520 15026
rect 22468 14962 22520 14968
rect 22652 15020 22704 15026
rect 22652 14962 22704 14968
rect 21916 13932 21968 13938
rect 21916 13874 21968 13880
rect 22192 13932 22244 13938
rect 22192 13874 22244 13880
rect 20996 13864 21048 13870
rect 20996 13806 21048 13812
rect 22204 13818 22232 13874
rect 25424 13870 25452 16050
rect 26148 15904 26200 15910
rect 26148 15846 26200 15852
rect 26160 15706 26188 15846
rect 26148 15700 26200 15706
rect 26148 15642 26200 15648
rect 26620 15502 26648 16526
rect 26976 16448 27028 16454
rect 26976 16390 27028 16396
rect 26988 16114 27016 16390
rect 26976 16108 27028 16114
rect 26976 16050 27028 16056
rect 27620 15904 27672 15910
rect 27620 15846 27672 15852
rect 26608 15496 26660 15502
rect 26608 15438 26660 15444
rect 27160 15360 27212 15366
rect 27160 15302 27212 15308
rect 26516 14408 26568 14414
rect 26516 14350 26568 14356
rect 26528 14074 26556 14350
rect 26516 14068 26568 14074
rect 26516 14010 26568 14016
rect 25504 13932 25556 13938
rect 25504 13874 25556 13880
rect 25412 13864 25464 13870
rect 22100 13796 22152 13802
rect 22204 13790 22416 13818
rect 25412 13806 25464 13812
rect 22100 13738 22152 13744
rect 22008 13728 22060 13734
rect 22008 13670 22060 13676
rect 21548 13320 21600 13326
rect 21548 13262 21600 13268
rect 21180 12844 21232 12850
rect 21180 12786 21232 12792
rect 20720 12640 20772 12646
rect 20720 12582 20772 12588
rect 20628 12436 20680 12442
rect 20628 12378 20680 12384
rect 20640 12170 20668 12378
rect 20260 12164 20312 12170
rect 20260 12106 20312 12112
rect 20628 12164 20680 12170
rect 20628 12106 20680 12112
rect 20272 11898 20300 12106
rect 19708 11892 19760 11898
rect 19708 11834 19760 11840
rect 20260 11892 20312 11898
rect 20260 11834 20312 11840
rect 20272 11694 20300 11834
rect 20260 11688 20312 11694
rect 20260 11630 20312 11636
rect 20640 11354 20668 12106
rect 20732 11830 20760 12582
rect 20996 12232 21048 12238
rect 20996 12174 21048 12180
rect 20720 11824 20772 11830
rect 20720 11766 20772 11772
rect 21008 11694 21036 12174
rect 20996 11688 21048 11694
rect 20996 11630 21048 11636
rect 21192 11354 21220 12786
rect 21560 12238 21588 13262
rect 21824 13252 21876 13258
rect 21824 13194 21876 13200
rect 21836 12986 21864 13194
rect 21824 12980 21876 12986
rect 21824 12922 21876 12928
rect 22020 12850 22048 13670
rect 22008 12844 22060 12850
rect 22008 12786 22060 12792
rect 21548 12232 21600 12238
rect 21548 12174 21600 12180
rect 21824 12232 21876 12238
rect 21824 12174 21876 12180
rect 21456 11892 21508 11898
rect 21456 11834 21508 11840
rect 20444 11348 20496 11354
rect 20444 11290 20496 11296
rect 20628 11348 20680 11354
rect 20628 11290 20680 11296
rect 21180 11348 21232 11354
rect 21180 11290 21232 11296
rect 19524 11144 19576 11150
rect 19524 11086 19576 11092
rect 19536 10674 19564 11086
rect 19524 10668 19576 10674
rect 19524 10610 19576 10616
rect 19536 10130 19564 10610
rect 20076 10600 20128 10606
rect 20076 10542 20128 10548
rect 19524 10124 19576 10130
rect 19524 10066 19576 10072
rect 20088 9722 20116 10542
rect 20456 10062 20484 11290
rect 20536 11144 20588 11150
rect 20640 11132 20668 11290
rect 20588 11104 20668 11132
rect 20536 11086 20588 11092
rect 21468 10742 21496 11834
rect 21548 11620 21600 11626
rect 21548 11562 21600 11568
rect 21560 11150 21588 11562
rect 21548 11144 21600 11150
rect 21548 11086 21600 11092
rect 21456 10736 21508 10742
rect 21456 10678 21508 10684
rect 20444 10056 20496 10062
rect 20444 9998 20496 10004
rect 20352 9988 20404 9994
rect 20352 9930 20404 9936
rect 20720 9988 20772 9994
rect 20720 9930 20772 9936
rect 20076 9716 20128 9722
rect 20076 9658 20128 9664
rect 19800 9648 19852 9654
rect 19800 9590 19852 9596
rect 19812 9178 19840 9590
rect 20364 9586 20392 9930
rect 20732 9586 20760 9930
rect 20904 9920 20956 9926
rect 20904 9862 20956 9868
rect 20260 9580 20312 9586
rect 20260 9522 20312 9528
rect 20352 9580 20404 9586
rect 20352 9522 20404 9528
rect 20720 9580 20772 9586
rect 20720 9522 20772 9528
rect 19800 9172 19852 9178
rect 19800 9114 19852 9120
rect 19708 8560 19760 8566
rect 19708 8502 19760 8508
rect 19432 8424 19484 8430
rect 19432 8366 19484 8372
rect 19444 7886 19472 8366
rect 19524 8288 19576 8294
rect 19524 8230 19576 8236
rect 18788 7880 18840 7886
rect 18788 7822 18840 7828
rect 18880 7880 18932 7886
rect 18880 7822 18932 7828
rect 19064 7880 19116 7886
rect 19064 7822 19116 7828
rect 19432 7880 19484 7886
rect 19432 7822 19484 7828
rect 18420 7472 18472 7478
rect 18420 7414 18472 7420
rect 18512 7404 18564 7410
rect 18512 7346 18564 7352
rect 18696 7404 18748 7410
rect 18696 7346 18748 7352
rect 18328 6928 18380 6934
rect 18328 6870 18380 6876
rect 18236 6724 18288 6730
rect 18236 6666 18288 6672
rect 17776 5568 17828 5574
rect 17776 5510 17828 5516
rect 17960 5296 18012 5302
rect 17960 5238 18012 5244
rect 17684 5092 17736 5098
rect 17684 5034 17736 5040
rect 17972 4146 18000 5238
rect 18052 5228 18104 5234
rect 18052 5170 18104 5176
rect 18064 4826 18092 5170
rect 18052 4820 18104 4826
rect 18052 4762 18104 4768
rect 18248 4729 18276 6666
rect 18234 4720 18290 4729
rect 18234 4655 18290 4664
rect 17960 4140 18012 4146
rect 17960 4082 18012 4088
rect 17406 3975 17462 3984
rect 17592 4004 17644 4010
rect 17592 3946 17644 3952
rect 17604 3738 17632 3946
rect 17972 3738 18000 4082
rect 18340 3942 18368 6870
rect 18524 6322 18552 7346
rect 18604 7336 18656 7342
rect 18604 7278 18656 7284
rect 18616 6798 18644 7278
rect 18604 6792 18656 6798
rect 18604 6734 18656 6740
rect 18512 6316 18564 6322
rect 18512 6258 18564 6264
rect 18524 5370 18552 6258
rect 18708 6254 18736 7346
rect 18800 6866 18828 7822
rect 18788 6860 18840 6866
rect 18788 6802 18840 6808
rect 18892 6798 18920 7822
rect 18972 7812 19024 7818
rect 18972 7754 19024 7760
rect 19156 7812 19208 7818
rect 19156 7754 19208 7760
rect 18984 7426 19012 7754
rect 19168 7478 19196 7754
rect 19248 7744 19300 7750
rect 19248 7686 19300 7692
rect 19260 7478 19288 7686
rect 19444 7546 19472 7822
rect 19432 7540 19484 7546
rect 19432 7482 19484 7488
rect 19536 7478 19564 8230
rect 19720 8090 19748 8502
rect 19812 8362 19840 9114
rect 20076 8968 20128 8974
rect 20076 8910 20128 8916
rect 19892 8832 19944 8838
rect 19892 8774 19944 8780
rect 19800 8356 19852 8362
rect 19800 8298 19852 8304
rect 19904 8294 19932 8774
rect 20088 8498 20116 8910
rect 20168 8560 20220 8566
rect 20168 8502 20220 8508
rect 20076 8492 20128 8498
rect 20076 8434 20128 8440
rect 20180 8430 20208 8502
rect 20272 8430 20300 9522
rect 20364 8974 20392 9522
rect 20444 9512 20496 9518
rect 20444 9454 20496 9460
rect 20352 8968 20404 8974
rect 20352 8910 20404 8916
rect 20352 8560 20404 8566
rect 20352 8502 20404 8508
rect 20456 8514 20484 9454
rect 20732 9042 20760 9522
rect 20916 9178 20944 9862
rect 21180 9580 21232 9586
rect 21180 9522 21232 9528
rect 20904 9172 20956 9178
rect 20904 9114 20956 9120
rect 21192 9042 21220 9522
rect 20720 9036 20772 9042
rect 20720 8978 20772 8984
rect 21180 9036 21232 9042
rect 21180 8978 21232 8984
rect 20536 8968 20588 8974
rect 20536 8910 20588 8916
rect 20548 8634 20576 8910
rect 21088 8900 21140 8906
rect 21088 8842 21140 8848
rect 20812 8832 20864 8838
rect 20812 8774 20864 8780
rect 20536 8628 20588 8634
rect 20536 8570 20588 8576
rect 20824 8514 20852 8774
rect 21100 8634 21128 8842
rect 21088 8628 21140 8634
rect 21088 8570 21140 8576
rect 20168 8424 20220 8430
rect 20168 8366 20220 8372
rect 20260 8424 20312 8430
rect 20260 8366 20312 8372
rect 19892 8288 19944 8294
rect 19892 8230 19944 8236
rect 20260 8288 20312 8294
rect 20260 8230 20312 8236
rect 19708 8084 19760 8090
rect 19708 8026 19760 8032
rect 20272 7954 20300 8230
rect 20260 7948 20312 7954
rect 20260 7890 20312 7896
rect 20364 7886 20392 8502
rect 20456 8498 20576 8514
rect 20456 8492 20588 8498
rect 20456 8486 20536 8492
rect 20824 8486 21128 8514
rect 20536 8434 20588 8440
rect 21100 8430 21128 8486
rect 21088 8424 21140 8430
rect 21088 8366 21140 8372
rect 20352 7880 20404 7886
rect 20352 7822 20404 7828
rect 19156 7472 19208 7478
rect 18984 7398 19104 7426
rect 19156 7414 19208 7420
rect 19248 7472 19300 7478
rect 19248 7414 19300 7420
rect 19524 7472 19576 7478
rect 19524 7414 19576 7420
rect 19076 7002 19104 7398
rect 19064 6996 19116 7002
rect 19064 6938 19116 6944
rect 18880 6792 18932 6798
rect 18880 6734 18932 6740
rect 19168 6730 19196 7414
rect 21192 7206 21220 8978
rect 21468 7478 21496 10678
rect 21548 10464 21600 10470
rect 21548 10406 21600 10412
rect 21560 9382 21588 10406
rect 21836 9994 21864 12174
rect 21916 11212 21968 11218
rect 21916 11154 21968 11160
rect 21928 10470 21956 11154
rect 21916 10464 21968 10470
rect 21916 10406 21968 10412
rect 21824 9988 21876 9994
rect 21824 9930 21876 9936
rect 21548 9376 21600 9382
rect 21548 9318 21600 9324
rect 21836 8634 21864 9930
rect 21824 8628 21876 8634
rect 21824 8570 21876 8576
rect 22112 7886 22140 13738
rect 22192 13184 22244 13190
rect 22192 13126 22244 13132
rect 22204 12238 22232 13126
rect 22284 12640 22336 12646
rect 22284 12582 22336 12588
rect 22192 12232 22244 12238
rect 22192 12174 22244 12180
rect 22192 12096 22244 12102
rect 22192 12038 22244 12044
rect 22204 11642 22232 12038
rect 22296 11762 22324 12582
rect 22388 12306 22416 13790
rect 24860 13728 24912 13734
rect 24860 13670 24912 13676
rect 23204 13252 23256 13258
rect 23204 13194 23256 13200
rect 22560 12844 22612 12850
rect 22560 12786 22612 12792
rect 22376 12300 22428 12306
rect 22376 12242 22428 12248
rect 22468 12164 22520 12170
rect 22468 12106 22520 12112
rect 22284 11756 22336 11762
rect 22284 11698 22336 11704
rect 22376 11756 22428 11762
rect 22376 11698 22428 11704
rect 22204 11614 22324 11642
rect 22192 11280 22244 11286
rect 22192 11222 22244 11228
rect 22204 10674 22232 11222
rect 22296 11014 22324 11614
rect 22388 11354 22416 11698
rect 22376 11348 22428 11354
rect 22376 11290 22428 11296
rect 22480 11218 22508 12106
rect 22572 11558 22600 12786
rect 22652 12776 22704 12782
rect 22652 12718 22704 12724
rect 22664 11898 22692 12718
rect 22744 12708 22796 12714
rect 22744 12650 22796 12656
rect 22756 12170 22784 12650
rect 23216 12186 23244 13194
rect 23388 13184 23440 13190
rect 23388 13126 23440 13132
rect 23400 12918 23428 13126
rect 23388 12912 23440 12918
rect 23388 12854 23440 12860
rect 23296 12844 23348 12850
rect 23296 12786 23348 12792
rect 23308 12442 23336 12786
rect 24216 12776 24268 12782
rect 24216 12718 24268 12724
rect 23480 12640 23532 12646
rect 23480 12582 23532 12588
rect 23296 12436 23348 12442
rect 23296 12378 23348 12384
rect 22744 12164 22796 12170
rect 23216 12158 23428 12186
rect 22744 12106 22796 12112
rect 23400 12102 23428 12158
rect 23388 12096 23440 12102
rect 23388 12038 23440 12044
rect 22652 11892 22704 11898
rect 22652 11834 22704 11840
rect 22664 11626 22692 11834
rect 23400 11830 23428 12038
rect 23388 11824 23440 11830
rect 23388 11766 23440 11772
rect 22652 11620 22704 11626
rect 22652 11562 22704 11568
rect 22560 11552 22612 11558
rect 22560 11494 22612 11500
rect 22468 11212 22520 11218
rect 22468 11154 22520 11160
rect 22284 11008 22336 11014
rect 22284 10950 22336 10956
rect 22296 10742 22324 10950
rect 22480 10810 22508 11154
rect 23400 11082 23428 11766
rect 23388 11076 23440 11082
rect 23388 11018 23440 11024
rect 23112 11008 23164 11014
rect 23112 10950 23164 10956
rect 22468 10804 22520 10810
rect 22468 10746 22520 10752
rect 22284 10736 22336 10742
rect 22284 10678 22336 10684
rect 23124 10674 23152 10950
rect 23492 10674 23520 12582
rect 24228 12102 24256 12718
rect 24676 12640 24728 12646
rect 24676 12582 24728 12588
rect 24400 12300 24452 12306
rect 24400 12242 24452 12248
rect 24216 12096 24268 12102
rect 24216 12038 24268 12044
rect 23940 11076 23992 11082
rect 23940 11018 23992 11024
rect 23952 10810 23980 11018
rect 23940 10804 23992 10810
rect 23940 10746 23992 10752
rect 24228 10742 24256 12038
rect 24412 11762 24440 12242
rect 24400 11756 24452 11762
rect 24400 11698 24452 11704
rect 24412 11218 24440 11698
rect 24400 11212 24452 11218
rect 24400 11154 24452 11160
rect 24216 10736 24268 10742
rect 24216 10678 24268 10684
rect 22192 10668 22244 10674
rect 22192 10610 22244 10616
rect 22560 10668 22612 10674
rect 22560 10610 22612 10616
rect 23112 10668 23164 10674
rect 23112 10610 23164 10616
rect 23480 10668 23532 10674
rect 23480 10610 23532 10616
rect 24584 10668 24636 10674
rect 24584 10610 24636 10616
rect 22572 10554 22600 10610
rect 22572 10526 22692 10554
rect 22664 9654 22692 10526
rect 24596 10062 24624 10610
rect 22744 10056 22796 10062
rect 22744 9998 22796 10004
rect 24584 10056 24636 10062
rect 24584 9998 24636 10004
rect 22756 9654 22784 9998
rect 22652 9648 22704 9654
rect 22652 9590 22704 9596
rect 22744 9648 22796 9654
rect 22744 9590 22796 9596
rect 22664 9042 22692 9590
rect 23664 9580 23716 9586
rect 23664 9522 23716 9528
rect 22652 9036 22704 9042
rect 22652 8978 22704 8984
rect 22284 8968 22336 8974
rect 22284 8910 22336 8916
rect 22296 8498 22324 8910
rect 22744 8832 22796 8838
rect 22744 8774 22796 8780
rect 22756 8634 22784 8774
rect 22744 8628 22796 8634
rect 22744 8570 22796 8576
rect 22284 8492 22336 8498
rect 22284 8434 22336 8440
rect 22100 7880 22152 7886
rect 22100 7822 22152 7828
rect 22112 7546 22140 7822
rect 22100 7540 22152 7546
rect 22100 7482 22152 7488
rect 21456 7472 21508 7478
rect 21456 7414 21508 7420
rect 21180 7200 21232 7206
rect 21180 7142 21232 7148
rect 19156 6724 19208 6730
rect 19156 6666 19208 6672
rect 19800 6656 19852 6662
rect 19800 6598 19852 6604
rect 18696 6248 18748 6254
rect 18696 6190 18748 6196
rect 19064 6248 19116 6254
rect 19064 6190 19116 6196
rect 18512 5364 18564 5370
rect 18512 5306 18564 5312
rect 18708 5358 19012 5386
rect 19076 5370 19104 6190
rect 18510 4856 18566 4865
rect 18510 4791 18512 4800
rect 18564 4791 18566 4800
rect 18512 4762 18564 4768
rect 18524 4078 18552 4762
rect 18708 4758 18736 5358
rect 18788 5228 18840 5234
rect 18788 5170 18840 5176
rect 18880 5228 18932 5234
rect 18880 5170 18932 5176
rect 18696 4752 18748 4758
rect 18696 4694 18748 4700
rect 18800 4486 18828 5170
rect 18892 5030 18920 5170
rect 18984 5030 19012 5358
rect 19064 5364 19116 5370
rect 19064 5306 19116 5312
rect 19432 5364 19484 5370
rect 19432 5306 19484 5312
rect 19444 5166 19472 5306
rect 19812 5302 19840 6598
rect 20444 6384 20496 6390
rect 20444 6326 20496 6332
rect 20456 5370 20484 6326
rect 21192 6254 21220 7142
rect 21180 6248 21232 6254
rect 21180 6190 21232 6196
rect 21192 5710 21220 6190
rect 21180 5704 21232 5710
rect 21180 5646 21232 5652
rect 20444 5364 20496 5370
rect 20444 5306 20496 5312
rect 19524 5296 19576 5302
rect 19524 5238 19576 5244
rect 19800 5296 19852 5302
rect 19800 5238 19852 5244
rect 19432 5160 19484 5166
rect 19432 5102 19484 5108
rect 18880 5024 18932 5030
rect 18880 4966 18932 4972
rect 18972 5024 19024 5030
rect 18972 4966 19024 4972
rect 18788 4480 18840 4486
rect 18788 4422 18840 4428
rect 18892 4214 18920 4966
rect 18880 4208 18932 4214
rect 18880 4150 18932 4156
rect 18512 4072 18564 4078
rect 18512 4014 18564 4020
rect 18328 3936 18380 3942
rect 18328 3878 18380 3884
rect 17592 3732 17644 3738
rect 17592 3674 17644 3680
rect 17960 3732 18012 3738
rect 17960 3674 18012 3680
rect 17408 3528 17460 3534
rect 17328 3488 17408 3516
rect 17408 3470 17460 3476
rect 17132 3460 17184 3466
rect 17132 3402 17184 3408
rect 17144 3058 17172 3402
rect 17132 3052 17184 3058
rect 17132 2994 17184 3000
rect 17040 2984 17092 2990
rect 17040 2926 17092 2932
rect 18340 2854 18368 3878
rect 18984 3194 19012 4966
rect 19444 4758 19472 5102
rect 19432 4752 19484 4758
rect 19062 4720 19118 4729
rect 19432 4694 19484 4700
rect 19062 4655 19118 4664
rect 19076 4622 19104 4655
rect 19064 4616 19116 4622
rect 19064 4558 19116 4564
rect 19248 4548 19300 4554
rect 19248 4490 19300 4496
rect 19260 3738 19288 4490
rect 19444 4078 19472 4694
rect 19536 4486 19564 5238
rect 19616 5092 19668 5098
rect 19616 5034 19668 5040
rect 19628 4622 19656 5034
rect 19812 4690 19840 5238
rect 20168 5092 20220 5098
rect 20168 5034 20220 5040
rect 19800 4684 19852 4690
rect 19800 4626 19852 4632
rect 19616 4616 19668 4622
rect 19616 4558 19668 4564
rect 19812 4570 19840 4626
rect 20180 4622 20208 5034
rect 20456 4622 20484 5306
rect 20168 4616 20220 4622
rect 19524 4480 19576 4486
rect 19628 4468 19656 4558
rect 19812 4542 19932 4570
rect 20168 4558 20220 4564
rect 20444 4616 20496 4622
rect 20444 4558 20496 4564
rect 19628 4440 19840 4468
rect 19524 4422 19576 4428
rect 19536 4282 19564 4422
rect 19524 4276 19576 4282
rect 19524 4218 19576 4224
rect 19432 4072 19484 4078
rect 19432 4014 19484 4020
rect 19248 3732 19300 3738
rect 19248 3674 19300 3680
rect 19340 3460 19392 3466
rect 19340 3402 19392 3408
rect 18972 3188 19024 3194
rect 18972 3130 19024 3136
rect 19352 3058 19380 3402
rect 19444 3398 19472 4014
rect 19432 3392 19484 3398
rect 19432 3334 19484 3340
rect 19536 3194 19564 4218
rect 19708 4208 19760 4214
rect 19708 4150 19760 4156
rect 19720 3602 19748 4150
rect 19812 3738 19840 4440
rect 19904 4146 19932 4542
rect 19984 4480 20036 4486
rect 19984 4422 20036 4428
rect 19892 4140 19944 4146
rect 19892 4082 19944 4088
rect 19800 3732 19852 3738
rect 19800 3674 19852 3680
rect 19812 3602 19840 3674
rect 19708 3596 19760 3602
rect 19708 3538 19760 3544
rect 19800 3596 19852 3602
rect 19800 3538 19852 3544
rect 19524 3188 19576 3194
rect 19524 3130 19576 3136
rect 19720 3074 19748 3538
rect 19904 3466 19932 4082
rect 19996 3942 20024 4422
rect 20180 4146 20208 4558
rect 20260 4480 20312 4486
rect 20260 4422 20312 4428
rect 20996 4480 21048 4486
rect 20996 4422 21048 4428
rect 20272 4146 20300 4422
rect 21008 4146 21036 4422
rect 20168 4140 20220 4146
rect 20168 4082 20220 4088
rect 20260 4140 20312 4146
rect 20260 4082 20312 4088
rect 20628 4140 20680 4146
rect 20628 4082 20680 4088
rect 20996 4140 21048 4146
rect 20996 4082 21048 4088
rect 19984 3936 20036 3942
rect 19984 3878 20036 3884
rect 19892 3460 19944 3466
rect 19892 3402 19944 3408
rect 19628 3058 19748 3074
rect 19996 3058 20024 3878
rect 20180 3534 20208 4082
rect 20536 3936 20588 3942
rect 20536 3878 20588 3884
rect 20548 3534 20576 3878
rect 20640 3738 20668 4082
rect 20628 3732 20680 3738
rect 20628 3674 20680 3680
rect 21008 3670 21036 4082
rect 20996 3664 21048 3670
rect 20996 3606 21048 3612
rect 20168 3528 20220 3534
rect 20168 3470 20220 3476
rect 20536 3528 20588 3534
rect 21192 3516 21220 5646
rect 21272 3528 21324 3534
rect 21192 3488 21272 3516
rect 20536 3470 20588 3476
rect 21272 3470 21324 3476
rect 20548 3126 20576 3470
rect 20536 3120 20588 3126
rect 20536 3062 20588 3068
rect 21284 3058 21312 3470
rect 19340 3052 19392 3058
rect 19340 2994 19392 3000
rect 19616 3052 19748 3058
rect 19668 3046 19748 3052
rect 19984 3052 20036 3058
rect 19616 2994 19668 3000
rect 19984 2994 20036 3000
rect 21272 3052 21324 3058
rect 21272 2994 21324 3000
rect 21468 2854 21496 7414
rect 22296 6458 22324 8434
rect 23676 8430 23704 9522
rect 24032 9036 24084 9042
rect 24032 8978 24084 8984
rect 23940 8492 23992 8498
rect 23940 8434 23992 8440
rect 23664 8424 23716 8430
rect 23664 8366 23716 8372
rect 23572 6724 23624 6730
rect 23572 6666 23624 6672
rect 23584 6458 23612 6666
rect 22284 6452 22336 6458
rect 22284 6394 22336 6400
rect 23572 6452 23624 6458
rect 23572 6394 23624 6400
rect 22560 6384 22612 6390
rect 22560 6326 22612 6332
rect 22572 5710 22600 6326
rect 23480 6180 23532 6186
rect 23480 6122 23532 6128
rect 23492 5710 23520 6122
rect 23676 5930 23704 8366
rect 23952 7818 23980 8434
rect 23940 7812 23992 7818
rect 23940 7754 23992 7760
rect 23848 7744 23900 7750
rect 23848 7686 23900 7692
rect 23860 6322 23888 7686
rect 23848 6316 23900 6322
rect 23848 6258 23900 6264
rect 23756 6112 23808 6118
rect 23756 6054 23808 6060
rect 23584 5902 23704 5930
rect 22560 5704 22612 5710
rect 22560 5646 22612 5652
rect 23480 5704 23532 5710
rect 23480 5646 23532 5652
rect 22284 5364 22336 5370
rect 22284 5306 22336 5312
rect 22296 5114 22324 5306
rect 22572 5302 22600 5646
rect 22560 5296 22612 5302
rect 22560 5238 22612 5244
rect 22204 5098 22324 5114
rect 22192 5092 22324 5098
rect 22244 5086 22324 5092
rect 22192 5034 22244 5040
rect 22572 4554 22600 5238
rect 23584 5166 23612 5902
rect 23768 5710 23796 6054
rect 23756 5704 23808 5710
rect 23756 5646 23808 5652
rect 23768 5370 23796 5646
rect 23756 5364 23808 5370
rect 23756 5306 23808 5312
rect 23860 5234 23888 6258
rect 23848 5228 23900 5234
rect 23848 5170 23900 5176
rect 23572 5160 23624 5166
rect 23952 5114 23980 7754
rect 24044 6322 24072 8978
rect 24688 8974 24716 12582
rect 24768 9988 24820 9994
rect 24768 9930 24820 9936
rect 24780 9586 24808 9930
rect 24768 9580 24820 9586
rect 24768 9522 24820 9528
rect 24308 8968 24360 8974
rect 24308 8910 24360 8916
rect 24676 8968 24728 8974
rect 24676 8910 24728 8916
rect 24124 8628 24176 8634
rect 24124 8570 24176 8576
rect 24136 8022 24164 8570
rect 24216 8424 24268 8430
rect 24216 8366 24268 8372
rect 24124 8016 24176 8022
rect 24124 7958 24176 7964
rect 24228 7970 24256 8366
rect 24320 8294 24348 8910
rect 24492 8900 24544 8906
rect 24492 8842 24544 8848
rect 24308 8288 24360 8294
rect 24308 8230 24360 8236
rect 24400 8288 24452 8294
rect 24400 8230 24452 8236
rect 24320 8090 24348 8230
rect 24308 8084 24360 8090
rect 24308 8026 24360 8032
rect 24228 7942 24348 7970
rect 24320 7886 24348 7942
rect 24308 7880 24360 7886
rect 24308 7822 24360 7828
rect 24320 7546 24348 7822
rect 24308 7540 24360 7546
rect 24308 7482 24360 7488
rect 24216 6724 24268 6730
rect 24216 6666 24268 6672
rect 24124 6656 24176 6662
rect 24124 6598 24176 6604
rect 24136 6322 24164 6598
rect 24032 6316 24084 6322
rect 24032 6258 24084 6264
rect 24124 6316 24176 6322
rect 24124 6258 24176 6264
rect 24228 5846 24256 6666
rect 24216 5840 24268 5846
rect 24216 5782 24268 5788
rect 23572 5102 23624 5108
rect 23584 4690 23612 5102
rect 23860 5086 23980 5114
rect 23572 4684 23624 4690
rect 23572 4626 23624 4632
rect 22560 4548 22612 4554
rect 22560 4490 22612 4496
rect 22572 4282 22600 4490
rect 22560 4276 22612 4282
rect 22560 4218 22612 4224
rect 21548 3596 21600 3602
rect 21548 3538 21600 3544
rect 21560 3466 21588 3538
rect 22572 3466 22600 4218
rect 23584 4214 23612 4626
rect 23572 4208 23624 4214
rect 23572 4150 23624 4156
rect 23296 4072 23348 4078
rect 23296 4014 23348 4020
rect 23308 3534 23336 4014
rect 23584 3602 23612 4150
rect 23572 3596 23624 3602
rect 23572 3538 23624 3544
rect 22836 3528 22888 3534
rect 22836 3470 22888 3476
rect 23296 3528 23348 3534
rect 23296 3470 23348 3476
rect 23388 3528 23440 3534
rect 23388 3470 23440 3476
rect 21548 3460 21600 3466
rect 21548 3402 21600 3408
rect 22560 3460 22612 3466
rect 22560 3402 22612 3408
rect 14556 2848 14608 2854
rect 14556 2790 14608 2796
rect 18328 2848 18380 2854
rect 18328 2790 18380 2796
rect 21456 2848 21508 2854
rect 21456 2790 21508 2796
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 21560 2650 21588 3402
rect 22572 3126 22600 3402
rect 22560 3120 22612 3126
rect 22560 3062 22612 3068
rect 22192 2984 22244 2990
rect 22192 2926 22244 2932
rect 22204 2650 22232 2926
rect 22848 2650 22876 3470
rect 23400 2990 23428 3470
rect 23584 3058 23612 3538
rect 23860 3194 23888 5086
rect 23940 3460 23992 3466
rect 23940 3402 23992 3408
rect 23848 3188 23900 3194
rect 23848 3130 23900 3136
rect 23572 3052 23624 3058
rect 23572 2994 23624 3000
rect 23388 2984 23440 2990
rect 23388 2926 23440 2932
rect 23952 2854 23980 3402
rect 24320 3398 24348 7482
rect 24412 7410 24440 8230
rect 24504 7886 24532 8842
rect 24584 8832 24636 8838
rect 24584 8774 24636 8780
rect 24676 8832 24728 8838
rect 24676 8774 24728 8780
rect 24596 8634 24624 8774
rect 24584 8628 24636 8634
rect 24584 8570 24636 8576
rect 24688 8566 24716 8774
rect 24676 8560 24728 8566
rect 24676 8502 24728 8508
rect 24768 8424 24820 8430
rect 24768 8366 24820 8372
rect 24676 8356 24728 8362
rect 24676 8298 24728 8304
rect 24688 8022 24716 8298
rect 24676 8016 24728 8022
rect 24582 7984 24638 7993
rect 24676 7958 24728 7964
rect 24582 7919 24584 7928
rect 24636 7919 24638 7928
rect 24584 7890 24636 7896
rect 24492 7880 24544 7886
rect 24492 7822 24544 7828
rect 24688 7478 24716 7958
rect 24676 7472 24728 7478
rect 24676 7414 24728 7420
rect 24400 7404 24452 7410
rect 24400 7346 24452 7352
rect 24400 7200 24452 7206
rect 24400 7142 24452 7148
rect 24412 5778 24440 7142
rect 24584 6316 24636 6322
rect 24584 6258 24636 6264
rect 24596 5914 24624 6258
rect 24780 6186 24808 8366
rect 24872 7954 24900 13670
rect 25516 12170 25544 13874
rect 26528 13394 26556 14010
rect 27068 14000 27120 14006
rect 27068 13942 27120 13948
rect 26516 13388 26568 13394
rect 26516 13330 26568 13336
rect 26528 12850 26556 13330
rect 26976 13184 27028 13190
rect 26976 13126 27028 13132
rect 26792 12912 26844 12918
rect 26792 12854 26844 12860
rect 26516 12844 26568 12850
rect 26516 12786 26568 12792
rect 26608 12844 26660 12850
rect 26608 12786 26660 12792
rect 26528 12306 26556 12786
rect 26240 12300 26292 12306
rect 26240 12242 26292 12248
rect 26516 12300 26568 12306
rect 26516 12242 26568 12248
rect 25504 12164 25556 12170
rect 25504 12106 25556 12112
rect 25516 11898 25544 12106
rect 25504 11892 25556 11898
rect 25504 11834 25556 11840
rect 26252 11830 26280 12242
rect 26240 11824 26292 11830
rect 26240 11766 26292 11772
rect 25044 11552 25096 11558
rect 25044 11494 25096 11500
rect 25056 8974 25084 11494
rect 26252 11218 26280 11766
rect 26516 11552 26568 11558
rect 26516 11494 26568 11500
rect 26240 11212 26292 11218
rect 26240 11154 26292 11160
rect 26252 10742 26280 11154
rect 26240 10736 26292 10742
rect 26240 10678 26292 10684
rect 26424 10736 26476 10742
rect 26424 10678 26476 10684
rect 26252 10130 26280 10678
rect 26240 10124 26292 10130
rect 26240 10066 26292 10072
rect 26436 10062 26464 10678
rect 26424 10056 26476 10062
rect 26424 9998 26476 10004
rect 26332 9920 26384 9926
rect 26332 9862 26384 9868
rect 26344 9586 26372 9862
rect 26240 9580 26292 9586
rect 26240 9522 26292 9528
rect 26332 9580 26384 9586
rect 26332 9522 26384 9528
rect 25688 9444 25740 9450
rect 25688 9386 25740 9392
rect 25320 9104 25372 9110
rect 25320 9046 25372 9052
rect 25044 8968 25096 8974
rect 25044 8910 25096 8916
rect 25056 8566 25084 8910
rect 25228 8900 25280 8906
rect 25228 8842 25280 8848
rect 25044 8560 25096 8566
rect 25096 8508 25176 8514
rect 25044 8502 25176 8508
rect 25056 8486 25176 8502
rect 25240 8498 25268 8842
rect 25332 8498 25360 9046
rect 25700 8498 25728 9386
rect 25872 9376 25924 9382
rect 25872 9318 25924 9324
rect 25884 9042 25912 9318
rect 26252 9110 26280 9522
rect 26240 9104 26292 9110
rect 26240 9046 26292 9052
rect 25872 9036 25924 9042
rect 25872 8978 25924 8984
rect 26056 8968 26108 8974
rect 26056 8910 26108 8916
rect 26332 8968 26384 8974
rect 26332 8910 26384 8916
rect 26068 8616 26096 8910
rect 25976 8588 26096 8616
rect 25044 8424 25096 8430
rect 25044 8366 25096 8372
rect 24952 8356 25004 8362
rect 24952 8298 25004 8304
rect 24860 7948 24912 7954
rect 24860 7890 24912 7896
rect 24872 6458 24900 7890
rect 24860 6452 24912 6458
rect 24860 6394 24912 6400
rect 24768 6180 24820 6186
rect 24768 6122 24820 6128
rect 24584 5908 24636 5914
rect 24584 5850 24636 5856
rect 24872 5846 24900 6394
rect 24860 5840 24912 5846
rect 24860 5782 24912 5788
rect 24400 5772 24452 5778
rect 24400 5714 24452 5720
rect 24676 5704 24728 5710
rect 24676 5646 24728 5652
rect 24860 5704 24912 5710
rect 24860 5646 24912 5652
rect 24400 5568 24452 5574
rect 24400 5510 24452 5516
rect 24412 5302 24440 5510
rect 24688 5302 24716 5646
rect 24872 5370 24900 5646
rect 24860 5364 24912 5370
rect 24860 5306 24912 5312
rect 24400 5296 24452 5302
rect 24400 5238 24452 5244
rect 24676 5296 24728 5302
rect 24676 5238 24728 5244
rect 24964 5234 24992 8298
rect 25056 7993 25084 8366
rect 25042 7984 25098 7993
rect 25042 7919 25098 7928
rect 25148 7886 25176 8486
rect 25228 8492 25280 8498
rect 25228 8434 25280 8440
rect 25320 8492 25372 8498
rect 25320 8434 25372 8440
rect 25688 8492 25740 8498
rect 25688 8434 25740 8440
rect 25412 8424 25464 8430
rect 25412 8366 25464 8372
rect 25424 8090 25452 8366
rect 25412 8084 25464 8090
rect 25412 8026 25464 8032
rect 25228 7948 25280 7954
rect 25228 7890 25280 7896
rect 25136 7880 25188 7886
rect 25136 7822 25188 7828
rect 25240 7546 25268 7890
rect 25688 7812 25740 7818
rect 25688 7754 25740 7760
rect 25228 7540 25280 7546
rect 25228 7482 25280 7488
rect 25700 7478 25728 7754
rect 25688 7472 25740 7478
rect 25688 7414 25740 7420
rect 25504 7200 25556 7206
rect 25504 7142 25556 7148
rect 25044 6316 25096 6322
rect 25044 6258 25096 6264
rect 25056 5914 25084 6258
rect 25044 5908 25096 5914
rect 25044 5850 25096 5856
rect 25056 5710 25084 5850
rect 25044 5704 25096 5710
rect 25044 5646 25096 5652
rect 25412 5704 25464 5710
rect 25412 5646 25464 5652
rect 25056 5234 25084 5646
rect 24952 5228 25004 5234
rect 24952 5170 25004 5176
rect 25044 5228 25096 5234
rect 25044 5170 25096 5176
rect 24860 5160 24912 5166
rect 24860 5102 24912 5108
rect 24400 5024 24452 5030
rect 24400 4966 24452 4972
rect 24412 4758 24440 4966
rect 24872 4826 24900 5102
rect 24860 4820 24912 4826
rect 24860 4762 24912 4768
rect 24400 4752 24452 4758
rect 24400 4694 24452 4700
rect 25424 4078 25452 5646
rect 25516 5642 25544 7142
rect 25504 5636 25556 5642
rect 25504 5578 25556 5584
rect 25516 5234 25544 5578
rect 25976 5370 26004 8588
rect 26056 8492 26108 8498
rect 26056 8434 26108 8440
rect 26068 7546 26096 8434
rect 26344 8430 26372 8910
rect 26332 8424 26384 8430
rect 26332 8366 26384 8372
rect 26344 8090 26372 8366
rect 26528 8090 26556 11494
rect 26620 11218 26648 12786
rect 26608 11212 26660 11218
rect 26608 11154 26660 11160
rect 26804 10810 26832 12854
rect 26884 12640 26936 12646
rect 26884 12582 26936 12588
rect 26896 11762 26924 12582
rect 26884 11756 26936 11762
rect 26884 11698 26936 11704
rect 26792 10804 26844 10810
rect 26792 10746 26844 10752
rect 26988 10742 27016 13126
rect 27080 11558 27108 13942
rect 27172 12646 27200 15302
rect 27436 14272 27488 14278
rect 27436 14214 27488 14220
rect 27448 13938 27476 14214
rect 27528 14068 27580 14074
rect 27528 14010 27580 14016
rect 27436 13932 27488 13938
rect 27436 13874 27488 13880
rect 27344 13864 27396 13870
rect 27344 13806 27396 13812
rect 27160 12640 27212 12646
rect 27160 12582 27212 12588
rect 27172 12102 27200 12582
rect 27160 12096 27212 12102
rect 27160 12038 27212 12044
rect 27356 11898 27384 13806
rect 27436 12912 27488 12918
rect 27436 12854 27488 12860
rect 27344 11892 27396 11898
rect 27344 11834 27396 11840
rect 27160 11756 27212 11762
rect 27160 11698 27212 11704
rect 27068 11552 27120 11558
rect 27068 11494 27120 11500
rect 26976 10736 27028 10742
rect 26976 10678 27028 10684
rect 26792 9580 26844 9586
rect 26792 9522 26844 9528
rect 26700 9172 26752 9178
rect 26700 9114 26752 9120
rect 26608 8832 26660 8838
rect 26608 8774 26660 8780
rect 26332 8084 26384 8090
rect 26332 8026 26384 8032
rect 26516 8084 26568 8090
rect 26516 8026 26568 8032
rect 26620 7954 26648 8774
rect 26332 7948 26384 7954
rect 26332 7890 26384 7896
rect 26608 7948 26660 7954
rect 26608 7890 26660 7896
rect 26056 7540 26108 7546
rect 26056 7482 26108 7488
rect 26344 7410 26372 7890
rect 26516 7880 26568 7886
rect 26516 7822 26568 7828
rect 26332 7404 26384 7410
rect 26332 7346 26384 7352
rect 26424 7404 26476 7410
rect 26424 7346 26476 7352
rect 26240 7336 26292 7342
rect 26240 7278 26292 7284
rect 26252 6322 26280 7278
rect 26344 7274 26372 7346
rect 26332 7268 26384 7274
rect 26332 7210 26384 7216
rect 26240 6316 26292 6322
rect 26240 6258 26292 6264
rect 26240 6180 26292 6186
rect 26240 6122 26292 6128
rect 26148 6112 26200 6118
rect 26148 6054 26200 6060
rect 26160 5914 26188 6054
rect 26148 5908 26200 5914
rect 26148 5850 26200 5856
rect 26252 5642 26280 6122
rect 26240 5636 26292 5642
rect 26240 5578 26292 5584
rect 25964 5364 26016 5370
rect 25964 5306 26016 5312
rect 26252 5302 26280 5578
rect 26240 5296 26292 5302
rect 26240 5238 26292 5244
rect 25504 5228 25556 5234
rect 25504 5170 25556 5176
rect 25504 5024 25556 5030
rect 25504 4966 25556 4972
rect 25516 4826 25544 4966
rect 26252 4826 26280 5238
rect 26332 5024 26384 5030
rect 26332 4966 26384 4972
rect 25504 4820 25556 4826
rect 25504 4762 25556 4768
rect 25872 4820 25924 4826
rect 25872 4762 25924 4768
rect 26240 4820 26292 4826
rect 26240 4762 26292 4768
rect 25884 4146 25912 4762
rect 25964 4616 26016 4622
rect 25964 4558 26016 4564
rect 25976 4282 26004 4558
rect 26240 4480 26292 4486
rect 26240 4422 26292 4428
rect 26252 4282 26280 4422
rect 25964 4276 26016 4282
rect 25964 4218 26016 4224
rect 26240 4276 26292 4282
rect 26240 4218 26292 4224
rect 25872 4140 25924 4146
rect 25872 4082 25924 4088
rect 25964 4140 26016 4146
rect 25964 4082 26016 4088
rect 25412 4072 25464 4078
rect 25412 4014 25464 4020
rect 25596 4004 25648 4010
rect 25596 3946 25648 3952
rect 25320 3664 25372 3670
rect 25320 3606 25372 3612
rect 25332 3534 25360 3606
rect 25320 3528 25372 3534
rect 25320 3470 25372 3476
rect 24308 3392 24360 3398
rect 24308 3334 24360 3340
rect 24400 3392 24452 3398
rect 24400 3334 24452 3340
rect 24412 3126 24440 3334
rect 25332 3194 25360 3470
rect 25608 3466 25636 3946
rect 25688 3936 25740 3942
rect 25688 3878 25740 3884
rect 25700 3466 25728 3878
rect 25976 3670 26004 4082
rect 25964 3664 26016 3670
rect 25964 3606 26016 3612
rect 25596 3460 25648 3466
rect 25596 3402 25648 3408
rect 25688 3460 25740 3466
rect 25688 3402 25740 3408
rect 25320 3188 25372 3194
rect 25320 3130 25372 3136
rect 24400 3120 24452 3126
rect 24400 3062 24452 3068
rect 25700 2990 25728 3402
rect 25976 3058 26004 3606
rect 26252 3534 26280 4218
rect 26344 3738 26372 4966
rect 26332 3732 26384 3738
rect 26332 3674 26384 3680
rect 26240 3528 26292 3534
rect 26240 3470 26292 3476
rect 26252 3194 26280 3470
rect 26436 3194 26464 7346
rect 26528 5914 26556 7822
rect 26712 6730 26740 9114
rect 26804 9042 26832 9522
rect 26884 9512 26936 9518
rect 26884 9454 26936 9460
rect 26988 9466 27016 10678
rect 26896 9178 26924 9454
rect 26988 9438 27108 9466
rect 27080 9382 27108 9438
rect 26976 9376 27028 9382
rect 26976 9318 27028 9324
rect 27068 9376 27120 9382
rect 27068 9318 27120 9324
rect 26884 9172 26936 9178
rect 26884 9114 26936 9120
rect 26896 9042 26924 9114
rect 26792 9036 26844 9042
rect 26792 8978 26844 8984
rect 26884 9036 26936 9042
rect 26884 8978 26936 8984
rect 26988 8974 27016 9318
rect 27068 9104 27120 9110
rect 27068 9046 27120 9052
rect 27080 8974 27108 9046
rect 26976 8968 27028 8974
rect 26976 8910 27028 8916
rect 27068 8968 27120 8974
rect 27068 8910 27120 8916
rect 26884 8084 26936 8090
rect 26884 8026 26936 8032
rect 26792 8016 26844 8022
rect 26792 7958 26844 7964
rect 26700 6724 26752 6730
rect 26700 6666 26752 6672
rect 26608 6656 26660 6662
rect 26608 6598 26660 6604
rect 26516 5908 26568 5914
rect 26516 5850 26568 5856
rect 26516 5568 26568 5574
rect 26516 5510 26568 5516
rect 26528 5234 26556 5510
rect 26516 5228 26568 5234
rect 26516 5170 26568 5176
rect 26620 4622 26648 6598
rect 26804 6322 26832 7958
rect 26792 6316 26844 6322
rect 26792 6258 26844 6264
rect 26700 5908 26752 5914
rect 26700 5850 26752 5856
rect 26712 4690 26740 5850
rect 26804 5166 26832 6258
rect 26792 5160 26844 5166
rect 26792 5102 26844 5108
rect 26700 4684 26752 4690
rect 26700 4626 26752 4632
rect 26608 4616 26660 4622
rect 26608 4558 26660 4564
rect 26620 4214 26648 4558
rect 26804 4282 26832 5102
rect 26792 4276 26844 4282
rect 26792 4218 26844 4224
rect 26608 4208 26660 4214
rect 26608 4150 26660 4156
rect 26516 4072 26568 4078
rect 26516 4014 26568 4020
rect 26528 3738 26556 4014
rect 26516 3732 26568 3738
rect 26516 3674 26568 3680
rect 26528 3466 26556 3674
rect 26896 3670 26924 8026
rect 27172 6458 27200 11698
rect 27448 11694 27476 12854
rect 27540 12782 27568 14010
rect 27632 13802 27660 15846
rect 27804 15496 27856 15502
rect 27804 15438 27856 15444
rect 27816 15065 27844 15438
rect 27896 15428 27948 15434
rect 27896 15370 27948 15376
rect 27908 15094 27936 15370
rect 27896 15088 27948 15094
rect 27802 15056 27858 15065
rect 27896 15030 27948 15036
rect 27802 14991 27858 15000
rect 28000 14482 28028 20198
rect 28276 20058 28304 21422
rect 28368 20466 28396 22646
rect 28448 21956 28500 21962
rect 28448 21898 28500 21904
rect 28356 20460 28408 20466
rect 28356 20402 28408 20408
rect 28460 20330 28488 21898
rect 28448 20324 28500 20330
rect 28448 20266 28500 20272
rect 28264 20052 28316 20058
rect 28264 19994 28316 20000
rect 28460 19854 28488 20266
rect 28080 19848 28132 19854
rect 28080 19790 28132 19796
rect 28448 19848 28500 19854
rect 28448 19790 28500 19796
rect 28092 17270 28120 19790
rect 28264 17536 28316 17542
rect 28264 17478 28316 17484
rect 28080 17264 28132 17270
rect 28080 17206 28132 17212
rect 28092 15162 28120 17206
rect 28276 16658 28304 17478
rect 28264 16652 28316 16658
rect 28264 16594 28316 16600
rect 28356 16108 28408 16114
rect 28356 16050 28408 16056
rect 28368 15745 28396 16050
rect 28354 15736 28410 15745
rect 28354 15671 28410 15680
rect 28172 15428 28224 15434
rect 28172 15370 28224 15376
rect 28080 15156 28132 15162
rect 28080 15098 28132 15104
rect 27988 14476 28040 14482
rect 27988 14418 28040 14424
rect 28092 14346 28120 15098
rect 28080 14340 28132 14346
rect 28080 14282 28132 14288
rect 27988 13932 28040 13938
rect 27988 13874 28040 13880
rect 27620 13796 27672 13802
rect 27620 13738 27672 13744
rect 27632 13410 27660 13738
rect 28000 13705 28028 13874
rect 27986 13696 28042 13705
rect 27986 13631 28042 13640
rect 27632 13394 27844 13410
rect 27632 13388 27856 13394
rect 27632 13382 27804 13388
rect 27804 13330 27856 13336
rect 27804 13252 27856 13258
rect 27804 13194 27856 13200
rect 27528 12776 27580 12782
rect 27528 12718 27580 12724
rect 27816 12434 27844 13194
rect 28080 12844 28132 12850
rect 28080 12786 28132 12792
rect 27816 12406 27936 12434
rect 27908 12170 27936 12406
rect 28092 12345 28120 12786
rect 28184 12434 28212 15370
rect 28262 14376 28318 14385
rect 28262 14311 28318 14320
rect 28276 14074 28304 14311
rect 28264 14068 28316 14074
rect 28264 14010 28316 14016
rect 28354 13016 28410 13025
rect 28354 12951 28410 12960
rect 28368 12850 28396 12951
rect 28356 12844 28408 12850
rect 28356 12786 28408 12792
rect 28184 12406 28304 12434
rect 28078 12336 28134 12345
rect 28078 12271 28134 12280
rect 27896 12164 27948 12170
rect 27896 12106 27948 12112
rect 27908 11830 27936 12106
rect 28172 12096 28224 12102
rect 28172 12038 28224 12044
rect 27896 11824 27948 11830
rect 27896 11766 27948 11772
rect 27436 11688 27488 11694
rect 27436 11630 27488 11636
rect 27344 11552 27396 11558
rect 27344 11494 27396 11500
rect 27252 10600 27304 10606
rect 27252 10542 27304 10548
rect 27264 6730 27292 10542
rect 27356 10130 27384 11494
rect 27908 11082 27936 11766
rect 28080 11212 28132 11218
rect 28080 11154 28132 11160
rect 27896 11076 27948 11082
rect 27896 11018 27948 11024
rect 27528 10668 27580 10674
rect 27528 10610 27580 10616
rect 27436 10464 27488 10470
rect 27436 10406 27488 10412
rect 27344 10124 27396 10130
rect 27344 10066 27396 10072
rect 27448 9722 27476 10406
rect 27540 9926 27568 10610
rect 27908 10470 27936 11018
rect 27896 10464 27948 10470
rect 27896 10406 27948 10412
rect 27908 10062 27936 10406
rect 27896 10056 27948 10062
rect 27896 9998 27948 10004
rect 27528 9920 27580 9926
rect 27528 9862 27580 9868
rect 27436 9716 27488 9722
rect 27436 9658 27488 9664
rect 27448 9382 27476 9658
rect 27540 9586 27568 9862
rect 28092 9586 28120 11154
rect 28184 9586 28212 12038
rect 27528 9580 27580 9586
rect 27528 9522 27580 9528
rect 28080 9580 28132 9586
rect 28080 9522 28132 9528
rect 28172 9580 28224 9586
rect 28172 9522 28224 9528
rect 27436 9376 27488 9382
rect 27436 9318 27488 9324
rect 27448 8974 27476 9318
rect 27436 8968 27488 8974
rect 27436 8910 27488 8916
rect 28092 8906 28120 9522
rect 28184 9110 28212 9522
rect 28172 9104 28224 9110
rect 28172 9046 28224 9052
rect 28080 8900 28132 8906
rect 28080 8842 28132 8848
rect 27528 7744 27580 7750
rect 27528 7686 27580 7692
rect 27540 7002 27568 7686
rect 27896 7200 27948 7206
rect 27896 7142 27948 7148
rect 27528 6996 27580 7002
rect 27528 6938 27580 6944
rect 27252 6724 27304 6730
rect 27252 6666 27304 6672
rect 27160 6452 27212 6458
rect 27160 6394 27212 6400
rect 27264 5642 27292 6666
rect 27540 6118 27568 6938
rect 27620 6316 27672 6322
rect 27620 6258 27672 6264
rect 27528 6112 27580 6118
rect 27528 6054 27580 6060
rect 27252 5636 27304 5642
rect 27252 5578 27304 5584
rect 27264 4554 27292 5578
rect 27632 5370 27660 6258
rect 27908 6186 27936 7142
rect 28276 6882 28304 12406
rect 28356 11756 28408 11762
rect 28356 11698 28408 11704
rect 28368 11665 28396 11698
rect 28354 11656 28410 11665
rect 28354 11591 28410 11600
rect 28356 7880 28408 7886
rect 28356 7822 28408 7828
rect 28368 7585 28396 7822
rect 28354 7576 28410 7585
rect 28354 7511 28410 7520
rect 28356 7404 28408 7410
rect 28356 7346 28408 7352
rect 28368 6905 28396 7346
rect 28184 6854 28304 6882
rect 28354 6896 28410 6905
rect 27988 6248 28040 6254
rect 27988 6190 28040 6196
rect 27896 6180 27948 6186
rect 27896 6122 27948 6128
rect 27620 5364 27672 5370
rect 27620 5306 27672 5312
rect 27252 4548 27304 4554
rect 27252 4490 27304 4496
rect 27264 4010 27292 4490
rect 27620 4140 27672 4146
rect 27620 4082 27672 4088
rect 27712 4140 27764 4146
rect 27712 4082 27764 4088
rect 27252 4004 27304 4010
rect 27172 3964 27252 3992
rect 26884 3664 26936 3670
rect 26884 3606 26936 3612
rect 26516 3460 26568 3466
rect 26516 3402 26568 3408
rect 26240 3188 26292 3194
rect 26240 3130 26292 3136
rect 26424 3188 26476 3194
rect 26424 3130 26476 3136
rect 25964 3052 26016 3058
rect 25964 2994 26016 3000
rect 25688 2984 25740 2990
rect 25688 2926 25740 2932
rect 26528 2854 26556 3402
rect 27172 3398 27200 3964
rect 27252 3946 27304 3952
rect 27436 4004 27488 4010
rect 27436 3946 27488 3952
rect 27448 3466 27476 3946
rect 27526 3496 27582 3505
rect 27436 3460 27488 3466
rect 27526 3431 27582 3440
rect 27436 3402 27488 3408
rect 27160 3392 27212 3398
rect 27160 3334 27212 3340
rect 27540 3058 27568 3431
rect 27528 3052 27580 3058
rect 27528 2994 27580 3000
rect 27632 2922 27660 4082
rect 27724 3194 27752 4082
rect 27908 3466 27936 6122
rect 28000 5778 28028 6190
rect 27988 5772 28040 5778
rect 27988 5714 28040 5720
rect 27988 5364 28040 5370
rect 27988 5306 28040 5312
rect 28000 4690 28028 5306
rect 27988 4684 28040 4690
rect 27988 4626 28040 4632
rect 28184 4010 28212 6854
rect 28354 6831 28410 6840
rect 28264 6792 28316 6798
rect 28264 6734 28316 6740
rect 28276 5710 28304 6734
rect 28356 6316 28408 6322
rect 28356 6258 28408 6264
rect 28368 6225 28396 6258
rect 28354 6216 28410 6225
rect 28354 6151 28410 6160
rect 28264 5704 28316 5710
rect 28264 5646 28316 5652
rect 28276 4622 28304 5646
rect 28354 5536 28410 5545
rect 28354 5471 28410 5480
rect 28368 5234 28396 5471
rect 28356 5228 28408 5234
rect 28356 5170 28408 5176
rect 28264 4616 28316 4622
rect 28264 4558 28316 4564
rect 28172 4004 28224 4010
rect 28172 3946 28224 3952
rect 27896 3460 27948 3466
rect 27896 3402 27948 3408
rect 28184 3233 28212 3946
rect 28276 3602 28304 4558
rect 28264 3596 28316 3602
rect 28264 3538 28316 3544
rect 28170 3224 28226 3233
rect 27712 3188 27764 3194
rect 28170 3159 28226 3168
rect 27712 3130 27764 3136
rect 28184 3126 28212 3159
rect 28172 3120 28224 3126
rect 28172 3062 28224 3068
rect 27620 2916 27672 2922
rect 27620 2858 27672 2864
rect 23940 2848 23992 2854
rect 23940 2790 23992 2796
rect 26516 2848 26568 2854
rect 26516 2790 26568 2796
rect 23952 2650 23980 2790
rect 21548 2644 21600 2650
rect 21548 2586 21600 2592
rect 22192 2644 22244 2650
rect 22192 2586 22244 2592
rect 22836 2644 22888 2650
rect 22836 2586 22888 2592
rect 23940 2644 23992 2650
rect 23940 2586 23992 2592
rect 21272 2440 21324 2446
rect 21272 2382 21324 2388
rect 21916 2440 21968 2446
rect 21916 2382 21968 2388
rect 22560 2440 22612 2446
rect 22560 2382 22612 2388
rect 23204 2440 23256 2446
rect 23204 2382 23256 2388
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 21284 800 21312 2382
rect 21928 800 21956 2382
rect 22572 800 22600 2382
rect 23216 800 23244 2382
rect 21270 0 21326 800
rect 21914 0 21970 800
rect 22558 0 22614 800
rect 23202 0 23258 800
<< via2 >>
rect 4880 29402 4936 29404
rect 4960 29402 5016 29404
rect 5040 29402 5096 29404
rect 5120 29402 5176 29404
rect 4880 29350 4926 29402
rect 4926 29350 4936 29402
rect 4960 29350 4990 29402
rect 4990 29350 5002 29402
rect 5002 29350 5016 29402
rect 5040 29350 5054 29402
rect 5054 29350 5066 29402
rect 5066 29350 5096 29402
rect 5120 29350 5130 29402
rect 5130 29350 5176 29402
rect 4880 29348 4936 29350
rect 4960 29348 5016 29350
rect 5040 29348 5096 29350
rect 5120 29348 5176 29350
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4880 28314 4936 28316
rect 4960 28314 5016 28316
rect 5040 28314 5096 28316
rect 5120 28314 5176 28316
rect 4880 28262 4926 28314
rect 4926 28262 4936 28314
rect 4960 28262 4990 28314
rect 4990 28262 5002 28314
rect 5002 28262 5016 28314
rect 5040 28262 5054 28314
rect 5054 28262 5066 28314
rect 5066 28262 5096 28314
rect 5120 28262 5130 28314
rect 5130 28262 5176 28314
rect 4880 28260 4936 28262
rect 4960 28260 5016 28262
rect 5040 28260 5096 28262
rect 5120 28260 5176 28262
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4880 27226 4936 27228
rect 4960 27226 5016 27228
rect 5040 27226 5096 27228
rect 5120 27226 5176 27228
rect 4880 27174 4926 27226
rect 4926 27174 4936 27226
rect 4960 27174 4990 27226
rect 4990 27174 5002 27226
rect 5002 27174 5016 27226
rect 5040 27174 5054 27226
rect 5054 27174 5066 27226
rect 5066 27174 5096 27226
rect 5120 27174 5130 27226
rect 5130 27174 5176 27226
rect 4880 27172 4936 27174
rect 4960 27172 5016 27174
rect 5040 27172 5096 27174
rect 5120 27172 5176 27174
rect 110 26968 166 27024
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4880 26138 4936 26140
rect 4960 26138 5016 26140
rect 5040 26138 5096 26140
rect 5120 26138 5176 26140
rect 4880 26086 4926 26138
rect 4926 26086 4936 26138
rect 4960 26086 4990 26138
rect 4990 26086 5002 26138
rect 5002 26086 5016 26138
rect 5040 26086 5054 26138
rect 5054 26086 5066 26138
rect 5066 26086 5096 26138
rect 5120 26086 5130 26138
rect 5130 26086 5176 26138
rect 4880 26084 4936 26086
rect 4960 26084 5016 26086
rect 5040 26084 5096 26086
rect 5120 26084 5176 26086
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4880 25050 4936 25052
rect 4960 25050 5016 25052
rect 5040 25050 5096 25052
rect 5120 25050 5176 25052
rect 4880 24998 4926 25050
rect 4926 24998 4936 25050
rect 4960 24998 4990 25050
rect 4990 24998 5002 25050
rect 5002 24998 5016 25050
rect 5040 24998 5054 25050
rect 5054 24998 5066 25050
rect 5066 24998 5096 25050
rect 5120 24998 5130 25050
rect 5130 24998 5176 25050
rect 4880 24996 4936 24998
rect 4960 24996 5016 24998
rect 5040 24996 5096 24998
rect 5120 24996 5176 24998
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4880 23962 4936 23964
rect 4960 23962 5016 23964
rect 5040 23962 5096 23964
rect 5120 23962 5176 23964
rect 4880 23910 4926 23962
rect 4926 23910 4936 23962
rect 4960 23910 4990 23962
rect 4990 23910 5002 23962
rect 5002 23910 5016 23962
rect 5040 23910 5054 23962
rect 5054 23910 5066 23962
rect 5066 23910 5096 23962
rect 5120 23910 5130 23962
rect 5130 23910 5176 23962
rect 4880 23908 4936 23910
rect 4960 23908 5016 23910
rect 5040 23908 5096 23910
rect 5120 23908 5176 23910
rect 4880 22874 4936 22876
rect 4960 22874 5016 22876
rect 5040 22874 5096 22876
rect 5120 22874 5176 22876
rect 4880 22822 4926 22874
rect 4926 22822 4936 22874
rect 4960 22822 4990 22874
rect 4990 22822 5002 22874
rect 5002 22822 5016 22874
rect 5040 22822 5054 22874
rect 5054 22822 5066 22874
rect 5066 22822 5096 22874
rect 5120 22822 5130 22874
rect 5130 22822 5176 22874
rect 4880 22820 4936 22822
rect 4960 22820 5016 22822
rect 5040 22820 5096 22822
rect 5120 22820 5176 22822
rect 11702 24132 11758 24168
rect 11702 24112 11704 24132
rect 11704 24112 11756 24132
rect 11756 24112 11758 24132
rect 5814 21936 5870 21992
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4880 21786 4936 21788
rect 4960 21786 5016 21788
rect 5040 21786 5096 21788
rect 5120 21786 5176 21788
rect 4880 21734 4926 21786
rect 4926 21734 4936 21786
rect 4960 21734 4990 21786
rect 4990 21734 5002 21786
rect 5002 21734 5016 21786
rect 5040 21734 5054 21786
rect 5054 21734 5066 21786
rect 5066 21734 5096 21786
rect 5120 21734 5130 21786
rect 5130 21734 5176 21786
rect 4880 21732 4936 21734
rect 4960 21732 5016 21734
rect 5040 21732 5096 21734
rect 5120 21732 5176 21734
rect 4880 20698 4936 20700
rect 4960 20698 5016 20700
rect 5040 20698 5096 20700
rect 5120 20698 5176 20700
rect 4880 20646 4926 20698
rect 4926 20646 4936 20698
rect 4960 20646 4990 20698
rect 4990 20646 5002 20698
rect 5002 20646 5016 20698
rect 5040 20646 5054 20698
rect 5054 20646 5066 20698
rect 5066 20646 5096 20698
rect 5120 20646 5130 20698
rect 5130 20646 5176 20698
rect 4880 20644 4936 20646
rect 4960 20644 5016 20646
rect 5040 20644 5096 20646
rect 5120 20644 5176 20646
rect 4880 19610 4936 19612
rect 4960 19610 5016 19612
rect 5040 19610 5096 19612
rect 5120 19610 5176 19612
rect 4880 19558 4926 19610
rect 4926 19558 4936 19610
rect 4960 19558 4990 19610
rect 4990 19558 5002 19610
rect 5002 19558 5016 19610
rect 5040 19558 5054 19610
rect 5054 19558 5066 19610
rect 5066 19558 5096 19610
rect 5120 19558 5130 19610
rect 5130 19558 5176 19610
rect 4880 19556 4936 19558
rect 4960 19556 5016 19558
rect 5040 19556 5096 19558
rect 5120 19556 5176 19558
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 5262 19372 5318 19408
rect 5262 19352 5264 19372
rect 5264 19352 5316 19372
rect 5316 19352 5318 19372
rect 4880 18522 4936 18524
rect 4960 18522 5016 18524
rect 5040 18522 5096 18524
rect 5120 18522 5176 18524
rect 4880 18470 4926 18522
rect 4926 18470 4936 18522
rect 4960 18470 4990 18522
rect 4990 18470 5002 18522
rect 5002 18470 5016 18522
rect 5040 18470 5054 18522
rect 5054 18470 5066 18522
rect 5066 18470 5096 18522
rect 5120 18470 5130 18522
rect 5130 18470 5176 18522
rect 4880 18468 4936 18470
rect 4960 18468 5016 18470
rect 5040 18468 5096 18470
rect 5120 18468 5176 18470
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 110 14320 166 14376
rect 4880 17434 4936 17436
rect 4960 17434 5016 17436
rect 5040 17434 5096 17436
rect 5120 17434 5176 17436
rect 4880 17382 4926 17434
rect 4926 17382 4936 17434
rect 4960 17382 4990 17434
rect 4990 17382 5002 17434
rect 5002 17382 5016 17434
rect 5040 17382 5054 17434
rect 5054 17382 5066 17434
rect 5066 17382 5096 17434
rect 5120 17382 5130 17434
rect 5130 17382 5176 17434
rect 4880 17380 4936 17382
rect 4960 17380 5016 17382
rect 5040 17380 5096 17382
rect 5120 17380 5176 17382
rect 4880 16346 4936 16348
rect 4960 16346 5016 16348
rect 5040 16346 5096 16348
rect 5120 16346 5176 16348
rect 4880 16294 4926 16346
rect 4926 16294 4936 16346
rect 4960 16294 4990 16346
rect 4990 16294 5002 16346
rect 5002 16294 5016 16346
rect 5040 16294 5054 16346
rect 5054 16294 5066 16346
rect 5066 16294 5096 16346
rect 5120 16294 5130 16346
rect 5130 16294 5176 16346
rect 4880 16292 4936 16294
rect 4960 16292 5016 16294
rect 5040 16292 5096 16294
rect 5120 16292 5176 16294
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 5446 14456 5502 14512
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 9586 20440 9642 20496
rect 8850 19352 8906 19408
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 4618 10648 4674 10704
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 8574 14456 8630 14512
rect 12622 24112 12678 24168
rect 12070 21972 12072 21992
rect 12072 21972 12124 21992
rect 12124 21972 12126 21992
rect 12070 21936 12126 21972
rect 9126 15020 9182 15056
rect 9126 15000 9128 15020
rect 9128 15000 9180 15020
rect 9180 15000 9182 15020
rect 9218 14900 9220 14920
rect 9220 14900 9272 14920
rect 9272 14900 9274 14920
rect 9218 14864 9274 14900
rect 9586 15020 9642 15056
rect 9586 15000 9588 15020
rect 9588 15000 9640 15020
rect 9640 15000 9642 15020
rect 10046 14864 10102 14920
rect 9862 11328 9918 11384
rect 8758 10684 8760 10704
rect 8760 10684 8812 10704
rect 8812 10684 8814 10704
rect 8758 10648 8814 10684
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 6550 8492 6606 8528
rect 6550 8472 6552 8492
rect 6552 8472 6604 8492
rect 6604 8472 6606 8492
rect 7286 8492 7342 8528
rect 7286 8472 7288 8492
rect 7288 8472 7340 8492
rect 7340 8472 7342 8492
rect 6826 8336 6882 8392
rect 7194 8336 7250 8392
rect 7654 8336 7710 8392
rect 6918 5480 6974 5536
rect 6090 4684 6146 4720
rect 6090 4664 6092 4684
rect 6092 4664 6144 4684
rect 6144 4664 6146 4684
rect 9678 7928 9734 7984
rect 9954 7928 10010 7984
rect 9954 7792 10010 7848
rect 9678 7692 9680 7712
rect 9680 7692 9732 7712
rect 9732 7692 9734 7712
rect 9678 7656 9734 7692
rect 7102 4664 7158 4720
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 7286 4140 7342 4176
rect 7286 4120 7288 4140
rect 7288 4120 7340 4140
rect 7340 4120 7342 4140
rect 8482 4684 8538 4720
rect 8482 4664 8484 4684
rect 8484 4664 8536 4684
rect 8536 4664 8538 4684
rect 8666 4564 8668 4584
rect 8668 4564 8720 4584
rect 8720 4564 8722 4584
rect 8666 4528 8722 4564
rect 9494 4664 9550 4720
rect 9862 4528 9918 4584
rect 13358 24112 13414 24168
rect 13082 20440 13138 20496
rect 15290 20440 15346 20496
rect 10414 7948 10470 7984
rect 10414 7928 10416 7948
rect 10416 7928 10468 7948
rect 10468 7928 10470 7948
rect 9954 4120 10010 4176
rect 10874 7812 10930 7848
rect 10874 7792 10876 7812
rect 10876 7792 10928 7812
rect 10928 7792 10930 7812
rect 12806 11348 12862 11384
rect 12806 11328 12808 11348
rect 12808 11328 12860 11348
rect 12860 11328 12862 11348
rect 11518 4664 11574 4720
rect 12162 4564 12164 4584
rect 12164 4564 12216 4584
rect 12216 4564 12218 4584
rect 12162 4528 12218 4564
rect 11978 4020 11980 4040
rect 11980 4020 12032 4040
rect 12032 4020 12034 4040
rect 11978 3984 12034 4020
rect 12346 3712 12402 3768
rect 15290 14340 15346 14376
rect 15290 14320 15292 14340
rect 15292 14320 15344 14340
rect 15344 14320 15346 14340
rect 13726 12416 13782 12472
rect 19706 19372 19762 19408
rect 19706 19352 19708 19372
rect 19708 19352 19760 19372
rect 19760 19352 19762 19372
rect 15474 12416 15530 12472
rect 12990 5888 13046 5944
rect 13358 4548 13414 4584
rect 13358 4528 13360 4548
rect 13360 4528 13412 4548
rect 13412 4528 13414 4548
rect 13358 4004 13414 4040
rect 13358 3984 13360 4004
rect 13360 3984 13412 4004
rect 13412 3984 13414 4004
rect 13726 3732 13782 3768
rect 13726 3712 13728 3732
rect 13728 3712 13780 3732
rect 13780 3712 13782 3732
rect 15474 7792 15530 7848
rect 15750 8372 15752 8392
rect 15752 8372 15804 8392
rect 15804 8372 15806 8392
rect 15750 8336 15806 8372
rect 15750 6060 15752 6080
rect 15752 6060 15804 6080
rect 15804 6060 15806 6080
rect 15750 6024 15806 6060
rect 15382 4936 15438 4992
rect 15842 5228 15898 5264
rect 15842 5208 15844 5228
rect 15844 5208 15896 5228
rect 15896 5208 15898 5228
rect 14462 3168 14518 3224
rect 16118 5480 16174 5536
rect 16026 4800 16082 4856
rect 16210 3984 16266 4040
rect 16118 3848 16174 3904
rect 16946 5752 17002 5808
rect 16578 5228 16634 5264
rect 16578 5208 16580 5228
rect 16580 5208 16632 5228
rect 16632 5208 16634 5228
rect 17038 4936 17094 4992
rect 17222 5908 17278 5944
rect 17222 5888 17224 5908
rect 17224 5888 17276 5908
rect 17276 5888 17278 5908
rect 17222 5752 17278 5808
rect 17498 6024 17554 6080
rect 17498 4936 17554 4992
rect 17406 3984 17462 4040
rect 22282 19372 22338 19408
rect 22282 19352 22284 19372
rect 22284 19352 22336 19372
rect 22336 19352 22338 19372
rect 23754 19372 23810 19408
rect 23754 19352 23756 19372
rect 23756 19352 23808 19372
rect 23808 19352 23810 19372
rect 18234 4664 18290 4720
rect 18510 4820 18566 4856
rect 18510 4800 18512 4820
rect 18512 4800 18564 4820
rect 18564 4800 18566 4820
rect 19062 4664 19118 4720
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 24582 7948 24638 7984
rect 24582 7928 24584 7948
rect 24584 7928 24636 7948
rect 24636 7928 24638 7948
rect 25042 7928 25098 7984
rect 27802 15000 27858 15056
rect 28354 15680 28410 15736
rect 27986 13640 28042 13696
rect 28262 14320 28318 14376
rect 28354 12960 28410 13016
rect 28078 12280 28134 12336
rect 28354 11600 28410 11656
rect 28354 7520 28410 7576
rect 27526 3440 27582 3496
rect 28354 6840 28410 6896
rect 28354 6160 28410 6216
rect 28354 5480 28410 5536
rect 28170 3168 28226 3224
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
<< metal3 >>
rect 4870 29408 5186 29409
rect 4870 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5186 29408
rect 4870 29343 5186 29344
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 4870 28320 5186 28321
rect 4870 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5186 28320
rect 4870 28255 5186 28256
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 0 27298 800 27328
rect 0 27238 1042 27298
rect 0 27208 800 27238
rect 105 27026 171 27029
rect 982 27026 1042 27238
rect 4870 27232 5186 27233
rect 4870 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5186 27232
rect 4870 27167 5186 27168
rect 105 27024 1042 27026
rect 105 26968 110 27024
rect 166 26968 1042 27024
rect 105 26966 1042 26968
rect 105 26963 171 26966
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 4870 26144 5186 26145
rect 4870 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5186 26144
rect 4870 26079 5186 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 4870 25056 5186 25057
rect 4870 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5186 25056
rect 4870 24991 5186 24992
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 11697 24170 11763 24173
rect 12617 24170 12683 24173
rect 13353 24170 13419 24173
rect 11697 24168 13419 24170
rect 11697 24112 11702 24168
rect 11758 24112 12622 24168
rect 12678 24112 13358 24168
rect 13414 24112 13419 24168
rect 11697 24110 13419 24112
rect 11697 24107 11763 24110
rect 12617 24107 12683 24110
rect 13353 24107 13419 24110
rect 4870 23968 5186 23969
rect 4870 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5186 23968
rect 4870 23903 5186 23904
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 4870 22880 5186 22881
rect 4870 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5186 22880
rect 4870 22815 5186 22816
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 5809 21994 5875 21997
rect 12065 21994 12131 21997
rect 5809 21992 12131 21994
rect 5809 21936 5814 21992
rect 5870 21936 12070 21992
rect 12126 21936 12131 21992
rect 5809 21934 12131 21936
rect 5809 21931 5875 21934
rect 12065 21931 12131 21934
rect 4870 21792 5186 21793
rect 4870 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5186 21792
rect 4870 21727 5186 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 4870 20704 5186 20705
rect 4870 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5186 20704
rect 4870 20639 5186 20640
rect 9581 20498 9647 20501
rect 13077 20498 13143 20501
rect 15285 20498 15351 20501
rect 9581 20496 15351 20498
rect 9581 20440 9586 20496
rect 9642 20440 13082 20496
rect 13138 20440 15290 20496
rect 15346 20440 15351 20496
rect 9581 20438 15351 20440
rect 9581 20435 9647 20438
rect 13077 20435 13143 20438
rect 15285 20435 15351 20438
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 4870 19616 5186 19617
rect 4870 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5186 19616
rect 4870 19551 5186 19552
rect 5257 19410 5323 19413
rect 8845 19410 8911 19413
rect 5257 19408 8911 19410
rect 5257 19352 5262 19408
rect 5318 19352 8850 19408
rect 8906 19352 8911 19408
rect 5257 19350 8911 19352
rect 5257 19347 5323 19350
rect 8845 19347 8911 19350
rect 19701 19410 19767 19413
rect 22277 19410 22343 19413
rect 23749 19410 23815 19413
rect 19701 19408 23815 19410
rect 19701 19352 19706 19408
rect 19762 19352 22282 19408
rect 22338 19352 23754 19408
rect 23810 19352 23815 19408
rect 19701 19350 23815 19352
rect 19701 19347 19767 19350
rect 22277 19347 22343 19350
rect 23749 19347 23815 19350
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 4870 18528 5186 18529
rect 4870 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5186 18528
rect 4870 18463 5186 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 4870 17440 5186 17441
rect 4870 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5186 17440
rect 4870 17375 5186 17376
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 4870 16352 5186 16353
rect 4870 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5186 16352
rect 4870 16287 5186 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 28349 15738 28415 15741
rect 29064 15738 29864 15768
rect 28349 15736 29864 15738
rect 28349 15680 28354 15736
rect 28410 15680 29864 15736
rect 28349 15678 29864 15680
rect 28349 15675 28415 15678
rect 29064 15648 29864 15678
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 9121 15058 9187 15061
rect 9581 15058 9647 15061
rect 9121 15056 9647 15058
rect 9121 15000 9126 15056
rect 9182 15000 9586 15056
rect 9642 15000 9647 15056
rect 9121 14998 9647 15000
rect 9121 14995 9187 14998
rect 9581 14995 9647 14998
rect 27797 15058 27863 15061
rect 29064 15058 29864 15088
rect 27797 15056 29864 15058
rect 27797 15000 27802 15056
rect 27858 15000 29864 15056
rect 27797 14998 29864 15000
rect 27797 14995 27863 14998
rect 29064 14968 29864 14998
rect 9213 14922 9279 14925
rect 10041 14922 10107 14925
rect 9213 14920 10107 14922
rect 9213 14864 9218 14920
rect 9274 14864 10046 14920
rect 10102 14864 10107 14920
rect 9213 14862 10107 14864
rect 9213 14859 9279 14862
rect 10041 14859 10107 14862
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 5441 14514 5507 14517
rect 8569 14514 8635 14517
rect 5441 14512 8635 14514
rect 5441 14456 5446 14512
rect 5502 14456 8574 14512
rect 8630 14456 8635 14512
rect 5441 14454 8635 14456
rect 5441 14451 5507 14454
rect 8569 14451 8635 14454
rect 105 14378 171 14381
rect 15285 14378 15351 14381
rect 105 14376 15351 14378
rect 105 14320 110 14376
rect 166 14320 15290 14376
rect 15346 14320 15351 14376
rect 105 14318 15351 14320
rect 105 14315 171 14318
rect 15285 14315 15351 14318
rect 28257 14378 28323 14381
rect 29064 14378 29864 14408
rect 28257 14376 29864 14378
rect 28257 14320 28262 14376
rect 28318 14320 29864 14376
rect 28257 14318 29864 14320
rect 28257 14315 28323 14318
rect 29064 14288 29864 14318
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 27981 13698 28047 13701
rect 29064 13698 29864 13728
rect 27981 13696 29864 13698
rect 27981 13640 27986 13696
rect 28042 13640 29864 13696
rect 27981 13638 29864 13640
rect 27981 13635 28047 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 29064 13608 29864 13638
rect 4210 13567 4526 13568
rect 4870 13088 5186 13089
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 28349 13018 28415 13021
rect 29064 13018 29864 13048
rect 28349 13016 29864 13018
rect 28349 12960 28354 13016
rect 28410 12960 29864 13016
rect 28349 12958 29864 12960
rect 28349 12955 28415 12958
rect 29064 12928 29864 12958
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 13721 12474 13787 12477
rect 15469 12474 15535 12477
rect 13721 12472 15535 12474
rect 13721 12416 13726 12472
rect 13782 12416 15474 12472
rect 15530 12416 15535 12472
rect 13721 12414 15535 12416
rect 13721 12411 13787 12414
rect 15469 12411 15535 12414
rect 28073 12338 28139 12341
rect 29064 12338 29864 12368
rect 28073 12336 29864 12338
rect 28073 12280 28078 12336
rect 28134 12280 29864 12336
rect 28073 12278 29864 12280
rect 28073 12275 28139 12278
rect 29064 12248 29864 12278
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 28349 11658 28415 11661
rect 29064 11658 29864 11688
rect 28349 11656 29864 11658
rect 28349 11600 28354 11656
rect 28410 11600 29864 11656
rect 28349 11598 29864 11600
rect 28349 11595 28415 11598
rect 29064 11568 29864 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 9857 11386 9923 11389
rect 12801 11386 12867 11389
rect 9857 11384 12867 11386
rect 9857 11328 9862 11384
rect 9918 11328 12806 11384
rect 12862 11328 12867 11384
rect 9857 11326 12867 11328
rect 9857 11323 9923 11326
rect 12801 11323 12867 11326
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 4870 10847 5186 10848
rect 4613 10706 4679 10709
rect 8753 10706 8819 10709
rect 4613 10704 8819 10706
rect 4613 10648 4618 10704
rect 4674 10648 8758 10704
rect 8814 10648 8819 10704
rect 4613 10646 8819 10648
rect 4613 10643 4679 10646
rect 8753 10643 8819 10646
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 6545 8530 6611 8533
rect 7281 8530 7347 8533
rect 6545 8528 7347 8530
rect 6545 8472 6550 8528
rect 6606 8472 7286 8528
rect 7342 8472 7347 8528
rect 6545 8470 7347 8472
rect 6545 8467 6611 8470
rect 7281 8467 7347 8470
rect 6821 8394 6887 8397
rect 7189 8394 7255 8397
rect 7649 8394 7715 8397
rect 15745 8396 15811 8397
rect 6821 8392 7715 8394
rect 6821 8336 6826 8392
rect 6882 8336 7194 8392
rect 7250 8336 7654 8392
rect 7710 8336 7715 8392
rect 6821 8334 7715 8336
rect 6821 8331 6887 8334
rect 7189 8331 7255 8334
rect 7649 8331 7715 8334
rect 15694 8332 15700 8396
rect 15764 8394 15811 8396
rect 15764 8392 15856 8394
rect 15806 8336 15856 8392
rect 15764 8334 15856 8336
rect 15764 8332 15811 8334
rect 15745 8331 15811 8332
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 9673 7986 9739 7989
rect 9630 7984 9739 7986
rect 9630 7928 9678 7984
rect 9734 7928 9739 7984
rect 9630 7923 9739 7928
rect 9949 7986 10015 7989
rect 10409 7986 10475 7989
rect 9949 7984 10475 7986
rect 9949 7928 9954 7984
rect 10010 7928 10414 7984
rect 10470 7928 10475 7984
rect 9949 7926 10475 7928
rect 9949 7923 10015 7926
rect 10409 7923 10475 7926
rect 24577 7986 24643 7989
rect 25037 7986 25103 7989
rect 24577 7984 25103 7986
rect 24577 7928 24582 7984
rect 24638 7928 25042 7984
rect 25098 7928 25103 7984
rect 24577 7926 25103 7928
rect 24577 7923 24643 7926
rect 25037 7923 25103 7926
rect 9630 7717 9690 7923
rect 9949 7850 10015 7853
rect 10869 7850 10935 7853
rect 15469 7852 15535 7853
rect 15469 7850 15516 7852
rect 9949 7848 10935 7850
rect 9949 7792 9954 7848
rect 10010 7792 10874 7848
rect 10930 7792 10935 7848
rect 9949 7790 10935 7792
rect 15424 7848 15516 7850
rect 15424 7792 15474 7848
rect 15424 7790 15516 7792
rect 9949 7787 10015 7790
rect 10869 7787 10935 7790
rect 15469 7788 15516 7790
rect 15580 7788 15586 7852
rect 15469 7787 15535 7788
rect 9630 7712 9739 7717
rect 9630 7656 9678 7712
rect 9734 7656 9739 7712
rect 9630 7654 9739 7656
rect 9673 7651 9739 7654
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 28349 7578 28415 7581
rect 29064 7578 29864 7608
rect 28349 7576 29864 7578
rect 28349 7520 28354 7576
rect 28410 7520 29864 7576
rect 28349 7518 29864 7520
rect 28349 7515 28415 7518
rect 29064 7488 29864 7518
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 28349 6898 28415 6901
rect 29064 6898 29864 6928
rect 28349 6896 29864 6898
rect 28349 6840 28354 6896
rect 28410 6840 29864 6896
rect 28349 6838 29864 6840
rect 28349 6835 28415 6838
rect 29064 6808 29864 6838
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 28349 6218 28415 6221
rect 29064 6218 29864 6248
rect 28349 6216 29864 6218
rect 28349 6160 28354 6216
rect 28410 6160 29864 6216
rect 28349 6158 29864 6160
rect 28349 6155 28415 6158
rect 29064 6128 29864 6158
rect 15745 6082 15811 6085
rect 17493 6082 17559 6085
rect 15745 6080 17559 6082
rect 15745 6024 15750 6080
rect 15806 6024 17498 6080
rect 17554 6024 17559 6080
rect 15745 6022 17559 6024
rect 15745 6019 15811 6022
rect 17493 6019 17559 6022
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 12985 5946 13051 5949
rect 17217 5946 17283 5949
rect 12985 5944 17283 5946
rect 12985 5888 12990 5944
rect 13046 5888 17222 5944
rect 17278 5888 17283 5944
rect 12985 5886 17283 5888
rect 12985 5883 13051 5886
rect 17217 5883 17283 5886
rect 16941 5810 17007 5813
rect 17217 5810 17283 5813
rect 16941 5808 17283 5810
rect 16941 5752 16946 5808
rect 17002 5752 17222 5808
rect 17278 5752 17283 5808
rect 16941 5750 17283 5752
rect 16941 5747 17007 5750
rect 17217 5747 17283 5750
rect 6913 5538 6979 5541
rect 15694 5538 15700 5540
rect 6913 5536 15700 5538
rect 6913 5480 6918 5536
rect 6974 5480 15700 5536
rect 6913 5478 15700 5480
rect 6913 5475 6979 5478
rect 15694 5476 15700 5478
rect 15764 5538 15770 5540
rect 16113 5538 16179 5541
rect 15764 5536 16179 5538
rect 15764 5480 16118 5536
rect 16174 5480 16179 5536
rect 15764 5478 16179 5480
rect 15764 5476 15770 5478
rect 16113 5475 16179 5478
rect 28349 5538 28415 5541
rect 29064 5538 29864 5568
rect 28349 5536 29864 5538
rect 28349 5480 28354 5536
rect 28410 5480 29864 5536
rect 28349 5478 29864 5480
rect 28349 5475 28415 5478
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 29064 5448 29864 5478
rect 4870 5407 5186 5408
rect 15837 5266 15903 5269
rect 16573 5266 16639 5269
rect 15837 5264 16639 5266
rect 15837 5208 15842 5264
rect 15898 5208 16578 5264
rect 16634 5208 16639 5264
rect 15837 5206 16639 5208
rect 15837 5203 15903 5206
rect 16573 5203 16639 5206
rect 15377 4994 15443 4997
rect 17033 4994 17099 4997
rect 17493 4994 17559 4997
rect 15377 4992 17559 4994
rect 15377 4936 15382 4992
rect 15438 4936 17038 4992
rect 17094 4936 17498 4992
rect 17554 4936 17559 4992
rect 15377 4934 17559 4936
rect 15377 4931 15443 4934
rect 17033 4931 17099 4934
rect 17493 4931 17559 4934
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 16021 4858 16087 4861
rect 18505 4858 18571 4861
rect 16021 4856 18571 4858
rect 16021 4800 16026 4856
rect 16082 4800 18510 4856
rect 18566 4800 18571 4856
rect 16021 4798 18571 4800
rect 16021 4795 16087 4798
rect 18505 4795 18571 4798
rect 6085 4722 6151 4725
rect 7097 4722 7163 4725
rect 6085 4720 7163 4722
rect 6085 4664 6090 4720
rect 6146 4664 7102 4720
rect 7158 4664 7163 4720
rect 6085 4662 7163 4664
rect 6085 4659 6151 4662
rect 7097 4659 7163 4662
rect 8477 4722 8543 4725
rect 9489 4722 9555 4725
rect 11513 4722 11579 4725
rect 18229 4722 18295 4725
rect 19057 4722 19123 4725
rect 8477 4720 19123 4722
rect 8477 4664 8482 4720
rect 8538 4664 9494 4720
rect 9550 4664 11518 4720
rect 11574 4664 18234 4720
rect 18290 4664 19062 4720
rect 19118 4664 19123 4720
rect 8477 4662 19123 4664
rect 8477 4659 8543 4662
rect 9489 4659 9555 4662
rect 11513 4659 11579 4662
rect 18229 4659 18295 4662
rect 19057 4659 19123 4662
rect 8661 4586 8727 4589
rect 9857 4586 9923 4589
rect 8661 4584 9923 4586
rect 8661 4528 8666 4584
rect 8722 4528 9862 4584
rect 9918 4528 9923 4584
rect 8661 4526 9923 4528
rect 8661 4523 8727 4526
rect 9857 4523 9923 4526
rect 12157 4586 12223 4589
rect 13353 4586 13419 4589
rect 12157 4584 13419 4586
rect 12157 4528 12162 4584
rect 12218 4528 13358 4584
rect 13414 4528 13419 4584
rect 12157 4526 13419 4528
rect 12157 4523 12223 4526
rect 13353 4523 13419 4526
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 7281 4178 7347 4181
rect 9949 4178 10015 4181
rect 7281 4176 10015 4178
rect 7281 4120 7286 4176
rect 7342 4120 9954 4176
rect 10010 4120 10015 4176
rect 7281 4118 10015 4120
rect 7281 4115 7347 4118
rect 9949 4115 10015 4118
rect 11973 4042 12039 4045
rect 13353 4042 13419 4045
rect 11973 4040 13419 4042
rect 11973 3984 11978 4040
rect 12034 3984 13358 4040
rect 13414 3984 13419 4040
rect 11973 3982 13419 3984
rect 11973 3979 12039 3982
rect 13353 3979 13419 3982
rect 16205 4042 16271 4045
rect 17401 4042 17467 4045
rect 16205 4040 17467 4042
rect 16205 3984 16210 4040
rect 16266 3984 17406 4040
rect 17462 3984 17467 4040
rect 16205 3982 17467 3984
rect 16205 3979 16271 3982
rect 17401 3979 17467 3982
rect 15510 3844 15516 3908
rect 15580 3906 15586 3908
rect 16113 3906 16179 3909
rect 15580 3904 16179 3906
rect 15580 3848 16118 3904
rect 16174 3848 16179 3904
rect 15580 3846 16179 3848
rect 15580 3844 15586 3846
rect 16113 3843 16179 3846
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 12341 3770 12407 3773
rect 13721 3770 13787 3773
rect 12341 3768 13787 3770
rect 12341 3712 12346 3768
rect 12402 3712 13726 3768
rect 13782 3712 13787 3768
rect 12341 3710 13787 3712
rect 12341 3707 12407 3710
rect 13721 3707 13787 3710
rect 27521 3498 27587 3501
rect 29064 3498 29864 3528
rect 27521 3496 29864 3498
rect 27521 3440 27526 3496
rect 27582 3440 29864 3496
rect 27521 3438 29864 3440
rect 27521 3435 27587 3438
rect 29064 3408 29864 3438
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 14457 3226 14523 3229
rect 28165 3226 28231 3229
rect 14457 3224 28231 3226
rect 14457 3168 14462 3224
rect 14518 3168 28170 3224
rect 28226 3168 28231 3224
rect 14457 3166 28231 3168
rect 14457 3163 14523 3166
rect 28165 3163 28231 3166
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
<< via3 >>
rect 4876 29404 4940 29408
rect 4876 29348 4880 29404
rect 4880 29348 4936 29404
rect 4936 29348 4940 29404
rect 4876 29344 4940 29348
rect 4956 29404 5020 29408
rect 4956 29348 4960 29404
rect 4960 29348 5016 29404
rect 5016 29348 5020 29404
rect 4956 29344 5020 29348
rect 5036 29404 5100 29408
rect 5036 29348 5040 29404
rect 5040 29348 5096 29404
rect 5096 29348 5100 29404
rect 5036 29344 5100 29348
rect 5116 29404 5180 29408
rect 5116 29348 5120 29404
rect 5120 29348 5176 29404
rect 5176 29348 5180 29404
rect 5116 29344 5180 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 4876 28316 4940 28320
rect 4876 28260 4880 28316
rect 4880 28260 4936 28316
rect 4936 28260 4940 28316
rect 4876 28256 4940 28260
rect 4956 28316 5020 28320
rect 4956 28260 4960 28316
rect 4960 28260 5016 28316
rect 5016 28260 5020 28316
rect 4956 28256 5020 28260
rect 5036 28316 5100 28320
rect 5036 28260 5040 28316
rect 5040 28260 5096 28316
rect 5096 28260 5100 28316
rect 5036 28256 5100 28260
rect 5116 28316 5180 28320
rect 5116 28260 5120 28316
rect 5120 28260 5176 28316
rect 5176 28260 5180 28316
rect 5116 28256 5180 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 4876 27228 4940 27232
rect 4876 27172 4880 27228
rect 4880 27172 4936 27228
rect 4936 27172 4940 27228
rect 4876 27168 4940 27172
rect 4956 27228 5020 27232
rect 4956 27172 4960 27228
rect 4960 27172 5016 27228
rect 5016 27172 5020 27228
rect 4956 27168 5020 27172
rect 5036 27228 5100 27232
rect 5036 27172 5040 27228
rect 5040 27172 5096 27228
rect 5096 27172 5100 27228
rect 5036 27168 5100 27172
rect 5116 27228 5180 27232
rect 5116 27172 5120 27228
rect 5120 27172 5176 27228
rect 5176 27172 5180 27228
rect 5116 27168 5180 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 4876 26140 4940 26144
rect 4876 26084 4880 26140
rect 4880 26084 4936 26140
rect 4936 26084 4940 26140
rect 4876 26080 4940 26084
rect 4956 26140 5020 26144
rect 4956 26084 4960 26140
rect 4960 26084 5016 26140
rect 5016 26084 5020 26140
rect 4956 26080 5020 26084
rect 5036 26140 5100 26144
rect 5036 26084 5040 26140
rect 5040 26084 5096 26140
rect 5096 26084 5100 26140
rect 5036 26080 5100 26084
rect 5116 26140 5180 26144
rect 5116 26084 5120 26140
rect 5120 26084 5176 26140
rect 5176 26084 5180 26140
rect 5116 26080 5180 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 4876 25052 4940 25056
rect 4876 24996 4880 25052
rect 4880 24996 4936 25052
rect 4936 24996 4940 25052
rect 4876 24992 4940 24996
rect 4956 25052 5020 25056
rect 4956 24996 4960 25052
rect 4960 24996 5016 25052
rect 5016 24996 5020 25052
rect 4956 24992 5020 24996
rect 5036 25052 5100 25056
rect 5036 24996 5040 25052
rect 5040 24996 5096 25052
rect 5096 24996 5100 25052
rect 5036 24992 5100 24996
rect 5116 25052 5180 25056
rect 5116 24996 5120 25052
rect 5120 24996 5176 25052
rect 5176 24996 5180 25052
rect 5116 24992 5180 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 4876 23964 4940 23968
rect 4876 23908 4880 23964
rect 4880 23908 4936 23964
rect 4936 23908 4940 23964
rect 4876 23904 4940 23908
rect 4956 23964 5020 23968
rect 4956 23908 4960 23964
rect 4960 23908 5016 23964
rect 5016 23908 5020 23964
rect 4956 23904 5020 23908
rect 5036 23964 5100 23968
rect 5036 23908 5040 23964
rect 5040 23908 5096 23964
rect 5096 23908 5100 23964
rect 5036 23904 5100 23908
rect 5116 23964 5180 23968
rect 5116 23908 5120 23964
rect 5120 23908 5176 23964
rect 5176 23908 5180 23964
rect 5116 23904 5180 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 4876 22876 4940 22880
rect 4876 22820 4880 22876
rect 4880 22820 4936 22876
rect 4936 22820 4940 22876
rect 4876 22816 4940 22820
rect 4956 22876 5020 22880
rect 4956 22820 4960 22876
rect 4960 22820 5016 22876
rect 5016 22820 5020 22876
rect 4956 22816 5020 22820
rect 5036 22876 5100 22880
rect 5036 22820 5040 22876
rect 5040 22820 5096 22876
rect 5096 22820 5100 22876
rect 5036 22816 5100 22820
rect 5116 22876 5180 22880
rect 5116 22820 5120 22876
rect 5120 22820 5176 22876
rect 5176 22820 5180 22876
rect 5116 22816 5180 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 4876 21788 4940 21792
rect 4876 21732 4880 21788
rect 4880 21732 4936 21788
rect 4936 21732 4940 21788
rect 4876 21728 4940 21732
rect 4956 21788 5020 21792
rect 4956 21732 4960 21788
rect 4960 21732 5016 21788
rect 5016 21732 5020 21788
rect 4956 21728 5020 21732
rect 5036 21788 5100 21792
rect 5036 21732 5040 21788
rect 5040 21732 5096 21788
rect 5096 21732 5100 21788
rect 5036 21728 5100 21732
rect 5116 21788 5180 21792
rect 5116 21732 5120 21788
rect 5120 21732 5176 21788
rect 5176 21732 5180 21788
rect 5116 21728 5180 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 4876 20700 4940 20704
rect 4876 20644 4880 20700
rect 4880 20644 4936 20700
rect 4936 20644 4940 20700
rect 4876 20640 4940 20644
rect 4956 20700 5020 20704
rect 4956 20644 4960 20700
rect 4960 20644 5016 20700
rect 5016 20644 5020 20700
rect 4956 20640 5020 20644
rect 5036 20700 5100 20704
rect 5036 20644 5040 20700
rect 5040 20644 5096 20700
rect 5096 20644 5100 20700
rect 5036 20640 5100 20644
rect 5116 20700 5180 20704
rect 5116 20644 5120 20700
rect 5120 20644 5176 20700
rect 5176 20644 5180 20700
rect 5116 20640 5180 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 4876 19612 4940 19616
rect 4876 19556 4880 19612
rect 4880 19556 4936 19612
rect 4936 19556 4940 19612
rect 4876 19552 4940 19556
rect 4956 19612 5020 19616
rect 4956 19556 4960 19612
rect 4960 19556 5016 19612
rect 5016 19556 5020 19612
rect 4956 19552 5020 19556
rect 5036 19612 5100 19616
rect 5036 19556 5040 19612
rect 5040 19556 5096 19612
rect 5096 19556 5100 19612
rect 5036 19552 5100 19556
rect 5116 19612 5180 19616
rect 5116 19556 5120 19612
rect 5120 19556 5176 19612
rect 5176 19556 5180 19612
rect 5116 19552 5180 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 4876 18524 4940 18528
rect 4876 18468 4880 18524
rect 4880 18468 4936 18524
rect 4936 18468 4940 18524
rect 4876 18464 4940 18468
rect 4956 18524 5020 18528
rect 4956 18468 4960 18524
rect 4960 18468 5016 18524
rect 5016 18468 5020 18524
rect 4956 18464 5020 18468
rect 5036 18524 5100 18528
rect 5036 18468 5040 18524
rect 5040 18468 5096 18524
rect 5096 18468 5100 18524
rect 5036 18464 5100 18468
rect 5116 18524 5180 18528
rect 5116 18468 5120 18524
rect 5120 18468 5176 18524
rect 5176 18468 5180 18524
rect 5116 18464 5180 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 4876 17436 4940 17440
rect 4876 17380 4880 17436
rect 4880 17380 4936 17436
rect 4936 17380 4940 17436
rect 4876 17376 4940 17380
rect 4956 17436 5020 17440
rect 4956 17380 4960 17436
rect 4960 17380 5016 17436
rect 5016 17380 5020 17436
rect 4956 17376 5020 17380
rect 5036 17436 5100 17440
rect 5036 17380 5040 17436
rect 5040 17380 5096 17436
rect 5096 17380 5100 17436
rect 5036 17376 5100 17380
rect 5116 17436 5180 17440
rect 5116 17380 5120 17436
rect 5120 17380 5176 17436
rect 5176 17380 5180 17436
rect 5116 17376 5180 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 4876 16348 4940 16352
rect 4876 16292 4880 16348
rect 4880 16292 4936 16348
rect 4936 16292 4940 16348
rect 4876 16288 4940 16292
rect 4956 16348 5020 16352
rect 4956 16292 4960 16348
rect 4960 16292 5016 16348
rect 5016 16292 5020 16348
rect 4956 16288 5020 16292
rect 5036 16348 5100 16352
rect 5036 16292 5040 16348
rect 5040 16292 5096 16348
rect 5096 16292 5100 16348
rect 5036 16288 5100 16292
rect 5116 16348 5180 16352
rect 5116 16292 5120 16348
rect 5120 16292 5176 16348
rect 5176 16292 5180 16348
rect 5116 16288 5180 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 15700 8392 15764 8396
rect 15700 8336 15750 8392
rect 15750 8336 15764 8392
rect 15700 8332 15764 8336
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 15516 7848 15580 7852
rect 15516 7792 15530 7848
rect 15530 7792 15580 7848
rect 15516 7788 15580 7792
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 15700 5476 15764 5540
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 15516 3844 15580 3908
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
<< metal4 >>
rect 4208 28864 4528 29424
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 29408 5188 29424
rect 4868 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5188 29408
rect 4868 28320 5188 29344
rect 4868 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5188 28320
rect 4868 27232 5188 28256
rect 4868 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5188 27232
rect 4868 26144 5188 27168
rect 4868 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5188 26144
rect 4868 25056 5188 26080
rect 4868 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5188 25056
rect 4868 23968 5188 24992
rect 4868 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5188 23968
rect 4868 22880 5188 23904
rect 4868 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5188 22880
rect 4868 21792 5188 22816
rect 4868 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5188 21792
rect 4868 20704 5188 21728
rect 4868 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5188 20704
rect 4868 19616 5188 20640
rect 4868 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5188 19616
rect 4868 18528 5188 19552
rect 4868 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5188 18528
rect 4868 17440 5188 18464
rect 4868 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5188 17440
rect 4868 16352 5188 17376
rect 4868 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5188 16352
rect 4868 15264 5188 16288
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4868 13088 5188 14112
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4868 10912 5188 11936
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 15699 8396 15765 8397
rect 15699 8332 15700 8396
rect 15764 8332 15765 8396
rect 15699 8331 15765 8332
rect 15515 7852 15581 7853
rect 15515 7788 15516 7852
rect 15580 7788 15581 7852
rect 15515 7787 15581 7788
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 15518 3909 15578 7787
rect 15702 5541 15762 8331
rect 15699 5540 15765 5541
rect 15699 5476 15700 5540
rect 15764 5476 15765 5540
rect 15699 5475 15765 5476
rect 15515 3908 15581 3909
rect 15515 3844 15516 3908
rect 15580 3844 15581 3908
rect 15515 3843 15581 3844
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
use sky130_fd_sc_hd__inv_2  _0429_
timestamp 1
transform -1 0 18492 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0430_
timestamp 1
transform 1 0 16284 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0431_
timestamp 1
transform 1 0 14076 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0432_
timestamp 1
transform 1 0 8280 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0433_
timestamp 1
transform -1 0 8832 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0434_
timestamp 1
transform -1 0 27876 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0435_
timestamp 1
transform 1 0 26220 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0436_
timestamp 1
transform -1 0 25760 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0437_
timestamp 1
transform -1 0 25116 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0438_
timestamp 1
transform -1 0 22356 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0439_
timestamp 1
transform -1 0 22356 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0440_
timestamp 1
transform -1 0 22080 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0441_
timestamp 1
transform -1 0 22724 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0442_
timestamp 1
transform -1 0 26496 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0443_
timestamp 1
transform 1 0 25024 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0444_
timestamp 1
transform -1 0 24288 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0445_
timestamp 1
transform -1 0 26036 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0446_
timestamp 1
transform -1 0 25668 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0447_
timestamp 1
transform -1 0 25944 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _0448_
timestamp 1
transform -1 0 16744 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _0449_
timestamp 1
transform 1 0 14904 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0450_
timestamp 1
transform 1 0 10212 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0451_
timestamp 1
transform 1 0 11684 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0452_
timestamp 1
transform -1 0 13248 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0453_
timestamp 1
transform 1 0 16928 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0454_
timestamp 1
transform -1 0 18952 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o21bai_1  _0455_
timestamp 1
transform -1 0 19504 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0456_
timestamp 1
transform 1 0 15272 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0457_
timestamp 1
transform -1 0 16928 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0458_
timestamp 1
transform 1 0 14720 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0459_
timestamp 1
transform -1 0 17940 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_4  _0460_
timestamp 1
transform 1 0 19044 0 -1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_2  _0461_
timestamp 1
transform 1 0 7084 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _0462_
timestamp 1
transform -1 0 12604 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0463_
timestamp 1
transform -1 0 11408 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0464_
timestamp 1
transform 1 0 12328 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0465_
timestamp 1
transform -1 0 16100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0466_
timestamp 1
transform -1 0 11224 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0467_
timestamp 1
transform -1 0 10304 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0468_
timestamp 1
transform 1 0 18584 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _0469_
timestamp 1
transform -1 0 17112 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o21bai_4  _0470_
timestamp 1
transform 1 0 15272 0 1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__a22o_1  _0471_
timestamp 1
transform 1 0 9660 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0472_
timestamp 1
transform -1 0 10028 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0473_
timestamp 1
transform 1 0 9568 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _0474_
timestamp 1
transform 1 0 8280 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0475_
timestamp 1
transform -1 0 9476 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0476_
timestamp 1
transform -1 0 7820 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0477_
timestamp 1
transform -1 0 9568 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0478_
timestamp 1
transform -1 0 8464 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _0479_
timestamp 1
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _0480_
timestamp 1
transform -1 0 19964 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _0481_
timestamp 1
transform -1 0 20700 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0482_
timestamp 1
transform 1 0 19228 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_2  _0483_
timestamp 1
transform -1 0 19872 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0484_
timestamp 1
transform 1 0 11224 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_1  _0485_
timestamp 1
transform -1 0 20700 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0486_
timestamp 1
transform 1 0 18400 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0487_
timestamp 1
transform -1 0 14628 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0488_
timestamp 1
transform -1 0 13984 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0489_
timestamp 1
transform -1 0 12420 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0490_
timestamp 1
transform 1 0 17848 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_2  _0491_
timestamp 1
transform -1 0 17940 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0492_
timestamp 1
transform -1 0 13156 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0493_
timestamp 1
transform 1 0 16652 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_2  _0494_
timestamp 1
transform 1 0 16652 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0495_
timestamp 1
transform 1 0 10948 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0496_
timestamp 1
transform 1 0 18400 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0497_
timestamp 1
transform 1 0 19044 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0498_
timestamp 1
transform -1 0 18400 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0499_
timestamp 1
transform -1 0 11500 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0500_
timestamp 1
transform -1 0 11224 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0501_
timestamp 1
transform 1 0 10120 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _0502_
timestamp 1
transform -1 0 13340 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0503_
timestamp 1
transform 1 0 11868 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0504_
timestamp 1
transform 1 0 12972 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a311o_1  _0505_
timestamp 1
transform 1 0 12236 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o32a_2  _0506_
timestamp 1
transform -1 0 17480 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0507_
timestamp 1
transform -1 0 10948 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0508_
timestamp 1
transform -1 0 8648 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0509_
timestamp 1
transform -1 0 10028 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0510_
timestamp 1
transform 1 0 8648 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_2  _0511_
timestamp 1
transform 1 0 15640 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0512_
timestamp 1
transform -1 0 6256 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0513_
timestamp 1
transform 1 0 6256 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0514_
timestamp 1
transform 1 0 6716 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0515_
timestamp 1
transform 1 0 17112 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0516_
timestamp 1
transform 1 0 14996 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_2  _0517_
timestamp 1
transform -1 0 16376 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0518_
timestamp 1
transform 1 0 5796 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0519_
timestamp 1
transform 1 0 6348 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _0520_
timestamp 1
transform 1 0 8004 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0521_
timestamp 1
transform 1 0 8188 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0522_
timestamp 1
transform -1 0 7452 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0523_
timestamp 1
transform -1 0 6716 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0524_
timestamp 1
transform 1 0 7452 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_1  _0525_
timestamp 1
transform -1 0 16836 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0526_
timestamp 1
transform -1 0 16468 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0527_
timestamp 1
transform -1 0 8096 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0528_
timestamp 1
transform -1 0 7820 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0529_
timestamp 1
transform -1 0 6808 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _0530_
timestamp 1
transform 1 0 16376 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0531_
timestamp 1
transform 1 0 5888 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0532_
timestamp 1
transform -1 0 6164 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0533_
timestamp 1
transform -1 0 5520 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0534_
timestamp 1
transform 1 0 6348 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _0535_
timestamp 1
transform 1 0 17664 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0536_
timestamp 1
transform 1 0 16008 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0537_
timestamp 1
transform -1 0 17296 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0538_
timestamp 1
transform -1 0 6716 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0539_
timestamp 1
transform 1 0 7176 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0540_
timestamp 1
transform 1 0 6164 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0541_
timestamp 1
transform -1 0 15640 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_2  _0542_
timestamp 1
transform -1 0 16284 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0543_
timestamp 1
transform 1 0 6348 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0544_
timestamp 1
transform -1 0 7360 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0545_
timestamp 1
transform -1 0 7636 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0546_
timestamp 1
transform 1 0 7084 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0547_
timestamp 1
transform -1 0 7176 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0548_
timestamp 1
transform -1 0 6716 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0549_
timestamp 1
transform 1 0 6440 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _0550_
timestamp 1
transform -1 0 7452 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_2  _0551_
timestamp 1
transform -1 0 8096 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0552_
timestamp 1
transform 1 0 6532 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0553_
timestamp 1
transform 1 0 5520 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _0554_
timestamp 1
transform -1 0 7176 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _0555_
timestamp 1
transform 1 0 6992 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0556_
timestamp 1
transform 1 0 12696 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0557_
timestamp 1
transform 1 0 12144 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0558_
timestamp 1
transform 1 0 16008 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_4  _0559_
timestamp 1
transform -1 0 16468 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _0560_
timestamp 1
transform 1 0 13524 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _0561_
timestamp 1
transform 1 0 20792 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0562_
timestamp 1
transform 1 0 20976 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _0563_
timestamp 1
transform 1 0 21620 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0564_
timestamp 1
transform 1 0 23920 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _0565_
timestamp 1
transform 1 0 24656 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0566_
timestamp 1
transform 1 0 26956 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _0567_
timestamp 1
transform 1 0 26220 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0568_
timestamp 1
transform -1 0 28428 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0569_
timestamp 1
transform -1 0 27508 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0570_
timestamp 1
transform 1 0 26036 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0571_
timestamp 1
transform -1 0 27324 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0572_
timestamp 1
transform 1 0 27324 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0573_
timestamp 1
transform 1 0 25024 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0574_
timestamp 1
transform 1 0 26128 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0575_
timestamp 1
transform 1 0 25668 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0576_
timestamp 1
transform -1 0 25576 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0577_
timestamp 1
transform 1 0 26956 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _0578_
timestamp 1
transform -1 0 26496 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0579_
timestamp 1
transform 1 0 24748 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0580_
timestamp 1
transform -1 0 18308 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0581_
timestamp 1
transform 1 0 17848 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0582_
timestamp 1
transform -1 0 18860 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0583_
timestamp 1
transform -1 0 19504 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0584_
timestamp 1
transform 1 0 18400 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0585_
timestamp 1
transform -1 0 18952 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0586_
timestamp 1
transform 1 0 17572 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0587_
timestamp 1
transform -1 0 17940 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0588_
timestamp 1
transform -1 0 17388 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0589_
timestamp 1
transform -1 0 17296 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0590_
timestamp 1
transform 1 0 14260 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0591_
timestamp 1
transform 1 0 15364 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0592_
timestamp 1
transform 1 0 15916 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0593_
timestamp 1
transform -1 0 15456 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0594_
timestamp 1
transform -1 0 15364 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0595_
timestamp 1
transform 1 0 14720 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0596_
timestamp 1
transform 1 0 14628 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0597_
timestamp 1
transform -1 0 14720 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0598_
timestamp 1
transform -1 0 12972 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0599_
timestamp 1
transform -1 0 12604 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0600_
timestamp 1
transform 1 0 12604 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0601_
timestamp 1
transform -1 0 13708 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _0602_
timestamp 1
transform -1 0 13800 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a221oi_1  _0603_
timestamp 1
transform 1 0 12236 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0604_
timestamp 1
transform 1 0 12420 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0605_
timestamp 1
transform 1 0 18124 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0606_
timestamp 1
transform -1 0 19320 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0607_
timestamp 1
transform -1 0 19044 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0608_
timestamp 1
transform -1 0 19872 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0609_
timestamp 1
transform 1 0 20148 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0610_
timestamp 1
transform -1 0 20148 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0611_
timestamp 1
transform 1 0 19780 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0612_
timestamp 1
transform 1 0 20516 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0613_
timestamp 1
transform 1 0 20240 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0614_
timestamp 1
transform -1 0 20976 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0615_
timestamp 1
transform 1 0 20976 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0616_
timestamp 1
transform 1 0 19044 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0617_
timestamp 1
transform 1 0 20148 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0618_
timestamp 1
transform 1 0 19504 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0619_
timestamp 1
transform -1 0 17112 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0620_
timestamp 1
transform 1 0 17940 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0621_
timestamp 1
transform 1 0 18584 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0622_
timestamp 1
transform -1 0 18584 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0623_
timestamp 1
transform -1 0 17940 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0624_
timestamp 1
transform -1 0 16560 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0625_
timestamp 1
transform 1 0 15640 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0626_
timestamp 1
transform -1 0 16100 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0627_
timestamp 1
transform -1 0 14536 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0628_
timestamp 1
transform 1 0 14168 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0629_
timestamp 1
transform 1 0 14536 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0630_
timestamp 1
transform -1 0 13432 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0631_
timestamp 1
transform 1 0 12696 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0632_
timestamp 1
transform -1 0 13800 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0633_
timestamp 1
transform 1 0 14168 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0634_
timestamp 1
transform 1 0 13340 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0635_
timestamp 1
transform -1 0 13340 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0636_
timestamp 1
transform -1 0 13708 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0637_
timestamp 1
transform -1 0 11592 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0638_
timestamp 1
transform 1 0 12144 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0639_
timestamp 1
transform 1 0 12420 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0640_
timestamp 1
transform -1 0 13892 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0641_
timestamp 1
transform 1 0 11592 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0642_
timestamp 1
transform -1 0 13340 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0643_
timestamp 1
transform 1 0 11500 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0644_
timestamp 1
transform -1 0 10212 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0645_
timestamp 1
transform -1 0 8832 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0646_
timestamp 1
transform -1 0 8464 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0647_
timestamp 1
transform -1 0 9844 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _0648_
timestamp 1
transform -1 0 9292 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0649_
timestamp 1
transform 1 0 12144 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0650_
timestamp 1
transform -1 0 10304 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0651_
timestamp 1
transform 1 0 13616 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0652_
timestamp 1
transform 1 0 12512 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0653_
timestamp 1
transform 1 0 10764 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0654_
timestamp 1
transform 1 0 10948 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0655_
timestamp 1
transform 1 0 22540 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0656_
timestamp 1
transform 1 0 23092 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0657_
timestamp 1
transform 1 0 25852 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0658_
timestamp 1
transform 1 0 26404 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0659_
timestamp 1
transform 1 0 25484 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0660_
timestamp 1
transform -1 0 20332 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0661_
timestamp 1
transform -1 0 21804 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0662_
timestamp 1
transform 1 0 21252 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0663_
timestamp 1
transform 1 0 22080 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0664_
timestamp 1
transform 1 0 23000 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0665_
timestamp 1
transform 1 0 23644 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0666_
timestamp 1
transform 1 0 26312 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0667_
timestamp 1
transform 1 0 26956 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0668_
timestamp 1
transform -1 0 26496 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0669_
timestamp 1
transform 1 0 26956 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0670_
timestamp 1
transform -1 0 28428 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0671_
timestamp 1
transform -1 0 26680 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _0672_
timestamp 1
transform -1 0 25392 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0673_
timestamp 1
transform -1 0 24932 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0674_
timestamp 1
transform -1 0 25300 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0675_
timestamp 1
transform -1 0 25668 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0676_
timestamp 1
transform 1 0 24656 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0677_
timestamp 1
transform 1 0 25300 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0678_
timestamp 1
transform 1 0 27140 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and3_2  _0679_
timestamp 1
transform -1 0 24932 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0680_
timestamp 1
transform 1 0 17480 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0681_
timestamp 1
transform 1 0 17112 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0682_
timestamp 1
transform -1 0 18492 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _0683_
timestamp 1
transform 1 0 16836 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0684_
timestamp 1
transform 1 0 18216 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _0685_
timestamp 1
transform 1 0 17756 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0686_
timestamp 1
transform 1 0 19228 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _0687_
timestamp 1
transform 1 0 20240 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0688_
timestamp 1
transform 1 0 21804 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _0689_
timestamp 1
transform 1 0 21804 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0690_
timestamp 1
transform 1 0 23276 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _0691_
timestamp 1
transform 1 0 23460 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0692_
timestamp 1
transform 1 0 23552 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_1  _0693_
timestamp 1
transform 1 0 23920 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0694_
timestamp 1
transform -1 0 24932 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0695_
timestamp 1
transform -1 0 25852 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0696_
timestamp 1
transform -1 0 27692 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0697_
timestamp 1
transform 1 0 23092 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0698_
timestamp 1
transform -1 0 27508 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0699_
timestamp 1
transform 1 0 26956 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _0700_
timestamp 1
transform -1 0 27784 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0701_
timestamp 1
transform -1 0 11684 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0702_
timestamp 1
transform -1 0 11500 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _0703_
timestamp 1
transform 1 0 12604 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_1  _0704_
timestamp 1
transform -1 0 13892 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0705_
timestamp 1
transform -1 0 11500 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0706_
timestamp 1
transform -1 0 11040 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0707_
timestamp 1
transform 1 0 15456 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0708_
timestamp 1
transform 1 0 15732 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0709_
timestamp 1
transform 1 0 17112 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0710_
timestamp 1
transform 1 0 17388 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0711_
timestamp 1
transform 1 0 18676 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0712_
timestamp 1
transform -1 0 19504 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0713_
timestamp 1
transform 1 0 20332 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0714_
timestamp 1
transform 1 0 20792 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0715_
timestamp 1
transform -1 0 23736 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0716_
timestamp 1
transform 1 0 21896 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0717_
timestamp 1
transform 1 0 22172 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0718_
timestamp 1
transform 1 0 22172 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0719_
timestamp 1
transform -1 0 23184 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0720_
timestamp 1
transform 1 0 22172 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _0721_
timestamp 1
transform 1 0 18216 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0722_
timestamp 1
transform 1 0 19964 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0723_
timestamp 1
transform 1 0 20884 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0724_
timestamp 1
transform -1 0 22540 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0725_
timestamp 1
transform 1 0 21804 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0726_
timestamp 1
transform 1 0 21712 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0727_
timestamp 1
transform 1 0 23092 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0728_
timestamp 1
transform 1 0 22356 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0729_
timestamp 1
transform -1 0 24380 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0730_
timestamp 1
transform 1 0 21712 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0731_
timestamp 1
transform -1 0 22632 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0732_
timestamp 1
transform 1 0 20516 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0733_
timestamp 1
transform -1 0 20976 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0734_
timestamp 1
transform 1 0 18400 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0735_
timestamp 1
transform -1 0 19136 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0736_
timestamp 1
transform 1 0 17112 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0737_
timestamp 1
transform -1 0 17940 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0738_
timestamp 1
transform 1 0 15640 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0739_
timestamp 1
transform 1 0 15640 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0740_
timestamp 1
transform 1 0 15272 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0741_
timestamp 1
transform 1 0 15916 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0742_
timestamp 1
transform 1 0 15180 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0743_
timestamp 1
transform 1 0 15088 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0744_
timestamp 1
transform 1 0 13432 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0745_
timestamp 1
transform -1 0 13708 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0746_
timestamp 1
transform -1 0 13156 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0747_
timestamp 1
transform -1 0 12328 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0748_
timestamp 1
transform -1 0 11868 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0749_
timestamp 1
transform 1 0 10028 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0750_
timestamp 1
transform -1 0 12236 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0751_
timestamp 1
transform 1 0 9936 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0752_
timestamp 1
transform 1 0 14076 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0753_
timestamp 1
transform 1 0 19228 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0754_
timestamp 1
transform -1 0 20240 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0755_
timestamp 1
transform 1 0 20056 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0756_
timestamp 1
transform 1 0 21804 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0757_
timestamp 1
transform 1 0 23276 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0758_
timestamp 1
transform -1 0 25760 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0759_
timestamp 1
transform 1 0 26956 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0760_
timestamp 1
transform -1 0 27876 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _0761_
timestamp 1
transform 1 0 14076 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0762_
timestamp 1
transform -1 0 15364 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0763_
timestamp 1
transform -1 0 16744 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0764_
timestamp 1
transform -1 0 16376 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0765_
timestamp 1
transform 1 0 16652 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0766_
timestamp 1
transform -1 0 16560 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0767_
timestamp 1
transform -1 0 17756 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0768_
timestamp 1
transform -1 0 14444 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0769_
timestamp 1
transform 1 0 17756 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0770_
timestamp 1
transform -1 0 15640 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0771_
timestamp 1
transform 1 0 9568 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0772_
timestamp 1
transform -1 0 10120 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0773_
timestamp 1
transform -1 0 10856 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0774_
timestamp 1
transform 1 0 9108 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0775_
timestamp 1
transform -1 0 10764 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0776_
timestamp 1
transform 1 0 10856 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _0777_
timestamp 1
transform 1 0 9568 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0778_
timestamp 1
transform 1 0 11408 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0779_
timestamp 1
transform -1 0 12696 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0780_
timestamp 1
transform 1 0 12236 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0781_
timestamp 1
transform 1 0 13432 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0782_
timestamp 1
transform 1 0 11960 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0783_
timestamp 1
transform 1 0 13892 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0784_
timestamp 1
transform -1 0 13340 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0785_
timestamp 1
transform 1 0 12420 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__o211ai_1  _0786_
timestamp 1
transform -1 0 13892 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _0787_
timestamp 1
transform 1 0 11684 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0788_
timestamp 1
transform -1 0 11132 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _0789_
timestamp 1
transform -1 0 10028 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0790_
timestamp 1
transform 1 0 10028 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0791_
timestamp 1
transform 1 0 9016 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0792_
timestamp 1
transform 1 0 9108 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0793_
timestamp 1
transform 1 0 8740 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0794_
timestamp 1
transform -1 0 8740 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _0795_
timestamp 1
transform 1 0 6992 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0796_
timestamp 1
transform -1 0 8188 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0797_
timestamp 1
transform 1 0 6348 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0798_
timestamp 1
transform -1 0 7544 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _0799_
timestamp 1
transform 1 0 7360 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0800_
timestamp 1
transform -1 0 6532 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0801_
timestamp 1
transform 1 0 6532 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0802_
timestamp 1
transform -1 0 5796 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0803_
timestamp 1
transform 1 0 5612 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0804_
timestamp 1
transform 1 0 4692 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0805_
timestamp 1
transform -1 0 7084 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0806_
timestamp 1
transform 1 0 6624 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _0807_
timestamp 1
transform 1 0 6348 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0808_
timestamp 1
transform 1 0 5060 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0809_
timestamp 1
transform 1 0 7084 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0810_
timestamp 1
transform -1 0 6624 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0811_
timestamp 1
transform 1 0 4600 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0812_
timestamp 1
transform 1 0 4876 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__o21ba_1  _0813_
timestamp 1
transform 1 0 6348 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _0814_
timestamp 1
transform 1 0 4784 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0815_
timestamp 1
transform -1 0 6072 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0816_
timestamp 1
transform 1 0 4324 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__o21ba_2  _0817_
timestamp 1
transform 1 0 11408 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0818_
timestamp 1
transform 1 0 5888 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0819_
timestamp 1
transform -1 0 5888 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0820_
timestamp 1
transform 1 0 5244 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0821_
timestamp 1
transform -1 0 5888 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0822_
timestamp 1
transform -1 0 7268 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0823_
timestamp 1
transform -1 0 7820 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _0824_
timestamp 1
transform 1 0 6348 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0825_
timestamp 1
transform 1 0 5888 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0826_
timestamp 1
transform -1 0 8924 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0827_
timestamp 1
transform -1 0 8188 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0828_
timestamp 1
transform 1 0 10304 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0829_
timestamp 1
transform 1 0 8924 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0830_
timestamp 1
transform 1 0 8188 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0831_
timestamp 1
transform -1 0 10028 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o221ai_4  _0832_
timestamp 1
transform 1 0 8924 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__a32o_1  _0833_
timestamp 1
transform -1 0 9384 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0834_
timestamp 1
transform -1 0 9568 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0835_
timestamp 1
transform 1 0 8464 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0836_
timestamp 1
transform 1 0 9384 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _0837_
timestamp 1
transform 1 0 8188 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0838_
timestamp 1
transform -1 0 8188 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0839_
timestamp 1
transform 1 0 5428 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0840_
timestamp 1
transform -1 0 6808 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0841_
timestamp 1
transform -1 0 6072 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0842_
timestamp 1
transform 1 0 5612 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0843_
timestamp 1
transform -1 0 5520 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0844_
timestamp 1
transform 1 0 5152 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0845_
timestamp 1
transform -1 0 5612 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0846_
timestamp 1
transform 1 0 3772 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nor4_1  _0847_
timestamp 1
transform -1 0 5796 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0848_
timestamp 1
transform -1 0 6256 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0849_
timestamp 1
transform 1 0 4600 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0850_
timestamp 1
transform 1 0 4324 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _0851_
timestamp 1
transform 1 0 3956 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0852_
timestamp 1
transform -1 0 6164 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0853_
timestamp 1
transform -1 0 5888 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0854_
timestamp 1
transform -1 0 5428 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0855_
timestamp 1
transform -1 0 6072 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0856_
timestamp 1
transform 1 0 4232 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0857_
timestamp 1
transform -1 0 5612 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0858_
timestamp 1
transform -1 0 5520 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0859_
timestamp 1
transform -1 0 6900 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0860_
timestamp 1
transform -1 0 9476 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _0861_
timestamp 1
transform -1 0 6256 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0862_
timestamp 1
transform 1 0 6164 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_1  _0863_
timestamp 1
transform 1 0 6992 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0864_
timestamp 1
transform -1 0 8096 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0865_
timestamp 1
transform 1 0 8924 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0866_
timestamp 1
transform -1 0 8556 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0867_
timestamp 1
transform -1 0 9568 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0868_
timestamp 1
transform 1 0 8924 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0869_
timestamp 1
transform 1 0 9752 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0870_
timestamp 1
transform 1 0 26036 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0871_
timestamp 1
transform 1 0 26220 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0872_
timestamp 1
transform -1 0 26220 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0873_
timestamp 1
transform -1 0 24104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0874_
timestamp 1
transform 1 0 23736 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0875_
timestamp 1
transform 1 0 24380 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_1  _0876_
timestamp 1
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _0877_
timestamp 1
transform -1 0 26772 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0878_
timestamp 1
transform 1 0 25944 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0879_
timestamp 1
transform 1 0 25116 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _0880_
timestamp 1
transform -1 0 25024 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or4bb_1  _0881_
timestamp 1
transform 1 0 25668 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0882_
timestamp 1
transform 1 0 26404 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _0883_
timestamp 1
transform -1 0 26588 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _0884_
timestamp 1
transform -1 0 28244 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_1  _0885_
timestamp 1
transform 1 0 26312 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _0886_
timestamp 1
transform 1 0 25484 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _0887_
timestamp 1
transform 1 0 24380 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0888_
timestamp 1
transform 1 0 24840 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _0889_
timestamp 1
transform -1 0 27600 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_1  _0890_
timestamp 1
transform 1 0 26220 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0891_
timestamp 1
transform 1 0 25392 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0892_
timestamp 1
transform 1 0 25116 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _0893_
timestamp 1
transform 1 0 23276 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_1  _0894_
timestamp 1
transform 1 0 25576 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__o21a_1  _0895_
timestamp 1
transform 1 0 25668 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0896_
timestamp 1
transform 1 0 25576 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _0897_
timestamp 1
transform 1 0 23644 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _0898_
timestamp 1
transform 1 0 24104 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_1  _0899_
timestamp 1
transform -1 0 24748 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _0900_
timestamp 1
transform 1 0 24380 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dfstp_1  _0901_
timestamp 1
transform -1 0 13892 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0902_
timestamp 1
transform 1 0 12144 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0903_
timestamp 1
transform 1 0 9568 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0904_
timestamp 1
transform 1 0 14628 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0905_
timestamp 1
transform 1 0 11500 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0906_
timestamp 1
transform 1 0 24380 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0907_
timestamp 1
transform 1 0 25208 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0908_
timestamp 1
transform 1 0 26496 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0909_
timestamp 1
transform 1 0 17848 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0910_
timestamp 1
transform 1 0 19228 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0911_
timestamp 1
transform 1 0 19872 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0912_
timestamp 1
transform -1 0 23736 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0913_
timestamp 1
transform 1 0 20884 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0914_
timestamp 1
transform 1 0 19780 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0915_
timestamp 1
transform -1 0 18860 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0916_
timestamp 1
transform -1 0 18216 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0917_
timestamp 1
transform 1 0 15456 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0918_
timestamp 1
transform 1 0 12420 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0919_
timestamp 1
transform 1 0 12052 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0920_
timestamp 1
transform 1 0 13800 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0921_
timestamp 1
transform 1 0 11592 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0922_
timestamp 1
transform -1 0 13708 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0923_
timestamp 1
transform 1 0 9568 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  _0924__65
timestamp 1
transform -1 0 8556 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _0924_
timestamp 1
transform 1 0 8004 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0925_
timestamp 1
transform -1 0 9660 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0926_
timestamp 1
transform 1 0 6900 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0927_
timestamp 1
transform 1 0 8924 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0928_
timestamp 1
transform 1 0 10672 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0929_
timestamp 1
transform 1 0 11776 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0930_
timestamp 1
transform 1 0 10948 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  _0931__64
timestamp 1
transform -1 0 5152 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _0931_
timestamp 1
transform 1 0 4416 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  _0932__63
timestamp 1
transform -1 0 5796 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _0932_
timestamp 1
transform 1 0 5152 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0933_
timestamp 1
transform 1 0 15088 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0934_
timestamp 1
transform 1 0 16836 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0935_
timestamp 1
transform 1 0 19228 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0936_
timestamp 1
transform 1 0 20424 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0937_
timestamp 1
transform 1 0 21436 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0938_
timestamp 1
transform 1 0 21804 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0939_
timestamp 1
transform 1 0 22080 0 1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0940_
timestamp 1
transform 1 0 17848 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0941_
timestamp 1
transform 1 0 19872 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0942_
timestamp 1
transform 1 0 21528 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0943_
timestamp 1
transform 1 0 22448 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0944_
timestamp 1
transform -1 0 24288 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0945_
timestamp 1
transform -1 0 24472 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0946_
timestamp 1
transform -1 0 20976 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0947_
timestamp 1
transform -1 0 21068 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0948_
timestamp 1
transform -1 0 17940 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0949_
timestamp 1
transform 1 0 14720 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0950_
timestamp 1
transform 1 0 14720 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0951_
timestamp 1
transform 1 0 14444 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0952_
timestamp 1
transform -1 0 14260 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0953_
timestamp 1
transform -1 0 12788 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0954_
timestamp 1
transform 1 0 8924 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0955_
timestamp 1
transform 1 0 8924 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0956_
timestamp 1
transform 1 0 17204 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0957_
timestamp 1
transform 1 0 17296 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0958_
timestamp 1
transform 1 0 18124 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0959_
timestamp 1
transform 1 0 19872 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0960_
timestamp 1
transform 1 0 21712 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0961_
timestamp 1
transform 1 0 23460 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0962_
timestamp 1
transform 1 0 25024 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0963_
timestamp 1
transform 1 0 26128 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0964_
timestamp 1
transform 1 0 13800 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0965_
timestamp 1
transform 1 0 17572 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0966_
timestamp 1
transform 1 0 17296 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0967_
timestamp 1
transform 1 0 19228 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0968_
timestamp 1
transform 1 0 21068 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0969_
timestamp 1
transform 1 0 22724 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0970_
timestamp 1
transform -1 0 26312 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0971_
timestamp 1
transform 1 0 26312 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0972_
timestamp 1
transform 1 0 26496 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0973_
timestamp 1
transform 1 0 14720 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0974_
timestamp 1
transform 1 0 14168 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0975_
timestamp 1
transform 1 0 14444 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0976_
timestamp 1
transform 1 0 14260 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0977_
timestamp 1
transform 1 0 15180 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0978_
timestamp 1
transform 1 0 9016 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0979_
timestamp 1
transform 1 0 8740 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0980_
timestamp 1
transform 1 0 11868 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0981_
timestamp 1
transform 1 0 11960 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0982_
timestamp 1
transform -1 0 11224 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0983_
timestamp 1
transform 1 0 8188 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0984_
timestamp 1
transform -1 0 6624 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0985_
timestamp 1
transform 1 0 3312 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0986_
timestamp 1
transform 1 0 3220 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0987_
timestamp 1
transform 1 0 3036 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0988_
timestamp 1
transform 1 0 3312 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0989_
timestamp 1
transform 1 0 4416 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0990_
timestamp 1
transform 1 0 5060 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0991_
timestamp 1
transform 1 0 8556 0 -1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0992_
timestamp 1
transform 1 0 8924 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0993_
timestamp 1
transform 1 0 7544 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0994_
timestamp 1
transform -1 0 6256 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0995_
timestamp 1
transform 1 0 1840 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0996_
timestamp 1
transform 1 0 2116 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0997_
timestamp 1
transform 1 0 3588 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0998_
timestamp 1
transform -1 0 5888 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0999_
timestamp 1
transform 1 0 5980 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1000_
timestamp 1
transform 1 0 7820 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1001_
timestamp 1
transform 1 0 9568 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1002_
timestamp 1
transform -1 0 24288 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1003_
timestamp 1
transform 1 0 19228 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1004_
timestamp 1
transform 1 0 19872 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1005_
timestamp 1
transform -1 0 23644 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1006_
timestamp 1
transform 1 0 24012 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1007_
timestamp 1
transform -1 0 26220 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1008_
timestamp 1
transform 1 0 26496 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1009_
timestamp 1
transform 1 0 26496 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1010_
timestamp 1
transform 1 0 26496 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1011_
timestamp 1
transform -1 0 22908 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1012_
timestamp 1
transform 1 0 21160 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1013_
timestamp 1
transform 1 0 21804 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1014_
timestamp 1
transform -1 0 23644 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1015_
timestamp 1
transform 1 0 24104 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1016_
timestamp 1
transform 1 0 26496 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1017_
timestamp 1
transform 1 0 26496 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1018_
timestamp 1
transform 1 0 26220 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1019_
timestamp 1
transform 1 0 26312 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1020_
timestamp 1
transform -1 0 26864 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1021_
timestamp 1
transform -1 0 26496 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1022_
timestamp 1
transform 1 0 21252 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1023_
timestamp 1
transform 1 0 21804 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1024_
timestamp 1
transform 1 0 23644 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1025_
timestamp 1
transform 1 0 23000 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1026_
timestamp 1
transform -1 0 28336 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1027_
timestamp 1
transform -1 0 28336 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1028_
timestamp 1
transform -1 0 28336 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1029_
timestamp 1
transform -1 0 28336 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 1
transform 1 0 15272 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_clk
timestamp 1
transform 1 0 6992 0 -1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_clk
timestamp 1
transform -1 0 7820 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_clk
timestamp 1
transform -1 0 12604 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_clk
timestamp 1
transform 1 0 11960 0 -1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_clk
timestamp 1
transform 1 0 6900 0 1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_clk
timestamp 1
transform 1 0 7820 0 1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_clk
timestamp 1
transform 1 0 13432 0 -1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_clk
timestamp 1
transform -1 0 14168 0 -1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_clk
timestamp 1
transform -1 0 22816 0 -1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_clk
timestamp 1
transform -1 0 20516 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_clk
timestamp 1
transform 1 0 24564 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_clk
timestamp 1
transform 1 0 25208 0 -1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_clk
timestamp 1
transform 1 0 19320 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_clk
timestamp 1
transform 1 0 19044 0 -1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_clk
timestamp 1
transform 1 0 24288 0 -1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_clk
timestamp 1
transform 1 0 24380 0 1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_2  clkload0
timestamp 1
transform -1 0 6992 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkinvlp_4  clkload1
timestamp 1
transform 1 0 6808 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_4  clkload2
timestamp 1
transform 1 0 11592 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__clkinvlp_4  clkload3
timestamp 1
transform 1 0 13708 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__bufinv_16  clkload4
timestamp 1
transform -1 0 9108 0 -1 21760
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_2  clkload5
timestamp 1
transform 1 0 7268 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  clkload6
timestamp 1
transform -1 0 13432 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  clkload7
timestamp 1
transform 1 0 13340 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkinvlp_4  clkload8
timestamp 1
transform -1 0 21528 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  clkload9
timestamp 1
transform 1 0 19504 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkload10
timestamp 1
transform 1 0 24564 0 -1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__bufinv_16  clkload11
timestamp 1
transform -1 0 21528 0 -1 19584
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_4  clkload12
timestamp 1
transform 1 0 19228 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  clkload13
timestamp 1
transform 1 0 23184 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  clkload14
timestamp 1
transform -1 0 24932 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout17
timestamp 1
transform -1 0 13800 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout19
timestamp 1
transform 1 0 19320 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout20
timestamp 1
transform 1 0 17848 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout21
timestamp 1
transform -1 0 13892 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout22
timestamp 1
transform -1 0 19136 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout23
timestamp 1
transform -1 0 12420 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout24
timestamp 1
transform -1 0 13616 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout25
timestamp 1
transform 1 0 14628 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout26
timestamp 1
transform -1 0 12052 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout27
timestamp 1
transform -1 0 12420 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout28
timestamp 1
transform -1 0 11960 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout29
timestamp 1
transform 1 0 18492 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout30
timestamp 1
transform -1 0 17480 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout31
timestamp 1
transform -1 0 20516 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout32
timestamp 1
transform 1 0 19688 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout33
timestamp 1
transform 1 0 23736 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout34
timestamp 1
transform -1 0 20240 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout35
timestamp 1
transform -1 0 24748 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout36
timestamp 1
transform -1 0 21068 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout37
timestamp 1
transform 1 0 14076 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout38
timestamp 1
transform -1 0 12144 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout39
timestamp 1
transform -1 0 12236 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout40
timestamp 1
transform -1 0 11960 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout41
timestamp 1
transform -1 0 9844 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout42
timestamp 1
transform 1 0 11500 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout43
timestamp 1
transform -1 0 12512 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout44
timestamp 1
transform -1 0 15916 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout45
timestamp 1
transform -1 0 16284 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout46
timestamp 1
transform -1 0 13800 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout47
timestamp 1
transform -1 0 14628 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout48
timestamp 1
transform -1 0 9476 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout49
timestamp 1
transform -1 0 14260 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout50
timestamp 1
transform 1 0 15272 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout51
timestamp 1
transform -1 0 13156 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout52
timestamp 1
transform -1 0 25024 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout53
timestamp 1
transform 1 0 27692 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout54
timestamp 1
transform 1 0 27508 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout55
timestamp 1
transform -1 0 28336 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout56
timestamp 1
transform -1 0 21620 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout57
timestamp 1
transform 1 0 20700 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout58
timestamp 1
transform -1 0 28244 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout59
timestamp 1
transform 1 0 27876 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout60
timestamp 1
transform -1 0 28060 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout61
timestamp 1
transform -1 0 28244 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout62
timestamp 1
transform 1 0 27876 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3
timestamp 1636968456
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1636968456
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp 1
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1636968456
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1636968456
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp 1
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1636968456
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1636968456
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1636968456
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1636968456
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1636968456
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1636968456
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1636968456
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1636968456
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1636968456
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1636968456
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1636968456
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_209
timestamp 1
transform 1 0 20332 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_217
timestamp 1
transform 1 0 21068 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_230
timestamp 1
transform 1 0 22264 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_237
timestamp 1
transform 1 0 22908 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_244
timestamp 1
transform 1 0 23552 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1636968456
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1636968456
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1636968456
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_293
timestamp 1
transform 1 0 28060 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1636968456
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1636968456
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1636968456
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1636968456
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_64
timestamp 1636968456
transform 1 0 6992 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_76
timestamp 1
transform 1 0 8096 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_97
timestamp 1636968456
transform 1 0 10028 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_109
timestamp 1
transform 1 0 11132 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_113
timestamp 1
transform 1 0 11500 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_119
timestamp 1
transform 1 0 12052 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_138
timestamp 1
transform 1 0 13800 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_147
timestamp 1636968456
transform 1 0 14628 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_159
timestamp 1
transform 1 0 15732 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_175
timestamp 1636968456
transform 1 0 17204 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_187
timestamp 1
transform 1 0 18308 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_193
timestamp 1
transform 1 0 18860 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1636968456
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_265
timestamp 1
transform 1 0 25484 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_276
timestamp 1
transform 1 0 26496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_281
timestamp 1
transform 1 0 26956 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_296
timestamp 1
transform 1 0 28336 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1636968456
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1636968456
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_29
timestamp 1
transform 1 0 3772 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_37
timestamp 1
transform 1 0 4508 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_75
timestamp 1
transform 1 0 8004 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_85
timestamp 1
transform 1 0 8924 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_89
timestamp 1
transform 1 0 9292 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_117
timestamp 1
transform 1 0 11868 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_149
timestamp 1
transform 1 0 14812 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_183
timestamp 1
transform 1 0 17940 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_189
timestamp 1
transform 1 0 18492 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_213
timestamp 1
transform 1 0 20700 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_253
timestamp 1
transform 1 0 24380 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_260
timestamp 1
transform 1 0 25024 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_296
timestamp 1
transform 1 0 28336 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1636968456
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1636968456
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1636968456
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1636968456
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_70
timestamp 1
transform 1 0 7544 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_78
timestamp 1
transform 1 0 8280 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_97
timestamp 1
transform 1 0 10028 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_109
timestamp 1
transform 1 0 11132 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_113
timestamp 1
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_123
timestamp 1
transform 1 0 12420 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_147
timestamp 1636968456
transform 1 0 14628 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_159
timestamp 1
transform 1 0 15732 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_178
timestamp 1
transform 1 0 17480 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1636968456
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_237
timestamp 1
transform 1 0 22908 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_258
timestamp 1
transform 1 0 24840 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_295
timestamp 1
transform 1 0 28244 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1636968456
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1636968456
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_29
timestamp 1
transform 1 0 3772 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_37
timestamp 1
transform 1 0 4508 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_51
timestamp 1
transform 1 0 5796 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_63
timestamp 1
transform 1 0 6900 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_85
timestamp 1
transform 1 0 8924 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_107
timestamp 1
transform 1 0 10948 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_115
timestamp 1
transform 1 0 11684 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1636968456
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_153
timestamp 1
transform 1 0 15180 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_157
timestamp 1
transform 1 0 15548 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_176
timestamp 1
transform 1 0 17296 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_184
timestamp 1
transform 1 0 18032 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_211
timestamp 1
transform 1 0 20516 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1636968456
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_265
timestamp 1
transform 1 0 25484 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_269
timestamp 1
transform 1 0 25852 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_296
timestamp 1
transform 1 0 28336 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1636968456
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_15
timestamp 1
transform 1 0 2484 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_23
timestamp 1
transform 1 0 3220 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_44
timestamp 1
transform 1 0 5152 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_48
timestamp 1
transform 1 0 5520 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_95
timestamp 1636968456
transform 1 0 9844 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_107
timestamp 1
transform 1 0 10948 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1636968456
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_125
timestamp 1
transform 1 0 12604 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_131
timestamp 1636968456
transform 1 0 13156 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_143
timestamp 1
transform 1 0 14260 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_151
timestamp 1
transform 1 0 14996 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_176
timestamp 1
transform 1 0 17296 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_186
timestamp 1
transform 1 0 18216 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_206
timestamp 1636968456
transform 1 0 20056 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_218
timestamp 1
transform 1 0 21160 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1636968456
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_293
timestamp 1
transform 1 0 28060 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1636968456
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1636968456
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1636968456
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1636968456
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_66
timestamp 1636968456
transform 1 0 7176 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_78
timestamp 1
transform 1 0 8280 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1636968456
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1636968456
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1636968456
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1636968456
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_141
timestamp 1
transform 1 0 14076 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_147
timestamp 1
transform 1 0 14628 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_183
timestamp 1636968456
transform 1 0 17940 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1636968456
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_209
timestamp 1
transform 1 0 20332 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_217
timestamp 1
transform 1 0 21068 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_238
timestamp 1
transform 1 0 23000 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_249
timestamp 1
transform 1 0 24012 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_267
timestamp 1
transform 1 0 25668 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_296
timestamp 1
transform 1 0 28336 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1636968456
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1636968456
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1636968456
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1636968456
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1636968456
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1636968456
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1636968456
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1636968456
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_113
timestamp 1
transform 1 0 11500 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_136
timestamp 1636968456
transform 1 0 13616 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_148
timestamp 1
transform 1 0 14720 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_178
timestamp 1
transform 1 0 17480 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_182
timestamp 1
transform 1 0 17848 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_188
timestamp 1636968456
transform 1 0 18400 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_200
timestamp 1636968456
transform 1 0 19504 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_212
timestamp 1636968456
transform 1 0 20608 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_260
timestamp 1
transform 1 0 25024 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_268
timestamp 1
transform 1 0 25760 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_276
timestamp 1
transform 1 0 26496 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_281
timestamp 1
transform 1 0 26956 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_289
timestamp 1
transform 1 0 27692 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_293
timestamp 1
transform 1 0 28060 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1636968456
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1636968456
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1636968456
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1636968456
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1636968456
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1636968456
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_85
timestamp 1
transform 1 0 8924 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_91
timestamp 1
transform 1 0 9476 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_105
timestamp 1
transform 1 0 10764 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_137
timestamp 1
transform 1 0 13708 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_145
timestamp 1636968456
transform 1 0 14444 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_157
timestamp 1636968456
transform 1 0 15548 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_169
timestamp 1636968456
transform 1 0 16652 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_181
timestamp 1
transform 1 0 17756 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_187
timestamp 1
transform 1 0 18308 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1636968456
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1636968456
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1636968456
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1636968456
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_245
timestamp 1
transform 1 0 23644 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1636968456
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_265
timestamp 1
transform 1 0 25484 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_273
timestamp 1
transform 1 0 26220 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_296
timestamp 1
transform 1 0 28336 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1636968456
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_15
timestamp 1
transform 1 0 2484 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_52
timestamp 1
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_68
timestamp 1636968456
transform 1 0 7360 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_80
timestamp 1
transform 1 0 8464 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_113
timestamp 1
transform 1 0 11500 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_117
timestamp 1
transform 1 0 11868 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_133
timestamp 1636968456
transform 1 0 13340 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_145
timestamp 1636968456
transform 1 0 14444 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_157
timestamp 1
transform 1 0 15548 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_165
timestamp 1
transform 1 0 16284 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_169
timestamp 1
transform 1 0 16652 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_177
timestamp 1
transform 1 0 17388 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_200
timestamp 1
transform 1 0 19504 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1636968456
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1636968456
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_249
timestamp 1
transform 1 0 24012 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_257
timestamp 1
transform 1 0 24748 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_265
timestamp 1
transform 1 0 25484 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_278
timestamp 1
transform 1 0 26680 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1636968456
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_293
timestamp 1
transform 1 0 28060 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1636968456
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1636968456
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_29
timestamp 1
transform 1 0 3772 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_37
timestamp 1
transform 1 0 4508 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_71
timestamp 1636968456
transform 1 0 7636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_85
timestamp 1
transform 1 0 8924 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_113
timestamp 1636968456
transform 1 0 11500 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_125
timestamp 1636968456
transform 1 0 12604 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_137
timestamp 1
transform 1 0 13708 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_141
timestamp 1
transform 1 0 14076 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_147
timestamp 1
transform 1 0 14628 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_155
timestamp 1
transform 1 0 15364 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_167
timestamp 1
transform 1 0 16468 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_177
timestamp 1
transform 1 0 17388 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_181
timestamp 1
transform 1 0 17756 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_197
timestamp 1
transform 1 0 19228 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_204
timestamp 1636968456
transform 1 0 19872 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_216
timestamp 1636968456
transform 1 0 20976 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_228
timestamp 1636968456
transform 1 0 22080 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_240
timestamp 1
transform 1 0 23184 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_266
timestamp 1
transform 1 0 25576 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1636968456
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_289
timestamp 1
transform 1 0 27692 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_293
timestamp 1
transform 1 0 28060 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1636968456
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_15
timestamp 1
transform 1 0 2484 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_11_50
timestamp 1
transform 1 0 5704 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_11_68
timestamp 1
transform 1 0 7360 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_76
timestamp 1
transform 1 0 8096 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_81
timestamp 1
transform 1 0 8556 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_85
timestamp 1
transform 1 0 8924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_106
timestamp 1
transform 1 0 10856 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_11_113
timestamp 1
transform 1 0 11500 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_121
timestamp 1
transform 1 0 12236 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_164
timestamp 1
transform 1 0 16192 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_183
timestamp 1636968456
transform 1 0 17940 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_195
timestamp 1
transform 1 0 19044 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_199
timestamp 1
transform 1 0 19412 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_220
timestamp 1
transform 1 0 21344 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_246
timestamp 1
transform 1 0 23736 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_272
timestamp 1
transform 1 0 26128 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1636968456
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_293
timestamp 1
transform 1 0 28060 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1636968456
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1636968456
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1636968456
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_41
timestamp 1
transform 1 0 4876 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_51
timestamp 1
transform 1 0 5796 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_71
timestamp 1636968456
transform 1 0 7636 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_85
timestamp 1
transform 1 0 8924 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_91
timestamp 1
transform 1 0 9476 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_114
timestamp 1
transform 1 0 11592 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_118
timestamp 1
transform 1 0 11960 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_141
timestamp 1
transform 1 0 14076 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_156
timestamp 1636968456
transform 1 0 15456 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_168
timestamp 1
transform 1 0 16560 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_174
timestamp 1636968456
transform 1 0 17112 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_186
timestamp 1
transform 1 0 18216 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_197
timestamp 1
transform 1 0 19228 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_244
timestamp 1
transform 1 0 23552 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_248
timestamp 1
transform 1 0 23920 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_263
timestamp 1
transform 1 0 25300 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_279
timestamp 1
transform 1 0 26772 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_290
timestamp 1
transform 1 0 27784 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_296
timestamp 1
transform 1 0 28336 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1636968456
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1636968456
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1636968456
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1636968456
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_71
timestamp 1636968456
transform 1 0 7636 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_83
timestamp 1636968456
transform 1 0 8740 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_95
timestamp 1636968456
transform 1 0 9844 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_107
timestamp 1
transform 1 0 10948 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_113
timestamp 1
transform 1 0 11500 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_121
timestamp 1
transform 1 0 12236 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_125
timestamp 1
transform 1 0 12604 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1636968456
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_187
timestamp 1
transform 1 0 18308 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_214
timestamp 1
transform 1 0 20792 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_222
timestamp 1
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_236
timestamp 1636968456
transform 1 0 22816 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_248
timestamp 1
transform 1 0 23920 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_254
timestamp 1
transform 1 0 24472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_266
timestamp 1
transform 1 0 25576 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_270
timestamp 1
transform 1 0 25944 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_295
timestamp 1
transform 1 0 28244 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1636968456
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1636968456
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1636968456
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_41
timestamp 1
transform 1 0 4876 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_48
timestamp 1
transform 1 0 5520 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_56
timestamp 1
transform 1 0 6256 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_76
timestamp 1
transform 1 0 8096 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_105
timestamp 1
transform 1 0 10764 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_113
timestamp 1
transform 1 0 11500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_125
timestamp 1636968456
transform 1 0 12604 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_137
timestamp 1
transform 1 0 13708 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_146
timestamp 1636968456
transform 1 0 14536 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_193
timestamp 1
transform 1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_197
timestamp 1
transform 1 0 19228 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_216
timestamp 1636968456
transform 1 0 20976 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_228
timestamp 1636968456
transform 1 0 22080 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_240
timestamp 1636968456
transform 1 0 23184 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_266
timestamp 1
transform 1 0 25576 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_272
timestamp 1
transform 1 0 26128 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_296
timestamp 1
transform 1 0 28336 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1636968456
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1636968456
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1636968456
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_39
timestamp 1
transform 1 0 4692 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_95
timestamp 1
transform 1 0 9844 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_102
timestamp 1
transform 1 0 10488 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_113
timestamp 1
transform 1 0 11500 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_121
timestamp 1
transform 1 0 12236 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_128
timestamp 1
transform 1 0 12880 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_138
timestamp 1636968456
transform 1 0 13800 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_150
timestamp 1
transform 1 0 14904 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_15_169
timestamp 1
transform 1 0 16652 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_193
timestamp 1
transform 1 0 18860 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_201
timestamp 1
transform 1 0 19596 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_225
timestamp 1
transform 1 0 21804 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_253
timestamp 1
transform 1 0 24380 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_261
timestamp 1
transform 1 0 25116 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_281
timestamp 1
transform 1 0 26956 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_287
timestamp 1
transform 1 0 27508 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_295
timestamp 1
transform 1 0 28244 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1636968456
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1636968456
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_29
timestamp 1
transform 1 0 3772 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_44
timestamp 1
transform 1 0 5152 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_76
timestamp 1
transform 1 0 8096 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_148
timestamp 1
transform 1 0 14720 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_176
timestamp 1636968456
transform 1 0 17296 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_188
timestamp 1
transform 1 0 18400 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_197
timestamp 1
transform 1 0 19228 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_219
timestamp 1
transform 1 0 21252 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_223
timestamp 1
transform 1 0 21620 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1636968456
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_265
timestamp 1
transform 1 0 25484 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_273
timestamp 1
transform 1 0 26220 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_294
timestamp 1
transform 1 0 28152 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1636968456
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_15
timestamp 1
transform 1 0 2484 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_23
timestamp 1
transform 1 0 3220 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_57
timestamp 1
transform 1 0 6348 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_61
timestamp 1
transform 1 0 6716 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_73
timestamp 1
transform 1 0 7820 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_77
timestamp 1
transform 1 0 8188 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_81
timestamp 1
transform 1 0 8556 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_89
timestamp 1
transform 1 0 9292 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_113
timestamp 1
transform 1 0 11500 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_117
timestamp 1
transform 1 0 11868 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_143
timestamp 1636968456
transform 1 0 14260 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_155
timestamp 1636968456
transform 1 0 15364 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1636968456
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_181
timestamp 1
transform 1 0 17756 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_187
timestamp 1
transform 1 0 18308 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_216
timestamp 1
transform 1 0 20976 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_225
timestamp 1
transform 1 0 21804 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_254
timestamp 1
transform 1 0 24472 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_17_286
timestamp 1
transform 1 0 27416 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1636968456
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1636968456
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1636968456
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_41
timestamp 1
transform 1 0 4876 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_55
timestamp 1636968456
transform 1 0 6164 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_67
timestamp 1636968456
transform 1 0 7268 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_79
timestamp 1
transform 1 0 8372 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1636968456
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_103
timestamp 1
transform 1 0 10580 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_117
timestamp 1
transform 1 0 11868 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_141
timestamp 1
transform 1 0 14076 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_149
timestamp 1636968456
transform 1 0 14812 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_161
timestamp 1636968456
transform 1 0 15916 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_173
timestamp 1636968456
transform 1 0 17020 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_185
timestamp 1
transform 1 0 18124 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_189
timestamp 1
transform 1 0 18492 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_217
timestamp 1
transform 1 0 21068 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_223
timestamp 1
transform 1 0 21620 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1636968456
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_265
timestamp 1
transform 1 0 25484 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_293
timestamp 1
transform 1 0 28060 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1636968456
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1636968456
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1636968456
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1636968456
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1636968456
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1636968456
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1636968456
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1636968456
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_113
timestamp 1
transform 1 0 11500 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_118
timestamp 1
transform 1 0 11960 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_129
timestamp 1
transform 1 0 12972 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_133
timestamp 1
transform 1 0 13340 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_169
timestamp 1
transform 1 0 16652 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_173
timestamp 1
transform 1 0 17020 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_182
timestamp 1636968456
transform 1 0 17848 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_216
timestamp 1
transform 1 0 20976 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_245
timestamp 1
transform 1 0 23644 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_254
timestamp 1
transform 1 0 24472 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_276
timestamp 1
transform 1 0 26496 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_287
timestamp 1
transform 1 0 27508 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1636968456
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1636968456
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1636968456
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_41
timestamp 1
transform 1 0 4876 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_63
timestamp 1636968456
transform 1 0 6900 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_75
timestamp 1
transform 1 0 8004 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1636968456
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1636968456
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1636968456
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1636968456
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1636968456
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_153
timestamp 1
transform 1 0 15180 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_162
timestamp 1
transform 1 0 16008 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_183
timestamp 1636968456
transform 1 0 17940 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1636968456
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1636968456
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_221
timestamp 1
transform 1 0 21436 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_250
timestamp 1
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1636968456
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_265
timestamp 1
transform 1 0 25484 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_273
timestamp 1
transform 1 0 26220 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_296
timestamp 1
transform 1 0 28336 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1636968456
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1636968456
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_27
timestamp 1
transform 1 0 3588 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_35
timestamp 1
transform 1 0 4324 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_65
timestamp 1
transform 1 0 7084 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_73
timestamp 1
transform 1 0 7820 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_21_104
timestamp 1
transform 1 0 10672 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_21_113
timestamp 1
transform 1 0 11500 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_119
timestamp 1
transform 1 0 12052 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_137
timestamp 1
transform 1 0 13708 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_145
timestamp 1
transform 1 0 14444 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_183
timestamp 1
transform 1 0 17940 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_191
timestamp 1
transform 1 0 18676 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_198
timestamp 1
transform 1 0 19320 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_212
timestamp 1636968456
transform 1 0 20608 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_233
timestamp 1636968456
transform 1 0 22540 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_245
timestamp 1
transform 1 0 23644 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_249
timestamp 1
transform 1 0 24012 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_270
timestamp 1
transform 1 0 25944 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_278
timestamp 1
transform 1 0 26680 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_281
timestamp 1
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1636968456
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1636968456
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1636968456
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_41
timestamp 1
transform 1 0 4876 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_73
timestamp 1
transform 1 0 7820 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_105
timestamp 1
transform 1 0 10764 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1636968456
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_153
timestamp 1
transform 1 0 15180 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_174
timestamp 1
transform 1 0 17112 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_182
timestamp 1
transform 1 0 17848 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_188
timestamp 1
transform 1 0 18400 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_218
timestamp 1636968456
transform 1 0 21160 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_230
timestamp 1636968456
transform 1 0 22264 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_242
timestamp 1
transform 1 0 23368 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1636968456
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_265
timestamp 1
transform 1 0 25484 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_273
timestamp 1
transform 1 0 26220 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_296
timestamp 1
transform 1 0 28336 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1636968456
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1636968456
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1636968456
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1636968456
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_57
timestamp 1
transform 1 0 6348 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_61
timestamp 1
transform 1 0 6716 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_67
timestamp 1636968456
transform 1 0 7268 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_98
timestamp 1636968456
transform 1 0 10120 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_113
timestamp 1
transform 1 0 11500 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_143
timestamp 1636968456
transform 1 0 14260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_155
timestamp 1
transform 1 0 15364 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_164
timestamp 1
transform 1 0 16192 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_177
timestamp 1
transform 1 0 17388 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_181
timestamp 1
transform 1 0 17756 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_203
timestamp 1
transform 1 0 19780 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_225
timestamp 1
transform 1 0 21804 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_235
timestamp 1636968456
transform 1 0 22724 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_247
timestamp 1636968456
transform 1 0 23828 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_259
timestamp 1636968456
transform 1 0 24932 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_271
timestamp 1
transform 1 0 26036 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_281
timestamp 1
transform 1 0 26956 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_293
timestamp 1
transform 1 0 28060 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1636968456
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1636968456
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1636968456
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1636968456
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1636968456
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1636968456
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_106
timestamp 1
transform 1 0 10856 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_114
timestamp 1
transform 1 0 11592 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_122
timestamp 1
transform 1 0 12328 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_126
timestamp 1
transform 1 0 12696 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_137
timestamp 1
transform 1 0 13708 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1636968456
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_167
timestamp 1636968456
transform 1 0 16468 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_179
timestamp 1
transform 1 0 17572 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_185
timestamp 1
transform 1 0 18124 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_219
timestamp 1
transform 1 0 21252 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_273
timestamp 1636968456
transform 1 0 26220 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_285
timestamp 1
transform 1 0 27324 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_295
timestamp 1
transform 1 0 28244 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1636968456
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1636968456
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_27
timestamp 1
transform 1 0 3588 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1636968456
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_69
timestamp 1
transform 1 0 7452 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_80
timestamp 1
transform 1 0 8464 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_97
timestamp 1636968456
transform 1 0 10028 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_109
timestamp 1
transform 1 0 11132 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_121
timestamp 1
transform 1 0 12236 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_131
timestamp 1
transform 1 0 13156 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_142
timestamp 1
transform 1 0 14168 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_177
timestamp 1
transform 1 0 17388 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_181
timestamp 1
transform 1 0 17756 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_210
timestamp 1
transform 1 0 20424 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_214
timestamp 1
transform 1 0 20792 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_221
timestamp 1
transform 1 0 21436 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_245
timestamp 1636968456
transform 1 0 23644 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_257
timestamp 1
transform 1 0 24748 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_278
timestamp 1
transform 1 0 26680 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1636968456
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_293
timestamp 1
transform 1 0 28060 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1636968456
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1636968456
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1636968456
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_41
timestamp 1
transform 1 0 4876 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_47
timestamp 1
transform 1 0 5428 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_62
timestamp 1636968456
transform 1 0 6808 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_74
timestamp 1
transform 1 0 7912 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_85
timestamp 1
transform 1 0 8924 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_91
timestamp 1636968456
transform 1 0 9476 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_103
timestamp 1
transform 1 0 10580 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_141
timestamp 1
transform 1 0 14076 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1636968456
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1636968456
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_193
timestamp 1
transform 1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1636968456
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1636968456
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_221
timestamp 1
transform 1 0 21436 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_235
timestamp 1
transform 1 0 22724 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_247
timestamp 1
transform 1 0 23828 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_253
timestamp 1
transform 1 0 24380 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_292
timestamp 1
transform 1 0 27968 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_296
timestamp 1
transform 1 0 28336 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1636968456
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1636968456
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1636968456
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_39
timestamp 1
transform 1 0 4692 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_43
timestamp 1
transform 1 0 5060 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_65
timestamp 1636968456
transform 1 0 7084 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_77
timestamp 1
transform 1 0 8188 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_100
timestamp 1636968456
transform 1 0 10304 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_113
timestamp 1
transform 1 0 11500 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_143
timestamp 1
transform 1 0 14260 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_151
timestamp 1
transform 1 0 14996 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_158
timestamp 1
transform 1 0 15640 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_183
timestamp 1
transform 1 0 17940 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_200
timestamp 1
transform 1 0 19504 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_214
timestamp 1
transform 1 0 20792 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_225
timestamp 1
transform 1 0 21804 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_234
timestamp 1
transform 1 0 22632 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_240
timestamp 1636968456
transform 1 0 23184 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_252
timestamp 1
transform 1 0 24288 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_260
timestamp 1
transform 1 0 25024 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_267
timestamp 1636968456
transform 1 0 25668 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_281
timestamp 1
transform 1 0 26956 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_295
timestamp 1
transform 1 0 28244 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_3
timestamp 1
transform 1 0 1380 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_7
timestamp 1
transform 1 0 1748 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_54
timestamp 1
transform 1 0 6072 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_58
timestamp 1
transform 1 0 6440 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_66
timestamp 1636968456
transform 1 0 7176 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_78
timestamp 1
transform 1 0 8280 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_85
timestamp 1
transform 1 0 8924 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_89
timestamp 1
transform 1 0 9292 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_113
timestamp 1636968456
transform 1 0 11500 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_125
timestamp 1636968456
transform 1 0 12604 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_137
timestamp 1
transform 1 0 13708 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1636968456
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_153
timestamp 1
transform 1 0 15180 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_161
timestamp 1
transform 1 0 15916 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_169
timestamp 1
transform 1 0 16652 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_217
timestamp 1
transform 1 0 21068 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_246
timestamp 1
transform 1 0 23736 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_270
timestamp 1
transform 1 0 25944 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_296
timestamp 1
transform 1 0 28336 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_3
timestamp 1
transform 1 0 1380 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1636968456
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_69
timestamp 1
transform 1 0 7452 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_108
timestamp 1
transform 1 0 11040 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_123
timestamp 1636968456
transform 1 0 12420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_135
timestamp 1
transform 1 0 13524 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_158
timestamp 1
transform 1 0 15640 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_165
timestamp 1
transform 1 0 16284 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_169
timestamp 1
transform 1 0 16652 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_173
timestamp 1
transform 1 0 17020 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_179
timestamp 1
transform 1 0 17572 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_196
timestamp 1
transform 1 0 19136 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_202
timestamp 1
transform 1 0 19688 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_208
timestamp 1
transform 1 0 20240 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_220
timestamp 1
transform 1 0 21344 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_225
timestamp 1
transform 1 0 21804 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_232
timestamp 1
transform 1 0 22448 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_250
timestamp 1
transform 1 0 24104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_259
timestamp 1
transform 1 0 24932 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_269
timestamp 1
transform 1 0 25852 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_277
timestamp 1
transform 1 0 26588 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1636968456
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_293
timestamp 1
transform 1 0 28060 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1636968456
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1636968456
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_29
timestamp 1
transform 1 0 3772 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_33
timestamp 1
transform 1 0 4140 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_42
timestamp 1
transform 1 0 4968 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_59
timestamp 1636968456
transform 1 0 6532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_71
timestamp 1636968456
transform 1 0 7636 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_95
timestamp 1636968456
transform 1 0 9844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_107
timestamp 1
transform 1 0 10948 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_151
timestamp 1
transform 1 0 14996 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_180
timestamp 1
transform 1 0 17664 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_197
timestamp 1
transform 1 0 19228 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_209
timestamp 1
transform 1 0 20332 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_238
timestamp 1
transform 1 0 23000 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_249
timestamp 1
transform 1 0 24012 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_253
timestamp 1
transform 1 0 24380 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_259
timestamp 1636968456
transform 1 0 24932 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_271
timestamp 1
transform 1 0 26036 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_292
timestamp 1
transform 1 0 27968 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_296
timestamp 1
transform 1 0 28336 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1636968456
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1636968456
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1636968456
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1636968456
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_69
timestamp 1
transform 1 0 7452 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_90
timestamp 1636968456
transform 1 0 9384 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_102
timestamp 1
transform 1 0 10488 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_108
timestamp 1
transform 1 0 11040 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_113
timestamp 1
transform 1 0 11500 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_139
timestamp 1636968456
transform 1 0 13892 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_151
timestamp 1
transform 1 0 14996 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_160
timestamp 1
transform 1 0 15824 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_165
timestamp 1
transform 1 0 16284 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_194
timestamp 1
transform 1 0 18952 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_249
timestamp 1
transform 1 0 24012 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_263
timestamp 1636968456
transform 1 0 25300 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_275
timestamp 1
transform 1 0 26404 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_281
timestamp 1
transform 1 0 26956 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1636968456
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1636968456
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1636968456
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1636968456
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_53
timestamp 1
transform 1 0 5980 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_61
timestamp 1
transform 1 0 6716 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_70
timestamp 1
transform 1 0 7544 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_91
timestamp 1636968456
transform 1 0 9476 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_103
timestamp 1
transform 1 0 10580 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_111
timestamp 1
transform 1 0 11316 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_120
timestamp 1
transform 1 0 12144 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_144
timestamp 1636968456
transform 1 0 14352 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_156
timestamp 1
transform 1 0 15456 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_161
timestamp 1
transform 1 0 15916 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_169
timestamp 1
transform 1 0 16652 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_178
timestamp 1
transform 1 0 17480 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_205
timestamp 1
transform 1 0 19964 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_215
timestamp 1
transform 1 0 20884 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_223
timestamp 1
transform 1 0 21620 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_232
timestamp 1
transform 1 0 22448 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_259
timestamp 1
transform 1 0 24932 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_280
timestamp 1
transform 1 0 26864 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1636968456
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1636968456
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_57
timestamp 1
transform 1 0 6348 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_63
timestamp 1
transform 1 0 6900 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_71
timestamp 1
transform 1 0 7636 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_93
timestamp 1
transform 1 0 9660 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_101
timestamp 1
transform 1 0 10396 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_109
timestamp 1
transform 1 0 11132 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_33_113
timestamp 1
transform 1 0 11500 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_119
timestamp 1
transform 1 0 12052 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_124
timestamp 1
transform 1 0 12512 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_145
timestamp 1
transform 1 0 14444 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_169
timestamp 1
transform 1 0 16652 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_173
timestamp 1
transform 1 0 17020 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_181
timestamp 1
transform 1 0 17756 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_205
timestamp 1636968456
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_235
timestamp 1
transform 1 0 22724 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_33_263
timestamp 1
transform 1 0 25300 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_271
timestamp 1
transform 1 0 26036 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1636968456
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1636968456
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1636968456
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_41
timestamp 1
transform 1 0 4876 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_49
timestamp 1
transform 1 0 5612 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_62
timestamp 1
transform 1 0 6808 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_74
timestamp 1
transform 1 0 7912 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_129
timestamp 1
transform 1 0 12972 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_137
timestamp 1
transform 1 0 13708 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_141
timestamp 1
transform 1 0 14076 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_163
timestamp 1636968456
transform 1 0 16100 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_175
timestamp 1
transform 1 0 17204 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_184
timestamp 1636968456
transform 1 0 18032 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_203
timestamp 1
transform 1 0 19780 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_264
timestamp 1636968456
transform 1 0 25392 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_296
timestamp 1
transform 1 0 28336 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1636968456
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1636968456
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_27
timestamp 1
transform 1 0 3588 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_33
timestamp 1
transform 1 0 4140 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_57
timestamp 1
transform 1 0 6348 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_91
timestamp 1
transform 1 0 9476 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_139
timestamp 1
transform 1 0 13892 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1636968456
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1636968456
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_193
timestamp 1
transform 1 0 18860 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_234
timestamp 1
transform 1 0 22632 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_255
timestamp 1
transform 1 0 24564 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_276
timestamp 1
transform 1 0 26496 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1636968456
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1636968456
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_29
timestamp 1
transform 1 0 3772 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_52
timestamp 1
transform 1 0 5888 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_92
timestamp 1636968456
transform 1 0 9568 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_104
timestamp 1
transform 1 0 10672 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_108
timestamp 1
transform 1 0 11040 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_115
timestamp 1
transform 1 0 11684 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_141
timestamp 1
transform 1 0 14076 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_170
timestamp 1
transform 1 0 16744 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_237
timestamp 1
transform 1 0 22908 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_253
timestamp 1
transform 1 0 24380 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_294
timestamp 1
transform 1 0 28152 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1636968456
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1636968456
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1636968456
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1636968456
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_57
timestamp 1
transform 1 0 6348 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_65
timestamp 1
transform 1 0 7084 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_71
timestamp 1
transform 1 0 7636 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_76
timestamp 1636968456
transform 1 0 8096 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_88
timestamp 1636968456
transform 1 0 9200 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_100
timestamp 1636968456
transform 1 0 10304 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_113
timestamp 1
transform 1 0 11500 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_121
timestamp 1
transform 1 0 12236 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_129
timestamp 1
transform 1 0 12972 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_166
timestamp 1
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_177
timestamp 1636968456
transform 1 0 17388 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_189
timestamp 1636968456
transform 1 0 18492 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_201
timestamp 1
transform 1 0 19596 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_211
timestamp 1636968456
transform 1 0 20516 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_233
timestamp 1
transform 1 0 22540 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_239
timestamp 1
transform 1 0 23092 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1636968456
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1636968456
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1636968456
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1636968456
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1636968456
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1636968456
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1636968456
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_97
timestamp 1
transform 1 0 10028 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_105
timestamp 1
transform 1 0 10764 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_112
timestamp 1636968456
transform 1 0 11408 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_124
timestamp 1636968456
transform 1 0 12512 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_136
timestamp 1
transform 1 0 13616 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_141
timestamp 1
transform 1 0 14076 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_149
timestamp 1
transform 1 0 14812 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_155
timestamp 1
transform 1 0 15364 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_167
timestamp 1
transform 1 0 16468 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_197
timestamp 1
transform 1 0 19228 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_208
timestamp 1636968456
transform 1 0 20240 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_220
timestamp 1
transform 1 0 21344 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_232
timestamp 1636968456
transform 1 0 22448 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_244
timestamp 1
transform 1 0 23552 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1636968456
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_265
timestamp 1
transform 1 0 25484 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_296
timestamp 1
transform 1 0 28336 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1636968456
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1636968456
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1636968456
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1636968456
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1636968456
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1636968456
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_81
timestamp 1
transform 1 0 8556 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_89
timestamp 1636968456
transform 1 0 9292 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_101
timestamp 1
transform 1 0 10396 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_113
timestamp 1
transform 1 0 11500 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_123
timestamp 1636968456
transform 1 0 12420 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_135
timestamp 1636968456
transform 1 0 13524 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_147
timestamp 1
transform 1 0 14628 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp 1
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_172
timestamp 1
transform 1 0 16928 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_178
timestamp 1
transform 1 0 17480 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_225
timestamp 1
transform 1 0 21804 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_39_231
timestamp 1
transform 1 0 22356 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_235
timestamp 1636968456
transform 1 0 22724 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_247
timestamp 1636968456
transform 1 0 23828 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_259
timestamp 1
transform 1 0 24932 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_39_268
timestamp 1
transform 1 0 25760 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_274
timestamp 1
transform 1 0 26312 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_281
timestamp 1
transform 1 0 26956 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1636968456
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1636968456
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1636968456
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1636968456
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_53
timestamp 1
transform 1 0 5980 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_61
timestamp 1
transform 1 0 6716 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_105
timestamp 1
transform 1 0 10764 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_132
timestamp 1
transform 1 0 13248 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_170
timestamp 1
transform 1 0 16744 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1636968456
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_272
timestamp 1
transform 1 0 26128 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_296
timestamp 1
transform 1 0 28336 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1636968456
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1636968456
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_27
timestamp 1
transform 1 0 3588 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_35
timestamp 1
transform 1 0 4324 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_57
timestamp 1
transform 1 0 6348 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_70
timestamp 1
transform 1 0 7544 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_41_93
timestamp 1
transform 1 0 9660 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_108
timestamp 1
transform 1 0 11040 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_140
timestamp 1
transform 1 0 13984 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_185
timestamp 1
transform 1 0 18124 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_189
timestamp 1
transform 1 0 18492 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_198
timestamp 1
transform 1 0 19320 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_241
timestamp 1636968456
transform 1 0 23276 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_253
timestamp 1
transform 1 0 24380 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_257
timestamp 1
transform 1 0 24748 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_278
timestamp 1
transform 1 0 26680 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_284
timestamp 1
transform 1 0 27232 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_291
timestamp 1
transform 1 0 27876 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1636968456
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1636968456
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1636968456
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_64
timestamp 1
transform 1 0 6992 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_130
timestamp 1
transform 1 0 13064 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_141
timestamp 1
transform 1 0 14076 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_173
timestamp 1636968456
transform 1 0 17020 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_185
timestamp 1
transform 1 0 18124 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_193
timestamp 1
transform 1 0 18860 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_217
timestamp 1
transform 1 0 21068 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_222
timestamp 1
transform 1 0 21528 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_244
timestamp 1
transform 1 0 23552 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_284
timestamp 1636968456
transform 1 0 27232 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_296
timestamp 1
transform 1 0 28336 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1636968456
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1636968456
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1636968456
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_39
timestamp 1
transform 1 0 4692 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_47
timestamp 1
transform 1 0 5428 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1636968456
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_69
timestamp 1
transform 1 0 7452 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_75
timestamp 1
transform 1 0 8004 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_80
timestamp 1
transform 1 0 8464 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_88
timestamp 1
transform 1 0 9200 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_95
timestamp 1636968456
transform 1 0 9844 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_107
timestamp 1
transform 1 0 10948 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_121
timestamp 1636968456
transform 1 0 12236 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_133
timestamp 1636968456
transform 1 0 13340 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_145
timestamp 1
transform 1 0 14444 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_153
timestamp 1
transform 1 0 15180 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_166
timestamp 1
transform 1 0 16376 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_177
timestamp 1636968456
transform 1 0 17388 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_189
timestamp 1636968456
transform 1 0 18492 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_201
timestamp 1
transform 1 0 19596 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_43_209
timestamp 1
transform 1 0 20332 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_220
timestamp 1
transform 1 0 21344 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_245
timestamp 1
transform 1 0 23644 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_269
timestamp 1
transform 1 0 25852 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_277
timestamp 1
transform 1 0 26588 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1636968456
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_293
timestamp 1
transform 1 0 28060 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1636968456
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1636968456
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1636968456
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1636968456
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1636968456
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1636968456
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1636968456
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1636968456
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1636968456
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1636968456
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1636968456
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1636968456
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1636968456
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1636968456
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1636968456
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1636968456
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1636968456
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_233
timestamp 1636968456
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1636968456
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1636968456
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1636968456
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_289
timestamp 1
transform 1 0 27692 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1636968456
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1636968456
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1636968456
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1636968456
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1636968456
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1636968456
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1636968456
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1636968456
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1636968456
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1636968456
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1636968456
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1636968456
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1636968456
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1636968456
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1636968456
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_205
timestamp 1636968456
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1636968456
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1636968456
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1636968456
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1636968456
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1636968456
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_293
timestamp 1
transform 1 0 28060 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1636968456
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1636968456
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1636968456
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1636968456
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1636968456
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1636968456
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1636968456
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1636968456
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1636968456
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1636968456
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1636968456
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1636968456
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_165
timestamp 1636968456
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_177
timestamp 1636968456
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1636968456
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1636968456
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1636968456
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_233
timestamp 1636968456
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1636968456
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1636968456
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_277
timestamp 1636968456
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_289
timestamp 1
transform 1 0 27692 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1636968456
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1636968456
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1636968456
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1636968456
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1636968456
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1636968456
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1636968456
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1636968456
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1636968456
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1636968456
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1636968456
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1636968456
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1636968456
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1636968456
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_193
timestamp 1636968456
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_205
timestamp 1636968456
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1636968456
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 1636968456
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_249
timestamp 1636968456
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_261
timestamp 1636968456
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1636968456
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_293
timestamp 1
transform 1 0 28060 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1636968456
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1636968456
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1636968456
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1636968456
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1636968456
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1636968456
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1636968456
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1636968456
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1636968456
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1636968456
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1636968456
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1636968456
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_165
timestamp 1636968456
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_177
timestamp 1636968456
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1636968456
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1636968456
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_221
timestamp 1636968456
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_233
timestamp 1636968456
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1636968456
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1636968456
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1636968456
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_289
timestamp 1
transform 1 0 27692 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1636968456
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1636968456
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_27
timestamp 1
transform 1 0 3588 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_29
timestamp 1636968456
transform 1 0 3772 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_41
timestamp 1636968456
transform 1 0 4876 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_53
timestamp 1
transform 1 0 5980 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1636968456
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1636968456
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_81
timestamp 1
transform 1 0 8556 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_85
timestamp 1636968456
transform 1 0 8924 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_97
timestamp 1636968456
transform 1 0 10028 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_109
timestamp 1
transform 1 0 11132 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1636968456
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1636968456
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_137
timestamp 1
transform 1 0 13708 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_141
timestamp 1636968456
transform 1 0 14076 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_153
timestamp 1636968456
transform 1 0 15180 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_165
timestamp 1
transform 1 0 16284 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1636968456
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1636968456
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_193
timestamp 1
transform 1 0 18860 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_197
timestamp 1636968456
transform 1 0 19228 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_209
timestamp 1636968456
transform 1 0 20332 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_221
timestamp 1
transform 1 0 21436 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1636968456
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1636968456
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_249
timestamp 1
transform 1 0 24012 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_253
timestamp 1636968456
transform 1 0 24380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_265
timestamp 1636968456
transform 1 0 25484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_277
timestamp 1
transform 1 0 26588 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1636968456
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_293
timestamp 1
transform 1 0 28060 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 1
transform -1 0 26496 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1
transform 1 0 25484 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1
transform -1 0 28428 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1
transform -1 0 28428 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1
transform 1 0 26128 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1
transform -1 0 27692 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1
transform 1 0 21988 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1
transform -1 0 22540 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1
transform 1 0 23552 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1
transform -1 0 23920 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1
transform -1 0 21620 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1
transform -1 0 20516 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1
transform -1 0 20976 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1
transform -1 0 19320 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1
transform 1 0 11408 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1
transform 1 0 16652 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1
transform -1 0 16376 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1
transform 1 0 19504 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1
transform -1 0 20792 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1
transform -1 0 20424 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1
transform -1 0 9660 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1
transform -1 0 8464 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1
transform -1 0 15916 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1
transform 1 0 14444 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1
transform 1 0 12788 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1
transform -1 0 17388 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1
transform 1 0 16652 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1
transform -1 0 24104 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1
transform -1 0 11500 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1
transform 1 0 23092 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1
transform -1 0 22080 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1
transform -1 0 24472 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1
transform -1 0 11316 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1
transform 1 0 22356 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1
transform -1 0 17388 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1
transform -1 0 17388 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1
transform 1 0 19688 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 1
transform -1 0 19688 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1
transform 1 0 11500 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 1
transform -1 0 19964 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 1
transform 1 0 14168 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1
transform 1 0 14812 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1
transform 1 0 22908 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 1
transform -1 0 23552 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 1
transform 1 0 16836 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 1
transform -1 0 12236 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1
transform -1 0 14168 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 1
transform -1 0 20608 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 1
transform 1 0 16652 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 1
transform -1 0 16376 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 1
transform -1 0 17388 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 1
transform 1 0 23644 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 1
transform -1 0 10764 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 1
transform 1 0 12788 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 1
transform 1 0 25116 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 1
transform 1 0 26220 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 1
transform -1 0 22540 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp 1
transform -1 0 21344 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp 1
transform -1 0 27784 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold60
timestamp 1
transform -1 0 23092 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp 1
transform -1 0 5888 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold62
timestamp 1
transform -1 0 11040 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold63
timestamp 1
transform -1 0 11592 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold64
timestamp 1
transform -1 0 23000 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold65
timestamp 1
transform -1 0 13984 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold66
timestamp 1
transform -1 0 18952 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold67
timestamp 1
transform -1 0 23460 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold68
timestamp 1
transform -1 0 7452 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold69
timestamp 1
transform -1 0 8832 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold70
timestamp 1
transform -1 0 5980 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold71
timestamp 1
transform -1 0 17664 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold72
timestamp 1
transform -1 0 14812 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold73
timestamp 1
transform -1 0 5796 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold74
timestamp 1
transform -1 0 20792 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold75
timestamp 1
transform -1 0 23828 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold76
timestamp 1
transform 1 0 16744 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold77
timestamp 1
transform 1 0 27692 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold78
timestamp 1
transform 1 0 6624 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold79
timestamp 1
transform -1 0 4968 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold80
timestamp 1
transform -1 0 15824 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold81
timestamp 1
transform -1 0 23276 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold82
timestamp 1
transform -1 0 19136 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold83
timestamp 1
transform 1 0 23276 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold84
timestamp 1
transform 1 0 17480 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1
transform 1 0 28152 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1
transform 1 0 28152 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1
transform 1 0 28152 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1
transform 1 0 28152 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1
transform 1 0 28152 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1
transform 1 0 28152 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1
transform 1 0 27600 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1
transform 1 0 28152 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1
transform 1 0 27876 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1
transform 1 0 27784 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1
transform -1 0 21620 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1
transform -1 0 22264 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1
transform -1 0 23552 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1
transform -1 0 22908 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1
transform -1 0 27784 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  max_cap18
timestamp 1
transform 1 0 6256 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 1
transform 1 0 28060 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_50
timestamp 1
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1
transform -1 0 28704 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_51
timestamp 1
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1
transform -1 0 28704 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_52
timestamp 1
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1
transform -1 0 28704 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_53
timestamp 1
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1
transform -1 0 28704 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_54
timestamp 1
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1
transform -1 0 28704 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_55
timestamp 1
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1
transform -1 0 28704 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_56
timestamp 1
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1
transform -1 0 28704 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_57
timestamp 1
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1
transform -1 0 28704 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_58
timestamp 1
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1
transform -1 0 28704 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_59
timestamp 1
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1
transform -1 0 28704 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_60
timestamp 1
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1
transform -1 0 28704 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_61
timestamp 1
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1
transform -1 0 28704 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_62
timestamp 1
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1
transform -1 0 28704 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_63
timestamp 1
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1
transform -1 0 28704 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_64
timestamp 1
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1
transform -1 0 28704 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_65
timestamp 1
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1
transform -1 0 28704 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_66
timestamp 1
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1
transform -1 0 28704 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_67
timestamp 1
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1
transform -1 0 28704 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_68
timestamp 1
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1
transform -1 0 28704 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_69
timestamp 1
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1
transform -1 0 28704 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_70
timestamp 1
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1
transform -1 0 28704 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_71
timestamp 1
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1
transform -1 0 28704 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_72
timestamp 1
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1
transform -1 0 28704 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_73
timestamp 1
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1
transform -1 0 28704 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_74
timestamp 1
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1
transform -1 0 28704 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_75
timestamp 1
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1
transform -1 0 28704 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_76
timestamp 1
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1
transform -1 0 28704 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_77
timestamp 1
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1
transform -1 0 28704 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_78
timestamp 1
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1
transform -1 0 28704 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_79
timestamp 1
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1
transform -1 0 28704 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_80
timestamp 1
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1
transform -1 0 28704 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_81
timestamp 1
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1
transform -1 0 28704 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_82
timestamp 1
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1
transform -1 0 28704 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_83
timestamp 1
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1
transform -1 0 28704 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_84
timestamp 1
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 1
transform -1 0 28704 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_85
timestamp 1
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 1
transform -1 0 28704 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_86
timestamp 1
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 1
transform -1 0 28704 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_87
timestamp 1
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 1
transform -1 0 28704 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_88
timestamp 1
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 1
transform -1 0 28704 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_89
timestamp 1
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 1
transform -1 0 28704 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_90
timestamp 1
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 1
transform -1 0 28704 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_91
timestamp 1
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp 1
transform -1 0 28704 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Left_92
timestamp 1
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Right_42
timestamp 1
transform -1 0 28704 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Left_93
timestamp 1
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Right_43
timestamp 1
transform -1 0 28704 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Left_94
timestamp 1
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Right_44
timestamp 1
transform -1 0 28704 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Left_95
timestamp 1
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Right_45
timestamp 1
transform -1 0 28704 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Left_96
timestamp 1
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Right_46
timestamp 1
transform -1 0 28704 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Left_97
timestamp 1
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Right_47
timestamp 1
transform -1 0 28704 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Left_98
timestamp 1
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Right_48
timestamp 1
transform -1 0 28704 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Left_99
timestamp 1
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Right_49
timestamp 1
transform -1 0 28704 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_100
timestamp 1
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_101
timestamp 1
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_102
timestamp 1
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_103
timestamp 1
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_104
timestamp 1
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_105
timestamp 1
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_106
timestamp 1
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_107
timestamp 1
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_108
timestamp 1
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_109
timestamp 1
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_110
timestamp 1
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_111
timestamp 1
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_112
timestamp 1
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_113
timestamp 1
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_114
timestamp 1
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_115
timestamp 1
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_116
timestamp 1
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_117
timestamp 1
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_118
timestamp 1
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_119
timestamp 1
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_120
timestamp 1
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_121
timestamp 1
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_122
timestamp 1
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_123
timestamp 1
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_124
timestamp 1
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_125
timestamp 1
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_126
timestamp 1
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_127
timestamp 1
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_128
timestamp 1
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_129
timestamp 1
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_130
timestamp 1
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_131
timestamp 1
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_132
timestamp 1
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_133
timestamp 1
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_134
timestamp 1
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_135
timestamp 1
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_136
timestamp 1
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_137
timestamp 1
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_138
timestamp 1
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_139
timestamp 1
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_140
timestamp 1
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_141
timestamp 1
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_142
timestamp 1
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_143
timestamp 1
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_144
timestamp 1
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_145
timestamp 1
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_146
timestamp 1
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_147
timestamp 1
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_148
timestamp 1
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_149
timestamp 1
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_150
timestamp 1
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_151
timestamp 1
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_152
timestamp 1
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_153
timestamp 1
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_154
timestamp 1
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_155
timestamp 1
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_156
timestamp 1
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_157
timestamp 1
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_158
timestamp 1
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_159
timestamp 1
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_160
timestamp 1
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_161
timestamp 1
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_162
timestamp 1
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_163
timestamp 1
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_164
timestamp 1
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_165
timestamp 1
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_166
timestamp 1
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_167
timestamp 1
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_168
timestamp 1
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_169
timestamp 1
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_170
timestamp 1
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_171
timestamp 1
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_172
timestamp 1
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_173
timestamp 1
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_174
timestamp 1
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_175
timestamp 1
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_176
timestamp 1
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_177
timestamp 1
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_178
timestamp 1
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_179
timestamp 1
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_180
timestamp 1
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_181
timestamp 1
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_182
timestamp 1
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_183
timestamp 1
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_184
timestamp 1
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_185
timestamp 1
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_186
timestamp 1
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_187
timestamp 1
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_188
timestamp 1
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_189
timestamp 1
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_190
timestamp 1
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_191
timestamp 1
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_192
timestamp 1
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_193
timestamp 1
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_194
timestamp 1
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_195
timestamp 1
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_196
timestamp 1
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_197
timestamp 1
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_198
timestamp 1
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_199
timestamp 1
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_200
timestamp 1
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_201
timestamp 1
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_202
timestamp 1
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_203
timestamp 1
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_204
timestamp 1
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_205
timestamp 1
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_206
timestamp 1
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_207
timestamp 1
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_208
timestamp 1
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_209
timestamp 1
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_210
timestamp 1
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_211
timestamp 1
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_212
timestamp 1
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_213
timestamp 1
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_214
timestamp 1
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_215
timestamp 1
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_216
timestamp 1
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_217
timestamp 1
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_218
timestamp 1
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_219
timestamp 1
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_220
timestamp 1
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_221
timestamp 1
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_222
timestamp 1
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_223
timestamp 1
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_224
timestamp 1
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_225
timestamp 1
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_226
timestamp 1
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_227
timestamp 1
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_228
timestamp 1
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_229
timestamp 1
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_230
timestamp 1
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_231
timestamp 1
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_232
timestamp 1
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_233
timestamp 1
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_234
timestamp 1
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_235
timestamp 1
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_236
timestamp 1
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_237
timestamp 1
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_238
timestamp 1
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_239
timestamp 1
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_240
timestamp 1
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_241
timestamp 1
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_242
timestamp 1
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_243
timestamp 1
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_244
timestamp 1
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_245
timestamp 1
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_246
timestamp 1
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_247
timestamp 1
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_248
timestamp 1
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_249
timestamp 1
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_250
timestamp 1
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_251
timestamp 1
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_252
timestamp 1
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_253
timestamp 1
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_254
timestamp 1
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_255
timestamp 1
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_256
timestamp 1
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_257
timestamp 1
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_258
timestamp 1
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_259
timestamp 1
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_260
timestamp 1
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_261
timestamp 1
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_262
timestamp 1
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_263
timestamp 1
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_264
timestamp 1
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_265
timestamp 1
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_266
timestamp 1
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_267
timestamp 1
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_268
timestamp 1
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_269
timestamp 1
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_270
timestamp 1
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_271
timestamp 1
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_272
timestamp 1
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_273
timestamp 1
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_274
timestamp 1
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_275
timestamp 1
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_276
timestamp 1
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_277
timestamp 1
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_278
timestamp 1
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_279
timestamp 1
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_280
timestamp 1
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_281
timestamp 1
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_282
timestamp 1
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_283
timestamp 1
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_284
timestamp 1
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_285
timestamp 1
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_286
timestamp 1
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_287
timestamp 1
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_288
timestamp 1
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_289
timestamp 1
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_290
timestamp 1
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_291
timestamp 1
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_292
timestamp 1
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_293
timestamp 1
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_294
timestamp 1
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_295
timestamp 1
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_296
timestamp 1
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_297
timestamp 1
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_298
timestamp 1
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_299
timestamp 1
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_300
timestamp 1
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_301
timestamp 1
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_302
timestamp 1
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_303
timestamp 1
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_304
timestamp 1
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_305
timestamp 1
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_306
timestamp 1
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_307
timestamp 1
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_308
timestamp 1
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_309
timestamp 1
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_310
timestamp 1
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_311
timestamp 1
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_312
timestamp 1
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_313
timestamp 1
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_314
timestamp 1
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_315
timestamp 1
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_316
timestamp 1
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_317
timestamp 1
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_318
timestamp 1
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_319
timestamp 1
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_320
timestamp 1
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_321
timestamp 1
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_322
timestamp 1
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_323
timestamp 1
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_324
timestamp 1
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_325
timestamp 1
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_326
timestamp 1
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_327
timestamp 1
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_328
timestamp 1
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_329
timestamp 1
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_330
timestamp 1
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_331
timestamp 1
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_332
timestamp 1
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_333
timestamp 1
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_334
timestamp 1
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_335
timestamp 1
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_336
timestamp 1
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_337
timestamp 1
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_338
timestamp 1
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_339
timestamp 1
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_340
timestamp 1
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_341
timestamp 1
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_342
timestamp 1
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_343
timestamp 1
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_344
timestamp 1
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_345
timestamp 1
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_346
timestamp 1
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_347
timestamp 1
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_348
timestamp 1
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_349
timestamp 1
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_350
timestamp 1
transform 1 0 3680 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_351
timestamp 1
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_352
timestamp 1
transform 1 0 8832 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_353
timestamp 1
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_354
timestamp 1
transform 1 0 13984 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_355
timestamp 1
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_356
timestamp 1
transform 1 0 19136 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_357
timestamp 1
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_358
timestamp 1
transform 1 0 24288 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_359
timestamp 1
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
<< labels >>
flabel metal4 s 4868 2128 5188 29424 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4208 2128 4528 29424 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 27208 800 27328 0 FreeSans 480 0 0 0 clk
port 2 nsew signal input
flabel metal3 s 29064 15648 29864 15768 0 FreeSans 480 0 0 0 keypad_i[0]
port 3 nsew signal input
flabel metal3 s 29064 7488 29864 7608 0 FreeSans 480 0 0 0 keypad_i[10]
port 4 nsew signal input
flabel metal3 s 29064 6808 29864 6928 0 FreeSans 480 0 0 0 keypad_i[11]
port 5 nsew signal input
flabel metal3 s 29064 5448 29864 5568 0 FreeSans 480 0 0 0 keypad_i[12]
port 6 nsew signal input
flabel metal3 s 29064 6128 29864 6248 0 FreeSans 480 0 0 0 keypad_i[13]
port 7 nsew signal input
flabel metal3 s 29064 11568 29864 11688 0 FreeSans 480 0 0 0 keypad_i[1]
port 8 nsew signal input
flabel metal3 s 29064 14968 29864 15088 0 FreeSans 480 0 0 0 keypad_i[2]
port 9 nsew signal input
flabel metal3 s 29064 12928 29864 13048 0 FreeSans 480 0 0 0 keypad_i[3]
port 10 nsew signal input
flabel metal3 s 29064 12248 29864 12368 0 FreeSans 480 0 0 0 keypad_i[4]
port 11 nsew signal input
flabel metal3 s 29064 13608 29864 13728 0 FreeSans 480 0 0 0 keypad_i[5]
port 12 nsew signal input
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 keypad_i[6]
port 13 nsew signal input
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 keypad_i[7]
port 14 nsew signal input
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 keypad_i[8]
port 15 nsew signal input
flabel metal2 s 22558 0 22614 800 0 FreeSans 224 90 0 0 keypad_i[9]
port 16 nsew signal input
flabel metal3 s 29064 3408 29864 3528 0 FreeSans 480 0 0 0 n_rst
port 17 nsew signal input
flabel metal3 s 29064 14288 29864 14408 0 FreeSans 480 0 0 0 pwm
port 18 nsew signal output
rlabel metal1 14904 29376 14904 29376 0 VGND
rlabel metal1 14904 28832 14904 28832 0 VPWR
rlabel metal2 11822 21726 11822 21726 0 _0000_
rlabel metal1 13524 19346 13524 19346 0 _0001_
rlabel metal2 12466 21522 12466 21522 0 _0002_
rlabel metal1 15456 20366 15456 20366 0 _0003_
rlabel metal1 15594 18394 15594 18394 0 _0004_
rlabel metal2 17434 17442 17434 17442 0 _0005_
rlabel metal2 19458 17374 19458 17374 0 _0006_
rlabel metal2 20838 18530 20838 18530 0 _0007_
rlabel metal2 21758 17884 21758 17884 0 _0008_
rlabel metal1 22172 16150 22172 16150 0 _0009_
rlabel metal1 22310 15130 22310 15130 0 _0010_
rlabel metal2 18262 15844 18262 15844 0 _0011_
rlabel metal1 20562 14926 20562 14926 0 _0012_
rlabel metal2 21850 13090 21850 13090 0 _0013_
rlabel metal1 22954 12682 22954 12682 0 _0014_
rlabel metal1 24150 10778 24150 10778 0 _0015_
rlabel metal1 23368 11662 23368 11662 0 _0016_
rlabel metal1 20838 12614 20838 12614 0 _0017_
rlabel metal1 19918 12274 19918 12274 0 _0018_
rlabel metal2 17618 13532 17618 13532 0 _0019_
rlabel metal1 15364 13838 15364 13838 0 _0020_
rlabel metal1 15502 15674 15502 15674 0 _0021_
rlabel metal2 14766 16796 14766 16796 0 _0022_
rlabel metal1 13800 15674 13800 15674 0 _0023_
rlabel metal2 12466 16082 12466 16082 0 _0024_
rlabel metal2 9246 11628 9246 11628 0 _0025_
rlabel metal1 9614 10098 9614 10098 0 _0026_
rlabel metal2 14122 18394 14122 18394 0 _0027_
rlabel metal1 19228 24378 19228 24378 0 _0028_
rlabel metal2 20194 24004 20194 24004 0 _0029_
rlabel metal1 20240 21658 20240 21658 0 _0030_
rlabel metal1 22126 21658 22126 21658 0 _0031_
rlabel metal1 23644 22542 23644 22542 0 _0032_
rlabel metal1 25668 21658 25668 21658 0 _0033_
rlabel metal1 27324 20570 27324 20570 0 _0034_
rlabel metal1 28060 20026 28060 20026 0 _0035_
rlabel metal2 14858 21148 14858 21148 0 _0036_
rlabel metal1 15548 22066 15548 22066 0 _0037_
rlabel metal1 15594 24718 15594 24718 0 _0038_
rlabel metal2 14398 24956 14398 24956 0 _0039_
rlabel metal1 16238 25772 16238 25772 0 _0040_
rlabel metal2 9338 8670 9338 8670 0 _0041_
rlabel metal1 9338 6970 9338 6970 0 _0042_
rlabel metal1 12236 6426 12236 6426 0 _0043_
rlabel metal2 12282 3298 12282 3298 0 _0044_
rlabel metal2 10902 3740 10902 3740 0 _0045_
rlabel metal1 8648 3094 8648 3094 0 _0046_
rlabel metal1 6863 3706 6863 3706 0 _0047_
rlabel metal1 4186 4794 4186 4794 0 _0048_
rlabel metal1 4324 7310 4324 7310 0 _0049_
rlabel metal1 4140 8398 4140 8398 0 _0050_
rlabel metal1 4002 11322 4002 11322 0 _0051_
rlabel metal2 4738 14110 4738 14110 0 _0052_
rlabel metal1 5520 13226 5520 13226 0 _0053_
rlabel metal1 8832 13974 8832 13974 0 _0054_
rlabel metal1 9108 17306 9108 17306 0 _0055_
rlabel metal2 7590 18802 7590 18802 0 _0056_
rlabel metal1 5980 16150 5980 16150 0 _0057_
rlabel metal1 2990 17714 2990 17714 0 _0058_
rlabel metal1 3220 18190 3220 18190 0 _0059_
rlabel metal1 4692 20366 4692 20366 0 _0060_
rlabel metal1 5244 21658 5244 21658 0 _0061_
rlabel metal1 6532 21114 6532 21114 0 _0062_
rlabel metal1 8050 20026 8050 20026 0 _0063_
rlabel metal1 10120 20570 10120 20570 0 _0064_
rlabel metal1 22678 4658 22678 4658 0 _0065_
rlabel metal1 22402 5746 22402 5746 0 _0066_
rlabel metal1 22908 6222 22908 6222 0 _0067_
rlabel metal1 23874 5270 23874 5270 0 _0068_
rlabel metal1 17526 4794 17526 4794 0 _0069_
rlabel metal2 15318 5372 15318 5372 0 _0070_
rlabel metal1 13570 19856 13570 19856 0 _0071_
rlabel metal1 10856 18258 10856 18258 0 _0072_
rlabel metal1 7958 21454 7958 21454 0 _0073_
rlabel metal1 27370 22474 27370 22474 0 _0074_
rlabel metal1 26542 22576 26542 22576 0 _0075_
rlabel metal1 25346 23494 25346 23494 0 _0076_
rlabel metal1 24932 24786 24932 24786 0 _0077_
rlabel metal2 22126 22882 22126 22882 0 _0078_
rlabel metal1 21597 23698 21597 23698 0 _0079_
rlabel metal1 21620 24242 21620 24242 0 _0080_
rlabel metal1 24104 23834 24104 23834 0 _0081_
rlabel metal2 26358 9724 26358 9724 0 _0082_
rlabel metal1 25070 8874 25070 8874 0 _0083_
rlabel metal1 24472 8874 24472 8874 0 _0084_
rlabel metal1 26036 5882 26036 5882 0 _0085_
rlabel metal1 25392 17646 25392 17646 0 _0086_
rlabel metal2 25806 16864 25806 16864 0 _0087_
rlabel metal2 15870 23698 15870 23698 0 _0088_
rlabel metal1 15410 20910 15410 20910 0 _0089_
rlabel metal2 9890 24174 9890 24174 0 _0090_
rlabel via1 13010 24106 13010 24106 0 _0091_
rlabel metal1 12558 18836 12558 18836 0 _0092_
rlabel metal1 17066 5644 17066 5644 0 _0093_
rlabel via2 18538 4811 18538 4811 0 _0094_
rlabel metal1 17020 3502 17020 3502 0 _0095_
rlabel via2 15778 6069 15778 6069 0 _0096_
rlabel metal2 16790 3604 16790 3604 0 _0097_
rlabel metal2 14766 6052 14766 6052 0 _0098_
rlabel metal1 15410 3536 15410 3536 0 _0099_
rlabel metal1 12558 12784 12558 12784 0 _0100_
rlabel metal2 13478 24276 13478 24276 0 _0101_
rlabel metal1 11638 18938 11638 18938 0 _0102_
rlabel viali 12558 19827 12558 19827 0 _0103_
rlabel metal1 14398 18870 14398 18870 0 _0104_
rlabel metal2 10258 17340 10258 17340 0 _0105_
rlabel metal1 9706 17612 9706 17612 0 _0106_
rlabel metal1 16054 4046 16054 4046 0 _0107_
rlabel metal1 16192 5678 16192 5678 0 _0108_
rlabel metal1 12742 12920 12742 12920 0 _0109_
rlabel metal2 9798 15232 9798 15232 0 _0110_
rlabel metal1 9437 16558 9437 16558 0 _0111_
rlabel metal1 9522 16048 9522 16048 0 _0112_
rlabel metal1 6762 17204 6762 17204 0 _0113_
rlabel metal1 9016 16422 9016 16422 0 _0114_
rlabel metal1 7636 14994 7636 14994 0 _0115_
rlabel metal1 9430 14790 9430 14790 0 _0116_
rlabel metal2 6946 16694 6946 16694 0 _0117_
rlabel metal1 15962 4182 15962 4182 0 _0118_
rlabel metal2 19550 3808 19550 3808 0 _0119_
rlabel metal1 18400 5202 18400 5202 0 _0120_
rlabel metal2 19274 4114 19274 4114 0 _0121_
rlabel metal1 19596 4522 19596 4522 0 _0122_
rlabel metal2 12926 4301 12926 4301 0 _0123_
rlabel metal1 18906 4012 18906 4012 0 _0124_
rlabel metal1 18998 6970 18998 6970 0 _0125_
rlabel metal1 13478 4012 13478 4012 0 _0126_
rlabel metal2 12834 3774 12834 3774 0 _0127_
rlabel metal2 13478 3740 13478 3740 0 _0128_
rlabel metal1 17066 5066 17066 5066 0 _0129_
rlabel metal2 13018 6256 13018 6256 0 _0130_
rlabel metal2 13018 4828 13018 4828 0 _0131_
rlabel metal2 17250 5559 17250 5559 0 _0132_
rlabel metal1 16422 5542 16422 5542 0 _0133_
rlabel metal2 11546 6834 11546 6834 0 _0134_
rlabel metal1 18446 6290 18446 6290 0 _0135_
rlabel metal1 18170 6256 18170 6256 0 _0136_
rlabel metal1 12144 7854 12144 7854 0 _0137_
rlabel metal1 9154 7990 9154 7990 0 _0138_
rlabel metal2 9338 7684 9338 7684 0 _0139_
rlabel metal2 10534 7344 10534 7344 0 _0140_
rlabel metal2 12558 7004 12558 7004 0 _0141_
rlabel metal1 11960 6154 11960 6154 0 _0142_
rlabel via2 13386 4539 13386 4539 0 _0143_
rlabel metal1 8970 4454 8970 4454 0 _0144_
rlabel metal1 17434 4114 17434 4114 0 _0145_
rlabel metal1 7866 4556 7866 4556 0 _0146_
rlabel metal1 8142 5066 8142 5066 0 _0147_
rlabel metal1 8510 4148 8510 4148 0 _0148_
rlabel metal1 9614 5066 9614 5066 0 _0149_
rlabel metal2 16146 5151 16146 5151 0 _0150_
rlabel metal1 6670 5746 6670 5746 0 _0151_
rlabel metal2 6670 5440 6670 5440 0 _0152_
rlabel metal1 7038 5168 7038 5168 0 _0153_
rlabel metal1 16238 3706 16238 3706 0 _0154_
rlabel metal1 15778 3502 15778 3502 0 _0155_
rlabel metal1 15686 3638 15686 3638 0 _0156_
rlabel metal1 6256 4794 6256 4794 0 _0157_
rlabel metal2 7038 3774 7038 3774 0 _0158_
rlabel metal1 8004 4998 8004 4998 0 _0159_
rlabel metal1 7912 4726 7912 4726 0 _0160_
rlabel metal1 6670 5236 6670 5236 0 _0161_
rlabel metal1 7682 5134 7682 5134 0 _0162_
rlabel metal1 7038 7888 7038 7888 0 _0163_
rlabel metal2 16422 5542 16422 5542 0 _0164_
rlabel metal1 14306 11152 14306 11152 0 _0165_
rlabel metal1 6762 11220 6762 11220 0 _0166_
rlabel metal1 7038 11730 7038 11730 0 _0167_
rlabel metal1 6026 11050 6026 11050 0 _0168_
rlabel metal1 15364 7922 15364 7922 0 _0169_
rlabel metal2 6302 10608 6302 10608 0 _0170_
rlabel metal1 5750 10030 5750 10030 0 _0171_
rlabel metal1 6256 10642 6256 10642 0 _0172_
rlabel metal2 7222 10268 7222 10268 0 _0173_
rlabel metal1 17480 4250 17480 4250 0 _0174_
rlabel metal1 16790 4250 16790 4250 0 _0175_
rlabel metal1 8418 8942 8418 8942 0 _0176_
rlabel metal2 7314 9724 7314 9724 0 _0177_
rlabel metal1 6578 8874 6578 8874 0 _0178_
rlabel metal2 6394 8330 6394 8330 0 _0179_
rlabel metal1 15686 5100 15686 5100 0 _0180_
rlabel metal2 15594 6902 15594 6902 0 _0181_
rlabel metal1 7084 8874 7084 8874 0 _0182_
rlabel metal1 7452 7854 7452 7854 0 _0183_
rlabel metal1 7176 8058 7176 8058 0 _0184_
rlabel metal1 7728 9690 7728 9690 0 _0185_
rlabel metal1 7038 9588 7038 9588 0 _0186_
rlabel metal1 6808 10098 6808 10098 0 _0187_
rlabel metal2 6946 10285 6946 10285 0 _0188_
rlabel metal1 7452 9962 7452 9962 0 _0189_
rlabel metal1 7038 14960 7038 14960 0 _0190_
rlabel metal1 6164 17102 6164 17102 0 _0191_
rlabel metal2 6670 17850 6670 17850 0 _0192_
rlabel metal1 7038 17850 7038 17850 0 _0193_
rlabel metal2 12742 21386 12742 21386 0 _0194_
rlabel metal1 12650 20876 12650 20876 0 _0195_
rlabel metal1 16330 21998 16330 21998 0 _0196_
rlabel metal1 20148 21454 20148 21454 0 _0197_
rlabel metal2 21022 23868 21022 23868 0 _0198_
rlabel metal2 21666 23290 21666 23290 0 _0199_
rlabel metal2 23966 22780 23966 22780 0 _0200_
rlabel metal1 24656 22610 24656 22610 0 _0201_
rlabel metal1 26036 22474 26036 22474 0 _0202_
rlabel metal2 28198 20910 28198 20910 0 _0203_
rlabel metal1 27324 22678 27324 22678 0 _0204_
rlabel metal1 27646 9350 27646 9350 0 _0205_
rlabel metal2 25898 9180 25898 9180 0 _0206_
rlabel metal1 26956 9486 26956 9486 0 _0207_
rlabel via1 26358 7922 26358 7922 0 _0208_
rlabel metal1 25898 7786 25898 7786 0 _0209_
rlabel metal2 25530 6392 25530 6392 0 _0210_
rlabel metal1 26634 7344 26634 7344 0 _0211_
rlabel metal1 25530 3434 25530 3434 0 _0212_
rlabel metal1 26634 5134 26634 5134 0 _0213_
rlabel metal1 25392 6290 25392 6290 0 _0214_
rlabel metal1 17802 6834 17802 6834 0 _0215_
rlabel metal2 19274 7582 19274 7582 0 _0216_
rlabel metal1 19458 7276 19458 7276 0 _0217_
rlabel metal1 18446 7242 18446 7242 0 _0218_
rlabel metal1 18262 6970 18262 6970 0 _0219_
rlabel metal1 17802 7412 17802 7412 0 _0220_
rlabel metal1 17756 7514 17756 7514 0 _0221_
rlabel metal2 17342 8058 17342 8058 0 _0222_
rlabel metal1 16514 7854 16514 7854 0 _0223_
rlabel metal1 16514 8058 16514 8058 0 _0224_
rlabel metal2 14950 8058 14950 8058 0 _0225_
rlabel metal2 16146 8058 16146 8058 0 _0226_
rlabel metal2 15962 8534 15962 8534 0 _0227_
rlabel metal1 15042 7820 15042 7820 0 _0228_
rlabel metal1 14904 8602 14904 8602 0 _0229_
rlabel metal1 14812 8058 14812 8058 0 _0230_
rlabel metal2 14674 9894 14674 9894 0 _0231_
rlabel metal1 13892 10574 13892 10574 0 _0232_
rlabel metal1 12650 12614 12650 12614 0 _0233_
rlabel metal2 13202 11934 13202 11934 0 _0234_
rlabel metal2 13018 11900 13018 11900 0 _0235_
rlabel metal1 13524 10574 13524 10574 0 _0236_
rlabel metal1 13018 10710 13018 10710 0 _0237_
rlabel metal1 12972 11186 12972 11186 0 _0238_
rlabel metal1 13432 12818 13432 12818 0 _0239_
rlabel metal2 18998 14178 18998 14178 0 _0240_
rlabel metal1 19780 8058 19780 8058 0 _0241_
rlabel metal2 20378 9758 20378 9758 0 _0242_
rlabel metal1 20010 9146 20010 9146 0 _0243_
rlabel metal1 20792 9146 20792 9146 0 _0244_
rlabel metal1 20838 8534 20838 8534 0 _0245_
rlabel metal2 16882 9520 16882 9520 0 _0246_
rlabel metal1 20056 9350 20056 9350 0 _0247_
rlabel metal2 16698 9962 16698 9962 0 _0248_
rlabel metal1 18400 9418 18400 9418 0 _0249_
rlabel metal1 18078 9622 18078 9622 0 _0250_
rlabel metal2 14306 11118 14306 11118 0 _0251_
rlabel metal2 15686 10336 15686 10336 0 _0252_
rlabel metal1 14076 10234 14076 10234 0 _0253_
rlabel metal1 14536 9554 14536 9554 0 _0254_
rlabel metal1 12926 9622 12926 9622 0 _0255_
rlabel metal1 13478 13702 13478 13702 0 _0256_
rlabel metal1 14030 12342 14030 12342 0 _0257_
rlabel metal1 12466 14008 12466 14008 0 _0258_
rlabel metal1 12926 13906 12926 13906 0 _0259_
rlabel metal1 12098 14042 12098 14042 0 _0260_
rlabel metal2 12834 14110 12834 14110 0 _0261_
rlabel metal2 13110 10880 13110 10880 0 _0262_
rlabel metal1 9154 25398 9154 25398 0 _0263_
rlabel metal2 8602 25670 8602 25670 0 _0264_
rlabel metal1 9522 23698 9522 23698 0 _0265_
rlabel metal1 11178 23834 11178 23834 0 _0266_
rlabel metal2 13662 24922 13662 24922 0 _0267_
rlabel metal2 11178 23290 11178 23290 0 _0268_
rlabel metal1 22540 24922 22540 24922 0 _0269_
rlabel metal2 23782 25126 23782 25126 0 _0270_
rlabel via1 26174 24021 26174 24021 0 _0271_
rlabel metal1 27462 23698 27462 23698 0 _0272_
rlabel metal2 21298 24820 21298 24820 0 _0273_
rlabel metal2 23046 24956 23046 24956 0 _0274_
rlabel metal2 26358 24956 26358 24956 0 _0275_
rlabel metal1 26726 24378 26726 24378 0 _0276_
rlabel metal1 26082 16014 26082 16014 0 _0277_
rlabel via1 17983 19822 17983 19822 0 _0278_
rlabel metal1 19642 19754 19642 19754 0 _0279_
rlabel metal1 24978 16558 24978 16558 0 _0280_
rlabel metal2 25070 16864 25070 16864 0 _0281_
rlabel viali 21850 19346 21850 19346 0 _0282_
rlabel via1 18280 19822 18280 19822 0 _0283_
rlabel metal1 17894 19210 17894 19210 0 _0284_
rlabel metal1 18906 18870 18906 18870 0 _0285_
rlabel via1 21942 19346 21942 19346 0 _0286_
rlabel viali 23414 19346 23414 19346 0 _0287_
rlabel metal2 24058 18938 24058 18938 0 _0288_
rlabel metal1 24794 17782 24794 17782 0 _0289_
rlabel metal1 25024 17850 25024 17850 0 _0290_
rlabel metal2 27186 9078 27186 9078 0 _0291_
rlabel metal1 24840 3706 24840 3706 0 _0292_
rlabel metal1 26956 12614 26956 12614 0 _0293_
rlabel metal2 27370 12852 27370 12852 0 _0294_
rlabel metal1 14490 19176 14490 19176 0 _0295_
rlabel metal2 12650 18428 12650 18428 0 _0296_
rlabel metal1 13478 18598 13478 18598 0 _0297_
rlabel via1 17350 18326 17350 18326 0 _0298_
rlabel metal1 14076 16558 14076 16558 0 _0299_
rlabel metal1 15916 17850 15916 17850 0 _0300_
rlabel metal1 17572 17170 17572 17170 0 _0301_
rlabel metal2 19274 17340 19274 17340 0 _0302_
rlabel metal1 20884 18258 20884 18258 0 _0303_
rlabel metal1 22724 17850 22724 17850 0 _0304_
rlabel metal1 22494 16558 22494 16558 0 _0305_
rlabel metal1 22448 14994 22448 14994 0 _0306_
rlabel metal2 20654 15878 20654 15878 0 _0307_
rlabel metal2 22034 13260 22034 13260 0 _0308_
rlabel metal1 22862 12410 22862 12410 0 _0309_
rlabel metal1 24150 10574 24150 10574 0 _0310_
rlabel metal2 22402 11526 22402 11526 0 _0311_
rlabel metal1 20976 12818 20976 12818 0 _0312_
rlabel metal1 18998 11866 18998 11866 0 _0313_
rlabel metal1 17756 12954 17756 12954 0 _0314_
rlabel metal1 16100 12954 16100 12954 0 _0315_
rlabel metal2 15962 14484 15962 14484 0 _0316_
rlabel metal2 15870 16388 15870 16388 0 _0317_
rlabel metal2 13478 15674 13478 15674 0 _0318_
rlabel metal2 12558 15674 12558 15674 0 _0319_
rlabel metal1 10258 12240 10258 12240 0 _0320_
rlabel metal1 10856 10642 10856 10642 0 _0321_
rlabel metal1 15364 23222 15364 23222 0 _0322_
rlabel metal1 16284 24786 16284 24786 0 _0323_
rlabel metal2 16790 24310 16790 24310 0 _0324_
rlabel metal1 17158 24650 17158 24650 0 _0325_
rlabel metal1 17756 24650 17756 24650 0 _0326_
rlabel metal1 10304 8942 10304 8942 0 _0327_
rlabel metal1 10350 8058 10350 8058 0 _0328_
rlabel metal2 10718 6970 10718 6970 0 _0329_
rlabel metal1 10074 6630 10074 6630 0 _0330_
rlabel metal1 9934 6766 9934 6766 0 _0331_
rlabel metal2 12466 7004 12466 7004 0 _0332_
rlabel metal2 12742 6868 12742 6868 0 _0333_
rlabel metal2 13938 4454 13938 4454 0 _0334_
rlabel metal2 13018 4318 13018 4318 0 _0335_
rlabel metal1 13386 4114 13386 4114 0 _0336_
rlabel metal2 12926 3536 12926 3536 0 _0337_
rlabel metal1 11914 4080 11914 4080 0 _0338_
rlabel metal1 11178 4046 11178 4046 0 _0339_
rlabel metal1 9706 4522 9706 4522 0 _0340_
rlabel metal1 9936 4794 9936 4794 0 _0341_
rlabel metal1 9246 4794 9246 4794 0 _0342_
rlabel metal1 9200 4250 9200 4250 0 _0343_
rlabel metal1 8234 4590 8234 4590 0 _0344_
rlabel metal1 6946 4726 6946 4726 0 _0345_
rlabel metal1 6762 3944 6762 3944 0 _0346_
rlabel metal1 7268 3502 7268 3502 0 _0347_
rlabel metal2 7682 3706 7682 3706 0 _0348_
rlabel metal1 6026 4794 6026 4794 0 _0349_
rlabel metal1 6670 4794 6670 4794 0 _0350_
rlabel metal1 4922 4556 4922 4556 0 _0351_
rlabel metal2 5014 4828 5014 4828 0 _0352_
rlabel metal1 7130 7412 7130 7412 0 _0353_
rlabel metal2 6670 7548 6670 7548 0 _0354_
rlabel metal1 5980 7514 5980 7514 0 _0355_
rlabel metal1 6854 7514 6854 7514 0 _0356_
rlabel metal1 4830 7888 4830 7888 0 _0357_
rlabel metal1 5290 8058 5290 8058 0 _0358_
rlabel metal1 5106 10540 5106 10540 0 _0359_
rlabel metal1 5612 10574 5612 10574 0 _0360_
rlabel metal1 5152 10778 5152 10778 0 _0361_
rlabel metal1 7038 14314 7038 14314 0 _0362_
rlabel metal2 5750 11356 5750 11356 0 _0363_
rlabel metal1 5428 11322 5428 11322 0 _0364_
rlabel metal1 5888 14382 5888 14382 0 _0365_
rlabel metal1 9890 15436 9890 15436 0 _0366_
rlabel metal1 6762 13906 6762 13906 0 _0367_
rlabel metal2 6394 14144 6394 14144 0 _0368_
rlabel metal1 9614 14858 9614 14858 0 _0369_
rlabel metal1 9246 14416 9246 14416 0 _0370_
rlabel metal1 9154 14314 9154 14314 0 _0371_
rlabel metal2 8234 14450 8234 14450 0 _0372_
rlabel metal1 9522 16150 9522 16150 0 _0373_
rlabel metal2 9154 15878 9154 15878 0 _0374_
rlabel metal1 9430 16218 9430 16218 0 _0375_
rlabel metal2 8418 18020 8418 18020 0 _0376_
rlabel metal1 9062 17850 9062 17850 0 _0377_
rlabel metal1 8142 18326 8142 18326 0 _0378_
rlabel metal2 6486 16796 6486 16796 0 _0379_
rlabel metal1 5980 16558 5980 16558 0 _0380_
rlabel metal2 6026 18292 6026 18292 0 _0381_
rlabel metal1 5244 17170 5244 17170 0 _0382_
rlabel metal2 5290 17442 5290 17442 0 _0383_
rlabel metal1 4002 17714 4002 17714 0 _0384_
rlabel metal1 6118 18870 6118 18870 0 _0385_
rlabel metal1 5014 18292 5014 18292 0 _0386_
rlabel metal1 4186 18292 4186 18292 0 _0387_
rlabel metal1 4508 17850 4508 17850 0 _0388_
rlabel metal1 5106 19414 5106 19414 0 _0389_
rlabel metal1 5198 19380 5198 19380 0 _0390_
rlabel metal1 5474 19278 5474 19278 0 _0391_
rlabel metal2 5382 21148 5382 21148 0 _0392_
rlabel metal1 5382 21114 5382 21114 0 _0393_
rlabel metal1 5934 21624 5934 21624 0 _0394_
rlabel metal1 6026 21556 6026 21556 0 _0395_
rlabel metal2 6210 21114 6210 21114 0 _0396_
rlabel metal1 7590 20026 7590 20026 0 _0397_
rlabel metal1 9108 19822 9108 19822 0 _0398_
rlabel metal1 8510 19856 8510 19856 0 _0399_
rlabel metal1 9062 21862 9062 21862 0 _0400_
rlabel metal2 9798 20604 9798 20604 0 _0401_
rlabel metal1 26358 7854 26358 7854 0 _0402_
rlabel metal2 26266 3978 26266 3978 0 _0403_
rlabel metal1 24242 7412 24242 7412 0 _0404_
rlabel metal1 24288 8602 24288 8602 0 _0405_
rlabel via2 24610 7939 24610 7939 0 _0406_
rlabel metal2 23874 7004 23874 7004 0 _0407_
rlabel metal1 25898 5134 25898 5134 0 _0408_
rlabel metal1 26036 4250 26036 4250 0 _0409_
rlabel metal1 25760 4794 25760 4794 0 _0410_
rlabel metal1 24932 5066 24932 5066 0 _0411_
rlabel metal2 25346 8772 25346 8772 0 _0412_
rlabel metal2 26450 5270 26450 5270 0 _0413_
rlabel via1 26082 7514 26082 7514 0 _0414_
rlabel metal1 25806 8432 25806 8432 0 _0415_
rlabel metal1 27094 9554 27094 9554 0 _0416_
rlabel metal2 25714 8942 25714 8942 0 _0417_
rlabel metal1 24886 5202 24886 5202 0 _0418_
rlabel metal1 24380 6154 24380 6154 0 _0419_
rlabel metal1 26864 8942 26864 8942 0 _0420_
rlabel metal1 23920 5814 23920 5814 0 _0421_
rlabel metal2 25438 4862 25438 4862 0 _0422_
rlabel metal1 24610 5610 24610 5610 0 _0423_
rlabel metal1 26404 3706 26404 3706 0 _0424_
rlabel metal1 25852 5338 25852 5338 0 _0425_
rlabel metal2 24058 7650 24058 7650 0 _0426_
rlabel metal2 24426 7820 24426 7820 0 _0427_
rlabel metal1 24610 5746 24610 5746 0 _0428_
rlabel metal3 575 26996 575 26996 0 clk
rlabel metal1 16514 14246 16514 14246 0 clknet_0_clk
rlabel metal1 6578 3468 6578 3468 0 clknet_4_0_0_clk
rlabel metal2 28290 4080 28290 4080 0 clknet_4_10_0_clk
rlabel metal2 26542 13702 26542 13702 0 clknet_4_11_0_clk
rlabel metal2 20470 19074 20470 19074 0 clknet_4_12_0_clk
rlabel metal1 20194 22066 20194 22066 0 clknet_4_13_0_clk
rlabel metal2 21850 15776 21850 15776 0 clknet_4_14_0_clk
rlabel metal1 23828 25806 23828 25806 0 clknet_4_15_0_clk
rlabel metal1 5244 13362 5244 13362 0 clknet_4_1_0_clk
rlabel via1 12006 3587 12006 3587 0 clknet_4_2_0_clk
rlabel metal1 13754 14926 13754 14926 0 clknet_4_3_0_clk
rlabel metal1 2162 18122 2162 18122 0 clknet_4_4_0_clk
rlabel metal1 9154 21930 9154 21930 0 clknet_4_5_0_clk
rlabel metal1 13616 16626 13616 16626 0 clknet_4_6_0_clk
rlabel metal1 13708 22066 13708 22066 0 clknet_4_7_0_clk
rlabel metal2 21298 3264 21298 3264 0 clknet_4_8_0_clk
rlabel metal1 18584 13362 18584 13362 0 clknet_4_9_0_clk
rlabel metal1 19366 13906 19366 13906 0 count\[0\]
rlabel metal1 14950 13226 14950 13226 0 count\[10\]
rlabel metal1 15502 12954 15502 12954 0 count\[11\]
rlabel metal1 13432 14246 13432 14246 0 count\[12\]
rlabel metal2 13018 15606 13018 15606 0 count\[13\]
rlabel metal1 12466 11084 12466 11084 0 count\[14\]
rlabel metal2 12282 10812 12282 10812 0 count\[15\]
rlabel metal1 19136 13702 19136 13702 0 count\[1\]
rlabel via1 20386 8534 20386 8534 0 count\[2\]
rlabel metal1 21298 9962 21298 9962 0 count\[3\]
rlabel metal1 18722 7854 18722 7854 0 count\[4\]
rlabel metal1 17618 8432 17618 8432 0 count\[5\]
rlabel metal2 17066 10846 17066 10846 0 count\[6\]
rlabel metal2 18538 10081 18538 10081 0 count\[7\]
rlabel metal1 16882 12750 16882 12750 0 count\[8\]
rlabel metal1 15180 12750 15180 12750 0 count\[9\]
rlabel metal2 21022 3876 21022 3876 0 freq_div.keycode\[0\]
rlabel metal1 23782 5882 23782 5882 0 freq_div.keycode\[1\]
rlabel metal2 23598 6562 23598 6562 0 freq_div.keycode\[2\]
rlabel metal2 20470 5474 20470 5474 0 freq_div.keycode\[3\]
rlabel metal1 27646 13158 27646 13158 0 keypad.keypad_reg\[0\]
rlabel metal1 26542 4590 26542 4590 0 keypad.keypad_reg\[10\]
rlabel metal1 26772 4046 26772 4046 0 keypad.keypad_reg\[11\]
rlabel metal2 26266 5882 26266 5882 0 keypad.keypad_reg\[12\]
rlabel metal2 26542 5372 26542 5372 0 keypad.keypad_reg\[13\]
rlabel metal1 27922 9894 27922 9894 0 keypad.keypad_reg\[1\]
rlabel metal2 28198 10812 28198 10812 0 keypad.keypad_reg\[2\]
rlabel metal1 28014 9554 28014 9554 0 keypad.keypad_reg\[3\]
rlabel metal2 25070 10234 25070 10234 0 keypad.keypad_reg\[4\]
rlabel metal1 24472 8942 24472 8942 0 keypad.keypad_reg\[5\]
rlabel metal1 24058 7854 24058 7854 0 keypad.keypad_reg\[6\]
rlabel metal1 23920 8466 23920 8466 0 keypad.keypad_reg\[7\]
rlabel metal1 26772 4114 26772 4114 0 keypad.keypad_reg\[8\]
rlabel metal1 25806 3978 25806 3978 0 keypad.keypad_reg\[9\]
rlabel metal1 25346 16082 25346 16082 0 keypad.modekey
rlabel metal1 24649 13702 24649 13702 0 keypad.n_modekey
rlabel metal2 28382 15895 28382 15895 0 keypad_i[0]
rlabel metal2 28382 7701 28382 7701 0 keypad_i[10]
rlabel metal2 28382 7123 28382 7123 0 keypad_i[11]
rlabel metal2 28382 5355 28382 5355 0 keypad_i[12]
rlabel metal2 28382 6239 28382 6239 0 keypad_i[13]
rlabel metal2 28382 11679 28382 11679 0 keypad_i[1]
rlabel metal2 27830 15249 27830 15249 0 keypad_i[2]
rlabel metal2 28382 12903 28382 12903 0 keypad_i[3]
rlabel metal3 28620 12308 28620 12308 0 keypad_i[4]
rlabel metal2 28014 13787 28014 13787 0 keypad_i[5]
rlabel metal2 21298 1588 21298 1588 0 keypad_i[6]
rlabel metal2 21942 1588 21942 1588 0 keypad_i[7]
rlabel metal2 23230 1588 23230 1588 0 keypad_i[8]
rlabel metal2 22586 1588 22586 1588 0 keypad_i[9]
rlabel metal1 27738 16558 27738 16558 0 mode\[1\]
rlabel metal2 27554 3247 27554 3247 0 n_rst
rlabel metal1 27554 13770 27554 13770 0 net1
rlabel metal1 27462 12750 27462 12750 0 net10
rlabel metal1 16422 14926 16422 14926 0 net100
rlabel metal1 16146 17102 16146 17102 0 net101
rlabel metal1 20424 12750 20424 12750 0 net102
rlabel metal1 18814 12274 18814 12274 0 net103
rlabel metal2 11822 15708 11822 15708 0 net104
rlabel metal1 18860 14382 18860 14382 0 net105
rlabel metal2 14398 21148 14398 21148 0 net106
rlabel metal2 15502 21284 15502 21284 0 net107
rlabel metal1 24242 4794 24242 4794 0 net108
rlabel metal1 21643 8534 21643 8534 0 net109
rlabel metal2 21574 3502 21574 3502 0 net11
rlabel metal1 17618 9622 17618 9622 0 net110
rlabel metal1 10442 24718 10442 24718 0 net111
rlabel metal1 12926 9520 12926 9520 0 net112
rlabel metal1 19320 13974 19320 13974 0 net113
rlabel metal2 16882 24140 16882 24140 0 net114
rlabel metal1 15502 22746 15502 22746 0 net115
rlabel metal2 16698 22202 16698 22202 0 net116
rlabel metal1 24610 5338 24610 5338 0 net117
rlabel metal1 9246 17204 9246 17204 0 net118
rlabel metal1 14122 19788 14122 19788 0 net119
rlabel metal1 22770 2958 22770 2958 0 net12
rlabel metal1 26082 24786 26082 24786 0 net120
rlabel metal1 26956 25262 26956 25262 0 net121
rlabel metal2 21758 24378 21758 24378 0 net122
rlabel metal1 20378 25874 20378 25874 0 net123
rlabel metal2 25898 24004 25898 24004 0 net124
rlabel metal1 22356 25262 22356 25262 0 net125
rlabel metal1 4968 11118 4968 11118 0 net126
rlabel metal2 10350 25364 10350 25364 0 net127
rlabel metal1 10856 8942 10856 8942 0 net128
rlabel metal1 21620 18394 21620 18394 0 net129
rlabel metal1 23736 2618 23736 2618 0 net13
rlabel metal1 13156 25262 13156 25262 0 net130
rlabel metal1 18032 17238 18032 17238 0 net131
rlabel metal1 22540 18326 22540 18326 0 net132
rlabel metal1 5566 14484 5566 14484 0 net133
rlabel metal2 8234 20298 8234 20298 0 net134
rlabel metal2 5474 7616 5474 7616 0 net135
rlabel metal1 16560 18394 16560 18394 0 net136
rlabel metal1 13478 3094 13478 3094 0 net137
rlabel metal2 5290 8704 5290 8704 0 net138
rlabel metal1 19596 17238 19596 17238 0 net139
rlabel metal1 23092 3502 23092 3502 0 net14
rlabel metal1 22862 16422 22862 16422 0 net140
rlabel metal2 17434 20400 17434 20400 0 net141
rlabel metal1 28244 22406 28244 22406 0 net142
rlabel metal1 7866 3502 7866 3502 0 net143
rlabel metal2 4554 18428 4554 18428 0 net144
rlabel metal2 14582 18938 14582 18938 0 net145
rlabel metal1 22402 19414 22402 19414 0 net146
rlabel metal1 18538 18938 18538 18938 0 net147
rlabel metal1 23828 18938 23828 18938 0 net148
rlabel metal1 18124 19482 18124 19482 0 net149
rlabel metal2 27738 3638 27738 3638 0 net15
rlabel metal1 28106 13872 28106 13872 0 net16
rlabel metal2 18170 14110 18170 14110 0 net17
rlabel metal2 6118 19142 6118 19142 0 net18
rlabel metal2 20010 14756 20010 14756 0 net19
rlabel metal1 27790 6970 27790 6970 0 net2
rlabel metal2 18170 18428 18170 18428 0 net20
rlabel metal1 17066 18258 17066 18258 0 net21
rlabel metal1 19734 12682 19734 12682 0 net22
rlabel metal2 19090 17510 19090 17510 0 net23
rlabel metal1 13156 6086 13156 6086 0 net24
rlabel metal1 14674 18938 14674 18938 0 net25
rlabel metal2 8602 14433 8602 14433 0 net26
rlabel metal1 11914 18224 11914 18224 0 net27
rlabel metal1 13064 18734 13064 18734 0 net28
rlabel metal1 18078 12886 18078 12886 0 net29
rlabel metal1 27370 6222 27370 6222 0 net3
rlabel metal1 17020 6358 17020 6358 0 net30
rlabel metal2 20286 4284 20286 4284 0 net31
rlabel metal1 15318 5338 15318 5338 0 net32
rlabel metal2 19826 5950 19826 5950 0 net33
rlabel metal2 20010 3740 20010 3740 0 net34
rlabel metal2 20194 4828 20194 4828 0 net35
rlabel metal2 16974 5440 16974 5440 0 net36
rlabel metal1 5888 5202 5888 5202 0 net37
rlabel metal1 12144 20910 12144 20910 0 net38
rlabel metal1 12558 6664 12558 6664 0 net39
rlabel metal1 27922 5338 27922 5338 0 net4
rlabel metal1 11592 12614 11592 12614 0 net40
rlabel via1 8865 16082 8865 16082 0 net41
rlabel metal1 12742 18632 12742 18632 0 net42
rlabel metal2 11638 19516 11638 19516 0 net43
rlabel metal1 20516 15402 20516 15402 0 net44
rlabel metal2 16054 19652 16054 19652 0 net45
rlabel metal2 13386 3332 13386 3332 0 net46
rlabel metal1 13202 3026 13202 3026 0 net47
rlabel via1 8970 19142 8970 19142 0 net48
rlabel metal2 12926 21726 12926 21726 0 net49
rlabel metal1 27876 6222 27876 6222 0 net5
rlabel metal2 15502 22168 15502 22168 0 net50
rlabel metal1 13018 15674 13018 15674 0 net51
rlabel metal2 22310 8704 22310 8704 0 net52
rlabel metal1 23145 13226 23145 13226 0 net53
rlabel metal1 26273 12886 26273 12886 0 net54
rlabel metal1 21443 7446 21443 7446 0 net55
rlabel metal2 20654 20672 20654 20672 0 net56
rlabel metal1 20983 17578 20983 17578 0 net57
rlabel metal1 26687 19754 26687 19754 0 net58
rlabel metal1 23828 25942 23828 25942 0 net59
rlabel metal1 27324 13974 27324 13974 0 net6
rlabel metal1 25491 25194 25491 25194 0 net60
rlabel metal1 20838 15368 20838 15368 0 net61
rlabel metal1 12558 15368 12558 15368 0 net62
rlabel metal1 5520 25194 5520 25194 0 net63
rlabel metal2 4738 25058 4738 25058 0 net64
rlabel metal2 8326 11118 8326 11118 0 net65
rlabel metal1 25576 21522 25576 21522 0 net66
rlabel metal1 26091 22202 26091 22202 0 net67
rlabel metal2 27738 19584 27738 19584 0 net68
rlabel metal2 26818 21182 26818 21182 0 net69
rlabel metal2 27186 13974 27186 13974 0 net7
rlabel metal1 27094 20434 27094 20434 0 net70
rlabel metal1 26811 22202 26811 22202 0 net71
rlabel metal1 22448 20570 22448 20570 0 net72
rlabel metal1 21613 22202 21613 22202 0 net73
rlabel metal1 23966 21114 23966 21114 0 net74
rlabel metal1 23138 22406 23138 22406 0 net75
rlabel metal1 20700 21522 20700 21522 0 net76
rlabel via1 19543 22202 19543 22202 0 net77
rlabel metal1 19964 23766 19964 23766 0 net78
rlabel metal2 17894 24174 17894 24174 0 net79
rlabel metal1 27416 12818 27416 12818 0 net8
rlabel metal1 12558 20944 12558 20944 0 net80
rlabel metal1 16376 25942 16376 25942 0 net81
rlabel metal2 15502 25500 15502 25500 0 net82
rlabel metal1 20010 23290 20010 23290 0 net83
rlabel metal1 19504 24106 19504 24106 0 net84
rlabel metal1 19320 15538 19320 15538 0 net85
rlabel metal2 8970 25636 8970 25636 0 net86
rlabel metal2 7222 24616 7222 24616 0 net87
rlabel metal1 14720 23834 14720 23834 0 net88
rlabel metal2 14582 24616 14582 24616 0 net89
rlabel metal1 27462 12920 27462 12920 0 net9
rlabel metal2 13202 15980 13202 15980 0 net90
rlabel metal1 16560 15538 16560 15538 0 net91
rlabel metal1 17388 13838 17388 13838 0 net92
rlabel metal1 22310 12852 22310 12852 0 net93
rlabel metal2 10810 11764 10810 11764 0 net94
rlabel metal1 23828 10574 23828 10574 0 net95
rlabel metal2 21390 15844 21390 15844 0 net96
rlabel metal1 23690 12750 23690 12750 0 net97
rlabel metal1 10534 10574 10534 10574 0 net98
rlabel metal1 22678 12614 22678 12614 0 net99
rlabel metal2 18262 14756 18262 14756 0 oscill.n_count\[0\]
rlabel metal2 12374 9180 12374 9180 0 oscill.n_count\[10\]
rlabel metal1 14030 12410 14030 12410 0 oscill.n_count\[11\]
rlabel metal1 11684 14314 11684 14314 0 oscill.n_count\[12\]
rlabel metal1 13432 14518 13432 14518 0 oscill.n_count\[13\]
rlabel metal1 12880 11322 12880 11322 0 oscill.n_count\[14\]
rlabel metal1 19274 14450 19274 14450 0 oscill.n_count\[1\]
rlabel metal1 19872 7446 19872 7446 0 oscill.n_count\[2\]
rlabel metal2 21114 8449 21114 8449 0 oscill.n_count\[3\]
rlabel via1 21117 8602 21117 8602 0 oscill.n_count\[4\]
rlabel metal2 20102 10132 20102 10132 0 oscill.n_count\[5\]
rlabel metal1 18584 10234 18584 10234 0 oscill.n_count\[6\]
rlabel metal2 17894 9690 17894 9690 0 oscill.n_count\[7\]
rlabel metal1 15640 10778 15640 10778 0 oscill.n_count\[8\]
rlabel metal1 12742 8568 12742 8568 0 oscill.n_count\[9\]
rlabel metal2 28290 14195 28290 14195 0 pwm
rlabel metal1 27370 13906 27370 13906 0 pwm1
rlabel metal1 19964 24038 19964 24038 0 pwm_counter.active_sample\[0\]
rlabel metal1 19596 23698 19596 23698 0 pwm_counter.active_sample\[1\]
rlabel metal2 21022 21760 21022 21760 0 pwm_counter.active_sample\[2\]
rlabel metal2 22862 22338 22862 22338 0 pwm_counter.active_sample\[3\]
rlabel via1 24610 22678 24610 22678 0 pwm_counter.active_sample\[4\]
rlabel metal1 25254 21420 25254 21420 0 pwm_counter.active_sample\[5\]
rlabel metal1 27324 21590 27324 21590 0 pwm_counter.active_sample\[6\]
rlabel metal1 27278 22610 27278 22610 0 pwm_counter.active_sample\[7\]
rlabel viali 22778 24854 22778 24854 0 pwm_counter.count\[0\]
rlabel metal1 21114 25466 21114 25466 0 pwm_counter.count\[1\]
rlabel metal1 22586 24786 22586 24786 0 pwm_counter.count\[2\]
rlabel metal2 22954 25466 22954 25466 0 pwm_counter.count\[3\]
rlabel metal1 25944 24582 25944 24582 0 pwm_counter.count\[4\]
rlabel metal2 25162 24956 25162 24956 0 pwm_counter.count\[5\]
rlabel metal1 25806 24140 25806 24140 0 pwm_counter.count\[6\]
rlabel metal1 27830 23630 27830 23630 0 pwm_counter.count\[7\]
rlabel metal1 24702 24174 24702 24174 0 pwm_counter.n_count\[0\]
rlabel metal2 19550 25500 19550 25500 0 pwm_counter.n_count\[1\]
rlabel metal1 20792 24718 20792 24718 0 pwm_counter.n_count\[2\]
rlabel metal1 23230 24922 23230 24922 0 pwm_counter.n_count\[3\]
rlabel metal1 24242 25466 24242 25466 0 pwm_counter.n_count\[4\]
rlabel metal1 26496 25194 26496 25194 0 pwm_counter.n_count\[5\]
rlabel metal2 26818 24412 26818 24412 0 pwm_counter.n_count\[6\]
rlabel metal1 26864 23154 26864 23154 0 pwm_counter.n_count\[7\]
rlabel metal1 27416 14450 27416 14450 0 pwm_counter.n_pwm
rlabel metal1 19918 23222 19918 23222 0 pwm_counter.sample\[0\]
rlabel metal1 19228 21862 19228 21862 0 pwm_counter.sample\[1\]
rlabel metal1 20700 20570 20700 20570 0 pwm_counter.sample\[2\]
rlabel metal1 21850 20434 21850 20434 0 pwm_counter.sample\[3\]
rlabel metal1 23552 20978 23552 20978 0 pwm_counter.sample\[4\]
rlabel metal1 25806 20570 25806 20570 0 pwm_counter.sample\[5\]
rlabel metal1 26772 20026 26772 20026 0 pwm_counter.sample\[6\]
rlabel metal2 27922 19108 27922 19108 0 pwm_counter.sample\[7\]
rlabel metal1 8280 25262 8280 25262 0 sample_rate.count\[0\]
rlabel metal2 8786 24820 8786 24820 0 sample_rate.count\[1\]
rlabel metal1 10672 24786 10672 24786 0 sample_rate.count\[2\]
rlabel metal1 11454 23630 11454 23630 0 sample_rate.count\[3\]
rlabel metal1 13708 24582 13708 24582 0 sample_rate.count\[4\]
rlabel metal1 12190 24038 12190 24038 0 sample_rate.count\[5\]
rlabel metal1 7130 24752 7130 24752 0 sample_rate.count\[6\]
rlabel metal1 7130 24854 7130 24854 0 sample_rate.count\[7\]
rlabel metal1 9430 24718 9430 24718 0 sample_rate.n_count\[0\]
rlabel metal2 8418 25500 8418 25500 0 sample_rate.n_count\[1\]
rlabel metal2 9246 23970 9246 23970 0 sample_rate.n_count\[2\]
rlabel metal1 10626 24922 10626 24922 0 sample_rate.n_count\[3\]
rlabel metal2 12558 24922 12558 24922 0 sample_rate.n_count\[4\]
rlabel metal1 11316 23290 11316 23290 0 sample_rate.n_count\[5\]
rlabel metal1 25668 15946 25668 15946 0 state_machine.fsmState\[0\]
rlabel metal1 27278 16422 27278 16422 0 state_machine.fsmState\[1\]
rlabel metal2 24702 15912 24702 15912 0 state_machine.nextState\[0\]
rlabel metal1 25438 16218 25438 16218 0 state_machine.nextState\[1\]
rlabel metal1 27002 16762 27002 16762 0 state_machine.nextState\[2\]
rlabel metal1 16652 19890 16652 19890 0 waveshape.scaled_count\[0\]
rlabel metal1 17342 19278 17342 19278 0 waveshape.scaled_count\[1\]
rlabel metal1 18538 18802 18538 18802 0 waveshape.scaled_count\[2\]
rlabel metal1 20010 19890 20010 19890 0 waveshape.scaled_count\[3\]
rlabel metal1 23184 18802 23184 18802 0 waveshape.scaled_count\[4\]
rlabel metal1 22816 17510 22816 17510 0 waveshape.scaled_count\[5\]
rlabel metal2 23966 18700 23966 18700 0 waveshape.scaled_count\[6\]
rlabel metal2 17066 19856 17066 19856 0 waveshape.scaled_count\[7\]
rlabel metal1 22770 13158 22770 13158 0 waveshape.seq_div.dividend\[10\]
rlabel metal1 24288 12750 24288 12750 0 waveshape.seq_div.dividend\[11\]
rlabel metal1 22816 10982 22816 10982 0 waveshape.seq_div.dividend\[12\]
rlabel metal2 21574 11356 21574 11356 0 waveshape.seq_div.dividend\[13\]
rlabel metal1 19458 11866 19458 11866 0 waveshape.seq_div.dividend\[14\]
rlabel metal1 18607 12818 18607 12818 0 waveshape.seq_div.dividend\[15\]
rlabel metal1 16376 13498 16376 13498 0 waveshape.seq_div.dividend\[16\]
rlabel metal2 16514 14518 16514 14518 0 waveshape.seq_div.dividend\[17\]
rlabel metal1 16882 16014 16882 16014 0 waveshape.seq_div.dividend\[18\]
rlabel metal1 16146 16422 16146 16422 0 waveshape.seq_div.dividend\[19\]
rlabel metal2 12834 16762 12834 16762 0 waveshape.seq_div.dividend\[20\]
rlabel metal1 11500 16014 11500 16014 0 waveshape.seq_div.dividend\[21\]
rlabel metal1 11040 11186 11040 11186 0 waveshape.seq_div.dividend\[22\]
rlabel metal1 10350 9894 10350 9894 0 waveshape.seq_div.dividend\[23\]
rlabel metal1 10902 8602 10902 8602 0 waveshape.seq_div.dividend\[24\]
rlabel metal1 11500 7378 11500 7378 0 waveshape.seq_div.dividend\[25\]
rlabel metal1 12834 5202 12834 5202 0 waveshape.seq_div.dividend\[26\]
rlabel via2 13754 3723 13754 3723 0 waveshape.seq_div.dividend\[27\]
rlabel metal1 11086 4114 11086 4114 0 waveshape.seq_div.dividend\[28\]
rlabel metal1 9154 4080 9154 4080 0 waveshape.seq_div.dividend\[29\]
rlabel metal2 5842 3876 5842 3876 0 waveshape.seq_div.dividend\[30\]
rlabel metal2 6486 6494 6486 6494 0 waveshape.seq_div.dividend\[31\]
rlabel metal1 5474 7854 5474 7854 0 waveshape.seq_div.dividend\[32\]
rlabel metal2 5658 8738 5658 8738 0 waveshape.seq_div.dividend\[33\]
rlabel metal2 5842 11424 5842 11424 0 waveshape.seq_div.dividend\[34\]
rlabel metal1 6210 14008 6210 14008 0 waveshape.seq_div.dividend\[35\]
rlabel metal1 7452 13906 7452 13906 0 waveshape.seq_div.dividend\[36\]
rlabel metal2 10074 15266 10074 15266 0 waveshape.seq_div.dividend\[37\]
rlabel metal1 9752 18054 9752 18054 0 waveshape.seq_div.dividend\[38\]
rlabel metal2 8418 16252 8418 16252 0 waveshape.seq_div.dividend\[39\]
rlabel metal1 5014 16626 5014 16626 0 waveshape.seq_div.dividend\[40\]
rlabel metal1 4278 17612 4278 17612 0 waveshape.seq_div.dividend\[41\]
rlabel metal2 4830 18564 4830 18564 0 waveshape.seq_div.dividend\[42\]
rlabel metal2 5658 18700 5658 18700 0 waveshape.seq_div.dividend\[43\]
rlabel metal1 6854 21352 6854 21352 0 waveshape.seq_div.dividend\[44\]
rlabel metal1 8786 19788 8786 19788 0 waveshape.seq_div.dividend\[45\]
rlabel metal2 7314 20128 7314 20128 0 waveshape.seq_div.dividend\[46\]
rlabel metal2 12926 21114 12926 21114 0 waveshape.seq_div.dividend\[47\]
rlabel metal1 19964 16014 19964 16014 0 waveshape.seq_div.dividend\[8\]
rlabel metal1 21804 15130 21804 15130 0 waveshape.seq_div.dividend\[9\]
rlabel metal1 15640 21658 15640 21658 0 waveshape.seq_div.n\[0\]
rlabel metal1 16008 21930 16008 21930 0 waveshape.seq_div.n\[1\]
rlabel metal1 16468 24650 16468 24650 0 waveshape.seq_div.n\[2\]
rlabel metal1 17848 24786 17848 24786 0 waveshape.seq_div.n\[3\]
rlabel metal2 16974 24752 16974 24752 0 waveshape.seq_div.n\[4\]
rlabel metal1 13340 18734 13340 18734 0 waveshape.seq_div.state\[0\]
rlabel metal1 14536 21862 14536 21862 0 waveshape.seq_div.state\[1\]
rlabel metal1 11408 20978 11408 20978 0 waveshape.seq_div.state\[2\]
rlabel metal2 16238 19788 16238 19788 0 waveshape.seq_div.state\[3\]
rlabel metal1 13202 21386 13202 21386 0 waveshape.seq_div.state\[4\]
rlabel metal2 17526 22066 17526 22066 0 waveshape.shaper.n_sample\[0\]
rlabel metal1 17710 20026 17710 20026 0 waveshape.shaper.n_sample\[1\]
rlabel metal2 18906 19924 18906 19924 0 waveshape.shaper.n_sample\[2\]
rlabel metal1 20056 20026 20056 20026 0 waveshape.shaper.n_sample\[3\]
rlabel metal1 22402 19482 22402 19482 0 waveshape.shaper.n_sample\[4\]
rlabel metal1 23874 19482 23874 19482 0 waveshape.shaper.n_sample\[5\]
rlabel metal1 24794 19754 24794 19754 0 waveshape.shaper.n_sample\[6\]
rlabel metal2 25806 18530 25806 18530 0 waveshape.shaper.n_sample\[7\]
<< properties >>
string FIXED_BBOX 0 0 29864 32008
<< end >>
