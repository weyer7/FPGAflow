VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fpga
  CLASS BLOCK ;
  FOREIGN fpga ;
  ORIGIN -15.000 -15.000 ;
  SIZE 435.000 BY 429.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 198.630 440.000 198.910 444.000 ;
    END
  END clk
  PIN config_data_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 15.000 225.840 19.000 226.440 ;
    END
  END config_data_in
  PIN config_data_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 236.040 450.000 236.640 ;
    END
  END config_data_out
  PIN config_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.860700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 182.530 440.000 182.810 444.000 ;
    END
  END config_en
  PIN io_east_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 151.040 450.000 151.640 ;
    END
  END io_east_in[0]
  PIN io_east_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 205.440 450.000 206.040 ;
    END
  END io_east_in[10]
  PIN io_east_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 212.240 450.000 212.840 ;
    END
  END io_east_in[11]
  PIN io_east_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 215.640 450.000 216.240 ;
    END
  END io_east_in[12]
  PIN io_east_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 219.040 450.000 219.640 ;
    END
  END io_east_in[13]
  PIN io_east_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.090 15.000 15.370 19.000 ;
    END
  END io_east_in[14]
  PIN io_east_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.310 15.000 18.590 19.000 ;
    END
  END io_east_in[15]
  PIN io_east_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 334.640 450.000 335.240 ;
    END
  END io_east_in[16]
  PIN io_east_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 338.040 450.000 338.640 ;
    END
  END io_east_in[17]
  PIN io_east_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 344.840 450.000 345.440 ;
    END
  END io_east_in[18]
  PIN io_east_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 351.640 450.000 352.240 ;
    END
  END io_east_in[19]
  PIN io_east_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 157.840 450.000 158.440 ;
    END
  END io_east_in[1]
  PIN io_east_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 355.040 450.000 355.640 ;
    END
  END io_east_in[20]
  PIN io_east_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 361.840 450.000 362.440 ;
    END
  END io_east_in[21]
  PIN io_east_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 365.240 450.000 365.840 ;
    END
  END io_east_in[22]
  PIN io_east_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 372.040 450.000 372.640 ;
    END
  END io_east_in[23]
  PIN io_east_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 378.840 450.000 379.440 ;
    END
  END io_east_in[24]
  PIN io_east_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 382.240 450.000 382.840 ;
    END
  END io_east_in[25]
  PIN io_east_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 389.040 450.000 389.640 ;
    END
  END io_east_in[26]
  PIN io_east_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 392.440 450.000 393.040 ;
    END
  END io_east_in[27]
  PIN io_east_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 399.240 450.000 399.840 ;
    END
  END io_east_in[28]
  PIN io_east_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 406.040 450.000 406.640 ;
    END
  END io_east_in[29]
  PIN io_east_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 161.240 450.000 161.840 ;
    END
  END io_east_in[2]
  PIN io_east_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.530 15.000 21.810 19.000 ;
    END
  END io_east_in[30]
  PIN io_east_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.750 15.000 25.030 19.000 ;
    END
  END io_east_in[31]
  PIN io_east_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 168.040 450.000 168.640 ;
    END
  END io_east_in[3]
  PIN io_east_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 174.840 450.000 175.440 ;
    END
  END io_east_in[4]
  PIN io_east_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 178.240 450.000 178.840 ;
    END
  END io_east_in[5]
  PIN io_east_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 185.040 450.000 185.640 ;
    END
  END io_east_in[6]
  PIN io_east_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 188.440 450.000 189.040 ;
    END
  END io_east_in[7]
  PIN io_east_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 195.240 450.000 195.840 ;
    END
  END io_east_in[8]
  PIN io_east_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 202.040 450.000 202.640 ;
    END
  END io_east_in[9]
  PIN io_east_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 76.240 450.000 76.840 ;
    END
  END io_east_out[0]
  PIN io_east_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 130.640 450.000 131.240 ;
    END
  END io_east_out[10]
  PIN io_east_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 134.040 450.000 134.640 ;
    END
  END io_east_out[11]
  PIN io_east_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 140.840 450.000 141.440 ;
    END
  END io_east_out[12]
  PIN io_east_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 147.640 450.000 148.240 ;
    END
  END io_east_out[13]
  PIN io_east_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.830 440.000 231.110 444.000 ;
    END
  END io_east_out[14]
  PIN io_east_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.150 440.000 250.430 444.000 ;
    END
  END io_east_out[15]
  PIN io_east_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 256.440 450.000 257.040 ;
    END
  END io_east_out[16]
  PIN io_east_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 263.240 450.000 263.840 ;
    END
  END io_east_out[17]
  PIN io_east_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 270.040 450.000 270.640 ;
    END
  END io_east_out[18]
  PIN io_east_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 273.440 450.000 274.040 ;
    END
  END io_east_out[19]
  PIN io_east_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 79.640 450.000 80.240 ;
    END
  END io_east_out[1]
  PIN io_east_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 280.240 450.000 280.840 ;
    END
  END io_east_out[20]
  PIN io_east_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 283.640 450.000 284.240 ;
    END
  END io_east_out[21]
  PIN io_east_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 290.440 450.000 291.040 ;
    END
  END io_east_out[22]
  PIN io_east_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 297.240 450.000 297.840 ;
    END
  END io_east_out[23]
  PIN io_east_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 300.640 450.000 301.240 ;
    END
  END io_east_out[24]
  PIN io_east_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 307.440 450.000 308.040 ;
    END
  END io_east_out[25]
  PIN io_east_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 310.840 450.000 311.440 ;
    END
  END io_east_out[26]
  PIN io_east_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 317.640 450.000 318.240 ;
    END
  END io_east_out[27]
  PIN io_east_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 324.440 450.000 325.040 ;
    END
  END io_east_out[28]
  PIN io_east_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 327.840 450.000 328.440 ;
    END
  END io_east_out[29]
  PIN io_east_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 86.440 450.000 87.040 ;
    END
  END io_east_out[2]
  PIN io_east_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.270 440.000 237.550 444.000 ;
    END
  END io_east_out[30]
  PIN io_east_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.290 440.000 208.570 444.000 ;
    END
  END io_east_out[31]
  PIN io_east_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 93.240 450.000 93.840 ;
    END
  END io_east_out[3]
  PIN io_east_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 96.640 450.000 97.240 ;
    END
  END io_east_out[4]
  PIN io_east_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 103.440 450.000 104.040 ;
    END
  END io_east_out[5]
  PIN io_east_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 106.840 450.000 107.440 ;
    END
  END io_east_out[6]
  PIN io_east_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 113.640 450.000 114.240 ;
    END
  END io_east_out[7]
  PIN io_east_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 120.440 450.000 121.040 ;
    END
  END io_east_out[8]
  PIN io_east_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 123.840 450.000 124.440 ;
    END
  END io_east_out[9]
  PIN io_north_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 76.270 440.000 76.550 444.000 ;
    END
  END io_north_in[0]
  PIN io_north_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 131.010 440.000 131.290 444.000 ;
    END
  END io_north_in[10]
  PIN io_north_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 134.230 440.000 134.510 444.000 ;
    END
  END io_north_in[11]
  PIN io_north_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 140.670 440.000 140.950 444.000 ;
    END
  END io_north_in[12]
  PIN io_north_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 147.110 440.000 147.390 444.000 ;
    END
  END io_north_in[13]
  PIN io_north_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.970 15.000 28.250 19.000 ;
    END
  END io_north_in[14]
  PIN io_north_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.190 15.000 31.470 19.000 ;
    END
  END io_north_in[15]
  PIN io_north_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 263.030 440.000 263.310 444.000 ;
    END
  END io_north_in[16]
  PIN io_north_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 266.250 440.000 266.530 444.000 ;
    END
  END io_north_in[17]
  PIN io_north_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 272.690 440.000 272.970 444.000 ;
    END
  END io_north_in[18]
  PIN io_north_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 279.130 440.000 279.410 444.000 ;
    END
  END io_north_in[19]
  PIN io_north_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 79.490 440.000 79.770 444.000 ;
    END
  END io_north_in[1]
  PIN io_north_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 285.570 440.000 285.850 444.000 ;
    END
  END io_north_in[20]
  PIN io_north_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 288.790 440.000 289.070 444.000 ;
    END
  END io_north_in[21]
  PIN io_north_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 295.230 440.000 295.510 444.000 ;
    END
  END io_north_in[22]
  PIN io_north_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 301.670 440.000 301.950 444.000 ;
    END
  END io_north_in[23]
  PIN io_north_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 304.890 440.000 305.170 444.000 ;
    END
  END io_north_in[24]
  PIN io_north_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 311.330 440.000 311.610 444.000 ;
    END
  END io_north_in[25]
  PIN io_north_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 317.770 440.000 318.050 444.000 ;
    END
  END io_north_in[26]
  PIN io_north_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 324.210 440.000 324.490 444.000 ;
    END
  END io_north_in[27]
  PIN io_north_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 327.430 440.000 327.710 444.000 ;
    END
  END io_north_in[28]
  PIN io_north_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 333.870 440.000 334.150 444.000 ;
    END
  END io_north_in[29]
  PIN io_north_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 85.930 440.000 86.210 444.000 ;
    END
  END io_north_in[2]
  PIN io_north_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.410 15.000 34.690 19.000 ;
    END
  END io_north_in[30]
  PIN io_north_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.630 15.000 37.910 19.000 ;
    END
  END io_north_in[31]
  PIN io_north_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 92.370 440.000 92.650 444.000 ;
    END
  END io_north_in[3]
  PIN io_north_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 95.590 440.000 95.870 444.000 ;
    END
  END io_north_in[4]
  PIN io_north_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 102.030 440.000 102.310 444.000 ;
    END
  END io_north_in[5]
  PIN io_north_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 108.470 440.000 108.750 444.000 ;
    END
  END io_north_in[6]
  PIN io_north_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 114.910 440.000 115.190 444.000 ;
    END
  END io_north_in[7]
  PIN io_north_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 118.130 440.000 118.410 444.000 ;
    END
  END io_north_in[8]
  PIN io_north_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 124.570 440.000 124.850 444.000 ;
    END
  END io_north_in[9]
  PIN io_north_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 153.550 440.000 153.830 444.000 ;
    END
  END io_north_out[0]
  PIN io_north_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 205.070 440.000 205.350 444.000 ;
    END
  END io_north_out[10]
  PIN io_north_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 211.510 440.000 211.790 444.000 ;
    END
  END io_north_out[11]
  PIN io_north_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 217.950 440.000 218.230 444.000 ;
    END
  END io_north_out[12]
  PIN io_north_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 221.170 440.000 221.450 444.000 ;
    END
  END io_north_out[13]
  PIN io_north_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.710 440.000 243.990 444.000 ;
    END
  END io_north_out[14]
  PIN io_north_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 239.440 450.000 240.040 ;
    END
  END io_north_out[15]
  PIN io_north_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 340.310 440.000 340.590 444.000 ;
    END
  END io_north_out[16]
  PIN io_north_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 343.530 440.000 343.810 444.000 ;
    END
  END io_north_out[17]
  PIN io_north_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 349.970 440.000 350.250 444.000 ;
    END
  END io_north_out[18]
  PIN io_north_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 356.410 440.000 356.690 444.000 ;
    END
  END io_north_out[19]
  PIN io_north_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 156.770 440.000 157.050 444.000 ;
    END
  END io_north_out[1]
  PIN io_north_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 362.850 440.000 363.130 444.000 ;
    END
  END io_north_out[20]
  PIN io_north_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 366.070 440.000 366.350 444.000 ;
    END
  END io_north_out[21]
  PIN io_north_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 372.510 440.000 372.790 444.000 ;
    END
  END io_north_out[22]
  PIN io_north_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 378.950 440.000 379.230 444.000 ;
    END
  END io_north_out[23]
  PIN io_north_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 382.170 440.000 382.450 444.000 ;
    END
  END io_north_out[24]
  PIN io_north_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 388.610 440.000 388.890 444.000 ;
    END
  END io_north_out[25]
  PIN io_north_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 395.050 440.000 395.330 444.000 ;
    END
  END io_north_out[26]
  PIN io_north_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 401.490 440.000 401.770 444.000 ;
    END
  END io_north_out[27]
  PIN io_north_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 404.710 440.000 404.990 444.000 ;
    END
  END io_north_out[28]
  PIN io_north_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 411.150 440.000 411.430 444.000 ;
    END
  END io_north_out[29]
  PIN io_north_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 163.210 440.000 163.490 444.000 ;
    END
  END io_north_out[2]
  PIN io_north_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 222.440 450.000 223.040 ;
    END
  END io_north_out[30]
  PIN io_north_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.730 440.000 215.010 444.000 ;
    END
  END io_north_out[31]
  PIN io_north_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 169.650 440.000 169.930 444.000 ;
    END
  END io_north_out[3]
  PIN io_north_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 172.870 440.000 173.150 444.000 ;
    END
  END io_north_out[4]
  PIN io_north_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 179.310 440.000 179.590 444.000 ;
    END
  END io_north_out[5]
  PIN io_north_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 185.750 440.000 186.030 444.000 ;
    END
  END io_north_out[6]
  PIN io_north_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 192.190 440.000 192.470 444.000 ;
    END
  END io_north_out[7]
  PIN io_north_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 195.410 440.000 195.690 444.000 ;
    END
  END io_north_out[8]
  PIN io_north_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 201.850 440.000 202.130 444.000 ;
    END
  END io_north_out[9]
  PIN io_south_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 153.550 15.000 153.830 19.000 ;
    END
  END io_south_in[0]
  PIN io_south_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 208.290 15.000 208.570 19.000 ;
    END
  END io_south_in[10]
  PIN io_south_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 211.510 15.000 211.790 19.000 ;
    END
  END io_south_in[11]
  PIN io_south_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 217.950 15.000 218.230 19.000 ;
    END
  END io_south_in[12]
  PIN io_south_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 224.390 15.000 224.670 19.000 ;
    END
  END io_south_in[13]
  PIN io_south_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.850 15.000 41.130 19.000 ;
    END
  END io_south_in[14]
  PIN io_south_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.070 15.000 44.350 19.000 ;
    END
  END io_south_in[15]
  PIN io_south_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 340.310 15.000 340.590 19.000 ;
    END
  END io_south_in[16]
  PIN io_south_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 343.530 15.000 343.810 19.000 ;
    END
  END io_south_in[17]
  PIN io_south_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 349.970 15.000 350.250 19.000 ;
    END
  END io_south_in[18]
  PIN io_south_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 356.410 15.000 356.690 19.000 ;
    END
  END io_south_in[19]
  PIN io_south_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 156.770 15.000 157.050 19.000 ;
    END
  END io_south_in[1]
  PIN io_south_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 362.850 15.000 363.130 19.000 ;
    END
  END io_south_in[20]
  PIN io_south_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 366.070 15.000 366.350 19.000 ;
    END
  END io_south_in[21]
  PIN io_south_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 372.510 15.000 372.790 19.000 ;
    END
  END io_south_in[22]
  PIN io_south_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 378.950 15.000 379.230 19.000 ;
    END
  END io_south_in[23]
  PIN io_south_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 382.170 15.000 382.450 19.000 ;
    END
  END io_south_in[24]
  PIN io_south_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 388.610 15.000 388.890 19.000 ;
    END
  END io_south_in[25]
  PIN io_south_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 395.050 15.000 395.330 19.000 ;
    END
  END io_south_in[26]
  PIN io_south_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 401.490 15.000 401.770 19.000 ;
    END
  END io_south_in[27]
  PIN io_south_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 404.710 15.000 404.990 19.000 ;
    END
  END io_south_in[28]
  PIN io_south_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 52.440 450.000 53.040 ;
    END
  END io_south_in[29]
  PIN io_south_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 163.210 15.000 163.490 19.000 ;
    END
  END io_south_in[2]
  PIN io_south_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.290 15.000 47.570 19.000 ;
    END
  END io_south_in[30]
  PIN io_south_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.510 15.000 50.790 19.000 ;
    END
  END io_south_in[31]
  PIN io_south_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 169.650 15.000 169.930 19.000 ;
    END
  END io_south_in[3]
  PIN io_south_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 172.870 15.000 173.150 19.000 ;
    END
  END io_south_in[4]
  PIN io_south_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 179.310 15.000 179.590 19.000 ;
    END
  END io_south_in[5]
  PIN io_south_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 185.750 15.000 186.030 19.000 ;
    END
  END io_south_in[6]
  PIN io_south_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 192.190 15.000 192.470 19.000 ;
    END
  END io_south_in[7]
  PIN io_south_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 195.410 15.000 195.690 19.000 ;
    END
  END io_south_in[8]
  PIN io_south_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 201.850 15.000 202.130 19.000 ;
    END
  END io_south_in[9]
  PIN io_south_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 76.270 15.000 76.550 19.000 ;
    END
  END io_south_out[0]
  PIN io_south_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 131.010 15.000 131.290 19.000 ;
    END
  END io_south_out[10]
  PIN io_south_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 134.230 15.000 134.510 19.000 ;
    END
  END io_south_out[11]
  PIN io_south_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 140.670 15.000 140.950 19.000 ;
    END
  END io_south_out[12]
  PIN io_south_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 147.110 15.000 147.390 19.000 ;
    END
  END io_south_out[13]
  PIN io_south_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.390 440.000 224.670 444.000 ;
    END
  END io_south_out[14]
  PIN io_south_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.930 440.000 247.210 444.000 ;
    END
  END io_south_out[15]
  PIN io_south_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 263.030 15.000 263.310 19.000 ;
    END
  END io_south_out[16]
  PIN io_south_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 266.250 15.000 266.530 19.000 ;
    END
  END io_south_out[17]
  PIN io_south_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 272.690 15.000 272.970 19.000 ;
    END
  END io_south_out[18]
  PIN io_south_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 279.130 15.000 279.410 19.000 ;
    END
  END io_south_out[19]
  PIN io_south_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 79.490 15.000 79.770 19.000 ;
    END
  END io_south_out[1]
  PIN io_south_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 285.570 15.000 285.850 19.000 ;
    END
  END io_south_out[20]
  PIN io_south_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 288.790 15.000 289.070 19.000 ;
    END
  END io_south_out[21]
  PIN io_south_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 295.230 15.000 295.510 19.000 ;
    END
  END io_south_out[22]
  PIN io_south_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 301.670 15.000 301.950 19.000 ;
    END
  END io_south_out[23]
  PIN io_south_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 304.890 15.000 305.170 19.000 ;
    END
  END io_south_out[24]
  PIN io_south_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 311.330 15.000 311.610 19.000 ;
    END
  END io_south_out[25]
  PIN io_south_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 317.770 15.000 318.050 19.000 ;
    END
  END io_south_out[26]
  PIN io_south_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 324.210 15.000 324.490 19.000 ;
    END
  END io_south_out[27]
  PIN io_south_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 327.430 15.000 327.710 19.000 ;
    END
  END io_south_out[28]
  PIN io_south_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 333.870 15.000 334.150 19.000 ;
    END
  END io_south_out[29]
  PIN io_south_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 85.930 15.000 86.210 19.000 ;
    END
  END io_south_out[2]
  PIN io_south_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 225.840 450.000 226.440 ;
    END
  END io_south_out[30]
  PIN io_south_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 232.640 450.000 233.240 ;
    END
  END io_south_out[31]
  PIN io_south_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 92.370 15.000 92.650 19.000 ;
    END
  END io_south_out[3]
  PIN io_south_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 95.590 15.000 95.870 19.000 ;
    END
  END io_south_out[4]
  PIN io_south_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 102.030 15.000 102.310 19.000 ;
    END
  END io_south_out[5]
  PIN io_south_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 108.470 15.000 108.750 19.000 ;
    END
  END io_south_out[6]
  PIN io_south_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 114.910 15.000 115.190 19.000 ;
    END
  END io_south_out[7]
  PIN io_south_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 118.130 15.000 118.410 19.000 ;
    END
  END io_south_out[8]
  PIN io_south_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 124.570 15.000 124.850 19.000 ;
    END
  END io_south_out[9]
  PIN io_west_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 15.000 76.240 19.000 76.840 ;
    END
  END io_west_in[0]
  PIN io_west_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 15.000 130.640 19.000 131.240 ;
    END
  END io_west_in[10]
  PIN io_west_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 15.000 134.040 19.000 134.640 ;
    END
  END io_west_in[11]
  PIN io_west_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 15.000 140.840 19.000 141.440 ;
    END
  END io_west_in[12]
  PIN io_west_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 15.000 147.640 19.000 148.240 ;
    END
  END io_west_in[13]
  PIN io_west_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.730 15.000 54.010 19.000 ;
    END
  END io_west_in[14]
  PIN io_west_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.950 15.000 57.230 19.000 ;
    END
  END io_west_in[15]
  PIN io_west_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 15.000 256.440 19.000 257.040 ;
    END
  END io_west_in[16]
  PIN io_west_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 15.000 263.240 19.000 263.840 ;
    END
  END io_west_in[17]
  PIN io_west_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 15.000 270.040 19.000 270.640 ;
    END
  END io_west_in[18]
  PIN io_west_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 15.000 273.440 19.000 274.040 ;
    END
  END io_west_in[19]
  PIN io_west_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 15.000 79.640 19.000 80.240 ;
    END
  END io_west_in[1]
  PIN io_west_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 15.000 280.240 19.000 280.840 ;
    END
  END io_west_in[20]
  PIN io_west_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 15.000 283.640 19.000 284.240 ;
    END
  END io_west_in[21]
  PIN io_west_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 15.000 290.440 19.000 291.040 ;
    END
  END io_west_in[22]
  PIN io_west_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 15.000 297.240 19.000 297.840 ;
    END
  END io_west_in[23]
  PIN io_west_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 15.000 300.640 19.000 301.240 ;
    END
  END io_west_in[24]
  PIN io_west_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 15.000 307.440 19.000 308.040 ;
    END
  END io_west_in[25]
  PIN io_west_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 15.000 310.840 19.000 311.440 ;
    END
  END io_west_in[26]
  PIN io_west_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 15.000 317.640 19.000 318.240 ;
    END
  END io_west_in[27]
  PIN io_west_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 15.000 324.440 19.000 325.040 ;
    END
  END io_west_in[28]
  PIN io_west_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 15.000 327.840 19.000 328.440 ;
    END
  END io_west_in[29]
  PIN io_west_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 15.000 86.440 19.000 87.040 ;
    END
  END io_west_in[2]
  PIN io_west_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.170 15.000 60.450 19.000 ;
    END
  END io_west_in[30]
  PIN io_west_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.390 15.000 63.670 19.000 ;
    END
  END io_west_in[31]
  PIN io_west_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 15.000 93.240 19.000 93.840 ;
    END
  END io_west_in[3]
  PIN io_west_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 15.000 96.640 19.000 97.240 ;
    END
  END io_west_in[4]
  PIN io_west_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 15.000 103.440 19.000 104.040 ;
    END
  END io_west_in[5]
  PIN io_west_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 15.000 106.840 19.000 107.440 ;
    END
  END io_west_in[6]
  PIN io_west_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 15.000 113.640 19.000 114.240 ;
    END
  END io_west_in[7]
  PIN io_west_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 15.000 120.440 19.000 121.040 ;
    END
  END io_west_in[8]
  PIN io_west_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 15.000 123.840 19.000 124.440 ;
    END
  END io_west_in[9]
  PIN io_west_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 15.000 151.040 19.000 151.640 ;
    END
  END io_west_out[0]
  PIN io_west_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 15.000 205.440 19.000 206.040 ;
    END
  END io_west_out[10]
  PIN io_west_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 15.000 212.240 19.000 212.840 ;
    END
  END io_west_out[11]
  PIN io_west_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 15.000 215.640 19.000 216.240 ;
    END
  END io_west_out[12]
  PIN io_west_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 15.000 222.440 19.000 223.040 ;
    END
  END io_west_out[13]
  PIN io_west_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.610 440.000 227.890 444.000 ;
    END
  END io_west_out[14]
  PIN io_west_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 242.840 450.000 243.440 ;
    END
  END io_west_out[15]
  PIN io_west_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 15.000 334.640 19.000 335.240 ;
    END
  END io_west_out[16]
  PIN io_west_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 15.000 338.040 19.000 338.640 ;
    END
  END io_west_out[17]
  PIN io_west_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 15.000 344.840 19.000 345.440 ;
    END
  END io_west_out[18]
  PIN io_west_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 15.000 351.640 19.000 352.240 ;
    END
  END io_west_out[19]
  PIN io_west_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 15.000 157.840 19.000 158.440 ;
    END
  END io_west_out[1]
  PIN io_west_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 15.000 355.040 19.000 355.640 ;
    END
  END io_west_out[20]
  PIN io_west_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 15.000 361.840 19.000 362.440 ;
    END
  END io_west_out[21]
  PIN io_west_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 15.000 365.240 19.000 365.840 ;
    END
  END io_west_out[22]
  PIN io_west_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 15.000 372.040 19.000 372.640 ;
    END
  END io_west_out[23]
  PIN io_west_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 15.000 378.840 19.000 379.440 ;
    END
  END io_west_out[24]
  PIN io_west_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 15.000 382.240 19.000 382.840 ;
    END
  END io_west_out[25]
  PIN io_west_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 15.000 389.040 19.000 389.640 ;
    END
  END io_west_out[26]
  PIN io_west_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 15.000 392.440 19.000 393.040 ;
    END
  END io_west_out[27]
  PIN io_west_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 15.000 399.240 19.000 399.840 ;
    END
  END io_west_out[28]
  PIN io_west_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 15.000 406.040 19.000 406.640 ;
    END
  END io_west_out[29]
  PIN io_west_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 15.000 161.240 19.000 161.840 ;
    END
  END io_west_out[2]
  PIN io_west_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.050 440.000 234.330 444.000 ;
    END
  END io_west_out[30]
  PIN io_west_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.490 440.000 240.770 444.000 ;
    END
  END io_west_out[31]
  PIN io_west_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 15.000 168.040 19.000 168.640 ;
    END
  END io_west_out[3]
  PIN io_west_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 15.000 174.840 19.000 175.440 ;
    END
  END io_west_out[4]
  PIN io_west_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 15.000 178.240 19.000 178.840 ;
    END
  END io_west_out[5]
  PIN io_west_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 15.000 185.040 19.000 185.640 ;
    END
  END io_west_out[6]
  PIN io_west_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 15.000 188.440 19.000 189.040 ;
    END
  END io_west_out[7]
  PIN io_west_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 15.000 195.240 19.000 195.840 ;
    END
  END io_west_out[8]
  PIN io_west_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 15.000 202.040 19.000 202.640 ;
    END
  END io_west_out[9]
  PIN le_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 62.640 450.000 63.240 ;
    END
  END le_clk
  PIN le_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 66.040 450.000 66.640 ;
    END
  END le_en
  PIN le_nrst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 72.840 450.000 73.440 ;
    END
  END le_nrst
  PIN nrst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.860700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 188.970 440.000 189.250 444.000 ;
    END
  END nrst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 16.780 16.880 18.380 445.520 ;
    END
    PORT
      LAYER met5 ;
        RECT 16.780 16.880 450.580 18.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 16.780 443.920 450.580 445.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 448.980 16.880 450.580 445.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 88.580 13.580 90.180 50.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 88.580 405.145 90.180 448.820 ;
    END
    PORT
      LAYER met4 ;
        RECT 180.580 13.580 182.180 50.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 180.580 405.145 182.180 448.820 ;
    END
    PORT
      LAYER met4 ;
        RECT 272.580 13.580 274.180 50.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 272.580 405.145 274.180 448.820 ;
    END
    PORT
      LAYER met4 ;
        RECT 364.580 13.580 366.180 50.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 364.580 405.145 366.180 448.820 ;
    END
    PORT
      LAYER met5 ;
        RECT 13.480 88.680 453.880 90.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 13.480 180.680 453.880 182.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 13.480 272.680 453.880 274.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 13.480 364.680 453.880 366.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 29.380 35.120 30.980 424.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 432.340 35.120 433.940 424.560 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 13.480 13.580 15.080 448.820 ;
    END
    PORT
      LAYER met5 ;
        RECT 13.480 13.580 453.880 15.180 ;
    END
    PORT
      LAYER met5 ;
        RECT 13.480 447.220 453.880 448.820 ;
    END
    PORT
      LAYER met4 ;
        RECT 452.280 13.580 453.880 448.820 ;
    END
    PORT
      LAYER met4 ;
        RECT 91.880 13.580 93.480 50.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 91.880 405.145 93.480 448.820 ;
    END
    PORT
      LAYER met4 ;
        RECT 183.880 13.580 185.480 50.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 183.880 405.145 185.480 448.820 ;
    END
    PORT
      LAYER met4 ;
        RECT 275.880 13.580 277.480 50.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 275.880 405.145 277.480 448.820 ;
    END
    PORT
      LAYER met4 ;
        RECT 367.880 13.580 369.480 50.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 367.880 405.145 369.480 448.820 ;
    END
    PORT
      LAYER met5 ;
        RECT 13.480 91.980 453.880 93.580 ;
    END
    PORT
      LAYER met5 ;
        RECT 13.480 183.980 453.880 185.580 ;
    END
    PORT
      LAYER met5 ;
        RECT 13.480 275.980 453.880 277.580 ;
    END
    PORT
      LAYER met5 ;
        RECT 13.480 367.980 453.880 369.580 ;
    END
    PORT
      LAYER met4 ;
        RECT 33.060 35.120 34.660 424.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 436.020 35.120 437.620 424.560 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 24.190 24.395 443.170 438.005 ;
      LAYER li1 ;
        RECT 24.380 24.395 442.980 438.005 ;
      LAYER met1 ;
        RECT 19.670 24.240 443.650 438.600 ;
      LAYER met2 ;
        RECT 19.690 439.720 75.990 440.410 ;
        RECT 76.830 439.720 79.210 440.410 ;
        RECT 80.050 439.720 85.650 440.410 ;
        RECT 86.490 439.720 92.090 440.410 ;
        RECT 92.930 439.720 95.310 440.410 ;
        RECT 96.150 439.720 101.750 440.410 ;
        RECT 102.590 439.720 108.190 440.410 ;
        RECT 109.030 439.720 114.630 440.410 ;
        RECT 115.470 439.720 117.850 440.410 ;
        RECT 118.690 439.720 124.290 440.410 ;
        RECT 125.130 439.720 130.730 440.410 ;
        RECT 131.570 439.720 133.950 440.410 ;
        RECT 134.790 439.720 140.390 440.410 ;
        RECT 141.230 439.720 146.830 440.410 ;
        RECT 147.670 439.720 153.270 440.410 ;
        RECT 154.110 439.720 156.490 440.410 ;
        RECT 157.330 439.720 162.930 440.410 ;
        RECT 163.770 439.720 169.370 440.410 ;
        RECT 170.210 439.720 172.590 440.410 ;
        RECT 173.430 439.720 179.030 440.410 ;
        RECT 179.870 439.720 182.250 440.410 ;
        RECT 183.090 439.720 185.470 440.410 ;
        RECT 186.310 439.720 188.690 440.410 ;
        RECT 189.530 439.720 191.910 440.410 ;
        RECT 192.750 439.720 195.130 440.410 ;
        RECT 195.970 439.720 198.350 440.410 ;
        RECT 199.190 439.720 201.570 440.410 ;
        RECT 202.410 439.720 204.790 440.410 ;
        RECT 205.630 439.720 208.010 440.410 ;
        RECT 208.850 439.720 211.230 440.410 ;
        RECT 212.070 439.720 214.450 440.410 ;
        RECT 215.290 439.720 217.670 440.410 ;
        RECT 218.510 439.720 220.890 440.410 ;
        RECT 221.730 439.720 224.110 440.410 ;
        RECT 224.950 439.720 227.330 440.410 ;
        RECT 228.170 439.720 230.550 440.410 ;
        RECT 231.390 439.720 233.770 440.410 ;
        RECT 234.610 439.720 236.990 440.410 ;
        RECT 237.830 439.720 240.210 440.410 ;
        RECT 241.050 439.720 243.430 440.410 ;
        RECT 244.270 439.720 246.650 440.410 ;
        RECT 247.490 439.720 249.870 440.410 ;
        RECT 250.710 439.720 262.750 440.410 ;
        RECT 263.590 439.720 265.970 440.410 ;
        RECT 266.810 439.720 272.410 440.410 ;
        RECT 273.250 439.720 278.850 440.410 ;
        RECT 279.690 439.720 285.290 440.410 ;
        RECT 286.130 439.720 288.510 440.410 ;
        RECT 289.350 439.720 294.950 440.410 ;
        RECT 295.790 439.720 301.390 440.410 ;
        RECT 302.230 439.720 304.610 440.410 ;
        RECT 305.450 439.720 311.050 440.410 ;
        RECT 311.890 439.720 317.490 440.410 ;
        RECT 318.330 439.720 323.930 440.410 ;
        RECT 324.770 439.720 327.150 440.410 ;
        RECT 327.990 439.720 333.590 440.410 ;
        RECT 334.430 439.720 340.030 440.410 ;
        RECT 340.870 439.720 343.250 440.410 ;
        RECT 344.090 439.720 349.690 440.410 ;
        RECT 350.530 439.720 356.130 440.410 ;
        RECT 356.970 439.720 362.570 440.410 ;
        RECT 363.410 439.720 365.790 440.410 ;
        RECT 366.630 439.720 372.230 440.410 ;
        RECT 373.070 439.720 378.670 440.410 ;
        RECT 379.510 439.720 381.890 440.410 ;
        RECT 382.730 439.720 388.330 440.410 ;
        RECT 389.170 439.720 394.770 440.410 ;
        RECT 395.610 439.720 401.210 440.410 ;
        RECT 402.050 439.720 404.430 440.410 ;
        RECT 405.270 439.720 410.870 440.410 ;
        RECT 411.710 439.720 443.630 440.410 ;
        RECT 19.690 19.280 443.630 439.720 ;
        RECT 19.690 18.670 21.250 19.280 ;
        RECT 22.090 18.670 24.470 19.280 ;
        RECT 25.310 18.670 27.690 19.280 ;
        RECT 28.530 18.670 30.910 19.280 ;
        RECT 31.750 18.670 34.130 19.280 ;
        RECT 34.970 18.670 37.350 19.280 ;
        RECT 38.190 18.670 40.570 19.280 ;
        RECT 41.410 18.670 43.790 19.280 ;
        RECT 44.630 18.670 47.010 19.280 ;
        RECT 47.850 18.670 50.230 19.280 ;
        RECT 51.070 18.670 53.450 19.280 ;
        RECT 54.290 18.670 56.670 19.280 ;
        RECT 57.510 18.670 59.890 19.280 ;
        RECT 60.730 18.670 63.110 19.280 ;
        RECT 63.950 18.670 75.990 19.280 ;
        RECT 76.830 18.670 79.210 19.280 ;
        RECT 80.050 18.670 85.650 19.280 ;
        RECT 86.490 18.670 92.090 19.280 ;
        RECT 92.930 18.670 95.310 19.280 ;
        RECT 96.150 18.670 101.750 19.280 ;
        RECT 102.590 18.670 108.190 19.280 ;
        RECT 109.030 18.670 114.630 19.280 ;
        RECT 115.470 18.670 117.850 19.280 ;
        RECT 118.690 18.670 124.290 19.280 ;
        RECT 125.130 18.670 130.730 19.280 ;
        RECT 131.570 18.670 133.950 19.280 ;
        RECT 134.790 18.670 140.390 19.280 ;
        RECT 141.230 18.670 146.830 19.280 ;
        RECT 147.670 18.670 153.270 19.280 ;
        RECT 154.110 18.670 156.490 19.280 ;
        RECT 157.330 18.670 162.930 19.280 ;
        RECT 163.770 18.670 169.370 19.280 ;
        RECT 170.210 18.670 172.590 19.280 ;
        RECT 173.430 18.670 179.030 19.280 ;
        RECT 179.870 18.670 185.470 19.280 ;
        RECT 186.310 18.670 191.910 19.280 ;
        RECT 192.750 18.670 195.130 19.280 ;
        RECT 195.970 18.670 201.570 19.280 ;
        RECT 202.410 18.670 208.010 19.280 ;
        RECT 208.850 18.670 211.230 19.280 ;
        RECT 212.070 18.670 217.670 19.280 ;
        RECT 218.510 18.670 224.110 19.280 ;
        RECT 224.950 18.670 262.750 19.280 ;
        RECT 263.590 18.670 265.970 19.280 ;
        RECT 266.810 18.670 272.410 19.280 ;
        RECT 273.250 18.670 278.850 19.280 ;
        RECT 279.690 18.670 285.290 19.280 ;
        RECT 286.130 18.670 288.510 19.280 ;
        RECT 289.350 18.670 294.950 19.280 ;
        RECT 295.790 18.670 301.390 19.280 ;
        RECT 302.230 18.670 304.610 19.280 ;
        RECT 305.450 18.670 311.050 19.280 ;
        RECT 311.890 18.670 317.490 19.280 ;
        RECT 318.330 18.670 323.930 19.280 ;
        RECT 324.770 18.670 327.150 19.280 ;
        RECT 327.990 18.670 333.590 19.280 ;
        RECT 334.430 18.670 340.030 19.280 ;
        RECT 340.870 18.670 343.250 19.280 ;
        RECT 344.090 18.670 349.690 19.280 ;
        RECT 350.530 18.670 356.130 19.280 ;
        RECT 356.970 18.670 362.570 19.280 ;
        RECT 363.410 18.670 365.790 19.280 ;
        RECT 366.630 18.670 372.230 19.280 ;
        RECT 373.070 18.670 378.670 19.280 ;
        RECT 379.510 18.670 381.890 19.280 ;
        RECT 382.730 18.670 388.330 19.280 ;
        RECT 389.170 18.670 394.770 19.280 ;
        RECT 395.610 18.670 401.210 19.280 ;
        RECT 402.050 18.670 404.430 19.280 ;
        RECT 405.270 18.670 443.630 19.280 ;
      LAYER met3 ;
        RECT 19.000 407.040 446.000 438.085 ;
        RECT 19.400 405.640 445.600 407.040 ;
        RECT 19.000 400.240 446.000 405.640 ;
        RECT 19.400 398.840 445.600 400.240 ;
        RECT 19.000 393.440 446.000 398.840 ;
        RECT 19.400 392.040 445.600 393.440 ;
        RECT 19.000 390.040 446.000 392.040 ;
        RECT 19.400 388.640 445.600 390.040 ;
        RECT 19.000 383.240 446.000 388.640 ;
        RECT 19.400 381.840 445.600 383.240 ;
        RECT 19.000 379.840 446.000 381.840 ;
        RECT 19.400 378.440 445.600 379.840 ;
        RECT 19.000 373.040 446.000 378.440 ;
        RECT 19.400 371.640 445.600 373.040 ;
        RECT 19.000 366.240 446.000 371.640 ;
        RECT 19.400 364.840 445.600 366.240 ;
        RECT 19.000 362.840 446.000 364.840 ;
        RECT 19.400 361.440 445.600 362.840 ;
        RECT 19.000 356.040 446.000 361.440 ;
        RECT 19.400 354.640 445.600 356.040 ;
        RECT 19.000 352.640 446.000 354.640 ;
        RECT 19.400 351.240 445.600 352.640 ;
        RECT 19.000 345.840 446.000 351.240 ;
        RECT 19.400 344.440 445.600 345.840 ;
        RECT 19.000 339.040 446.000 344.440 ;
        RECT 19.400 337.640 445.600 339.040 ;
        RECT 19.000 335.640 446.000 337.640 ;
        RECT 19.400 334.240 445.600 335.640 ;
        RECT 19.000 328.840 446.000 334.240 ;
        RECT 19.400 327.440 445.600 328.840 ;
        RECT 19.000 325.440 446.000 327.440 ;
        RECT 19.400 324.040 445.600 325.440 ;
        RECT 19.000 318.640 446.000 324.040 ;
        RECT 19.400 317.240 445.600 318.640 ;
        RECT 19.000 311.840 446.000 317.240 ;
        RECT 19.400 310.440 445.600 311.840 ;
        RECT 19.000 308.440 446.000 310.440 ;
        RECT 19.400 307.040 445.600 308.440 ;
        RECT 19.000 301.640 446.000 307.040 ;
        RECT 19.400 300.240 445.600 301.640 ;
        RECT 19.000 298.240 446.000 300.240 ;
        RECT 19.400 296.840 445.600 298.240 ;
        RECT 19.000 291.440 446.000 296.840 ;
        RECT 19.400 290.040 445.600 291.440 ;
        RECT 19.000 284.640 446.000 290.040 ;
        RECT 19.400 283.240 445.600 284.640 ;
        RECT 19.000 281.240 446.000 283.240 ;
        RECT 19.400 279.840 445.600 281.240 ;
        RECT 19.000 274.440 446.000 279.840 ;
        RECT 19.400 273.040 445.600 274.440 ;
        RECT 19.000 271.040 446.000 273.040 ;
        RECT 19.400 269.640 445.600 271.040 ;
        RECT 19.000 264.240 446.000 269.640 ;
        RECT 19.400 262.840 445.600 264.240 ;
        RECT 19.000 257.440 446.000 262.840 ;
        RECT 19.400 256.040 445.600 257.440 ;
        RECT 19.000 243.840 446.000 256.040 ;
        RECT 19.000 242.440 445.600 243.840 ;
        RECT 19.000 240.440 446.000 242.440 ;
        RECT 19.000 239.040 445.600 240.440 ;
        RECT 19.000 237.040 446.000 239.040 ;
        RECT 19.000 235.640 445.600 237.040 ;
        RECT 19.000 233.640 446.000 235.640 ;
        RECT 19.000 232.240 445.600 233.640 ;
        RECT 19.000 226.840 446.000 232.240 ;
        RECT 19.400 225.440 445.600 226.840 ;
        RECT 19.000 223.440 446.000 225.440 ;
        RECT 19.400 222.040 445.600 223.440 ;
        RECT 19.000 220.040 446.000 222.040 ;
        RECT 19.000 218.640 445.600 220.040 ;
        RECT 19.000 216.640 446.000 218.640 ;
        RECT 19.400 215.240 445.600 216.640 ;
        RECT 19.000 213.240 446.000 215.240 ;
        RECT 19.400 211.840 445.600 213.240 ;
        RECT 19.000 206.440 446.000 211.840 ;
        RECT 19.400 205.040 445.600 206.440 ;
        RECT 19.000 203.040 446.000 205.040 ;
        RECT 19.400 201.640 445.600 203.040 ;
        RECT 19.000 196.240 446.000 201.640 ;
        RECT 19.400 194.840 445.600 196.240 ;
        RECT 19.000 189.440 446.000 194.840 ;
        RECT 19.400 188.040 445.600 189.440 ;
        RECT 19.000 186.040 446.000 188.040 ;
        RECT 19.400 184.640 445.600 186.040 ;
        RECT 19.000 179.240 446.000 184.640 ;
        RECT 19.400 177.840 445.600 179.240 ;
        RECT 19.000 175.840 446.000 177.840 ;
        RECT 19.400 174.440 445.600 175.840 ;
        RECT 19.000 169.040 446.000 174.440 ;
        RECT 19.400 167.640 445.600 169.040 ;
        RECT 19.000 162.240 446.000 167.640 ;
        RECT 19.400 160.840 445.600 162.240 ;
        RECT 19.000 158.840 446.000 160.840 ;
        RECT 19.400 157.440 445.600 158.840 ;
        RECT 19.000 152.040 446.000 157.440 ;
        RECT 19.400 150.640 445.600 152.040 ;
        RECT 19.000 148.640 446.000 150.640 ;
        RECT 19.400 147.240 445.600 148.640 ;
        RECT 19.000 141.840 446.000 147.240 ;
        RECT 19.400 140.440 445.600 141.840 ;
        RECT 19.000 135.040 446.000 140.440 ;
        RECT 19.400 133.640 445.600 135.040 ;
        RECT 19.000 131.640 446.000 133.640 ;
        RECT 19.400 130.240 445.600 131.640 ;
        RECT 19.000 124.840 446.000 130.240 ;
        RECT 19.400 123.440 445.600 124.840 ;
        RECT 19.000 121.440 446.000 123.440 ;
        RECT 19.400 120.040 445.600 121.440 ;
        RECT 19.000 114.640 446.000 120.040 ;
        RECT 19.400 113.240 445.600 114.640 ;
        RECT 19.000 107.840 446.000 113.240 ;
        RECT 19.400 106.440 445.600 107.840 ;
        RECT 19.000 104.440 446.000 106.440 ;
        RECT 19.400 103.040 445.600 104.440 ;
        RECT 19.000 97.640 446.000 103.040 ;
        RECT 19.400 96.240 445.600 97.640 ;
        RECT 19.000 94.240 446.000 96.240 ;
        RECT 19.400 92.840 445.600 94.240 ;
        RECT 19.000 87.440 446.000 92.840 ;
        RECT 19.400 86.040 445.600 87.440 ;
        RECT 19.000 80.640 446.000 86.040 ;
        RECT 19.400 79.240 445.600 80.640 ;
        RECT 19.000 77.240 446.000 79.240 ;
        RECT 19.400 75.840 445.600 77.240 ;
        RECT 19.000 73.840 446.000 75.840 ;
        RECT 19.000 72.440 445.600 73.840 ;
        RECT 19.000 67.040 446.000 72.440 ;
        RECT 19.000 65.640 445.600 67.040 ;
        RECT 19.000 63.640 446.000 65.640 ;
        RECT 19.000 62.240 445.600 63.640 ;
        RECT 19.000 53.440 446.000 62.240 ;
        RECT 19.000 52.040 445.600 53.440 ;
        RECT 19.000 24.315 446.000 52.040 ;
      LAYER met4 ;
        RECT 52.420 404.745 88.180 406.320 ;
        RECT 90.580 404.745 91.480 406.320 ;
        RECT 93.880 404.745 180.180 406.320 ;
        RECT 182.580 404.745 183.480 406.320 ;
        RECT 185.880 404.745 272.180 406.320 ;
        RECT 274.580 404.745 275.480 406.320 ;
        RECT 277.880 404.745 364.180 406.320 ;
        RECT 366.580 404.745 367.480 406.320 ;
        RECT 369.880 404.745 407.320 406.320 ;
        RECT 52.420 51.535 407.320 404.745 ;
      LAYER met5 ;
        RECT 52.420 371.180 412.960 404.540 ;
        RECT 52.420 279.180 412.960 363.080 ;
        RECT 52.420 187.180 412.960 271.080 ;
        RECT 52.420 95.180 412.960 179.080 ;
        RECT 52.420 54.640 412.960 87.080 ;
  END
END fpga
END LIBRARY

