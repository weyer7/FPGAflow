magic
tech sky130A
magscale 1 2
timestamp 1752769994
<< viali >>
rect 16553 87405 16587 87439
rect 34697 87405 34731 87439
rect 37759 87405 37793 87439
rect 39691 87405 39725 87439
rect 41137 87405 41171 87439
rect 42425 87405 42459 87439
rect 44357 87405 44391 87439
rect 54181 87405 54215 87439
rect 68829 87405 68863 87439
rect 76557 87405 76591 87439
rect 15289 87337 15323 87371
rect 16369 87337 16403 87371
rect 16737 87337 16771 87371
rect 17381 87337 17415 87371
rect 17565 87337 17599 87371
rect 18669 87337 18703 87371
rect 18853 87337 18887 87371
rect 19157 87337 19191 87371
rect 19497 87337 19531 87371
rect 20601 87337 20635 87371
rect 20785 87337 20819 87371
rect 21889 87337 21923 87371
rect 22073 87337 22107 87371
rect 23177 87337 23211 87371
rect 23361 87337 23395 87371
rect 23665 87337 23699 87371
rect 24005 87337 24039 87371
rect 25109 87337 25143 87371
rect 25293 87337 25327 87371
rect 26397 87337 26431 87371
rect 26581 87337 26615 87371
rect 26885 87337 26919 87371
rect 27225 87337 27259 87371
rect 28329 87337 28363 87371
rect 28513 87337 28547 87371
rect 29617 87337 29651 87371
rect 29801 87337 29835 87371
rect 30745 87337 30779 87371
rect 31641 87337 31675 87371
rect 32677 87337 32711 87371
rect 33965 87337 33999 87371
rect 34861 87337 34895 87371
rect 35934 87337 35968 87371
rect 37456 87337 37490 87371
rect 37590 87337 37624 87371
rect 38050 87337 38084 87371
rect 38473 87337 38507 87371
rect 39485 87337 39519 87371
rect 40405 87337 40439 87371
rect 41301 87337 41335 87371
rect 41761 87337 41795 87371
rect 42589 87337 42623 87371
rect 43049 87337 43083 87371
rect 43662 87337 43696 87371
rect 44521 87337 44555 87371
rect 44981 87337 45015 87371
rect 45625 87337 45659 87371
rect 46269 87337 46303 87371
rect 46913 87337 46947 87371
rect 47557 87337 47591 87371
rect 48201 87337 48235 87371
rect 48845 87337 48879 87371
rect 49489 87337 49523 87371
rect 50133 87337 50167 87371
rect 52641 87337 52675 87371
rect 53721 87337 53755 87371
rect 53997 87337 54031 87371
rect 54733 87337 54767 87371
rect 54917 87337 54951 87371
rect 56021 87337 56055 87371
rect 56205 87337 56239 87371
rect 57309 87337 57343 87371
rect 57493 87337 57527 87371
rect 57797 87337 57831 87371
rect 58137 87337 58171 87371
rect 59241 87337 59275 87371
rect 59425 87337 59459 87371
rect 60529 87337 60563 87371
rect 60713 87337 60747 87371
rect 61017 87337 61051 87371
rect 61357 87337 61391 87371
rect 62461 87337 62495 87371
rect 62645 87337 62679 87371
rect 63749 87337 63783 87371
rect 63933 87337 63967 87371
rect 65037 87337 65071 87371
rect 65221 87337 65255 87371
rect 65525 87337 65559 87371
rect 65865 87337 65899 87371
rect 66969 87337 67003 87371
rect 67153 87337 67187 87371
rect 68097 87337 68131 87371
rect 68993 87337 69027 87371
rect 70029 87337 70063 87371
rect 71317 87337 71351 87371
rect 72605 87337 72639 87371
rect 73501 87337 73535 87371
rect 74537 87337 74571 87371
rect 75825 87337 75859 87371
rect 76721 87337 76755 87371
rect 77757 87337 77791 87371
rect 79045 87337 79079 87371
rect 80370 87337 80404 87371
rect 81229 87337 81263 87371
rect 82265 87337 82299 87371
rect 36609 87269 36643 87303
rect 39369 87269 39403 87303
rect 39921 87269 39955 87303
rect 15541 87201 15575 87235
rect 16210 87201 16244 87235
rect 17222 87201 17256 87235
rect 18510 87201 18544 87235
rect 19359 87201 19393 87235
rect 20442 87201 20476 87235
rect 21730 87201 21764 87235
rect 23018 87201 23052 87235
rect 23867 87201 23901 87235
rect 24950 87201 24984 87235
rect 26237 87201 26271 87235
rect 27087 87201 27121 87235
rect 28169 87201 28203 87235
rect 29458 87201 29492 87235
rect 30951 87201 30985 87235
rect 31477 87201 31511 87235
rect 32883 87201 32917 87235
rect 34171 87201 34205 87235
rect 36103 87201 36137 87235
rect 38219 87201 38253 87235
rect 40611 87201 40645 87235
rect 43831 87201 43865 87235
rect 52893 87201 52927 87235
rect 53562 87201 53596 87235
rect 54574 87201 54608 87235
rect 55862 87201 55896 87235
rect 57150 87201 57184 87235
rect 57999 87201 58033 87235
rect 59082 87201 59116 87235
rect 60370 87201 60404 87235
rect 61219 87201 61253 87235
rect 62311 87201 62345 87235
rect 63589 87201 63623 87235
rect 64878 87201 64912 87235
rect 65727 87201 65761 87235
rect 66810 87201 66844 87235
rect 68303 87201 68337 87235
rect 70235 87201 70269 87235
rect 71523 87201 71557 87235
rect 72811 87201 72845 87235
rect 73337 87201 73371 87235
rect 74743 87201 74777 87235
rect 76031 87201 76065 87235
rect 77963 87201 77997 87235
rect 79251 87201 79285 87235
rect 80539 87201 80573 87235
rect 81065 87201 81099 87235
rect 82471 87201 82505 87235
rect 37621 86861 37655 86895
rect 38541 86861 38575 86895
rect 37805 86589 37839 86623
rect 45441 84685 45475 84719
rect 50317 84685 50351 84719
rect 12873 84617 12907 84651
rect 11769 84549 11803 84583
rect 45625 84549 45659 84583
rect 28881 84481 28915 84515
rect 30585 84481 30619 84515
rect 31089 84481 31123 84515
rect 41049 84481 41083 84515
rect 42773 84481 42807 84515
rect 42957 84481 42991 84515
rect 10665 84413 10699 84447
rect 13977 84413 14011 84447
rect 30905 84413 30939 84447
rect 40841 84413 40875 84447
rect 45809 84413 45843 84447
rect 45993 84413 46027 84447
rect 48109 84413 48143 84447
rect 49213 84413 49247 84447
rect 51421 84413 51455 84447
rect 5257 81285 5291 81319
rect 5421 81285 5455 81319
rect 87761 81285 87795 81319
rect 88221 81285 88255 81319
rect 88061 81217 88095 81251
rect 5421 80197 5455 80231
rect 87761 80197 87795 80231
rect 88221 80197 88255 80231
rect 88061 80129 88095 80163
rect 5257 80061 5291 80095
rect 88061 78701 88095 78735
rect 5421 78633 5455 78667
rect 87945 78633 87979 78667
rect 88221 78633 88255 78667
rect 5257 78497 5291 78531
rect 5421 78021 5455 78055
rect 87761 78021 87795 78055
rect 88221 78021 88255 78055
rect 88061 77953 88095 77987
rect 5257 77885 5291 77919
rect 5421 76933 5455 76967
rect 87761 76933 87795 76967
rect 5257 76797 5291 76831
rect 87577 76797 87611 76831
rect 88037 76797 88071 76831
rect 5421 75845 5455 75879
rect 87761 75845 87795 75879
rect 88221 75845 88255 75879
rect 5257 75777 5291 75811
rect 88057 75777 88091 75811
rect 87761 74825 87795 74859
rect 5257 74757 5291 74791
rect 5421 74757 5455 74791
rect 88057 74757 88091 74791
rect 88221 74757 88255 74791
rect 88062 73261 88096 73295
rect 5421 73193 5455 73227
rect 87945 73193 87979 73227
rect 88221 73193 88255 73227
rect 5257 73057 5291 73091
rect 5421 72581 5455 72615
rect 87761 72581 87795 72615
rect 88221 72581 88255 72615
rect 5257 72445 5291 72479
rect 88062 72445 88096 72479
rect 5421 71493 5455 71527
rect 87761 71493 87795 71527
rect 88221 71493 88255 71527
rect 88061 71425 88095 71459
rect 5257 71357 5291 71391
rect 5421 70405 5455 70439
rect 87761 70405 87795 70439
rect 88221 70405 88255 70439
rect 5257 70337 5291 70371
rect 88061 70337 88095 70371
rect 5421 69317 5455 69351
rect 87761 69317 87795 69351
rect 88221 69317 88255 69351
rect 5257 69249 5291 69283
rect 88062 69249 88096 69283
rect 88061 67821 88095 67855
rect 5421 67753 5455 67787
rect 87945 67753 87979 67787
rect 88221 67753 88255 67787
rect 5257 67617 5291 67651
rect 5421 67141 5455 67175
rect 87761 67141 87795 67175
rect 88221 67141 88255 67175
rect 88062 67073 88096 67107
rect 5257 67005 5291 67039
rect 5375 66121 5409 66155
rect 5173 66053 5207 66087
rect 5513 66053 5547 66087
rect 87969 66053 88003 66087
rect 88175 65917 88209 65951
rect 5375 65033 5409 65067
rect 5173 64965 5207 64999
rect 5513 64965 5547 64999
rect 87969 64965 88003 64999
rect 88175 64829 88209 64863
rect 7537 64557 7571 64591
rect 5173 63877 5207 63911
rect 5513 63877 5547 63911
rect 7401 63877 7435 63911
rect 87969 63877 88003 63911
rect 5375 63741 5409 63775
rect 6617 63741 6651 63775
rect 88175 63741 88209 63775
rect 7537 63469 7571 63503
rect 5173 62313 5207 62347
rect 5513 62313 5547 62347
rect 87969 62313 88003 62347
rect 5375 62177 5409 62211
rect 88175 62109 88209 62143
rect 5173 61701 5207 61735
rect 5513 61701 5547 61735
rect 87969 61701 88003 61735
rect 5375 61633 5409 61667
rect 88175 61565 88209 61599
rect 5173 60613 5207 60647
rect 5513 60613 5547 60647
rect 87969 60613 88003 60647
rect 5375 60545 5409 60579
rect 88175 60477 88209 60511
rect 5173 59525 5207 59559
rect 5513 59525 5547 59559
rect 87969 59525 88003 59559
rect 5375 59389 5409 59423
rect 88175 59389 88209 59423
rect 5173 58437 5207 58471
rect 5513 58437 5547 58471
rect 87969 58437 88003 58471
rect 5375 58301 5409 58335
rect 88175 58301 88209 58335
rect 5375 56941 5409 56975
rect 88175 56941 88209 56975
rect 5173 56873 5207 56907
rect 5513 56873 5547 56907
rect 87969 56873 88003 56907
rect 5375 56329 5409 56363
rect 5173 56261 5207 56295
rect 5513 56261 5547 56295
rect 87969 56261 88003 56295
rect 88175 56125 88209 56159
rect 5375 55241 5409 55275
rect 5173 55173 5207 55207
rect 5513 55173 5547 55207
rect 87969 55173 88003 55207
rect 88175 55037 88209 55071
rect 5375 54153 5409 54187
rect 5173 54085 5207 54119
rect 5513 54085 5547 54119
rect 87969 54085 88003 54119
rect 88175 53949 88209 53983
rect 5375 53065 5409 53099
rect 5173 52997 5207 53031
rect 5513 52997 5547 53031
rect 87969 52997 88003 53031
rect 88175 52861 88209 52895
rect 5375 51501 5409 51535
rect 5173 51433 5207 51467
rect 5513 51433 5547 51467
rect 87969 51433 88003 51467
rect 88175 51297 88209 51331
rect 85645 50685 85679 50719
rect 85645 49597 85679 49631
rect 88221 48645 88255 48679
rect 85645 48577 85679 48611
rect 88221 47965 88255 47999
rect 87969 47557 88003 47591
rect 88175 47421 88209 47455
rect 88221 46877 88255 46911
rect 7353 45517 7387 45551
rect 85829 45517 85863 45551
rect 7169 45449 7203 45483
rect 5173 45381 5207 45415
rect 5513 45381 5547 45415
rect 86013 45381 86047 45415
rect 88221 45381 88255 45415
rect 5375 45313 5409 45347
rect 85645 45245 85679 45279
rect 86197 45245 86231 45279
rect 7537 44973 7571 45007
rect 5421 44905 5455 44939
rect 5257 44701 5291 44735
rect 88221 44701 88255 44735
rect 88061 44361 88095 44395
rect 87761 44293 87795 44327
rect 88221 44293 88255 44327
rect 88061 43341 88095 43375
rect 5257 43205 5291 43239
rect 5421 43205 5455 43239
rect 87761 43205 87795 43239
rect 88221 43205 88255 43239
rect 5421 42729 5455 42763
rect 87945 42729 87979 42763
rect 88221 42729 88255 42763
rect 88061 42593 88095 42627
rect 5257 42525 5291 42559
rect 5257 41641 5291 41675
rect 5421 41641 5455 41675
rect 88061 41641 88095 41675
rect 88221 41641 88255 41675
rect 87945 41573 87979 41607
rect 5421 40553 5455 40587
rect 87945 40485 87979 40519
rect 88221 40485 88255 40519
rect 5257 40417 5291 40451
rect 88221 40077 88255 40111
rect 5421 39465 5455 39499
rect 87853 39465 87887 39499
rect 88221 39465 88255 39499
rect 88057 39329 88091 39363
rect 5257 39261 5291 39295
rect 88057 37901 88091 37935
rect 5257 37765 5291 37799
rect 5421 37765 5455 37799
rect 87761 37765 87795 37799
rect 88221 37765 88255 37799
rect 5421 37289 5455 37323
rect 87945 37289 87979 37323
rect 88221 37289 88255 37323
rect 88062 37153 88096 37187
rect 5257 37085 5291 37119
rect 5421 36201 5455 36235
rect 87945 36201 87979 36235
rect 88221 36201 88255 36235
rect 5257 36133 5291 36167
rect 88062 36133 88096 36167
rect 5421 35113 5455 35147
rect 87945 35113 87979 35147
rect 88221 35113 88255 35147
rect 5257 35045 5291 35079
rect 88062 34977 88096 35011
rect 5421 34025 5455 34059
rect 87945 34025 87979 34059
rect 88221 34025 88255 34059
rect 88061 33889 88095 33923
rect 5257 33821 5291 33855
rect 88062 32461 88096 32495
rect 5257 32325 5291 32359
rect 5421 32325 5455 32359
rect 87761 32325 87795 32359
rect 88221 32325 88255 32359
rect 5421 31849 5455 31883
rect 87945 31849 87979 31883
rect 88221 31849 88255 31883
rect 88061 31713 88095 31747
rect 5257 31645 5291 31679
rect 5421 30761 5455 30795
rect 87945 30761 87979 30795
rect 88221 30761 88255 30795
rect 5257 30625 5291 30659
rect 88062 30625 88096 30659
rect 5173 29673 5207 29707
rect 5513 29673 5547 29707
rect 87969 29673 88003 29707
rect 5375 29537 5409 29571
rect 88175 29469 88209 29503
rect 5173 28585 5207 28619
rect 5513 28585 5547 28619
rect 87969 28585 88003 28619
rect 5375 28449 5409 28483
rect 88175 28381 88209 28415
rect 5375 27021 5409 27055
rect 5173 26885 5207 26919
rect 5513 26885 5547 26919
rect 87969 26885 88003 26919
rect 88175 26749 88209 26783
rect 5173 26409 5207 26443
rect 5513 26409 5547 26443
rect 87969 26409 88003 26443
rect 5375 26273 5409 26307
rect 88175 26205 88209 26239
rect 5173 25321 5207 25355
rect 5513 25321 5547 25355
rect 87969 25321 88003 25355
rect 5375 25117 5409 25151
rect 88175 25117 88209 25151
rect 5173 24233 5207 24267
rect 5513 24233 5547 24267
rect 87969 24233 88003 24267
rect 5375 24097 5409 24131
rect 88175 24097 88209 24131
rect 5173 23145 5207 23179
rect 5513 23145 5547 23179
rect 87969 23145 88003 23179
rect 5375 23009 5409 23043
rect 88175 22941 88209 22975
rect 5375 21581 5409 21615
rect 5173 21445 5207 21479
rect 5513 21445 5547 21479
rect 87969 21445 88003 21479
rect 88175 21309 88209 21343
rect 5375 21037 5409 21071
rect 88175 21037 88209 21071
rect 5173 20969 5207 21003
rect 5513 20969 5547 21003
rect 87969 20969 88003 21003
rect 5173 19881 5207 19915
rect 5513 19881 5547 19915
rect 87969 19881 88003 19915
rect 5375 19745 5409 19779
rect 88175 19677 88209 19711
rect 5173 18793 5207 18827
rect 5513 18793 5547 18827
rect 87969 18793 88003 18827
rect 5375 18657 5409 18691
rect 88175 18657 88209 18691
rect 5173 17705 5207 17739
rect 5513 17705 5547 17739
rect 87969 17705 88003 17739
rect 5375 17569 5409 17603
rect 88175 17501 88209 17535
rect 5375 16141 5409 16175
rect 5173 16005 5207 16039
rect 5513 16005 5547 16039
rect 87969 16005 88003 16039
rect 88175 15869 88209 15903
rect 5375 15597 5409 15631
rect 88175 15597 88209 15631
rect 5173 15529 5207 15563
rect 5513 15529 5547 15563
rect 87969 15529 88003 15563
rect 87485 14985 87519 15019
rect 88221 14985 88255 15019
rect 87808 14917 87842 14951
rect 88037 14781 88071 14815
rect 85645 14237 85679 14271
rect 85645 13421 85679 13455
rect 87669 13421 87703 13455
rect 88226 13344 88260 13378
rect 87945 13285 87979 13319
rect 88221 12877 88255 12911
rect 87808 12741 87842 12775
rect 87485 12673 87519 12707
rect 88037 12673 88071 12707
rect 85645 12333 85679 12367
rect 88129 12333 88163 12367
rect 85645 11245 85679 11279
rect 87761 10565 87795 10599
rect 88221 10565 88255 10599
rect 88061 10497 88095 10531
rect 45441 7437 45475 7471
rect 45625 7437 45659 7471
rect 45809 7437 45843 7471
rect 45993 7437 46027 7471
rect 30745 5261 30779 5295
rect 31595 5261 31629 5295
rect 32678 5261 32712 5295
rect 33966 5261 34000 5295
rect 34815 5261 34849 5295
rect 35907 5261 35941 5295
rect 37186 5261 37220 5295
rect 38474 5261 38508 5295
rect 39323 5261 39357 5295
rect 40406 5261 40440 5295
rect 41693 5261 41727 5295
rect 42543 5261 42577 5295
rect 43635 5261 43669 5295
rect 44913 5261 44947 5295
rect 68097 5261 68131 5295
rect 68947 5261 68981 5295
rect 70030 5261 70064 5295
rect 71318 5261 71352 5295
rect 72606 5261 72640 5295
rect 73455 5261 73489 5295
rect 74538 5261 74572 5295
rect 75826 5261 75860 5295
rect 76675 5261 76709 5295
rect 77758 5261 77792 5295
rect 79045 5261 79079 5295
rect 80333 5261 80367 5295
rect 81183 5261 81217 5295
rect 15289 5125 15323 5159
rect 16185 5125 16219 5159
rect 17221 5125 17255 5159
rect 18509 5125 18543 5159
rect 19405 5125 19439 5159
rect 20478 5125 20512 5159
rect 21729 5125 21763 5159
rect 23017 5125 23051 5159
rect 23913 5125 23947 5159
rect 24949 5125 24983 5159
rect 26237 5125 26271 5159
rect 27133 5125 27167 5159
rect 28206 5125 28240 5159
rect 29457 5125 29491 5159
rect 30905 5125 30939 5159
rect 31089 5125 31123 5159
rect 31393 5125 31427 5159
rect 31733 5125 31767 5159
rect 32837 5125 32871 5159
rect 33021 5125 33055 5159
rect 34125 5125 34159 5159
rect 34309 5125 34343 5159
rect 34613 5125 34647 5159
rect 34953 5125 34987 5159
rect 36057 5125 36091 5159
rect 36241 5125 36275 5159
rect 37345 5125 37379 5159
rect 37529 5125 37563 5159
rect 38633 5125 38667 5159
rect 38817 5125 38851 5159
rect 39121 5125 39155 5159
rect 39461 5125 39495 5159
rect 40565 5125 40599 5159
rect 40749 5125 40783 5159
rect 41853 5125 41887 5159
rect 42037 5125 42071 5159
rect 42341 5125 42375 5159
rect 42681 5125 42715 5159
rect 43785 5125 43819 5159
rect 43969 5125 44003 5159
rect 45073 5125 45107 5159
rect 45257 5125 45291 5159
rect 52641 5125 52675 5159
rect 53537 5125 53571 5159
rect 54573 5125 54607 5159
rect 55861 5125 55895 5159
rect 57149 5125 57183 5159
rect 58045 5125 58079 5159
rect 59081 5125 59115 5159
rect 60369 5125 60403 5159
rect 61265 5125 61299 5159
rect 62338 5125 62372 5159
rect 63589 5125 63623 5159
rect 64877 5125 64911 5159
rect 65773 5125 65807 5159
rect 66809 5125 66843 5159
rect 68257 5125 68291 5159
rect 68441 5125 68475 5159
rect 68745 5125 68779 5159
rect 69085 5125 69119 5159
rect 70189 5125 70223 5159
rect 70373 5125 70407 5159
rect 71477 5125 71511 5159
rect 71661 5125 71695 5159
rect 72765 5125 72799 5159
rect 72949 5125 72983 5159
rect 73253 5125 73287 5159
rect 73593 5125 73627 5159
rect 74697 5125 74731 5159
rect 74881 5125 74915 5159
rect 75985 5125 76019 5159
rect 76169 5125 76203 5159
rect 76473 5125 76507 5159
rect 76813 5125 76847 5159
rect 77917 5125 77951 5159
rect 78101 5125 78135 5159
rect 79205 5125 79239 5159
rect 79389 5125 79423 5159
rect 80493 5125 80527 5159
rect 80677 5125 80711 5159
rect 80981 5125 81015 5159
rect 81321 5125 81355 5159
rect 15495 4989 15529 5023
rect 16021 4989 16055 5023
rect 17427 4989 17461 5023
rect 18715 4989 18749 5023
rect 19241 4989 19275 5023
rect 20647 4989 20681 5023
rect 21935 4989 21969 5023
rect 23223 4989 23257 5023
rect 23749 4989 23783 5023
rect 25155 4989 25189 5023
rect 26443 4989 26477 5023
rect 26969 4989 27003 5023
rect 28375 4989 28409 5023
rect 29663 4989 29697 5023
rect 52847 4989 52881 5023
rect 53373 4989 53407 5023
rect 54779 4989 54813 5023
rect 56067 4989 56101 5023
rect 57355 4989 57389 5023
rect 57881 4989 57915 5023
rect 59287 4989 59321 5023
rect 60575 4989 60609 5023
rect 61101 4989 61135 5023
rect 62507 4989 62541 5023
rect 63795 4989 63829 5023
rect 65083 4989 65117 5023
rect 65609 4989 65643 5023
rect 67015 4989 67049 5023
<< metal1 >>
rect 36502 87668 36508 87720
rect 36560 87708 36566 87720
rect 37514 87708 37520 87720
rect 36560 87680 37520 87708
rect 36560 87668 36566 87680
rect 37514 87668 37520 87680
rect 37572 87668 37578 87720
rect 4876 87610 88596 87632
rect 4876 87558 18382 87610
rect 18434 87558 18446 87610
rect 18498 87558 18510 87610
rect 18562 87558 18574 87610
rect 18626 87558 18638 87610
rect 18690 87558 36782 87610
rect 36834 87558 36846 87610
rect 36898 87558 36910 87610
rect 36962 87558 36974 87610
rect 37026 87558 37038 87610
rect 37090 87558 55182 87610
rect 55234 87558 55246 87610
rect 55298 87558 55310 87610
rect 55362 87558 55374 87610
rect 55426 87558 55438 87610
rect 55490 87558 73582 87610
rect 73634 87558 73646 87610
rect 73698 87558 73710 87610
rect 73762 87558 73774 87610
rect 73826 87558 73838 87610
rect 73890 87558 88596 87610
rect 4876 87536 88596 87558
rect 16541 87439 16599 87445
rect 16541 87436 16553 87439
rect 15728 87408 16553 87436
rect 15250 87328 15256 87380
rect 15308 87377 15314 87380
rect 15308 87371 15335 87377
rect 15323 87368 15335 87371
rect 15728 87368 15756 87408
rect 16541 87405 16553 87408
rect 16587 87405 16599 87439
rect 16541 87399 16599 87405
rect 34570 87396 34576 87448
rect 34628 87436 34634 87448
rect 34685 87439 34743 87445
rect 34685 87436 34697 87439
rect 34628 87408 34697 87436
rect 34628 87396 34634 87408
rect 34685 87405 34697 87408
rect 34731 87405 34743 87439
rect 34685 87399 34743 87405
rect 37146 87396 37152 87448
rect 37204 87436 37210 87448
rect 37747 87439 37805 87445
rect 37747 87436 37759 87439
rect 37204 87408 37759 87436
rect 37204 87396 37210 87408
rect 37747 87405 37759 87408
rect 37793 87405 37805 87439
rect 37747 87399 37805 87405
rect 39078 87396 39084 87448
rect 39136 87436 39142 87448
rect 39679 87439 39737 87445
rect 39679 87436 39691 87439
rect 39136 87408 39691 87436
rect 39136 87396 39142 87408
rect 39679 87405 39691 87408
rect 39725 87405 39737 87439
rect 39679 87399 39737 87405
rect 41010 87396 41016 87448
rect 41068 87436 41074 87448
rect 41125 87439 41183 87445
rect 41125 87436 41137 87439
rect 41068 87408 41137 87436
rect 41068 87396 41074 87408
rect 41125 87405 41137 87408
rect 41171 87405 41183 87439
rect 41125 87399 41183 87405
rect 42298 87396 42304 87448
rect 42356 87436 42362 87448
rect 42413 87439 42471 87445
rect 42413 87436 42425 87439
rect 42356 87408 42425 87436
rect 42356 87396 42362 87408
rect 42413 87405 42425 87408
rect 42459 87405 42471 87439
rect 42413 87399 42471 87405
rect 44230 87396 44236 87448
rect 44288 87436 44294 87448
rect 44345 87439 44403 87445
rect 44345 87436 44357 87439
rect 44288 87408 44357 87436
rect 44288 87396 44294 87408
rect 44345 87405 44357 87408
rect 44391 87405 44403 87439
rect 54169 87439 54227 87445
rect 54169 87436 54181 87439
rect 44345 87399 44403 87405
rect 53172 87408 54181 87436
rect 15323 87340 15756 87368
rect 15323 87337 15335 87340
rect 15308 87331 15335 87337
rect 15308 87328 15314 87331
rect 15894 87328 15900 87380
rect 15952 87368 15958 87380
rect 16357 87371 16415 87377
rect 16357 87368 16369 87371
rect 15952 87340 16369 87368
rect 15952 87328 15958 87340
rect 16357 87337 16369 87340
rect 16403 87368 16415 87371
rect 16725 87371 16783 87377
rect 16725 87368 16737 87371
rect 16403 87340 16737 87368
rect 16403 87337 16415 87340
rect 16357 87331 16415 87337
rect 16725 87337 16737 87340
rect 16771 87337 16783 87371
rect 16725 87331 16783 87337
rect 17182 87328 17188 87380
rect 17240 87368 17246 87380
rect 17369 87371 17427 87377
rect 17369 87368 17381 87371
rect 17240 87340 17381 87368
rect 17240 87328 17246 87340
rect 17369 87337 17381 87340
rect 17415 87368 17427 87371
rect 17553 87371 17611 87377
rect 17553 87368 17565 87371
rect 17415 87340 17565 87368
rect 17415 87337 17427 87340
rect 17369 87331 17427 87337
rect 17553 87337 17565 87340
rect 17599 87337 17611 87371
rect 17553 87331 17611 87337
rect 18657 87371 18715 87377
rect 18657 87337 18669 87371
rect 18703 87368 18715 87371
rect 18746 87368 18752 87380
rect 18703 87340 18752 87368
rect 18703 87337 18715 87340
rect 18657 87331 18715 87337
rect 18746 87328 18752 87340
rect 18804 87368 18810 87380
rect 18841 87371 18899 87377
rect 18841 87368 18853 87371
rect 18804 87340 18853 87368
rect 18804 87328 18810 87340
rect 18841 87337 18853 87340
rect 18887 87337 18899 87371
rect 18841 87331 18899 87337
rect 19114 87328 19120 87380
rect 19172 87377 19178 87380
rect 19172 87371 19203 87377
rect 19191 87368 19203 87371
rect 19485 87371 19543 87377
rect 19485 87368 19497 87371
rect 19191 87340 19497 87368
rect 19191 87337 19203 87340
rect 19172 87331 19203 87337
rect 19485 87337 19497 87340
rect 19531 87337 19543 87371
rect 19485 87331 19543 87337
rect 19172 87328 19178 87331
rect 20402 87328 20408 87380
rect 20460 87368 20466 87380
rect 20589 87371 20647 87377
rect 20589 87368 20601 87371
rect 20460 87340 20601 87368
rect 20460 87328 20466 87340
rect 20589 87337 20601 87340
rect 20635 87368 20647 87371
rect 20773 87371 20831 87377
rect 20773 87368 20785 87371
rect 20635 87340 20785 87368
rect 20635 87337 20647 87340
rect 20589 87331 20647 87337
rect 20773 87337 20785 87340
rect 20819 87337 20831 87371
rect 20773 87331 20831 87337
rect 21690 87328 21696 87380
rect 21748 87368 21754 87380
rect 21877 87371 21935 87377
rect 21877 87368 21889 87371
rect 21748 87340 21889 87368
rect 21748 87328 21754 87340
rect 21877 87337 21889 87340
rect 21923 87368 21935 87371
rect 22061 87371 22119 87377
rect 22061 87368 22073 87371
rect 21923 87340 22073 87368
rect 21923 87337 21935 87340
rect 21877 87331 21935 87337
rect 22061 87337 22073 87340
rect 22107 87337 22119 87371
rect 22061 87331 22119 87337
rect 22978 87328 22984 87380
rect 23036 87368 23042 87380
rect 23165 87371 23223 87377
rect 23165 87368 23177 87371
rect 23036 87340 23177 87368
rect 23036 87328 23042 87340
rect 23165 87337 23177 87340
rect 23211 87368 23223 87371
rect 23349 87371 23407 87377
rect 23349 87368 23361 87371
rect 23211 87340 23361 87368
rect 23211 87337 23223 87340
rect 23165 87331 23223 87337
rect 23349 87337 23361 87340
rect 23395 87337 23407 87371
rect 23349 87331 23407 87337
rect 23622 87328 23628 87380
rect 23680 87377 23686 87380
rect 23680 87371 23711 87377
rect 23699 87368 23711 87371
rect 23993 87371 24051 87377
rect 23993 87368 24005 87371
rect 23699 87340 24005 87368
rect 23699 87337 23711 87340
rect 23680 87331 23711 87337
rect 23993 87337 24005 87340
rect 24039 87337 24051 87371
rect 23993 87331 24051 87337
rect 23680 87328 23686 87331
rect 24910 87328 24916 87380
rect 24968 87368 24974 87380
rect 25097 87371 25155 87377
rect 25097 87368 25109 87371
rect 24968 87340 25109 87368
rect 24968 87328 24974 87340
rect 25097 87337 25109 87340
rect 25143 87368 25155 87371
rect 25281 87371 25339 87377
rect 25281 87368 25293 87371
rect 25143 87340 25293 87368
rect 25143 87337 25155 87340
rect 25097 87331 25155 87337
rect 25281 87337 25293 87340
rect 25327 87337 25339 87371
rect 25281 87331 25339 87337
rect 26198 87328 26204 87380
rect 26256 87368 26262 87380
rect 26385 87371 26443 87377
rect 26385 87368 26397 87371
rect 26256 87340 26397 87368
rect 26256 87328 26262 87340
rect 26385 87337 26397 87340
rect 26431 87368 26443 87371
rect 26569 87371 26627 87377
rect 26569 87368 26581 87371
rect 26431 87340 26581 87368
rect 26431 87337 26443 87340
rect 26385 87331 26443 87337
rect 26569 87337 26581 87340
rect 26615 87337 26627 87371
rect 26569 87331 26627 87337
rect 26842 87328 26848 87380
rect 26900 87377 26906 87380
rect 26900 87371 26931 87377
rect 26919 87368 26931 87371
rect 27213 87371 27271 87377
rect 27213 87368 27225 87371
rect 26919 87340 27225 87368
rect 26919 87337 26931 87340
rect 26900 87331 26931 87337
rect 27213 87337 27225 87340
rect 27259 87337 27271 87371
rect 27213 87331 27271 87337
rect 26900 87328 26906 87331
rect 28130 87328 28136 87380
rect 28188 87368 28194 87380
rect 28317 87371 28375 87377
rect 28317 87368 28329 87371
rect 28188 87340 28329 87368
rect 28188 87328 28194 87340
rect 28317 87337 28329 87340
rect 28363 87368 28375 87371
rect 28501 87371 28559 87377
rect 28501 87368 28513 87371
rect 28363 87340 28513 87368
rect 28363 87337 28375 87340
rect 28317 87331 28375 87337
rect 28501 87337 28513 87340
rect 28547 87337 28559 87371
rect 28501 87331 28559 87337
rect 29418 87328 29424 87380
rect 29476 87368 29482 87380
rect 29605 87371 29663 87377
rect 29605 87368 29617 87371
rect 29476 87340 29617 87368
rect 29476 87328 29482 87340
rect 29605 87337 29617 87340
rect 29651 87368 29663 87371
rect 29789 87371 29847 87377
rect 29789 87368 29801 87371
rect 29651 87340 29801 87368
rect 29651 87337 29663 87340
rect 29605 87331 29663 87337
rect 29789 87337 29801 87340
rect 29835 87337 29847 87371
rect 29789 87331 29847 87337
rect 30614 87328 30620 87380
rect 30672 87368 30678 87380
rect 30733 87371 30791 87377
rect 30733 87368 30745 87371
rect 30672 87340 30745 87368
rect 30672 87328 30678 87340
rect 30733 87337 30745 87340
rect 30779 87337 30791 87371
rect 30733 87331 30791 87337
rect 31534 87328 31540 87380
rect 31592 87368 31598 87380
rect 31629 87371 31687 87377
rect 31629 87368 31641 87371
rect 31592 87340 31641 87368
rect 31592 87328 31598 87340
rect 31629 87337 31641 87340
rect 31675 87337 31687 87371
rect 31629 87331 31687 87337
rect 32638 87328 32644 87380
rect 32696 87377 32702 87380
rect 32696 87371 32723 87377
rect 32711 87337 32723 87371
rect 32696 87331 32723 87337
rect 32696 87328 32702 87331
rect 33742 87328 33748 87380
rect 33800 87368 33806 87380
rect 33953 87371 34011 87377
rect 33953 87368 33965 87371
rect 33800 87340 33965 87368
rect 33800 87328 33806 87340
rect 33953 87337 33965 87340
rect 33999 87337 34011 87371
rect 33953 87331 34011 87337
rect 34846 87328 34852 87380
rect 34904 87328 34910 87380
rect 35950 87377 35956 87380
rect 35922 87371 35956 87377
rect 35922 87337 35934 87371
rect 35922 87331 35956 87337
rect 35950 87328 35956 87331
rect 36008 87328 36014 87380
rect 37422 87328 37428 87380
rect 37480 87377 37486 87380
rect 37606 87377 37612 87380
rect 37480 87371 37502 87377
rect 37490 87337 37502 87371
rect 37480 87331 37502 87337
rect 37578 87371 37612 87377
rect 37578 87337 37590 87371
rect 37578 87331 37612 87337
rect 37480 87328 37486 87331
rect 37606 87328 37612 87331
rect 37664 87328 37670 87380
rect 38038 87371 38096 87377
rect 38038 87337 38050 87371
rect 38084 87368 38096 87371
rect 38158 87368 38164 87380
rect 38084 87340 38164 87368
rect 38084 87337 38096 87340
rect 38038 87331 38096 87337
rect 38158 87328 38164 87340
rect 38216 87328 38222 87380
rect 38434 87328 38440 87380
rect 38492 87377 38498 87380
rect 38492 87371 38519 87377
rect 38507 87337 38519 87371
rect 38492 87331 38519 87337
rect 38492 87328 38498 87331
rect 39262 87328 39268 87380
rect 39320 87368 39326 87380
rect 39473 87371 39531 87377
rect 39473 87368 39485 87371
rect 39320 87340 39485 87368
rect 39320 87328 39326 87340
rect 39473 87337 39485 87340
rect 39519 87337 39531 87371
rect 39473 87331 39531 87337
rect 40366 87328 40372 87380
rect 40424 87377 40430 87380
rect 40424 87371 40451 87377
rect 40439 87337 40451 87371
rect 40424 87331 40451 87337
rect 41289 87371 41347 87377
rect 41289 87337 41301 87371
rect 41335 87368 41347 87371
rect 41470 87368 41476 87380
rect 41335 87340 41476 87368
rect 41335 87337 41347 87340
rect 41289 87331 41347 87337
rect 40424 87328 40430 87331
rect 41470 87328 41476 87340
rect 41528 87328 41534 87380
rect 41654 87328 41660 87380
rect 41712 87368 41718 87380
rect 41749 87371 41807 87377
rect 41749 87368 41761 87371
rect 41712 87340 41761 87368
rect 41712 87328 41718 87340
rect 41749 87337 41761 87340
rect 41795 87337 41807 87371
rect 41749 87331 41807 87337
rect 42574 87328 42580 87380
rect 42632 87328 42638 87380
rect 42942 87328 42948 87380
rect 43000 87368 43006 87380
rect 43678 87377 43684 87380
rect 43037 87371 43095 87377
rect 43037 87368 43049 87371
rect 43000 87340 43049 87368
rect 43000 87328 43006 87340
rect 43037 87337 43049 87340
rect 43083 87337 43095 87371
rect 43037 87331 43095 87337
rect 43650 87371 43684 87377
rect 43650 87337 43662 87371
rect 43650 87331 43684 87337
rect 43678 87328 43684 87331
rect 43736 87328 43742 87380
rect 44509 87371 44567 87377
rect 44509 87337 44521 87371
rect 44555 87368 44567 87371
rect 44782 87368 44788 87380
rect 44555 87340 44788 87368
rect 44555 87337 44567 87340
rect 44509 87331 44567 87337
rect 44782 87328 44788 87340
rect 44840 87328 44846 87380
rect 44874 87328 44880 87380
rect 44932 87368 44938 87380
rect 44969 87371 45027 87377
rect 44969 87368 44981 87371
rect 44932 87340 44981 87368
rect 44932 87328 44938 87340
rect 44969 87337 44981 87340
rect 45015 87337 45027 87371
rect 44969 87331 45027 87337
rect 45518 87328 45524 87380
rect 45576 87368 45582 87380
rect 45613 87371 45671 87377
rect 45613 87368 45625 87371
rect 45576 87340 45625 87368
rect 45576 87328 45582 87340
rect 45613 87337 45625 87340
rect 45659 87337 45671 87371
rect 45613 87331 45671 87337
rect 46162 87328 46168 87380
rect 46220 87368 46226 87380
rect 46257 87371 46315 87377
rect 46257 87368 46269 87371
rect 46220 87340 46269 87368
rect 46220 87328 46226 87340
rect 46257 87337 46269 87340
rect 46303 87337 46315 87371
rect 46257 87331 46315 87337
rect 46806 87328 46812 87380
rect 46864 87368 46870 87380
rect 46901 87371 46959 87377
rect 46901 87368 46913 87371
rect 46864 87340 46913 87368
rect 46864 87328 46870 87340
rect 46901 87337 46913 87340
rect 46947 87337 46959 87371
rect 46901 87331 46959 87337
rect 47450 87328 47456 87380
rect 47508 87368 47514 87380
rect 47545 87371 47603 87377
rect 47545 87368 47557 87371
rect 47508 87340 47557 87368
rect 47508 87328 47514 87340
rect 47545 87337 47557 87340
rect 47591 87337 47603 87371
rect 47545 87331 47603 87337
rect 48094 87328 48100 87380
rect 48152 87368 48158 87380
rect 48189 87371 48247 87377
rect 48189 87368 48201 87371
rect 48152 87340 48201 87368
rect 48152 87328 48158 87340
rect 48189 87337 48201 87340
rect 48235 87337 48247 87371
rect 48189 87331 48247 87337
rect 48738 87328 48744 87380
rect 48796 87368 48802 87380
rect 48833 87371 48891 87377
rect 48833 87368 48845 87371
rect 48796 87340 48845 87368
rect 48796 87328 48802 87340
rect 48833 87337 48845 87340
rect 48879 87337 48891 87371
rect 48833 87331 48891 87337
rect 49382 87328 49388 87380
rect 49440 87368 49446 87380
rect 49477 87371 49535 87377
rect 49477 87368 49489 87371
rect 49440 87340 49489 87368
rect 49440 87328 49446 87340
rect 49477 87337 49489 87340
rect 49523 87337 49535 87371
rect 49477 87331 49535 87337
rect 50026 87328 50032 87380
rect 50084 87368 50090 87380
rect 50121 87371 50179 87377
rect 50121 87368 50133 87371
rect 50084 87340 50133 87368
rect 50084 87328 50090 87340
rect 50121 87337 50133 87340
rect 50167 87337 50179 87371
rect 50121 87331 50179 87337
rect 52602 87328 52608 87380
rect 52660 87377 52666 87380
rect 52660 87371 52687 87377
rect 52675 87368 52687 87371
rect 53172 87368 53200 87408
rect 54169 87405 54181 87408
rect 54215 87405 54227 87439
rect 54169 87399 54227 87405
rect 68702 87396 68708 87448
rect 68760 87436 68766 87448
rect 68817 87439 68875 87445
rect 68817 87436 68829 87439
rect 68760 87408 68829 87436
rect 68760 87396 68766 87408
rect 68817 87405 68829 87408
rect 68863 87405 68875 87439
rect 68817 87399 68875 87405
rect 76430 87396 76436 87448
rect 76488 87436 76494 87448
rect 76545 87439 76603 87445
rect 76545 87436 76557 87439
rect 76488 87408 76557 87436
rect 76488 87396 76494 87408
rect 76545 87405 76557 87408
rect 76591 87405 76603 87439
rect 76545 87399 76603 87405
rect 52675 87340 53200 87368
rect 52675 87337 52687 87340
rect 52660 87331 52687 87337
rect 52660 87328 52666 87331
rect 53246 87328 53252 87380
rect 53304 87368 53310 87380
rect 53709 87371 53767 87377
rect 53709 87368 53721 87371
rect 53304 87340 53721 87368
rect 53304 87328 53310 87340
rect 53709 87337 53721 87340
rect 53755 87368 53767 87371
rect 53985 87371 54043 87377
rect 53985 87368 53997 87371
rect 53755 87340 53997 87368
rect 53755 87337 53767 87340
rect 53709 87331 53767 87337
rect 53985 87337 53997 87340
rect 54031 87337 54043 87371
rect 53985 87331 54043 87337
rect 54534 87328 54540 87380
rect 54592 87368 54598 87380
rect 54721 87371 54779 87377
rect 54721 87368 54733 87371
rect 54592 87340 54733 87368
rect 54592 87328 54598 87340
rect 54721 87337 54733 87340
rect 54767 87368 54779 87371
rect 54905 87371 54963 87377
rect 54905 87368 54917 87371
rect 54767 87340 54917 87368
rect 54767 87337 54779 87340
rect 54721 87331 54779 87337
rect 54905 87337 54917 87340
rect 54951 87337 54963 87371
rect 54905 87331 54963 87337
rect 55822 87328 55828 87380
rect 55880 87368 55886 87380
rect 56009 87371 56067 87377
rect 56009 87368 56021 87371
rect 55880 87340 56021 87368
rect 55880 87328 55886 87340
rect 56009 87337 56021 87340
rect 56055 87368 56067 87371
rect 56193 87371 56251 87377
rect 56193 87368 56205 87371
rect 56055 87340 56205 87368
rect 56055 87337 56067 87340
rect 56009 87331 56067 87337
rect 56193 87337 56205 87340
rect 56239 87337 56251 87371
rect 56193 87331 56251 87337
rect 57110 87328 57116 87380
rect 57168 87368 57174 87380
rect 57297 87371 57355 87377
rect 57297 87368 57309 87371
rect 57168 87340 57309 87368
rect 57168 87328 57174 87340
rect 57297 87337 57309 87340
rect 57343 87368 57355 87371
rect 57481 87371 57539 87377
rect 57481 87368 57493 87371
rect 57343 87340 57493 87368
rect 57343 87337 57355 87340
rect 57297 87331 57355 87337
rect 57481 87337 57493 87340
rect 57527 87337 57539 87371
rect 57481 87331 57539 87337
rect 57754 87328 57760 87380
rect 57812 87377 57818 87380
rect 57812 87371 57843 87377
rect 57831 87368 57843 87371
rect 58125 87371 58183 87377
rect 58125 87368 58137 87371
rect 57831 87340 58137 87368
rect 57831 87337 57843 87340
rect 57812 87331 57843 87337
rect 58125 87337 58137 87340
rect 58171 87337 58183 87371
rect 58125 87331 58183 87337
rect 57812 87328 57818 87331
rect 59042 87328 59048 87380
rect 59100 87368 59106 87380
rect 59229 87371 59287 87377
rect 59229 87368 59241 87371
rect 59100 87340 59241 87368
rect 59100 87328 59106 87340
rect 59229 87337 59241 87340
rect 59275 87368 59287 87371
rect 59413 87371 59471 87377
rect 59413 87368 59425 87371
rect 59275 87340 59425 87368
rect 59275 87337 59287 87340
rect 59229 87331 59287 87337
rect 59413 87337 59425 87340
rect 59459 87337 59471 87371
rect 59413 87331 59471 87337
rect 60330 87328 60336 87380
rect 60388 87368 60394 87380
rect 60517 87371 60575 87377
rect 60517 87368 60529 87371
rect 60388 87340 60529 87368
rect 60388 87328 60394 87340
rect 60517 87337 60529 87340
rect 60563 87368 60575 87371
rect 60701 87371 60759 87377
rect 60701 87368 60713 87371
rect 60563 87340 60713 87368
rect 60563 87337 60575 87340
rect 60517 87331 60575 87337
rect 60701 87337 60713 87340
rect 60747 87337 60759 87371
rect 60701 87331 60759 87337
rect 60974 87328 60980 87380
rect 61032 87377 61038 87380
rect 61032 87371 61063 87377
rect 61051 87368 61063 87371
rect 61345 87371 61403 87377
rect 61345 87368 61357 87371
rect 61051 87340 61357 87368
rect 61051 87337 61063 87340
rect 61032 87331 61063 87337
rect 61345 87337 61357 87340
rect 61391 87337 61403 87371
rect 61345 87331 61403 87337
rect 61032 87328 61038 87331
rect 62262 87328 62268 87380
rect 62320 87368 62326 87380
rect 62449 87371 62507 87377
rect 62449 87368 62461 87371
rect 62320 87340 62461 87368
rect 62320 87328 62326 87340
rect 62449 87337 62461 87340
rect 62495 87368 62507 87371
rect 62633 87371 62691 87377
rect 62633 87368 62645 87371
rect 62495 87340 62645 87368
rect 62495 87337 62507 87340
rect 62449 87331 62507 87337
rect 62633 87337 62645 87340
rect 62679 87337 62691 87371
rect 62633 87331 62691 87337
rect 63550 87328 63556 87380
rect 63608 87368 63614 87380
rect 63737 87371 63795 87377
rect 63737 87368 63749 87371
rect 63608 87340 63749 87368
rect 63608 87328 63614 87340
rect 63737 87337 63749 87340
rect 63783 87368 63795 87371
rect 63921 87371 63979 87377
rect 63921 87368 63933 87371
rect 63783 87340 63933 87368
rect 63783 87337 63795 87340
rect 63737 87331 63795 87337
rect 63921 87337 63933 87340
rect 63967 87337 63979 87371
rect 63921 87331 63979 87337
rect 64838 87328 64844 87380
rect 64896 87368 64902 87380
rect 65025 87371 65083 87377
rect 65025 87368 65037 87371
rect 64896 87340 65037 87368
rect 64896 87328 64902 87340
rect 65025 87337 65037 87340
rect 65071 87368 65083 87371
rect 65209 87371 65267 87377
rect 65209 87368 65221 87371
rect 65071 87340 65221 87368
rect 65071 87337 65083 87340
rect 65025 87331 65083 87337
rect 65209 87337 65221 87340
rect 65255 87337 65267 87371
rect 65209 87331 65267 87337
rect 65482 87328 65488 87380
rect 65540 87377 65546 87380
rect 65540 87371 65571 87377
rect 65559 87368 65571 87371
rect 65853 87371 65911 87377
rect 65853 87368 65865 87371
rect 65559 87340 65865 87368
rect 65559 87337 65571 87340
rect 65540 87331 65571 87337
rect 65853 87337 65865 87340
rect 65899 87337 65911 87371
rect 65853 87331 65911 87337
rect 65540 87328 65546 87331
rect 66770 87328 66776 87380
rect 66828 87368 66834 87380
rect 66957 87371 67015 87377
rect 66957 87368 66969 87371
rect 66828 87340 66969 87368
rect 66828 87328 66834 87340
rect 66957 87337 66969 87340
rect 67003 87368 67015 87371
rect 67141 87371 67199 87377
rect 67141 87368 67153 87371
rect 67003 87340 67153 87368
rect 67003 87337 67015 87340
rect 66957 87331 67015 87337
rect 67141 87337 67153 87340
rect 67187 87337 67199 87371
rect 67141 87331 67199 87337
rect 67874 87328 67880 87380
rect 67932 87368 67938 87380
rect 68085 87371 68143 87377
rect 68085 87368 68097 87371
rect 67932 87340 68097 87368
rect 67932 87328 67938 87340
rect 68085 87337 68097 87340
rect 68131 87337 68143 87371
rect 68085 87331 68143 87337
rect 68978 87328 68984 87380
rect 69036 87328 69042 87380
rect 69990 87328 69996 87380
rect 70048 87377 70054 87380
rect 70048 87371 70075 87377
rect 70063 87337 70075 87371
rect 70048 87331 70075 87337
rect 70048 87328 70054 87331
rect 71186 87328 71192 87380
rect 71244 87368 71250 87380
rect 71305 87371 71363 87377
rect 71305 87368 71317 87371
rect 71244 87340 71317 87368
rect 71244 87328 71250 87340
rect 71305 87337 71317 87340
rect 71351 87337 71363 87371
rect 71305 87331 71363 87337
rect 72290 87328 72296 87380
rect 72348 87368 72354 87380
rect 72593 87371 72651 87377
rect 72593 87368 72605 87371
rect 72348 87340 72605 87368
rect 72348 87328 72354 87340
rect 72593 87337 72605 87340
rect 72639 87337 72651 87371
rect 72593 87331 72651 87337
rect 73394 87328 73400 87380
rect 73452 87368 73458 87380
rect 73489 87371 73547 87377
rect 73489 87368 73501 87371
rect 73452 87340 73501 87368
rect 73452 87328 73458 87340
rect 73489 87337 73501 87340
rect 73535 87337 73547 87371
rect 73489 87331 73547 87337
rect 74498 87328 74504 87380
rect 74556 87377 74562 87380
rect 74556 87371 74583 87377
rect 74571 87337 74583 87371
rect 74556 87331 74583 87337
rect 74556 87328 74562 87331
rect 75602 87328 75608 87380
rect 75660 87368 75666 87380
rect 75813 87371 75871 87377
rect 75813 87368 75825 87371
rect 75660 87340 75825 87368
rect 75660 87328 75666 87340
rect 75813 87337 75825 87340
rect 75859 87337 75871 87371
rect 75813 87331 75871 87337
rect 76706 87328 76712 87380
rect 76764 87328 76770 87380
rect 77718 87328 77724 87380
rect 77776 87377 77782 87380
rect 77776 87371 77803 87377
rect 77791 87337 77803 87371
rect 77776 87331 77803 87337
rect 77776 87328 77782 87331
rect 78914 87328 78920 87380
rect 78972 87368 78978 87380
rect 80386 87377 80392 87380
rect 79033 87371 79091 87377
rect 79033 87368 79045 87371
rect 78972 87340 79045 87368
rect 78972 87328 78978 87340
rect 79033 87337 79045 87340
rect 79079 87337 79091 87371
rect 79033 87331 79091 87337
rect 80358 87371 80392 87377
rect 80358 87337 80370 87371
rect 80358 87331 80392 87337
rect 80386 87328 80392 87331
rect 80444 87328 80450 87380
rect 81122 87328 81128 87380
rect 81180 87368 81186 87380
rect 81217 87371 81275 87377
rect 81217 87368 81229 87371
rect 81180 87340 81229 87368
rect 81180 87328 81186 87340
rect 81217 87337 81229 87340
rect 81263 87337 81275 87371
rect 81217 87331 81275 87337
rect 82226 87328 82232 87380
rect 82284 87377 82290 87380
rect 82284 87371 82311 87377
rect 82299 87337 82311 87371
rect 82284 87331 82311 87337
rect 82284 87328 82290 87331
rect 36594 87260 36600 87312
rect 36652 87260 36658 87312
rect 39078 87260 39084 87312
rect 39136 87300 39142 87312
rect 39357 87303 39415 87309
rect 39357 87300 39369 87303
rect 39136 87272 39369 87300
rect 39136 87260 39142 87272
rect 39357 87269 39369 87272
rect 39403 87300 39415 87303
rect 39909 87303 39967 87309
rect 39909 87300 39921 87303
rect 39403 87272 39921 87300
rect 39403 87269 39415 87272
rect 39357 87263 39415 87269
rect 39909 87269 39921 87272
rect 39955 87269 39967 87303
rect 39909 87263 39967 87269
rect 15526 87192 15532 87244
rect 15584 87192 15590 87244
rect 16078 87192 16084 87244
rect 16136 87232 16142 87244
rect 16198 87235 16256 87241
rect 16198 87232 16210 87235
rect 16136 87204 16210 87232
rect 16136 87192 16142 87204
rect 16198 87201 16210 87204
rect 16244 87201 16256 87235
rect 16198 87195 16256 87201
rect 17182 87192 17188 87244
rect 17240 87241 17246 87244
rect 17240 87235 17268 87241
rect 17256 87201 17268 87235
rect 17240 87195 17268 87201
rect 17240 87192 17246 87195
rect 18286 87192 18292 87244
rect 18344 87232 18350 87244
rect 19390 87241 19396 87244
rect 18498 87235 18556 87241
rect 18498 87232 18510 87235
rect 18344 87204 18510 87232
rect 18344 87192 18350 87204
rect 18498 87201 18510 87204
rect 18544 87201 18556 87235
rect 18498 87195 18556 87201
rect 19347 87235 19396 87241
rect 19347 87201 19359 87235
rect 19393 87201 19396 87235
rect 19347 87195 19396 87201
rect 19390 87192 19396 87195
rect 19448 87192 19454 87244
rect 20402 87192 20408 87244
rect 20460 87241 20466 87244
rect 20460 87235 20488 87241
rect 20476 87201 20488 87235
rect 20460 87195 20488 87201
rect 20460 87192 20466 87195
rect 21598 87192 21604 87244
rect 21656 87232 21662 87244
rect 21718 87235 21776 87241
rect 21718 87232 21730 87235
rect 21656 87204 21730 87232
rect 21656 87192 21662 87204
rect 21718 87201 21730 87204
rect 21764 87201 21776 87235
rect 21718 87195 21776 87201
rect 22702 87192 22708 87244
rect 22760 87232 22766 87244
rect 23006 87235 23064 87241
rect 23006 87232 23018 87235
rect 22760 87204 23018 87232
rect 22760 87192 22766 87204
rect 23006 87201 23018 87204
rect 23052 87201 23064 87235
rect 23006 87195 23064 87201
rect 23806 87192 23812 87244
rect 23864 87241 23870 87244
rect 23864 87235 23913 87241
rect 23864 87201 23867 87235
rect 23901 87201 23913 87235
rect 23864 87195 23913 87201
rect 23864 87192 23870 87195
rect 24910 87192 24916 87244
rect 24968 87241 24974 87244
rect 24968 87235 24996 87241
rect 24984 87201 24996 87235
rect 24968 87195 24996 87201
rect 24968 87192 24974 87195
rect 26014 87192 26020 87244
rect 26072 87232 26078 87244
rect 27118 87241 27124 87244
rect 26225 87235 26283 87241
rect 26225 87232 26237 87235
rect 26072 87204 26237 87232
rect 26072 87192 26078 87204
rect 26225 87201 26237 87204
rect 26271 87201 26283 87235
rect 26225 87195 26283 87201
rect 27075 87235 27124 87241
rect 27075 87201 27087 87235
rect 27121 87201 27124 87235
rect 27075 87195 27124 87201
rect 27118 87192 27124 87195
rect 27176 87192 27182 87244
rect 28130 87192 28136 87244
rect 28188 87241 28194 87244
rect 28188 87235 28215 87241
rect 28203 87201 28215 87235
rect 28188 87195 28215 87201
rect 28188 87192 28194 87195
rect 29326 87192 29332 87244
rect 29384 87232 29390 87244
rect 29446 87235 29504 87241
rect 29446 87232 29458 87235
rect 29384 87204 29458 87232
rect 29384 87192 29390 87204
rect 29446 87201 29458 87204
rect 29492 87201 29504 87235
rect 29446 87195 29504 87201
rect 30706 87192 30712 87244
rect 30764 87232 30770 87244
rect 30939 87235 30997 87241
rect 30939 87232 30951 87235
rect 30764 87204 30951 87232
rect 30764 87192 30770 87204
rect 30939 87201 30951 87204
rect 30985 87201 30997 87235
rect 30939 87195 30997 87201
rect 31350 87192 31356 87244
rect 31408 87232 31414 87244
rect 31465 87235 31523 87241
rect 31465 87232 31477 87235
rect 31408 87204 31477 87232
rect 31408 87192 31414 87204
rect 31465 87201 31477 87204
rect 31511 87201 31523 87235
rect 31465 87195 31523 87201
rect 32730 87192 32736 87244
rect 32788 87232 32794 87244
rect 32871 87235 32929 87241
rect 32871 87232 32883 87235
rect 32788 87204 32883 87232
rect 32788 87192 32794 87204
rect 32871 87201 32883 87204
rect 32917 87201 32929 87235
rect 32871 87195 32929 87201
rect 33926 87192 33932 87244
rect 33984 87232 33990 87244
rect 34159 87235 34217 87241
rect 34159 87232 34171 87235
rect 33984 87204 34171 87232
rect 33984 87192 33990 87204
rect 34159 87201 34171 87204
rect 34205 87201 34217 87235
rect 34159 87195 34217 87201
rect 35858 87192 35864 87244
rect 35916 87232 35922 87244
rect 36091 87235 36149 87241
rect 36091 87232 36103 87235
rect 35916 87204 36103 87232
rect 35916 87192 35922 87204
rect 36091 87201 36103 87204
rect 36137 87201 36149 87235
rect 36091 87195 36149 87201
rect 38207 87235 38265 87241
rect 38207 87201 38219 87235
rect 38253 87232 38265 87235
rect 38342 87232 38348 87244
rect 38253 87204 38348 87232
rect 38253 87201 38265 87204
rect 38207 87195 38265 87201
rect 38342 87192 38348 87204
rect 38400 87192 38406 87244
rect 40458 87192 40464 87244
rect 40516 87232 40522 87244
rect 40599 87235 40657 87241
rect 40599 87232 40611 87235
rect 40516 87204 40611 87232
rect 40516 87192 40522 87204
rect 40599 87201 40611 87204
rect 40645 87201 40657 87235
rect 40599 87195 40657 87201
rect 43586 87192 43592 87244
rect 43644 87232 43650 87244
rect 43819 87235 43877 87241
rect 43819 87232 43831 87235
rect 43644 87204 43831 87232
rect 43644 87192 43650 87204
rect 43819 87201 43831 87204
rect 43865 87201 43877 87235
rect 43819 87195 43877 87201
rect 52878 87192 52884 87244
rect 52936 87192 52942 87244
rect 53522 87192 53528 87244
rect 53580 87241 53586 87244
rect 53580 87235 53608 87241
rect 53596 87201 53608 87235
rect 53580 87195 53608 87201
rect 53580 87192 53586 87195
rect 54442 87192 54448 87244
rect 54500 87232 54506 87244
rect 54562 87235 54620 87241
rect 54562 87232 54574 87235
rect 54500 87204 54574 87232
rect 54500 87192 54506 87204
rect 54562 87201 54574 87204
rect 54608 87201 54620 87235
rect 54562 87195 54620 87201
rect 55730 87192 55736 87244
rect 55788 87232 55794 87244
rect 55850 87235 55908 87241
rect 55850 87232 55862 87235
rect 55788 87204 55862 87232
rect 55788 87192 55794 87204
rect 55850 87201 55862 87204
rect 55896 87201 55908 87235
rect 55850 87195 55908 87201
rect 56834 87192 56840 87244
rect 56892 87232 56898 87244
rect 57138 87235 57196 87241
rect 57138 87232 57150 87235
rect 56892 87204 57150 87232
rect 56892 87192 56898 87204
rect 57138 87201 57150 87204
rect 57184 87201 57196 87235
rect 57138 87195 57196 87201
rect 57938 87192 57944 87244
rect 57996 87241 58002 87244
rect 57996 87235 58045 87241
rect 57996 87201 57999 87235
rect 58033 87201 58045 87235
rect 57996 87195 58045 87201
rect 57996 87192 58002 87195
rect 59042 87192 59048 87244
rect 59100 87241 59106 87244
rect 59100 87235 59128 87241
rect 59116 87201 59128 87235
rect 59100 87195 59128 87201
rect 59100 87192 59106 87195
rect 60146 87192 60152 87244
rect 60204 87232 60210 87244
rect 60358 87235 60416 87241
rect 60358 87232 60370 87235
rect 60204 87204 60370 87232
rect 60204 87192 60210 87204
rect 60358 87201 60370 87204
rect 60404 87201 60416 87235
rect 60358 87195 60416 87201
rect 61158 87192 61164 87244
rect 61216 87241 61222 87244
rect 61216 87235 61265 87241
rect 61216 87201 61219 87235
rect 61253 87201 61265 87235
rect 61216 87195 61265 87201
rect 62299 87235 62357 87241
rect 62299 87201 62311 87235
rect 62345 87232 62357 87235
rect 62446 87232 62452 87244
rect 62345 87204 62452 87232
rect 62345 87201 62357 87204
rect 62299 87195 62357 87201
rect 61216 87192 61222 87195
rect 62446 87192 62452 87204
rect 62504 87192 62510 87244
rect 63458 87192 63464 87244
rect 63516 87232 63522 87244
rect 63577 87235 63635 87241
rect 63577 87232 63589 87235
rect 63516 87204 63589 87232
rect 63516 87192 63522 87204
rect 63577 87201 63589 87204
rect 63623 87201 63635 87235
rect 63577 87195 63635 87201
rect 64562 87192 64568 87244
rect 64620 87232 64626 87244
rect 64866 87235 64924 87241
rect 64866 87232 64878 87235
rect 64620 87204 64878 87232
rect 64620 87192 64626 87204
rect 64866 87201 64878 87204
rect 64912 87201 64924 87235
rect 64866 87195 64924 87201
rect 65666 87192 65672 87244
rect 65724 87241 65730 87244
rect 65724 87235 65773 87241
rect 65724 87201 65727 87235
rect 65761 87201 65773 87235
rect 65724 87195 65773 87201
rect 65724 87192 65730 87195
rect 66770 87192 66776 87244
rect 66828 87241 66834 87244
rect 66828 87235 66856 87241
rect 66844 87201 66856 87235
rect 66828 87195 66856 87201
rect 66828 87192 66834 87195
rect 68058 87192 68064 87244
rect 68116 87232 68122 87244
rect 68291 87235 68349 87241
rect 68291 87232 68303 87235
rect 68116 87204 68303 87232
rect 68116 87192 68122 87204
rect 68291 87201 68303 87204
rect 68337 87201 68349 87235
rect 68291 87195 68349 87201
rect 70082 87192 70088 87244
rect 70140 87232 70146 87244
rect 70223 87235 70281 87241
rect 70223 87232 70235 87235
rect 70140 87204 70235 87232
rect 70140 87192 70146 87204
rect 70223 87201 70235 87204
rect 70269 87201 70281 87235
rect 70223 87195 70281 87201
rect 71278 87192 71284 87244
rect 71336 87232 71342 87244
rect 71511 87235 71569 87241
rect 71511 87232 71523 87235
rect 71336 87204 71523 87232
rect 71336 87192 71342 87204
rect 71511 87201 71523 87204
rect 71557 87201 71569 87235
rect 71511 87195 71569 87201
rect 72566 87192 72572 87244
rect 72624 87232 72630 87244
rect 72799 87235 72857 87241
rect 72799 87232 72811 87235
rect 72624 87204 72811 87232
rect 72624 87192 72630 87204
rect 72799 87201 72811 87204
rect 72845 87201 72857 87235
rect 72799 87195 72857 87201
rect 73210 87192 73216 87244
rect 73268 87232 73274 87244
rect 73325 87235 73383 87241
rect 73325 87232 73337 87235
rect 73268 87204 73337 87232
rect 73268 87192 73274 87204
rect 73325 87201 73337 87204
rect 73371 87201 73383 87235
rect 73325 87195 73383 87201
rect 74590 87192 74596 87244
rect 74648 87232 74654 87244
rect 74731 87235 74789 87241
rect 74731 87232 74743 87235
rect 74648 87204 74743 87232
rect 74648 87192 74654 87204
rect 74731 87201 74743 87204
rect 74777 87201 74789 87235
rect 74731 87195 74789 87201
rect 75786 87192 75792 87244
rect 75844 87232 75850 87244
rect 76019 87235 76077 87241
rect 76019 87232 76031 87235
rect 75844 87204 76031 87232
rect 75844 87192 75850 87204
rect 76019 87201 76031 87204
rect 76065 87201 76077 87235
rect 76019 87195 76077 87201
rect 77810 87192 77816 87244
rect 77868 87232 77874 87244
rect 77951 87235 78009 87241
rect 77951 87232 77963 87235
rect 77868 87204 77963 87232
rect 77868 87192 77874 87204
rect 77951 87201 77963 87204
rect 77997 87201 78009 87235
rect 77951 87195 78009 87201
rect 79006 87192 79012 87244
rect 79064 87232 79070 87244
rect 79239 87235 79297 87241
rect 79239 87232 79251 87235
rect 79064 87204 79251 87232
rect 79064 87192 79070 87204
rect 79239 87201 79251 87204
rect 79285 87201 79297 87235
rect 79239 87195 79297 87201
rect 80294 87192 80300 87244
rect 80352 87232 80358 87244
rect 80527 87235 80585 87241
rect 80527 87232 80539 87235
rect 80352 87204 80539 87232
rect 80352 87192 80358 87204
rect 80527 87201 80539 87204
rect 80573 87201 80585 87235
rect 80527 87195 80585 87201
rect 80938 87192 80944 87244
rect 80996 87232 81002 87244
rect 81053 87235 81111 87241
rect 81053 87232 81065 87235
rect 80996 87204 81065 87232
rect 80996 87192 81002 87204
rect 81053 87201 81065 87204
rect 81099 87201 81111 87235
rect 81053 87195 81111 87201
rect 82318 87192 82324 87244
rect 82376 87232 82382 87244
rect 82459 87235 82517 87241
rect 82459 87232 82471 87235
rect 82376 87204 82471 87232
rect 82376 87192 82382 87204
rect 82459 87201 82471 87204
rect 82505 87201 82517 87235
rect 82459 87195 82517 87201
rect 4876 87066 88596 87088
rect 4876 87014 17722 87066
rect 17774 87014 17786 87066
rect 17838 87014 17850 87066
rect 17902 87014 17914 87066
rect 17966 87014 17978 87066
rect 18030 87014 36122 87066
rect 36174 87014 36186 87066
rect 36238 87014 36250 87066
rect 36302 87014 36314 87066
rect 36366 87014 36378 87066
rect 36430 87014 54522 87066
rect 54574 87014 54586 87066
rect 54638 87014 54650 87066
rect 54702 87014 54714 87066
rect 54766 87014 54778 87066
rect 54830 87014 72922 87066
rect 72974 87014 72986 87066
rect 73038 87014 73050 87066
rect 73102 87014 73114 87066
rect 73166 87014 73178 87066
rect 73230 87014 88596 87066
rect 4876 86992 88596 87014
rect 37514 86852 37520 86904
rect 37572 86892 37578 86904
rect 37609 86895 37667 86901
rect 37609 86892 37621 86895
rect 37572 86864 37621 86892
rect 37572 86852 37578 86864
rect 37609 86861 37621 86864
rect 37655 86861 37667 86895
rect 37609 86855 37667 86861
rect 37790 86852 37796 86904
rect 37848 86892 37854 86904
rect 38434 86892 38440 86904
rect 37848 86864 38440 86892
rect 37848 86852 37854 86864
rect 38434 86852 38440 86864
rect 38492 86892 38498 86904
rect 38529 86895 38587 86901
rect 38529 86892 38541 86895
rect 38492 86864 38541 86892
rect 38492 86852 38498 86864
rect 38529 86861 38541 86864
rect 38575 86861 38587 86895
rect 38529 86855 38587 86861
rect 36594 86580 36600 86632
rect 36652 86620 36658 86632
rect 37793 86623 37851 86629
rect 37793 86620 37805 86623
rect 36652 86592 37805 86620
rect 36652 86580 36658 86592
rect 37793 86589 37805 86592
rect 37839 86620 37851 86623
rect 46990 86620 46996 86632
rect 37839 86592 46996 86620
rect 37839 86589 37851 86592
rect 37793 86583 37851 86589
rect 46990 86580 46996 86592
rect 47048 86620 47054 86632
rect 50302 86620 50308 86632
rect 47048 86592 50308 86620
rect 47048 86580 47054 86592
rect 50302 86580 50308 86592
rect 50360 86580 50366 86632
rect 4876 86522 88596 86544
rect 4876 86470 18382 86522
rect 18434 86470 18446 86522
rect 18498 86470 18510 86522
rect 18562 86470 18574 86522
rect 18626 86470 18638 86522
rect 18690 86470 36782 86522
rect 36834 86470 36846 86522
rect 36898 86470 36910 86522
rect 36962 86470 36974 86522
rect 37026 86470 37038 86522
rect 37090 86470 55182 86522
rect 55234 86470 55246 86522
rect 55298 86470 55310 86522
rect 55362 86470 55374 86522
rect 55426 86470 55438 86522
rect 55490 86470 73582 86522
rect 73634 86470 73646 86522
rect 73698 86470 73710 86522
rect 73762 86470 73774 86522
rect 73826 86470 73838 86522
rect 73890 86470 88596 86522
rect 4876 86448 88596 86470
rect 4876 85978 88596 86000
rect 4876 85926 17722 85978
rect 17774 85926 17786 85978
rect 17838 85926 17850 85978
rect 17902 85926 17914 85978
rect 17966 85926 17978 85978
rect 18030 85926 36122 85978
rect 36174 85926 36186 85978
rect 36238 85926 36250 85978
rect 36302 85926 36314 85978
rect 36366 85926 36378 85978
rect 36430 85926 54522 85978
rect 54574 85926 54586 85978
rect 54638 85926 54650 85978
rect 54702 85926 54714 85978
rect 54766 85926 54778 85978
rect 54830 85926 72922 85978
rect 72974 85926 72986 85978
rect 73038 85926 73050 85978
rect 73102 85926 73114 85978
rect 73166 85926 73178 85978
rect 73230 85926 88596 85978
rect 4876 85904 88596 85926
rect 4876 85434 88596 85456
rect 4876 85382 18382 85434
rect 18434 85382 18446 85434
rect 18498 85382 18510 85434
rect 18562 85382 18574 85434
rect 18626 85382 18638 85434
rect 18690 85382 36782 85434
rect 36834 85382 36846 85434
rect 36898 85382 36910 85434
rect 36962 85382 36974 85434
rect 37026 85382 37038 85434
rect 37090 85382 55182 85434
rect 55234 85382 55246 85434
rect 55298 85382 55310 85434
rect 55362 85382 55374 85434
rect 55426 85382 55438 85434
rect 55490 85382 73582 85434
rect 73634 85382 73646 85434
rect 73698 85382 73710 85434
rect 73762 85382 73774 85434
rect 73826 85382 73838 85434
rect 73890 85382 88596 85434
rect 4876 85360 88596 85382
rect 4876 84890 88596 84912
rect 4876 84838 5882 84890
rect 5934 84838 5946 84890
rect 5998 84838 6010 84890
rect 6062 84838 6074 84890
rect 6126 84838 6138 84890
rect 6190 84838 17722 84890
rect 17774 84838 17786 84890
rect 17838 84838 17850 84890
rect 17902 84838 17914 84890
rect 17966 84838 17978 84890
rect 18030 84838 36122 84890
rect 36174 84838 36186 84890
rect 36238 84838 36250 84890
rect 36302 84838 36314 84890
rect 36366 84838 36378 84890
rect 36430 84838 54522 84890
rect 54574 84838 54586 84890
rect 54638 84838 54650 84890
rect 54702 84838 54714 84890
rect 54766 84838 54778 84890
rect 54830 84838 72922 84890
rect 72974 84838 72986 84890
rect 73038 84838 73050 84890
rect 73102 84838 73114 84890
rect 73166 84838 73178 84890
rect 73230 84838 86474 84890
rect 86526 84838 86538 84890
rect 86590 84838 86602 84890
rect 86654 84838 86666 84890
rect 86718 84838 86730 84890
rect 86782 84838 88596 84890
rect 4876 84816 88596 84838
rect 45429 84719 45487 84725
rect 45429 84685 45441 84719
rect 45475 84716 45487 84719
rect 46162 84716 46168 84728
rect 45475 84688 46168 84716
rect 45475 84685 45487 84688
rect 45429 84679 45487 84685
rect 46162 84676 46168 84688
rect 46220 84716 46226 84728
rect 46220 84688 50256 84716
rect 46220 84676 46226 84688
rect 12766 84608 12772 84660
rect 12824 84648 12830 84660
rect 12861 84651 12919 84657
rect 12861 84648 12873 84651
rect 12824 84620 12873 84648
rect 12824 84608 12830 84620
rect 12861 84617 12873 84620
rect 12907 84648 12919 84651
rect 36594 84648 36600 84660
rect 12907 84620 36600 84648
rect 12907 84617 12919 84620
rect 12861 84611 12919 84617
rect 36594 84608 36600 84620
rect 36652 84608 36658 84660
rect 39078 84648 39084 84660
rect 38866 84620 39084 84648
rect 11662 84540 11668 84592
rect 11720 84580 11726 84592
rect 11757 84583 11815 84589
rect 11757 84580 11769 84583
rect 11720 84552 11769 84580
rect 11720 84540 11726 84552
rect 11757 84549 11769 84552
rect 11803 84580 11815 84583
rect 38866 84580 38894 84620
rect 39078 84608 39084 84620
rect 39136 84648 39142 84660
rect 49106 84648 49112 84660
rect 39136 84620 49112 84648
rect 39136 84608 39142 84620
rect 49106 84608 49112 84620
rect 49164 84608 49170 84660
rect 50228 84648 50256 84688
rect 50302 84676 50308 84728
rect 50360 84676 50366 84728
rect 51314 84648 51320 84660
rect 50228 84620 51320 84648
rect 51314 84608 51320 84620
rect 51372 84608 51378 84660
rect 11803 84552 38894 84580
rect 45613 84583 45671 84589
rect 11803 84549 11815 84552
rect 11757 84543 11815 84549
rect 45613 84549 45625 84583
rect 45659 84580 45671 84583
rect 46070 84580 46076 84592
rect 45659 84552 46076 84580
rect 45659 84549 45671 84552
rect 45613 84543 45671 84549
rect 46070 84540 46076 84552
rect 46128 84540 46134 84592
rect 7522 84472 7528 84524
rect 7580 84512 7586 84524
rect 28869 84515 28927 84521
rect 28869 84512 28881 84515
rect 7580 84484 28881 84512
rect 7580 84472 7586 84484
rect 28869 84481 28881 84484
rect 28915 84512 28927 84515
rect 30573 84515 30631 84521
rect 28915 84484 29234 84512
rect 28915 84481 28927 84484
rect 28869 84475 28927 84481
rect 10558 84404 10564 84456
rect 10616 84444 10622 84456
rect 10653 84447 10711 84453
rect 10653 84444 10665 84447
rect 10616 84416 10665 84444
rect 10616 84404 10622 84416
rect 10653 84413 10665 84416
rect 10699 84413 10711 84447
rect 10653 84407 10711 84413
rect 13870 84404 13876 84456
rect 13928 84444 13934 84456
rect 13965 84447 14023 84453
rect 13965 84444 13977 84447
rect 13928 84416 13977 84444
rect 13928 84404 13934 84416
rect 13965 84413 13977 84416
rect 14011 84413 14023 84447
rect 29206 84444 29234 84484
rect 30573 84481 30585 84515
rect 30619 84512 30631 84515
rect 31077 84515 31135 84521
rect 31077 84512 31089 84515
rect 30619 84484 31089 84512
rect 30619 84481 30631 84484
rect 30573 84475 30631 84481
rect 31077 84481 31089 84484
rect 31123 84512 31135 84515
rect 39722 84512 39728 84524
rect 31123 84484 39728 84512
rect 31123 84481 31135 84484
rect 31077 84475 31135 84481
rect 39722 84472 39728 84484
rect 39780 84472 39786 84524
rect 41037 84515 41095 84521
rect 41037 84512 41049 84515
rect 40844 84484 41049 84512
rect 40844 84453 40872 84484
rect 41037 84481 41049 84484
rect 41083 84481 41095 84515
rect 41037 84475 41095 84481
rect 42761 84515 42819 84521
rect 42761 84481 42773 84515
rect 42807 84512 42819 84515
rect 42945 84515 43003 84521
rect 42945 84512 42957 84515
rect 42807 84484 42957 84512
rect 42807 84481 42819 84484
rect 42761 84475 42819 84481
rect 42945 84481 42957 84484
rect 42991 84512 43003 84515
rect 42991 84484 48048 84512
rect 42991 84481 43003 84484
rect 42945 84475 43003 84481
rect 48020 84456 48048 84484
rect 30893 84447 30951 84453
rect 30893 84444 30905 84447
rect 29206 84416 30905 84444
rect 13965 84407 14023 84413
rect 30893 84413 30905 84416
rect 30939 84444 30951 84447
rect 40829 84447 40887 84453
rect 40829 84444 40841 84447
rect 30939 84416 40841 84444
rect 30939 84413 30951 84416
rect 30893 84407 30951 84413
rect 40829 84413 40841 84416
rect 40875 84413 40887 84447
rect 40829 84407 40887 84413
rect 45797 84447 45855 84453
rect 45797 84413 45809 84447
rect 45843 84444 45855 84447
rect 45886 84444 45892 84456
rect 45843 84416 45892 84444
rect 45843 84413 45855 84416
rect 45797 84407 45855 84413
rect 45886 84404 45892 84416
rect 45944 84404 45950 84456
rect 45978 84404 45984 84456
rect 46036 84404 46042 84456
rect 48002 84404 48008 84456
rect 48060 84444 48066 84456
rect 48097 84447 48155 84453
rect 48097 84444 48109 84447
rect 48060 84416 48109 84444
rect 48060 84404 48066 84416
rect 48097 84413 48109 84416
rect 48143 84413 48155 84447
rect 48097 84407 48155 84413
rect 49106 84404 49112 84456
rect 49164 84444 49170 84456
rect 49201 84447 49259 84453
rect 49201 84444 49213 84447
rect 49164 84416 49213 84444
rect 49164 84404 49170 84416
rect 49201 84413 49213 84416
rect 49247 84413 49259 84447
rect 49201 84407 49259 84413
rect 51314 84404 51320 84456
rect 51372 84444 51378 84456
rect 51409 84447 51467 84453
rect 51409 84444 51421 84447
rect 51372 84416 51421 84444
rect 51372 84404 51378 84416
rect 51409 84413 51421 84416
rect 51455 84413 51467 84447
rect 51409 84407 51467 84413
rect 4876 84346 88596 84368
rect 4876 84294 6618 84346
rect 6670 84294 6682 84346
rect 6734 84294 6746 84346
rect 6798 84294 6810 84346
rect 6862 84294 6874 84346
rect 6926 84294 18382 84346
rect 18434 84294 18446 84346
rect 18498 84294 18510 84346
rect 18562 84294 18574 84346
rect 18626 84294 18638 84346
rect 18690 84294 36782 84346
rect 36834 84294 36846 84346
rect 36898 84294 36910 84346
rect 36962 84294 36974 84346
rect 37026 84294 37038 84346
rect 37090 84294 55182 84346
rect 55234 84294 55246 84346
rect 55298 84294 55310 84346
rect 55362 84294 55374 84346
rect 55426 84294 55438 84346
rect 55490 84294 73582 84346
rect 73634 84294 73646 84346
rect 73698 84294 73710 84346
rect 73762 84294 73774 84346
rect 73826 84294 73838 84346
rect 73890 84294 87210 84346
rect 87262 84294 87274 84346
rect 87326 84294 87338 84346
rect 87390 84294 87402 84346
rect 87454 84294 87466 84346
rect 87518 84294 88596 84346
rect 4876 84272 88596 84294
rect 4876 83802 7912 83824
rect 4876 83750 5882 83802
rect 5934 83750 5946 83802
rect 5998 83750 6010 83802
rect 6062 83750 6074 83802
rect 6126 83750 6138 83802
rect 6190 83750 7912 83802
rect 4876 83728 7912 83750
rect 85284 83802 88596 83824
rect 85284 83750 86474 83802
rect 86526 83750 86538 83802
rect 86590 83750 86602 83802
rect 86654 83750 86666 83802
rect 86718 83750 86730 83802
rect 86782 83750 88596 83802
rect 85284 83728 88596 83750
rect 4876 83258 7912 83280
rect 4876 83206 6618 83258
rect 6670 83206 6682 83258
rect 6734 83206 6746 83258
rect 6798 83206 6810 83258
rect 6862 83206 6874 83258
rect 6926 83206 7912 83258
rect 4876 83184 7912 83206
rect 85284 83258 88596 83280
rect 85284 83206 87210 83258
rect 87262 83206 87274 83258
rect 87326 83206 87338 83258
rect 87390 83206 87402 83258
rect 87454 83206 87466 83258
rect 87518 83206 88596 83258
rect 85284 83184 88596 83206
rect 13870 83112 13876 83164
rect 13928 83152 13934 83164
rect 83238 83152 83244 83164
rect 13928 83124 83244 83152
rect 13928 83112 13934 83124
rect 83238 83112 83244 83124
rect 83296 83112 83302 83164
rect 9822 83044 9828 83096
rect 9880 83084 9886 83096
rect 12766 83084 12772 83096
rect 9880 83056 12772 83084
rect 9880 83044 9886 83056
rect 12766 83044 12772 83056
rect 12824 83044 12830 83096
rect 14974 82976 14980 83028
rect 15032 83016 15038 83028
rect 15526 83016 15532 83028
rect 15032 82988 15532 83016
rect 15032 82976 15038 82988
rect 15526 82976 15532 82988
rect 15584 82976 15590 83028
rect 37054 82976 37060 83028
rect 37112 83016 37118 83028
rect 37606 83016 37612 83028
rect 37112 82988 37612 83016
rect 37112 82976 37118 82988
rect 37606 82976 37612 82988
rect 37664 82976 37670 83028
rect 4876 82714 7912 82736
rect 4876 82662 5882 82714
rect 5934 82662 5946 82714
rect 5998 82662 6010 82714
rect 6062 82662 6074 82714
rect 6126 82662 6138 82714
rect 6190 82662 7912 82714
rect 4876 82640 7912 82662
rect 85284 82714 88596 82736
rect 85284 82662 86474 82714
rect 86526 82662 86538 82714
rect 86590 82662 86602 82714
rect 86654 82662 86666 82714
rect 86718 82662 86730 82714
rect 86782 82662 88596 82714
rect 85284 82640 88596 82662
rect 7614 82364 7620 82416
rect 7672 82404 7678 82416
rect 11662 82404 11668 82416
rect 7672 82376 11668 82404
rect 7672 82364 7678 82376
rect 11662 82364 11668 82376
rect 11720 82364 11726 82416
rect 7798 82296 7804 82348
rect 7856 82336 7862 82348
rect 10558 82336 10564 82348
rect 7856 82308 10564 82336
rect 7856 82296 7862 82308
rect 10558 82296 10564 82308
rect 10616 82296 10622 82348
rect 52372 82296 52378 82348
rect 52430 82336 52436 82348
rect 52878 82336 52884 82348
rect 52430 82308 52884 82336
rect 52430 82296 52436 82308
rect 52878 82296 52884 82308
rect 52936 82296 52942 82348
rect 79972 82296 79978 82348
rect 80030 82336 80036 82348
rect 80386 82336 80392 82348
rect 80030 82308 80392 82336
rect 80030 82296 80036 82308
rect 80386 82296 80392 82308
rect 80444 82296 80450 82348
rect 4876 82170 7912 82192
rect 4876 82118 6618 82170
rect 6670 82118 6682 82170
rect 6734 82118 6746 82170
rect 6798 82118 6810 82170
rect 6862 82118 6874 82170
rect 6926 82118 7912 82170
rect 4876 82096 7912 82118
rect 85284 82170 88596 82192
rect 85284 82118 87210 82170
rect 87262 82118 87274 82170
rect 87326 82118 87338 82170
rect 87390 82118 87402 82170
rect 87454 82118 87466 82170
rect 87518 82118 88596 82170
rect 85284 82096 88596 82118
rect 4876 81626 7912 81648
rect 4876 81574 5882 81626
rect 5934 81574 5946 81626
rect 5998 81574 6010 81626
rect 6062 81574 6074 81626
rect 6126 81574 6138 81626
rect 6190 81574 7912 81626
rect 4876 81552 7912 81574
rect 85284 81626 88596 81648
rect 85284 81574 86474 81626
rect 86526 81574 86538 81626
rect 86590 81574 86602 81626
rect 86654 81574 86666 81626
rect 86718 81574 86730 81626
rect 86782 81574 88596 81626
rect 85284 81552 88596 81574
rect 4118 81276 4124 81328
rect 4176 81316 4182 81328
rect 5245 81319 5303 81325
rect 5245 81316 5257 81319
rect 4176 81288 5257 81316
rect 4176 81276 4182 81288
rect 5245 81285 5257 81288
rect 5291 81285 5303 81319
rect 5245 81279 5303 81285
rect 5409 81319 5467 81325
rect 5409 81285 5421 81319
rect 5455 81316 5467 81319
rect 8534 81316 8540 81328
rect 5455 81288 8540 81316
rect 5455 81285 5467 81288
rect 5409 81279 5467 81285
rect 8534 81276 8540 81288
rect 8592 81276 8598 81328
rect 87749 81319 87807 81325
rect 87749 81285 87761 81319
rect 87795 81316 87807 81319
rect 88206 81316 88212 81328
rect 87795 81288 88212 81316
rect 87795 81285 87807 81288
rect 87749 81279 87807 81285
rect 88206 81276 88212 81288
rect 88264 81276 88270 81328
rect 84342 81208 84348 81260
rect 84400 81248 84406 81260
rect 88049 81251 88107 81257
rect 88049 81248 88061 81251
rect 84400 81220 88061 81248
rect 84400 81208 84406 81220
rect 88049 81217 88061 81220
rect 88095 81217 88107 81251
rect 88049 81211 88107 81217
rect 4876 81082 7912 81104
rect 4876 81030 6618 81082
rect 6670 81030 6682 81082
rect 6734 81030 6746 81082
rect 6798 81030 6810 81082
rect 6862 81030 6874 81082
rect 6926 81030 7912 81082
rect 4876 81008 7912 81030
rect 85284 81082 88596 81104
rect 85284 81030 87210 81082
rect 87262 81030 87274 81082
rect 87326 81030 87338 81082
rect 87390 81030 87402 81082
rect 87454 81030 87466 81082
rect 87518 81030 88596 81082
rect 85284 81008 88596 81030
rect 4876 80538 7912 80560
rect 4876 80486 5882 80538
rect 5934 80486 5946 80538
rect 5998 80486 6010 80538
rect 6062 80486 6074 80538
rect 6126 80486 6138 80538
rect 6190 80486 7912 80538
rect 4876 80464 7912 80486
rect 85284 80538 88596 80560
rect 85284 80486 86474 80538
rect 86526 80486 86538 80538
rect 86590 80486 86602 80538
rect 86654 80486 86666 80538
rect 86718 80486 86730 80538
rect 86782 80486 88596 80538
rect 85284 80464 88596 80486
rect 5409 80231 5467 80237
rect 5409 80197 5421 80231
rect 5455 80228 5467 80231
rect 8534 80228 8540 80240
rect 5455 80200 8540 80228
rect 5455 80197 5467 80200
rect 5409 80191 5467 80197
rect 8534 80188 8540 80200
rect 8592 80188 8598 80240
rect 87749 80231 87807 80237
rect 87749 80197 87761 80231
rect 87795 80228 87807 80231
rect 88206 80228 88212 80240
rect 87795 80200 88212 80228
rect 87795 80197 87807 80200
rect 87749 80191 87807 80197
rect 88206 80188 88212 80200
rect 88264 80188 88270 80240
rect 85814 80120 85820 80172
rect 85872 80160 85878 80172
rect 88049 80163 88107 80169
rect 88049 80160 88061 80163
rect 85872 80132 88061 80160
rect 85872 80120 85878 80132
rect 88049 80129 88061 80132
rect 88095 80129 88107 80163
rect 88049 80123 88107 80129
rect 4118 80052 4124 80104
rect 4176 80092 4182 80104
rect 5245 80095 5303 80101
rect 5245 80092 5257 80095
rect 4176 80064 5257 80092
rect 4176 80052 4182 80064
rect 5245 80061 5257 80064
rect 5291 80061 5303 80095
rect 5245 80055 5303 80061
rect 4876 79994 7912 80016
rect 4876 79942 6618 79994
rect 6670 79942 6682 79994
rect 6734 79942 6746 79994
rect 6798 79942 6810 79994
rect 6862 79942 6874 79994
rect 6926 79942 7912 79994
rect 4876 79920 7912 79942
rect 85284 79994 88596 80016
rect 85284 79942 87210 79994
rect 87262 79942 87274 79994
rect 87326 79942 87338 79994
rect 87390 79942 87402 79994
rect 87454 79942 87466 79994
rect 87518 79942 88596 79994
rect 85284 79920 88596 79942
rect 4876 79450 7912 79472
rect 4876 79398 5882 79450
rect 5934 79398 5946 79450
rect 5998 79398 6010 79450
rect 6062 79398 6074 79450
rect 6126 79398 6138 79450
rect 6190 79398 7912 79450
rect 4876 79376 7912 79398
rect 85284 79450 88596 79472
rect 85284 79398 86474 79450
rect 86526 79398 86538 79450
rect 86590 79398 86602 79450
rect 86654 79398 86666 79450
rect 86718 79398 86730 79450
rect 86782 79398 88596 79450
rect 85284 79376 88596 79398
rect 4876 78906 7912 78928
rect 4876 78854 6618 78906
rect 6670 78854 6682 78906
rect 6734 78854 6746 78906
rect 6798 78854 6810 78906
rect 6862 78854 6874 78906
rect 6926 78854 7912 78906
rect 4876 78832 7912 78854
rect 85284 78906 88596 78928
rect 85284 78854 87210 78906
rect 87262 78854 87274 78906
rect 87326 78854 87338 78906
rect 87390 78854 87402 78906
rect 87454 78854 87466 78906
rect 87518 78854 88596 78906
rect 85284 78832 88596 78854
rect 85814 78692 85820 78744
rect 85872 78732 85878 78744
rect 88049 78735 88107 78741
rect 88049 78732 88061 78735
rect 85872 78704 88061 78732
rect 85872 78692 85878 78704
rect 88049 78701 88061 78704
rect 88095 78701 88107 78735
rect 88049 78695 88107 78701
rect 5409 78667 5467 78673
rect 5409 78633 5421 78667
rect 5455 78664 5467 78667
rect 8534 78664 8540 78676
rect 5455 78636 8540 78664
rect 5455 78633 5467 78636
rect 5409 78627 5467 78633
rect 8534 78624 8540 78636
rect 8592 78624 8598 78676
rect 87933 78667 87991 78673
rect 87933 78633 87945 78667
rect 87979 78664 87991 78667
rect 88206 78664 88212 78676
rect 87979 78636 88212 78664
rect 87979 78633 87991 78636
rect 87933 78627 87991 78633
rect 88206 78624 88212 78636
rect 88264 78624 88270 78676
rect 4118 78488 4124 78540
rect 4176 78528 4182 78540
rect 5245 78531 5303 78537
rect 5245 78528 5257 78531
rect 4176 78500 5257 78528
rect 4176 78488 4182 78500
rect 5245 78497 5257 78500
rect 5291 78497 5303 78531
rect 5245 78491 5303 78497
rect 4876 78362 7912 78384
rect 4876 78310 5882 78362
rect 5934 78310 5946 78362
rect 5998 78310 6010 78362
rect 6062 78310 6074 78362
rect 6126 78310 6138 78362
rect 6190 78310 7912 78362
rect 4876 78288 7912 78310
rect 85284 78362 88596 78384
rect 85284 78310 86474 78362
rect 86526 78310 86538 78362
rect 86590 78310 86602 78362
rect 86654 78310 86666 78362
rect 86718 78310 86730 78362
rect 86782 78310 88596 78362
rect 85284 78288 88596 78310
rect 5409 78055 5467 78061
rect 5409 78021 5421 78055
rect 5455 78052 5467 78055
rect 8534 78052 8540 78064
rect 5455 78024 8540 78052
rect 5455 78021 5467 78024
rect 5409 78015 5467 78021
rect 8534 78012 8540 78024
rect 8592 78012 8598 78064
rect 87749 78055 87807 78061
rect 87749 78021 87761 78055
rect 87795 78052 87807 78055
rect 88206 78052 88212 78064
rect 87795 78024 88212 78052
rect 87795 78021 87807 78024
rect 87749 78015 87807 78021
rect 88206 78012 88212 78024
rect 88264 78012 88270 78064
rect 85814 77944 85820 77996
rect 85872 77984 85878 77996
rect 88049 77987 88107 77993
rect 88049 77984 88061 77987
rect 85872 77956 88061 77984
rect 85872 77944 85878 77956
rect 88049 77953 88061 77956
rect 88095 77953 88107 77987
rect 88049 77947 88107 77953
rect 4118 77876 4124 77928
rect 4176 77916 4182 77928
rect 5245 77919 5303 77925
rect 5245 77916 5257 77919
rect 4176 77888 5257 77916
rect 4176 77876 4182 77888
rect 5245 77885 5257 77888
rect 5291 77885 5303 77919
rect 5245 77879 5303 77885
rect 4876 77818 7912 77840
rect 4876 77766 6618 77818
rect 6670 77766 6682 77818
rect 6734 77766 6746 77818
rect 6798 77766 6810 77818
rect 6862 77766 6874 77818
rect 6926 77766 7912 77818
rect 4876 77744 7912 77766
rect 85284 77818 88596 77840
rect 85284 77766 87210 77818
rect 87262 77766 87274 77818
rect 87326 77766 87338 77818
rect 87390 77766 87402 77818
rect 87454 77766 87466 77818
rect 87518 77766 88596 77818
rect 85284 77744 88596 77766
rect 4876 77274 7912 77296
rect 4876 77222 5882 77274
rect 5934 77222 5946 77274
rect 5998 77222 6010 77274
rect 6062 77222 6074 77274
rect 6126 77222 6138 77274
rect 6190 77222 7912 77274
rect 4876 77200 7912 77222
rect 85284 77274 88596 77296
rect 85284 77222 86474 77274
rect 86526 77222 86538 77274
rect 86590 77222 86602 77274
rect 86654 77222 86666 77274
rect 86718 77222 86730 77274
rect 86782 77222 88596 77274
rect 85284 77200 88596 77222
rect 5409 76967 5467 76973
rect 5409 76933 5421 76967
rect 5455 76964 5467 76967
rect 8534 76964 8540 76976
rect 5455 76936 8540 76964
rect 5455 76933 5467 76936
rect 5409 76927 5467 76933
rect 8534 76924 8540 76936
rect 8592 76924 8598 76976
rect 87749 76967 87807 76973
rect 87749 76933 87761 76967
rect 87795 76964 87807 76967
rect 87795 76936 88068 76964
rect 87795 76933 87807 76936
rect 87749 76927 87807 76933
rect 88040 76840 88068 76936
rect 4210 76788 4216 76840
rect 4268 76828 4274 76840
rect 5245 76831 5303 76837
rect 5245 76828 5257 76831
rect 4268 76800 5257 76828
rect 4268 76788 4274 76800
rect 5245 76797 5257 76800
rect 5291 76797 5303 76831
rect 5245 76791 5303 76797
rect 85814 76788 85820 76840
rect 85872 76828 85878 76840
rect 87565 76831 87623 76837
rect 87565 76828 87577 76831
rect 85872 76800 87577 76828
rect 85872 76788 85878 76800
rect 87565 76797 87577 76800
rect 87611 76797 87623 76831
rect 87565 76791 87623 76797
rect 88022 76788 88028 76840
rect 88080 76788 88086 76840
rect 4876 76730 7912 76752
rect 4876 76678 6618 76730
rect 6670 76678 6682 76730
rect 6734 76678 6746 76730
rect 6798 76678 6810 76730
rect 6862 76678 6874 76730
rect 6926 76678 7912 76730
rect 4876 76656 7912 76678
rect 85284 76730 88596 76752
rect 85284 76678 87210 76730
rect 87262 76678 87274 76730
rect 87326 76678 87338 76730
rect 87390 76678 87402 76730
rect 87454 76678 87466 76730
rect 87518 76678 88596 76730
rect 85284 76656 88596 76678
rect 4876 76186 7912 76208
rect 4876 76134 5882 76186
rect 5934 76134 5946 76186
rect 5998 76134 6010 76186
rect 6062 76134 6074 76186
rect 6126 76134 6138 76186
rect 6190 76134 7912 76186
rect 4876 76112 7912 76134
rect 85284 76186 88596 76208
rect 85284 76134 86474 76186
rect 86526 76134 86538 76186
rect 86590 76134 86602 76186
rect 86654 76134 86666 76186
rect 86718 76134 86730 76186
rect 86782 76134 88596 76186
rect 85284 76112 88596 76134
rect 5409 75879 5467 75885
rect 5409 75845 5421 75879
rect 5455 75876 5467 75879
rect 8534 75876 8540 75888
rect 5455 75848 8540 75876
rect 5455 75845 5467 75848
rect 5409 75839 5467 75845
rect 8534 75836 8540 75848
rect 8592 75836 8598 75888
rect 87749 75879 87807 75885
rect 87749 75845 87761 75879
rect 87795 75876 87807 75879
rect 88206 75876 88212 75888
rect 87795 75848 88212 75876
rect 87795 75845 87807 75848
rect 87749 75839 87807 75845
rect 88206 75836 88212 75848
rect 88264 75836 88270 75888
rect 4118 75768 4124 75820
rect 4176 75808 4182 75820
rect 5245 75811 5303 75817
rect 5245 75808 5257 75811
rect 4176 75780 5257 75808
rect 4176 75768 4182 75780
rect 5245 75777 5257 75780
rect 5291 75777 5303 75811
rect 5245 75771 5303 75777
rect 85814 75768 85820 75820
rect 85872 75808 85878 75820
rect 88045 75811 88103 75817
rect 88045 75808 88057 75811
rect 85872 75780 88057 75808
rect 85872 75768 85878 75780
rect 88045 75777 88057 75780
rect 88091 75777 88103 75811
rect 88045 75771 88103 75777
rect 4876 75642 7912 75664
rect 4876 75590 6618 75642
rect 6670 75590 6682 75642
rect 6734 75590 6746 75642
rect 6798 75590 6810 75642
rect 6862 75590 6874 75642
rect 6926 75590 7912 75642
rect 4876 75568 7912 75590
rect 85284 75642 88596 75664
rect 85284 75590 87210 75642
rect 87262 75590 87274 75642
rect 87326 75590 87338 75642
rect 87390 75590 87402 75642
rect 87454 75590 87466 75642
rect 87518 75590 88596 75642
rect 85284 75568 88596 75590
rect 4876 75098 7912 75120
rect 4876 75046 5882 75098
rect 5934 75046 5946 75098
rect 5998 75046 6010 75098
rect 6062 75046 6074 75098
rect 6126 75046 6138 75098
rect 6190 75046 7912 75098
rect 4876 75024 7912 75046
rect 85284 75098 88596 75120
rect 85284 75046 86474 75098
rect 86526 75046 86538 75098
rect 86590 75046 86602 75098
rect 86654 75046 86666 75098
rect 86718 75046 86730 75098
rect 86782 75046 88596 75098
rect 85284 75024 88596 75046
rect 87749 74859 87807 74865
rect 87749 74825 87761 74859
rect 87795 74856 87807 74859
rect 87795 74828 88252 74856
rect 87795 74825 87807 74828
rect 87749 74819 87807 74825
rect 4118 74748 4124 74800
rect 4176 74788 4182 74800
rect 5245 74791 5303 74797
rect 5245 74788 5257 74791
rect 4176 74760 5257 74788
rect 4176 74748 4182 74760
rect 5245 74757 5257 74760
rect 5291 74757 5303 74791
rect 5245 74751 5303 74757
rect 5406 74748 5412 74800
rect 5464 74748 5470 74800
rect 84526 74748 84532 74800
rect 84584 74788 84590 74800
rect 88224 74797 88252 74828
rect 88045 74791 88103 74797
rect 88045 74788 88057 74791
rect 84584 74760 88057 74788
rect 84584 74748 84590 74760
rect 88045 74757 88057 74760
rect 88091 74757 88103 74791
rect 88045 74751 88103 74757
rect 88209 74791 88267 74797
rect 88209 74757 88221 74791
rect 88255 74788 88267 74791
rect 88574 74788 88580 74800
rect 88255 74760 88580 74788
rect 88255 74757 88267 74760
rect 88209 74751 88267 74757
rect 88574 74748 88580 74760
rect 88632 74748 88638 74800
rect 4876 74554 7912 74576
rect 4876 74502 6618 74554
rect 6670 74502 6682 74554
rect 6734 74502 6746 74554
rect 6798 74502 6810 74554
rect 6862 74502 6874 74554
rect 6926 74502 7912 74554
rect 4876 74480 7912 74502
rect 85284 74554 88596 74576
rect 85284 74502 87210 74554
rect 87262 74502 87274 74554
rect 87326 74502 87338 74554
rect 87390 74502 87402 74554
rect 87454 74502 87466 74554
rect 87518 74502 88596 74554
rect 85284 74480 88596 74502
rect 4876 74010 7912 74032
rect 4876 73958 5882 74010
rect 5934 73958 5946 74010
rect 5998 73958 6010 74010
rect 6062 73958 6074 74010
rect 6126 73958 6138 74010
rect 6190 73958 7912 74010
rect 4876 73936 7912 73958
rect 85284 74010 88596 74032
rect 85284 73958 86474 74010
rect 86526 73958 86538 74010
rect 86590 73958 86602 74010
rect 86654 73958 86666 74010
rect 86718 73958 86730 74010
rect 86782 73958 88596 74010
rect 85284 73936 88596 73958
rect 4876 73466 7912 73488
rect 4876 73414 6618 73466
rect 6670 73414 6682 73466
rect 6734 73414 6746 73466
rect 6798 73414 6810 73466
rect 6862 73414 6874 73466
rect 6926 73414 7912 73466
rect 4876 73392 7912 73414
rect 85284 73466 88596 73488
rect 85284 73414 87210 73466
rect 87262 73414 87274 73466
rect 87326 73414 87338 73466
rect 87390 73414 87402 73466
rect 87454 73414 87466 73466
rect 87518 73414 88596 73466
rect 85284 73392 88596 73414
rect 84802 73252 84808 73304
rect 84860 73292 84866 73304
rect 88050 73295 88108 73301
rect 88050 73292 88062 73295
rect 84860 73264 88062 73292
rect 84860 73252 84866 73264
rect 88050 73261 88062 73264
rect 88096 73261 88108 73295
rect 88050 73255 88108 73261
rect 5406 73184 5412 73236
rect 5464 73184 5470 73236
rect 87933 73227 87991 73233
rect 87933 73193 87945 73227
rect 87979 73224 87991 73227
rect 88206 73224 88212 73236
rect 87979 73196 88212 73224
rect 87979 73193 87991 73196
rect 87933 73187 87991 73193
rect 88206 73184 88212 73196
rect 88264 73184 88270 73236
rect 4118 73048 4124 73100
rect 4176 73088 4182 73100
rect 5245 73091 5303 73097
rect 5245 73088 5257 73091
rect 4176 73060 5257 73088
rect 4176 73048 4182 73060
rect 5245 73057 5257 73060
rect 5291 73057 5303 73091
rect 5245 73051 5303 73057
rect 4876 72922 7912 72944
rect 4876 72870 5882 72922
rect 5934 72870 5946 72922
rect 5998 72870 6010 72922
rect 6062 72870 6074 72922
rect 6126 72870 6138 72922
rect 6190 72870 7912 72922
rect 4876 72848 7912 72870
rect 85284 72922 88596 72944
rect 85284 72870 86474 72922
rect 86526 72870 86538 72922
rect 86590 72870 86602 72922
rect 86654 72870 86666 72922
rect 86718 72870 86730 72922
rect 86782 72870 88596 72922
rect 85284 72848 88596 72870
rect 5409 72615 5467 72621
rect 5409 72581 5421 72615
rect 5455 72612 5467 72615
rect 8534 72612 8540 72624
rect 5455 72584 8540 72612
rect 5455 72581 5467 72584
rect 5409 72575 5467 72581
rect 8534 72572 8540 72584
rect 8592 72572 8598 72624
rect 87749 72615 87807 72621
rect 87749 72581 87761 72615
rect 87795 72612 87807 72615
rect 88206 72612 88212 72624
rect 87795 72584 88212 72612
rect 87795 72581 87807 72584
rect 87749 72575 87807 72581
rect 88206 72572 88212 72584
rect 88264 72572 88270 72624
rect 4118 72436 4124 72488
rect 4176 72476 4182 72488
rect 5245 72479 5303 72485
rect 5245 72476 5257 72479
rect 4176 72448 5257 72476
rect 4176 72436 4182 72448
rect 5245 72445 5257 72448
rect 5291 72445 5303 72479
rect 5245 72439 5303 72445
rect 87838 72436 87844 72488
rect 87896 72476 87902 72488
rect 88050 72479 88108 72485
rect 88050 72476 88062 72479
rect 87896 72448 88062 72476
rect 87896 72436 87902 72448
rect 88050 72445 88062 72448
rect 88096 72445 88108 72479
rect 88050 72439 88108 72445
rect 4876 72378 7912 72400
rect 4876 72326 6618 72378
rect 6670 72326 6682 72378
rect 6734 72326 6746 72378
rect 6798 72326 6810 72378
rect 6862 72326 6874 72378
rect 6926 72326 7912 72378
rect 4876 72304 7912 72326
rect 85284 72378 88596 72400
rect 85284 72326 87210 72378
rect 87262 72326 87274 72378
rect 87326 72326 87338 72378
rect 87390 72326 87402 72378
rect 87454 72326 87466 72378
rect 87518 72326 88596 72378
rect 85284 72304 88596 72326
rect 4876 71834 7912 71856
rect 4876 71782 5882 71834
rect 5934 71782 5946 71834
rect 5998 71782 6010 71834
rect 6062 71782 6074 71834
rect 6126 71782 6138 71834
rect 6190 71782 7912 71834
rect 4876 71760 7912 71782
rect 85284 71834 88596 71856
rect 85284 71782 86474 71834
rect 86526 71782 86538 71834
rect 86590 71782 86602 71834
rect 86654 71782 86666 71834
rect 86718 71782 86730 71834
rect 86782 71782 88596 71834
rect 85284 71760 88596 71782
rect 5409 71527 5467 71533
rect 5409 71493 5421 71527
rect 5455 71524 5467 71527
rect 8534 71524 8540 71536
rect 5455 71496 8540 71524
rect 5455 71493 5467 71496
rect 5409 71487 5467 71493
rect 8534 71484 8540 71496
rect 8592 71484 8598 71536
rect 87749 71527 87807 71533
rect 87749 71493 87761 71527
rect 87795 71524 87807 71527
rect 88206 71524 88212 71536
rect 87795 71496 88212 71524
rect 87795 71493 87807 71496
rect 87749 71487 87807 71493
rect 88206 71484 88212 71496
rect 88264 71484 88270 71536
rect 85814 71416 85820 71468
rect 85872 71456 85878 71468
rect 88049 71459 88107 71465
rect 88049 71456 88061 71459
rect 85872 71428 88061 71456
rect 85872 71416 85878 71428
rect 88049 71425 88061 71428
rect 88095 71425 88107 71459
rect 88049 71419 88107 71425
rect 4210 71348 4216 71400
rect 4268 71388 4274 71400
rect 5245 71391 5303 71397
rect 5245 71388 5257 71391
rect 4268 71360 5257 71388
rect 4268 71348 4274 71360
rect 5245 71357 5257 71360
rect 5291 71357 5303 71391
rect 5245 71351 5303 71357
rect 4876 71290 7912 71312
rect 4876 71238 6618 71290
rect 6670 71238 6682 71290
rect 6734 71238 6746 71290
rect 6798 71238 6810 71290
rect 6862 71238 6874 71290
rect 6926 71238 7912 71290
rect 4876 71216 7912 71238
rect 85284 71290 88596 71312
rect 85284 71238 87210 71290
rect 87262 71238 87274 71290
rect 87326 71238 87338 71290
rect 87390 71238 87402 71290
rect 87454 71238 87466 71290
rect 87518 71238 88596 71290
rect 85284 71216 88596 71238
rect 4876 70746 7912 70768
rect 4876 70694 5882 70746
rect 5934 70694 5946 70746
rect 5998 70694 6010 70746
rect 6062 70694 6074 70746
rect 6126 70694 6138 70746
rect 6190 70694 7912 70746
rect 4876 70672 7912 70694
rect 85284 70746 88596 70768
rect 85284 70694 86474 70746
rect 86526 70694 86538 70746
rect 86590 70694 86602 70746
rect 86654 70694 86666 70746
rect 86718 70694 86730 70746
rect 86782 70694 88596 70746
rect 85284 70672 88596 70694
rect 5409 70439 5467 70445
rect 5409 70405 5421 70439
rect 5455 70436 5467 70439
rect 8534 70436 8540 70448
rect 5455 70408 8540 70436
rect 5455 70405 5467 70408
rect 5409 70399 5467 70405
rect 8534 70396 8540 70408
rect 8592 70396 8598 70448
rect 87749 70439 87807 70445
rect 87749 70405 87761 70439
rect 87795 70436 87807 70439
rect 88206 70436 88212 70448
rect 87795 70408 88212 70436
rect 87795 70405 87807 70408
rect 87749 70399 87807 70405
rect 88206 70396 88212 70408
rect 88264 70396 88270 70448
rect 4118 70328 4124 70380
rect 4176 70368 4182 70380
rect 5245 70371 5303 70377
rect 5245 70368 5257 70371
rect 4176 70340 5257 70368
rect 4176 70328 4182 70340
rect 5245 70337 5257 70340
rect 5291 70337 5303 70371
rect 5245 70331 5303 70337
rect 85814 70328 85820 70380
rect 85872 70368 85878 70380
rect 88049 70371 88107 70377
rect 88049 70368 88061 70371
rect 85872 70340 88061 70368
rect 85872 70328 85878 70340
rect 88049 70337 88061 70340
rect 88095 70337 88107 70371
rect 88049 70331 88107 70337
rect 4876 70202 7912 70224
rect 4876 70150 6618 70202
rect 6670 70150 6682 70202
rect 6734 70150 6746 70202
rect 6798 70150 6810 70202
rect 6862 70150 6874 70202
rect 6926 70150 7912 70202
rect 4876 70128 7912 70150
rect 85284 70202 88596 70224
rect 85284 70150 87210 70202
rect 87262 70150 87274 70202
rect 87326 70150 87338 70202
rect 87390 70150 87402 70202
rect 87454 70150 87466 70202
rect 87518 70150 88596 70202
rect 85284 70128 88596 70150
rect 4876 69658 7912 69680
rect 4876 69606 5882 69658
rect 5934 69606 5946 69658
rect 5998 69606 6010 69658
rect 6062 69606 6074 69658
rect 6126 69606 6138 69658
rect 6190 69606 7912 69658
rect 4876 69584 7912 69606
rect 85284 69658 88596 69680
rect 85284 69606 86474 69658
rect 86526 69606 86538 69658
rect 86590 69606 86602 69658
rect 86654 69606 86666 69658
rect 86718 69606 86730 69658
rect 86782 69606 88596 69658
rect 85284 69584 88596 69606
rect 5406 69308 5412 69360
rect 5464 69308 5470 69360
rect 87749 69351 87807 69357
rect 87749 69317 87761 69351
rect 87795 69348 87807 69351
rect 88209 69351 88267 69357
rect 88209 69348 88221 69351
rect 87795 69320 88221 69348
rect 87795 69317 87807 69320
rect 87749 69311 87807 69317
rect 88209 69317 88221 69320
rect 88255 69348 88267 69351
rect 88574 69348 88580 69360
rect 88255 69320 88580 69348
rect 88255 69317 88267 69320
rect 88209 69311 88267 69317
rect 88574 69308 88580 69320
rect 88632 69308 88638 69360
rect 4118 69240 4124 69292
rect 4176 69280 4182 69292
rect 5245 69283 5303 69289
rect 5245 69280 5257 69283
rect 4176 69252 5257 69280
rect 4176 69240 4182 69252
rect 5245 69249 5257 69252
rect 5291 69249 5303 69283
rect 5245 69243 5303 69249
rect 84802 69240 84808 69292
rect 84860 69280 84866 69292
rect 88050 69283 88108 69289
rect 88050 69280 88062 69283
rect 84860 69252 88062 69280
rect 84860 69240 84866 69252
rect 88050 69249 88062 69252
rect 88096 69249 88108 69283
rect 88050 69243 88108 69249
rect 4876 69114 7912 69136
rect 4876 69062 6618 69114
rect 6670 69062 6682 69114
rect 6734 69062 6746 69114
rect 6798 69062 6810 69114
rect 6862 69062 6874 69114
rect 6926 69062 7912 69114
rect 4876 69040 7912 69062
rect 85284 69114 88596 69136
rect 85284 69062 87210 69114
rect 87262 69062 87274 69114
rect 87326 69062 87338 69114
rect 87390 69062 87402 69114
rect 87454 69062 87466 69114
rect 87518 69062 88596 69114
rect 85284 69040 88596 69062
rect 4876 68570 7912 68592
rect 4876 68518 5882 68570
rect 5934 68518 5946 68570
rect 5998 68518 6010 68570
rect 6062 68518 6074 68570
rect 6126 68518 6138 68570
rect 6190 68518 7912 68570
rect 4876 68496 7912 68518
rect 85284 68570 88596 68592
rect 85284 68518 86474 68570
rect 86526 68518 86538 68570
rect 86590 68518 86602 68570
rect 86654 68518 86666 68570
rect 86718 68518 86730 68570
rect 86782 68518 88596 68570
rect 85284 68496 88596 68518
rect 4876 68026 7912 68048
rect 4876 67974 6618 68026
rect 6670 67974 6682 68026
rect 6734 67974 6746 68026
rect 6798 67974 6810 68026
rect 6862 67974 6874 68026
rect 6926 67974 7912 68026
rect 4876 67952 7912 67974
rect 85284 68026 88596 68048
rect 85284 67974 87210 68026
rect 87262 67974 87274 68026
rect 87326 67974 87338 68026
rect 87390 67974 87402 68026
rect 87454 67974 87466 68026
rect 87518 67974 88596 68026
rect 85284 67952 88596 67974
rect 85262 67812 85268 67864
rect 85320 67852 85326 67864
rect 88049 67855 88107 67861
rect 88049 67852 88061 67855
rect 85320 67824 88061 67852
rect 85320 67812 85326 67824
rect 88049 67821 88061 67824
rect 88095 67821 88107 67855
rect 88049 67815 88107 67821
rect 5406 67744 5412 67796
rect 5464 67744 5470 67796
rect 87933 67787 87991 67793
rect 87933 67753 87945 67787
rect 87979 67784 87991 67787
rect 88206 67784 88212 67796
rect 87979 67756 88212 67784
rect 87979 67753 87991 67756
rect 87933 67747 87991 67753
rect 88206 67744 88212 67756
rect 88264 67744 88270 67796
rect 4026 67608 4032 67660
rect 4084 67648 4090 67660
rect 5245 67651 5303 67657
rect 5245 67648 5257 67651
rect 4084 67620 5257 67648
rect 4084 67608 4090 67620
rect 5245 67617 5257 67620
rect 5291 67617 5303 67651
rect 5245 67611 5303 67617
rect 4876 67482 7912 67504
rect 4876 67430 5882 67482
rect 5934 67430 5946 67482
rect 5998 67430 6010 67482
rect 6062 67430 6074 67482
rect 6126 67430 6138 67482
rect 6190 67430 7912 67482
rect 4876 67408 7912 67430
rect 85284 67482 88596 67504
rect 85284 67430 86474 67482
rect 86526 67430 86538 67482
rect 86590 67430 86602 67482
rect 86654 67430 86666 67482
rect 86718 67430 86730 67482
rect 86782 67430 88596 67482
rect 85284 67408 88596 67430
rect 5409 67175 5467 67181
rect 5409 67141 5421 67175
rect 5455 67172 5467 67175
rect 8534 67172 8540 67184
rect 5455 67144 8540 67172
rect 5455 67141 5467 67144
rect 5409 67135 5467 67141
rect 8534 67132 8540 67144
rect 8592 67132 8598 67184
rect 87749 67175 87807 67181
rect 87749 67141 87761 67175
rect 87795 67172 87807 67175
rect 88206 67172 88212 67184
rect 87795 67144 88212 67172
rect 87795 67141 87807 67144
rect 87749 67135 87807 67141
rect 88206 67132 88212 67144
rect 88264 67132 88270 67184
rect 85814 67064 85820 67116
rect 85872 67104 85878 67116
rect 88050 67107 88108 67113
rect 88050 67104 88062 67107
rect 85872 67076 88062 67104
rect 85872 67064 85878 67076
rect 88050 67073 88062 67076
rect 88096 67073 88108 67107
rect 88050 67067 88108 67073
rect 4118 66996 4124 67048
rect 4176 67036 4182 67048
rect 5245 67039 5303 67045
rect 5245 67036 5257 67039
rect 4176 67008 5257 67036
rect 4176 66996 4182 67008
rect 5245 67005 5257 67008
rect 5291 67005 5303 67039
rect 5245 66999 5303 67005
rect 4876 66938 7912 66960
rect 4876 66886 6618 66938
rect 6670 66886 6682 66938
rect 6734 66886 6746 66938
rect 6798 66886 6810 66938
rect 6862 66886 6874 66938
rect 6926 66886 7912 66938
rect 4876 66864 7912 66886
rect 85284 66938 88596 66960
rect 85284 66886 87210 66938
rect 87262 66886 87274 66938
rect 87326 66886 87338 66938
rect 87390 66886 87402 66938
rect 87454 66886 87466 66938
rect 87518 66886 88596 66938
rect 85284 66864 88596 66886
rect 4876 66394 7912 66416
rect 4876 66342 5882 66394
rect 5934 66342 5946 66394
rect 5998 66342 6010 66394
rect 6062 66342 6074 66394
rect 6126 66342 6138 66394
rect 6190 66342 7912 66394
rect 4876 66320 7912 66342
rect 85284 66394 88596 66416
rect 85284 66342 86474 66394
rect 86526 66342 86538 66394
rect 86590 66342 86602 66394
rect 86654 66342 86666 66394
rect 86718 66342 86730 66394
rect 86782 66342 88596 66394
rect 85284 66320 88596 66342
rect 5363 66155 5421 66161
rect 5363 66121 5375 66155
rect 5409 66152 5421 66155
rect 8534 66152 8540 66164
rect 5409 66124 8540 66152
rect 5409 66121 5421 66124
rect 5363 66115 5421 66121
rect 8534 66112 8540 66124
rect 8592 66112 8598 66164
rect 4302 66044 4308 66096
rect 4360 66084 4366 66096
rect 5161 66087 5219 66093
rect 5161 66084 5173 66087
rect 4360 66056 5173 66084
rect 4360 66044 4366 66056
rect 5161 66053 5173 66056
rect 5207 66084 5219 66087
rect 5501 66087 5559 66093
rect 5501 66084 5513 66087
rect 5207 66056 5513 66084
rect 5207 66053 5219 66056
rect 5161 66047 5219 66053
rect 5501 66053 5513 66056
rect 5547 66053 5559 66087
rect 5501 66047 5559 66053
rect 85814 66044 85820 66096
rect 85872 66084 85878 66096
rect 87957 66087 88015 66093
rect 87957 66084 87969 66087
rect 85872 66056 87969 66084
rect 85872 66044 85878 66056
rect 87957 66053 87969 66056
rect 88003 66053 88015 66087
rect 87957 66047 88015 66053
rect 88206 65957 88212 65960
rect 88163 65951 88212 65957
rect 88163 65917 88175 65951
rect 88209 65917 88212 65951
rect 88163 65911 88212 65917
rect 88206 65908 88212 65911
rect 88264 65908 88270 65960
rect 4876 65850 7912 65872
rect 4876 65798 6618 65850
rect 6670 65798 6682 65850
rect 6734 65798 6746 65850
rect 6798 65798 6810 65850
rect 6862 65798 6874 65850
rect 6926 65798 7912 65850
rect 4876 65776 7912 65798
rect 85284 65850 88596 65872
rect 85284 65798 87210 65850
rect 87262 65798 87274 65850
rect 87326 65798 87338 65850
rect 87390 65798 87402 65850
rect 87454 65798 87466 65850
rect 87518 65798 88596 65850
rect 85284 65776 88596 65798
rect 4876 65306 7912 65328
rect 4876 65254 5882 65306
rect 5934 65254 5946 65306
rect 5998 65254 6010 65306
rect 6062 65254 6074 65306
rect 6126 65254 6138 65306
rect 6190 65254 7912 65306
rect 4876 65232 7912 65254
rect 85284 65306 88596 65328
rect 85284 65254 86474 65306
rect 86526 65254 86538 65306
rect 86590 65254 86602 65306
rect 86654 65254 86666 65306
rect 86718 65254 86730 65306
rect 86782 65254 88596 65306
rect 85284 65232 88596 65254
rect 5363 65067 5421 65073
rect 5363 65033 5375 65067
rect 5409 65064 5421 65067
rect 8534 65064 8540 65076
rect 5409 65036 8540 65064
rect 5409 65033 5421 65036
rect 5363 65027 5421 65033
rect 8534 65024 8540 65036
rect 8592 65024 8598 65076
rect 4302 64956 4308 65008
rect 4360 64996 4366 65008
rect 5161 64999 5219 65005
rect 5161 64996 5173 64999
rect 4360 64968 5173 64996
rect 4360 64956 4366 64968
rect 5161 64965 5173 64968
rect 5207 64996 5219 64999
rect 5501 64999 5559 65005
rect 5501 64996 5513 64999
rect 5207 64968 5513 64996
rect 5207 64965 5219 64968
rect 5161 64959 5219 64965
rect 5501 64965 5513 64968
rect 5547 64965 5559 64999
rect 5501 64959 5559 64965
rect 85814 64956 85820 65008
rect 85872 64996 85878 65008
rect 87957 64999 88015 65005
rect 87957 64996 87969 64999
rect 85872 64968 87969 64996
rect 85872 64956 85878 64968
rect 87957 64965 87969 64968
rect 88003 64965 88015 64999
rect 87957 64959 88015 64965
rect 88163 64863 88221 64869
rect 88163 64829 88175 64863
rect 88209 64860 88221 64863
rect 88390 64860 88396 64872
rect 88209 64832 88396 64860
rect 88209 64829 88221 64832
rect 88163 64823 88221 64829
rect 88390 64820 88396 64832
rect 88448 64820 88454 64872
rect 4876 64762 7912 64784
rect 4876 64710 6618 64762
rect 6670 64710 6682 64762
rect 6734 64710 6746 64762
rect 6798 64710 6810 64762
rect 6862 64710 6874 64762
rect 6926 64710 7912 64762
rect 4876 64688 7912 64710
rect 85284 64762 88596 64784
rect 85284 64710 87210 64762
rect 87262 64710 87274 64762
rect 87326 64710 87338 64762
rect 87390 64710 87402 64762
rect 87454 64710 87466 64762
rect 87518 64710 88596 64762
rect 85284 64688 88596 64710
rect 7522 64548 7528 64600
rect 7580 64548 7586 64600
rect 4876 64218 7912 64240
rect 4876 64166 5882 64218
rect 5934 64166 5946 64218
rect 5998 64166 6010 64218
rect 6062 64166 6074 64218
rect 6126 64166 6138 64218
rect 6190 64166 7912 64218
rect 4876 64144 7912 64166
rect 85284 64218 88596 64240
rect 85284 64166 86474 64218
rect 86526 64166 86538 64218
rect 86590 64166 86602 64218
rect 86654 64166 86666 64218
rect 86718 64166 86730 64218
rect 86782 64166 88596 64218
rect 85284 64144 88596 64166
rect 4302 63868 4308 63920
rect 4360 63908 4366 63920
rect 5161 63911 5219 63917
rect 5161 63908 5173 63911
rect 4360 63880 5173 63908
rect 4360 63868 4366 63880
rect 5161 63877 5173 63880
rect 5207 63908 5219 63911
rect 5501 63911 5559 63917
rect 5501 63908 5513 63911
rect 5207 63880 5513 63908
rect 5207 63877 5219 63880
rect 5161 63871 5219 63877
rect 5501 63877 5513 63880
rect 5547 63877 5559 63911
rect 5501 63871 5559 63877
rect 7389 63911 7447 63917
rect 7389 63877 7401 63911
rect 7435 63908 7447 63911
rect 7522 63908 7528 63920
rect 7435 63880 7528 63908
rect 7435 63877 7447 63880
rect 7389 63871 7447 63877
rect 7522 63868 7528 63880
rect 7580 63868 7586 63920
rect 84526 63868 84532 63920
rect 84584 63908 84590 63920
rect 87957 63911 88015 63917
rect 87957 63908 87969 63911
rect 84584 63880 87969 63908
rect 84584 63868 84590 63880
rect 87957 63877 87969 63880
rect 88003 63877 88015 63911
rect 87957 63871 88015 63877
rect 5363 63775 5421 63781
rect 5363 63741 5375 63775
rect 5409 63772 5421 63775
rect 5682 63772 5688 63784
rect 5409 63744 5688 63772
rect 5409 63741 5421 63744
rect 5363 63735 5421 63741
rect 5682 63732 5688 63744
rect 5740 63732 5746 63784
rect 6605 63775 6663 63781
rect 6605 63741 6617 63775
rect 6651 63772 6663 63775
rect 7798 63772 7804 63784
rect 6651 63744 7804 63772
rect 6651 63741 6663 63744
rect 6605 63735 6663 63741
rect 7798 63732 7804 63744
rect 7856 63732 7862 63784
rect 88163 63775 88221 63781
rect 88163 63741 88175 63775
rect 88209 63772 88221 63775
rect 88574 63772 88580 63784
rect 88209 63744 88580 63772
rect 88209 63741 88221 63744
rect 88163 63735 88221 63741
rect 88574 63732 88580 63744
rect 88632 63732 88638 63784
rect 4876 63674 7912 63696
rect 4876 63622 6618 63674
rect 6670 63622 6682 63674
rect 6734 63622 6746 63674
rect 6798 63622 6810 63674
rect 6862 63622 6874 63674
rect 6926 63622 7912 63674
rect 4876 63600 7912 63622
rect 85284 63674 88596 63696
rect 85284 63622 87210 63674
rect 87262 63622 87274 63674
rect 87326 63622 87338 63674
rect 87390 63622 87402 63674
rect 87454 63622 87466 63674
rect 87518 63622 88596 63674
rect 85284 63600 88596 63622
rect 7338 63460 7344 63512
rect 7396 63500 7402 63512
rect 7525 63503 7583 63509
rect 7525 63500 7537 63503
rect 7396 63472 7537 63500
rect 7396 63460 7402 63472
rect 7525 63469 7537 63472
rect 7571 63500 7583 63503
rect 7798 63500 7804 63512
rect 7571 63472 7804 63500
rect 7571 63469 7583 63472
rect 7525 63463 7583 63469
rect 7798 63460 7804 63472
rect 7856 63460 7862 63512
rect 4876 63130 7912 63152
rect 4876 63078 5882 63130
rect 5934 63078 5946 63130
rect 5998 63078 6010 63130
rect 6062 63078 6074 63130
rect 6126 63078 6138 63130
rect 6190 63078 7912 63130
rect 4876 63056 7912 63078
rect 85284 63130 88596 63152
rect 85284 63078 86474 63130
rect 86526 63078 86538 63130
rect 86590 63078 86602 63130
rect 86654 63078 86666 63130
rect 86718 63078 86730 63130
rect 86782 63078 88596 63130
rect 85284 63056 88596 63078
rect 4876 62586 7912 62608
rect 4876 62534 6618 62586
rect 6670 62534 6682 62586
rect 6734 62534 6746 62586
rect 6798 62534 6810 62586
rect 6862 62534 6874 62586
rect 6926 62534 7912 62586
rect 4876 62512 7912 62534
rect 85284 62586 88596 62608
rect 85284 62534 87210 62586
rect 87262 62534 87274 62586
rect 87326 62534 87338 62586
rect 87390 62534 87402 62586
rect 87454 62534 87466 62586
rect 87518 62534 88596 62586
rect 85284 62512 88596 62534
rect 4302 62304 4308 62356
rect 4360 62344 4366 62356
rect 5161 62347 5219 62353
rect 5161 62344 5173 62347
rect 4360 62316 5173 62344
rect 4360 62304 4366 62316
rect 5161 62313 5173 62316
rect 5207 62344 5219 62347
rect 5501 62347 5559 62353
rect 5501 62344 5513 62347
rect 5207 62316 5513 62344
rect 5207 62313 5219 62316
rect 5161 62307 5219 62313
rect 5501 62313 5513 62316
rect 5547 62313 5559 62347
rect 5501 62307 5559 62313
rect 84802 62304 84808 62356
rect 84860 62344 84866 62356
rect 87957 62347 88015 62353
rect 87957 62344 87969 62347
rect 84860 62316 87969 62344
rect 84860 62304 84866 62316
rect 87957 62313 87969 62316
rect 88003 62313 88015 62347
rect 87957 62307 88015 62313
rect 5363 62211 5421 62217
rect 5363 62177 5375 62211
rect 5409 62208 5421 62211
rect 5682 62208 5688 62220
rect 5409 62180 5688 62208
rect 5409 62177 5421 62180
rect 5363 62171 5421 62177
rect 5682 62168 5688 62180
rect 5740 62168 5746 62220
rect 88163 62143 88221 62149
rect 88163 62109 88175 62143
rect 88209 62140 88221 62143
rect 88390 62140 88396 62152
rect 88209 62112 88396 62140
rect 88209 62109 88221 62112
rect 88163 62103 88221 62109
rect 88390 62100 88396 62112
rect 88448 62100 88454 62152
rect 4876 62042 7912 62064
rect 4876 61990 5882 62042
rect 5934 61990 5946 62042
rect 5998 61990 6010 62042
rect 6062 61990 6074 62042
rect 6126 61990 6138 62042
rect 6190 61990 7912 62042
rect 4876 61968 7912 61990
rect 85284 62042 88596 62064
rect 85284 61990 86474 62042
rect 86526 61990 86538 62042
rect 86590 61990 86602 62042
rect 86654 61990 86666 62042
rect 86718 61990 86730 62042
rect 86782 61990 88596 62042
rect 85284 61968 88596 61990
rect 4302 61692 4308 61744
rect 4360 61732 4366 61744
rect 5161 61735 5219 61741
rect 5161 61732 5173 61735
rect 4360 61704 5173 61732
rect 4360 61692 4366 61704
rect 5161 61701 5173 61704
rect 5207 61732 5219 61735
rect 5501 61735 5559 61741
rect 5501 61732 5513 61735
rect 5207 61704 5513 61732
rect 5207 61701 5219 61704
rect 5161 61695 5219 61701
rect 5501 61701 5513 61704
rect 5547 61701 5559 61735
rect 5501 61695 5559 61701
rect 85814 61692 85820 61744
rect 85872 61732 85878 61744
rect 87957 61735 88015 61741
rect 87957 61732 87969 61735
rect 85872 61704 87969 61732
rect 85872 61692 85878 61704
rect 87957 61701 87969 61704
rect 88003 61701 88015 61735
rect 87957 61695 88015 61701
rect 5363 61667 5421 61673
rect 5363 61633 5375 61667
rect 5409 61664 5421 61667
rect 8534 61664 8540 61676
rect 5409 61636 8540 61664
rect 5409 61633 5421 61636
rect 5363 61627 5421 61633
rect 8534 61624 8540 61636
rect 8592 61624 8598 61676
rect 88206 61605 88212 61608
rect 88163 61599 88212 61605
rect 88163 61565 88175 61599
rect 88209 61565 88212 61599
rect 88163 61559 88212 61565
rect 88206 61556 88212 61559
rect 88264 61556 88270 61608
rect 4876 61498 7912 61520
rect 4876 61446 6618 61498
rect 6670 61446 6682 61498
rect 6734 61446 6746 61498
rect 6798 61446 6810 61498
rect 6862 61446 6874 61498
rect 6926 61446 7912 61498
rect 4876 61424 7912 61446
rect 85284 61498 88596 61520
rect 85284 61446 87210 61498
rect 87262 61446 87274 61498
rect 87326 61446 87338 61498
rect 87390 61446 87402 61498
rect 87454 61446 87466 61498
rect 87518 61446 88596 61498
rect 85284 61424 88596 61446
rect 4876 60954 7912 60976
rect 4876 60902 5882 60954
rect 5934 60902 5946 60954
rect 5998 60902 6010 60954
rect 6062 60902 6074 60954
rect 6126 60902 6138 60954
rect 6190 60902 7912 60954
rect 4876 60880 7912 60902
rect 85284 60954 88596 60976
rect 85284 60902 86474 60954
rect 86526 60902 86538 60954
rect 86590 60902 86602 60954
rect 86654 60902 86666 60954
rect 86718 60902 86730 60954
rect 86782 60902 88596 60954
rect 85284 60880 88596 60902
rect 4302 60604 4308 60656
rect 4360 60644 4366 60656
rect 5161 60647 5219 60653
rect 5161 60644 5173 60647
rect 4360 60616 5173 60644
rect 4360 60604 4366 60616
rect 5161 60613 5173 60616
rect 5207 60644 5219 60647
rect 5501 60647 5559 60653
rect 5501 60644 5513 60647
rect 5207 60616 5513 60644
rect 5207 60613 5219 60616
rect 5161 60607 5219 60613
rect 5501 60613 5513 60616
rect 5547 60613 5559 60647
rect 5501 60607 5559 60613
rect 85814 60604 85820 60656
rect 85872 60644 85878 60656
rect 87957 60647 88015 60653
rect 87957 60644 87969 60647
rect 85872 60616 87969 60644
rect 85872 60604 85878 60616
rect 87957 60613 87969 60616
rect 88003 60613 88015 60647
rect 87957 60607 88015 60613
rect 5363 60579 5421 60585
rect 5363 60545 5375 60579
rect 5409 60576 5421 60579
rect 8534 60576 8540 60588
rect 5409 60548 8540 60576
rect 5409 60545 5421 60548
rect 5363 60539 5421 60545
rect 8534 60536 8540 60548
rect 8592 60536 8598 60588
rect 88206 60517 88212 60520
rect 88163 60511 88212 60517
rect 88163 60477 88175 60511
rect 88209 60477 88212 60511
rect 88163 60471 88212 60477
rect 88206 60468 88212 60471
rect 88264 60468 88270 60520
rect 4876 60410 7912 60432
rect 4876 60358 6618 60410
rect 6670 60358 6682 60410
rect 6734 60358 6746 60410
rect 6798 60358 6810 60410
rect 6862 60358 6874 60410
rect 6926 60358 7912 60410
rect 4876 60336 7912 60358
rect 85284 60410 88596 60432
rect 85284 60358 87210 60410
rect 87262 60358 87274 60410
rect 87326 60358 87338 60410
rect 87390 60358 87402 60410
rect 87454 60358 87466 60410
rect 87518 60358 88596 60410
rect 85284 60336 88596 60358
rect 4876 59866 7912 59888
rect 4876 59814 5882 59866
rect 5934 59814 5946 59866
rect 5998 59814 6010 59866
rect 6062 59814 6074 59866
rect 6126 59814 6138 59866
rect 6190 59814 7912 59866
rect 4876 59792 7912 59814
rect 85284 59866 88596 59888
rect 85284 59814 86474 59866
rect 86526 59814 86538 59866
rect 86590 59814 86602 59866
rect 86654 59814 86666 59866
rect 86718 59814 86730 59866
rect 86782 59814 88596 59866
rect 85284 59792 88596 59814
rect 4302 59516 4308 59568
rect 4360 59556 4366 59568
rect 5161 59559 5219 59565
rect 5161 59556 5173 59559
rect 4360 59528 5173 59556
rect 4360 59516 4366 59528
rect 5161 59525 5173 59528
rect 5207 59556 5219 59559
rect 5501 59559 5559 59565
rect 5501 59556 5513 59559
rect 5207 59528 5513 59556
rect 5207 59525 5219 59528
rect 5161 59519 5219 59525
rect 5501 59525 5513 59528
rect 5547 59525 5559 59559
rect 5501 59519 5559 59525
rect 87470 59516 87476 59568
rect 87528 59556 87534 59568
rect 87957 59559 88015 59565
rect 87957 59556 87969 59559
rect 87528 59528 87969 59556
rect 87528 59516 87534 59528
rect 87957 59525 87969 59528
rect 88003 59525 88015 59559
rect 87957 59519 88015 59525
rect 8534 59488 8540 59500
rect 5240 59460 8540 59488
rect 5240 59420 5268 59460
rect 8534 59448 8540 59460
rect 8592 59448 8598 59500
rect 88206 59429 88212 59432
rect 5363 59423 5421 59429
rect 5363 59420 5375 59423
rect 5240 59392 5375 59420
rect 5363 59389 5375 59392
rect 5409 59389 5421 59423
rect 5363 59383 5421 59389
rect 88163 59423 88212 59429
rect 88163 59389 88175 59423
rect 88209 59389 88212 59423
rect 88163 59383 88212 59389
rect 88206 59380 88212 59383
rect 88264 59380 88270 59432
rect 4876 59322 7912 59344
rect 4876 59270 6618 59322
rect 6670 59270 6682 59322
rect 6734 59270 6746 59322
rect 6798 59270 6810 59322
rect 6862 59270 6874 59322
rect 6926 59270 7912 59322
rect 4876 59248 7912 59270
rect 85284 59322 88596 59344
rect 85284 59270 87210 59322
rect 87262 59270 87274 59322
rect 87326 59270 87338 59322
rect 87390 59270 87402 59322
rect 87454 59270 87466 59322
rect 87518 59270 88596 59322
rect 85284 59248 88596 59270
rect 4876 58778 7912 58800
rect 4876 58726 5882 58778
rect 5934 58726 5946 58778
rect 5998 58726 6010 58778
rect 6062 58726 6074 58778
rect 6126 58726 6138 58778
rect 6190 58726 7912 58778
rect 4876 58704 7912 58726
rect 85284 58778 88596 58800
rect 85284 58726 86474 58778
rect 86526 58726 86538 58778
rect 86590 58726 86602 58778
rect 86654 58726 86666 58778
rect 86718 58726 86730 58778
rect 86782 58726 88596 58778
rect 85284 58704 88596 58726
rect 4302 58428 4308 58480
rect 4360 58468 4366 58480
rect 5161 58471 5219 58477
rect 5161 58468 5173 58471
rect 4360 58440 5173 58468
rect 4360 58428 4366 58440
rect 5161 58437 5173 58440
rect 5207 58468 5219 58471
rect 5501 58471 5559 58477
rect 5501 58468 5513 58471
rect 5207 58440 5513 58468
rect 5207 58437 5219 58440
rect 5161 58431 5219 58437
rect 5501 58437 5513 58440
rect 5547 58437 5559 58471
rect 5501 58431 5559 58437
rect 85078 58428 85084 58480
rect 85136 58468 85142 58480
rect 87957 58471 88015 58477
rect 87957 58468 87969 58471
rect 85136 58440 87969 58468
rect 85136 58428 85142 58440
rect 87957 58437 87969 58440
rect 88003 58437 88015 58471
rect 87957 58431 88015 58437
rect 5406 58341 5412 58344
rect 5363 58335 5412 58341
rect 5363 58301 5375 58335
rect 5409 58301 5412 58335
rect 5363 58295 5412 58301
rect 5406 58292 5412 58295
rect 5464 58292 5470 58344
rect 88163 58335 88221 58341
rect 88163 58301 88175 58335
rect 88209 58332 88221 58335
rect 88574 58332 88580 58344
rect 88209 58304 88580 58332
rect 88209 58301 88221 58304
rect 88163 58295 88221 58301
rect 88574 58292 88580 58304
rect 88632 58292 88638 58344
rect 4876 58234 7912 58256
rect 4876 58182 6618 58234
rect 6670 58182 6682 58234
rect 6734 58182 6746 58234
rect 6798 58182 6810 58234
rect 6862 58182 6874 58234
rect 6926 58182 7912 58234
rect 4876 58160 7912 58182
rect 85284 58234 88596 58256
rect 85284 58182 87210 58234
rect 87262 58182 87274 58234
rect 87326 58182 87338 58234
rect 87390 58182 87402 58234
rect 87454 58182 87466 58234
rect 87518 58182 88596 58234
rect 85284 58160 88596 58182
rect 4876 57690 7912 57712
rect 4876 57638 5882 57690
rect 5934 57638 5946 57690
rect 5998 57638 6010 57690
rect 6062 57638 6074 57690
rect 6126 57638 6138 57690
rect 6190 57638 7912 57690
rect 4876 57616 7912 57638
rect 85284 57690 88596 57712
rect 85284 57638 86474 57690
rect 86526 57638 86538 57690
rect 86590 57638 86602 57690
rect 86654 57638 86666 57690
rect 86718 57638 86730 57690
rect 86782 57638 88596 57690
rect 85284 57616 88596 57638
rect 4876 57146 7912 57168
rect 4876 57094 6618 57146
rect 6670 57094 6682 57146
rect 6734 57094 6746 57146
rect 6798 57094 6810 57146
rect 6862 57094 6874 57146
rect 6926 57094 7912 57146
rect 4876 57072 7912 57094
rect 85284 57146 88596 57168
rect 85284 57094 87210 57146
rect 87262 57094 87274 57146
rect 87326 57094 87338 57146
rect 87390 57094 87402 57146
rect 87454 57094 87466 57146
rect 87518 57094 88596 57146
rect 85284 57072 88596 57094
rect 5363 56975 5421 56981
rect 5363 56941 5375 56975
rect 5409 56972 5421 56975
rect 9914 56972 9920 56984
rect 5409 56944 9920 56972
rect 5409 56941 5421 56944
rect 5363 56935 5421 56941
rect 9914 56932 9920 56944
rect 9972 56932 9978 56984
rect 88163 56975 88221 56981
rect 88163 56941 88175 56975
rect 88209 56972 88221 56975
rect 88574 56972 88580 56984
rect 88209 56944 88580 56972
rect 88209 56941 88221 56944
rect 88163 56935 88221 56941
rect 88574 56932 88580 56944
rect 88632 56932 88638 56984
rect 4302 56864 4308 56916
rect 4360 56904 4366 56916
rect 5161 56907 5219 56913
rect 5161 56904 5173 56907
rect 4360 56876 5173 56904
rect 4360 56864 4366 56876
rect 5161 56873 5173 56876
rect 5207 56904 5219 56907
rect 5501 56907 5559 56913
rect 5501 56904 5513 56907
rect 5207 56876 5513 56904
rect 5207 56873 5219 56876
rect 5161 56867 5219 56873
rect 5501 56873 5513 56876
rect 5547 56873 5559 56907
rect 5501 56867 5559 56873
rect 87562 56864 87568 56916
rect 87620 56904 87626 56916
rect 87957 56907 88015 56913
rect 87957 56904 87969 56907
rect 87620 56876 87969 56904
rect 87620 56864 87626 56876
rect 87957 56873 87969 56876
rect 88003 56873 88015 56907
rect 87957 56867 88015 56873
rect 4876 56602 7912 56624
rect 4876 56550 5882 56602
rect 5934 56550 5946 56602
rect 5998 56550 6010 56602
rect 6062 56550 6074 56602
rect 6126 56550 6138 56602
rect 6190 56550 7912 56602
rect 4876 56528 7912 56550
rect 85284 56602 88596 56624
rect 85284 56550 86474 56602
rect 86526 56550 86538 56602
rect 86590 56550 86602 56602
rect 86654 56550 86666 56602
rect 86718 56550 86730 56602
rect 86782 56550 88596 56602
rect 85284 56528 88596 56550
rect 5363 56363 5421 56369
rect 5363 56329 5375 56363
rect 5409 56360 5421 56363
rect 9914 56360 9920 56372
rect 5409 56332 9920 56360
rect 5409 56329 5421 56332
rect 5363 56323 5421 56329
rect 9914 56320 9920 56332
rect 9972 56320 9978 56372
rect 4302 56252 4308 56304
rect 4360 56292 4366 56304
rect 5161 56295 5219 56301
rect 5161 56292 5173 56295
rect 4360 56264 5173 56292
rect 4360 56252 4366 56264
rect 5161 56261 5173 56264
rect 5207 56292 5219 56295
rect 5501 56295 5559 56301
rect 5501 56292 5513 56295
rect 5207 56264 5513 56292
rect 5207 56261 5219 56264
rect 5161 56255 5219 56261
rect 5501 56261 5513 56264
rect 5547 56261 5559 56295
rect 5501 56255 5559 56261
rect 85814 56252 85820 56304
rect 85872 56292 85878 56304
rect 87957 56295 88015 56301
rect 87957 56292 87969 56295
rect 85872 56264 87969 56292
rect 85872 56252 85878 56264
rect 87957 56261 87969 56264
rect 88003 56261 88015 56295
rect 87957 56255 88015 56261
rect 88206 56165 88212 56168
rect 88163 56159 88212 56165
rect 88163 56125 88175 56159
rect 88209 56125 88212 56159
rect 88163 56119 88212 56125
rect 88206 56116 88212 56119
rect 88264 56116 88270 56168
rect 4876 56058 7912 56080
rect 4876 56006 6618 56058
rect 6670 56006 6682 56058
rect 6734 56006 6746 56058
rect 6798 56006 6810 56058
rect 6862 56006 6874 56058
rect 6926 56006 7912 56058
rect 4876 55984 7912 56006
rect 85284 56058 88596 56080
rect 85284 56006 87210 56058
rect 87262 56006 87274 56058
rect 87326 56006 87338 56058
rect 87390 56006 87402 56058
rect 87454 56006 87466 56058
rect 87518 56006 88596 56058
rect 85284 55984 88596 56006
rect 4876 55514 7912 55536
rect 4876 55462 5882 55514
rect 5934 55462 5946 55514
rect 5998 55462 6010 55514
rect 6062 55462 6074 55514
rect 6126 55462 6138 55514
rect 6190 55462 7912 55514
rect 4876 55440 7912 55462
rect 85284 55514 88596 55536
rect 85284 55462 86474 55514
rect 86526 55462 86538 55514
rect 86590 55462 86602 55514
rect 86654 55462 86666 55514
rect 86718 55462 86730 55514
rect 86782 55462 88596 55514
rect 85284 55440 88596 55462
rect 5363 55275 5421 55281
rect 5363 55241 5375 55275
rect 5409 55272 5421 55275
rect 8534 55272 8540 55284
rect 5409 55244 8540 55272
rect 5409 55241 5421 55244
rect 5363 55235 5421 55241
rect 8534 55232 8540 55244
rect 8592 55232 8598 55284
rect 4302 55164 4308 55216
rect 4360 55204 4366 55216
rect 5161 55207 5219 55213
rect 5161 55204 5173 55207
rect 4360 55176 5173 55204
rect 4360 55164 4366 55176
rect 5161 55173 5173 55176
rect 5207 55204 5219 55207
rect 5501 55207 5559 55213
rect 5501 55204 5513 55207
rect 5207 55176 5513 55204
rect 5207 55173 5219 55176
rect 5161 55167 5219 55173
rect 5501 55173 5513 55176
rect 5547 55173 5559 55207
rect 5501 55167 5559 55173
rect 85814 55164 85820 55216
rect 85872 55204 85878 55216
rect 87957 55207 88015 55213
rect 87957 55204 87969 55207
rect 85872 55176 87969 55204
rect 85872 55164 85878 55176
rect 87957 55173 87969 55176
rect 88003 55173 88015 55207
rect 87957 55167 88015 55173
rect 88206 55077 88212 55080
rect 88163 55071 88212 55077
rect 88163 55037 88175 55071
rect 88209 55037 88212 55071
rect 88163 55031 88212 55037
rect 88206 55028 88212 55031
rect 88264 55028 88270 55080
rect 4876 54970 7912 54992
rect 4876 54918 6618 54970
rect 6670 54918 6682 54970
rect 6734 54918 6746 54970
rect 6798 54918 6810 54970
rect 6862 54918 6874 54970
rect 6926 54918 7912 54970
rect 4876 54896 7912 54918
rect 85284 54970 88596 54992
rect 85284 54918 87210 54970
rect 87262 54918 87274 54970
rect 87326 54918 87338 54970
rect 87390 54918 87402 54970
rect 87454 54918 87466 54970
rect 87518 54918 88596 54970
rect 85284 54896 88596 54918
rect 4876 54426 7912 54448
rect 4876 54374 5882 54426
rect 5934 54374 5946 54426
rect 5998 54374 6010 54426
rect 6062 54374 6074 54426
rect 6126 54374 6138 54426
rect 6190 54374 7912 54426
rect 4876 54352 7912 54374
rect 85284 54426 88596 54448
rect 85284 54374 86474 54426
rect 86526 54374 86538 54426
rect 86590 54374 86602 54426
rect 86654 54374 86666 54426
rect 86718 54374 86730 54426
rect 86782 54374 88596 54426
rect 85284 54352 88596 54374
rect 5363 54187 5421 54193
rect 5363 54153 5375 54187
rect 5409 54184 5421 54187
rect 5682 54184 5688 54196
rect 5409 54156 5688 54184
rect 5409 54153 5421 54156
rect 5363 54147 5421 54153
rect 5682 54144 5688 54156
rect 5740 54144 5746 54196
rect 4302 54076 4308 54128
rect 4360 54116 4366 54128
rect 5161 54119 5219 54125
rect 5161 54116 5173 54119
rect 4360 54088 5173 54116
rect 4360 54076 4366 54088
rect 5161 54085 5173 54088
rect 5207 54116 5219 54119
rect 5501 54119 5559 54125
rect 5501 54116 5513 54119
rect 5207 54088 5513 54116
rect 5207 54085 5219 54088
rect 5161 54079 5219 54085
rect 5501 54085 5513 54088
rect 5547 54085 5559 54119
rect 5501 54079 5559 54085
rect 84526 54076 84532 54128
rect 84584 54116 84590 54128
rect 87957 54119 88015 54125
rect 87957 54116 87969 54119
rect 84584 54088 87969 54116
rect 84584 54076 84590 54088
rect 87957 54085 87969 54088
rect 88003 54085 88015 54119
rect 88206 54116 88212 54128
rect 87957 54079 88015 54085
rect 88178 54076 88212 54116
rect 88264 54076 88270 54128
rect 88178 53989 88206 54076
rect 88163 53983 88221 53989
rect 88163 53949 88175 53983
rect 88209 53949 88221 53983
rect 88163 53943 88221 53949
rect 4876 53882 7912 53904
rect 4876 53830 6618 53882
rect 6670 53830 6682 53882
rect 6734 53830 6746 53882
rect 6798 53830 6810 53882
rect 6862 53830 6874 53882
rect 6926 53830 7912 53882
rect 4876 53808 7912 53830
rect 85284 53882 88596 53904
rect 85284 53830 87210 53882
rect 87262 53830 87274 53882
rect 87326 53830 87338 53882
rect 87390 53830 87402 53882
rect 87454 53830 87466 53882
rect 87518 53830 88596 53882
rect 85284 53808 88596 53830
rect 4876 53338 7912 53360
rect 4876 53286 5882 53338
rect 5934 53286 5946 53338
rect 5998 53286 6010 53338
rect 6062 53286 6074 53338
rect 6126 53286 6138 53338
rect 6190 53286 7912 53338
rect 4876 53264 7912 53286
rect 85284 53338 88596 53360
rect 85284 53286 86474 53338
rect 86526 53286 86538 53338
rect 86590 53286 86602 53338
rect 86654 53286 86666 53338
rect 86718 53286 86730 53338
rect 86782 53286 88596 53338
rect 85284 53264 88596 53286
rect 5363 53099 5421 53105
rect 5363 53065 5375 53099
rect 5409 53096 5421 53099
rect 8534 53096 8540 53108
rect 5409 53068 8540 53096
rect 5409 53065 5421 53068
rect 5363 53059 5421 53065
rect 8534 53056 8540 53068
rect 8592 53056 8598 53108
rect 4302 52988 4308 53040
rect 4360 53028 4366 53040
rect 5161 53031 5219 53037
rect 5161 53028 5173 53031
rect 4360 53000 5173 53028
rect 4360 52988 4366 53000
rect 5161 52997 5173 53000
rect 5207 53028 5219 53031
rect 5501 53031 5559 53037
rect 5501 53028 5513 53031
rect 5207 53000 5513 53028
rect 5207 52997 5219 53000
rect 5161 52991 5219 52997
rect 5501 52997 5513 53000
rect 5547 52997 5559 53031
rect 5501 52991 5559 52997
rect 87562 52988 87568 53040
rect 87620 53028 87626 53040
rect 87957 53031 88015 53037
rect 87957 53028 87969 53031
rect 87620 53000 87969 53028
rect 87620 52988 87626 53000
rect 87957 52997 87969 53000
rect 88003 52997 88015 53031
rect 87957 52991 88015 52997
rect 88206 52901 88212 52904
rect 88163 52895 88212 52901
rect 88163 52861 88175 52895
rect 88209 52861 88212 52895
rect 88163 52855 88212 52861
rect 88206 52852 88212 52855
rect 88264 52852 88270 52904
rect 4876 52794 7912 52816
rect 4876 52742 6618 52794
rect 6670 52742 6682 52794
rect 6734 52742 6746 52794
rect 6798 52742 6810 52794
rect 6862 52742 6874 52794
rect 6926 52742 7912 52794
rect 4876 52720 7912 52742
rect 85284 52794 88596 52816
rect 85284 52742 87210 52794
rect 87262 52742 87274 52794
rect 87326 52742 87338 52794
rect 87390 52742 87402 52794
rect 87454 52742 87466 52794
rect 87518 52742 88596 52794
rect 85284 52720 88596 52742
rect 4876 52250 7912 52272
rect 4876 52198 5882 52250
rect 5934 52198 5946 52250
rect 5998 52198 6010 52250
rect 6062 52198 6074 52250
rect 6126 52198 6138 52250
rect 6190 52198 7912 52250
rect 4876 52176 7912 52198
rect 85284 52250 88596 52272
rect 85284 52198 86474 52250
rect 86526 52198 86538 52250
rect 86590 52198 86602 52250
rect 86654 52198 86666 52250
rect 86718 52198 86730 52250
rect 86782 52198 88596 52250
rect 85284 52176 88596 52198
rect 4876 51706 7912 51728
rect 4876 51654 6618 51706
rect 6670 51654 6682 51706
rect 6734 51654 6746 51706
rect 6798 51654 6810 51706
rect 6862 51654 6874 51706
rect 6926 51654 7912 51706
rect 4876 51632 7912 51654
rect 85284 51706 88596 51728
rect 85284 51654 87210 51706
rect 87262 51654 87274 51706
rect 87326 51654 87338 51706
rect 87390 51654 87402 51706
rect 87454 51654 87466 51706
rect 87518 51654 88596 51706
rect 85284 51632 88596 51654
rect 5363 51535 5421 51541
rect 5363 51501 5375 51535
rect 5409 51532 5421 51535
rect 8534 51532 8540 51544
rect 5409 51504 8540 51532
rect 5409 51501 5421 51504
rect 5363 51495 5421 51501
rect 8534 51492 8540 51504
rect 8592 51492 8598 51544
rect 4302 51424 4308 51476
rect 4360 51464 4366 51476
rect 5161 51467 5219 51473
rect 5161 51464 5173 51467
rect 4360 51436 5173 51464
rect 4360 51424 4366 51436
rect 5161 51433 5173 51436
rect 5207 51464 5219 51467
rect 5501 51467 5559 51473
rect 5501 51464 5513 51467
rect 5207 51436 5513 51464
rect 5207 51433 5219 51436
rect 5161 51427 5219 51433
rect 5501 51433 5513 51436
rect 5547 51433 5559 51467
rect 5501 51427 5559 51433
rect 87562 51424 87568 51476
rect 87620 51464 87626 51476
rect 87957 51467 88015 51473
rect 87957 51464 87969 51467
rect 87620 51436 87969 51464
rect 87620 51424 87626 51436
rect 87957 51433 87969 51436
rect 88003 51433 88015 51467
rect 87957 51427 88015 51433
rect 88206 51337 88212 51340
rect 88163 51331 88212 51337
rect 88163 51297 88175 51331
rect 88209 51297 88212 51331
rect 88163 51291 88212 51297
rect 88206 51288 88212 51291
rect 88264 51288 88270 51340
rect 4876 51162 7912 51184
rect 4876 51110 5882 51162
rect 5934 51110 5946 51162
rect 5998 51110 6010 51162
rect 6062 51110 6074 51162
rect 6126 51110 6138 51162
rect 6190 51110 7912 51162
rect 4876 51088 7912 51110
rect 85284 51162 88596 51184
rect 85284 51110 86474 51162
rect 86526 51110 86538 51162
rect 86590 51110 86602 51162
rect 86654 51110 86666 51162
rect 86718 51110 86730 51162
rect 86782 51110 88596 51162
rect 85284 51088 88596 51110
rect 85630 50676 85636 50728
rect 85688 50676 85694 50728
rect 4876 50618 7912 50640
rect 4876 50566 6618 50618
rect 6670 50566 6682 50618
rect 6734 50566 6746 50618
rect 6798 50566 6810 50618
rect 6862 50566 6874 50618
rect 6926 50566 7912 50618
rect 4876 50544 7912 50566
rect 85284 50618 88596 50640
rect 85284 50566 87210 50618
rect 87262 50566 87274 50618
rect 87326 50566 87338 50618
rect 87390 50566 87402 50618
rect 87454 50566 87466 50618
rect 87518 50566 88596 50618
rect 85284 50544 88596 50566
rect 4876 50074 7912 50096
rect 4876 50022 5882 50074
rect 5934 50022 5946 50074
rect 5998 50022 6010 50074
rect 6062 50022 6074 50074
rect 6126 50022 6138 50074
rect 6190 50022 7912 50074
rect 4876 50000 7912 50022
rect 85284 50074 88596 50096
rect 85284 50022 86474 50074
rect 86526 50022 86538 50074
rect 86590 50022 86602 50074
rect 86654 50022 86666 50074
rect 86718 50022 86730 50074
rect 86782 50022 88596 50074
rect 85284 50000 88596 50022
rect 85630 49588 85636 49640
rect 85688 49588 85694 49640
rect 4876 49530 7912 49552
rect 4876 49478 6618 49530
rect 6670 49478 6682 49530
rect 6734 49478 6746 49530
rect 6798 49478 6810 49530
rect 6862 49478 6874 49530
rect 6926 49478 7912 49530
rect 4876 49456 7912 49478
rect 85284 49530 88596 49552
rect 85284 49478 87210 49530
rect 87262 49478 87274 49530
rect 87326 49478 87338 49530
rect 87390 49478 87402 49530
rect 87454 49478 87466 49530
rect 87518 49478 88596 49530
rect 85284 49456 88596 49478
rect 4876 48986 7912 49008
rect 4876 48934 5882 48986
rect 5934 48934 5946 48986
rect 5998 48934 6010 48986
rect 6062 48934 6074 48986
rect 6126 48934 6138 48986
rect 6190 48934 7912 48986
rect 4876 48912 7912 48934
rect 85284 48986 88596 49008
rect 85284 48934 86474 48986
rect 86526 48934 86538 48986
rect 86590 48934 86602 48986
rect 86654 48934 86666 48986
rect 86718 48934 86730 48986
rect 86782 48934 88596 48986
rect 85284 48912 88596 48934
rect 88206 48636 88212 48688
rect 88264 48636 88270 48688
rect 85354 48568 85360 48620
rect 85412 48608 85418 48620
rect 85633 48611 85691 48617
rect 85633 48608 85645 48611
rect 85412 48580 85645 48608
rect 85412 48568 85418 48580
rect 85633 48577 85645 48580
rect 85679 48577 85691 48611
rect 85633 48571 85691 48577
rect 4876 48442 7912 48464
rect 4876 48390 6618 48442
rect 6670 48390 6682 48442
rect 6734 48390 6746 48442
rect 6798 48390 6810 48442
rect 6862 48390 6874 48442
rect 6926 48390 7912 48442
rect 4876 48368 7912 48390
rect 85284 48442 88596 48464
rect 85284 48390 87210 48442
rect 87262 48390 87274 48442
rect 87326 48390 87338 48442
rect 87390 48390 87402 48442
rect 87454 48390 87466 48442
rect 87518 48390 88596 48442
rect 85284 48368 88596 48390
rect 88206 47956 88212 48008
rect 88264 47956 88270 48008
rect 4876 47898 7912 47920
rect 4876 47846 5882 47898
rect 5934 47846 5946 47898
rect 5998 47846 6010 47898
rect 6062 47846 6074 47898
rect 6126 47846 6138 47898
rect 6190 47846 7912 47898
rect 4876 47824 7912 47846
rect 85284 47898 88596 47920
rect 85284 47846 86474 47898
rect 86526 47846 86538 47898
rect 86590 47846 86602 47898
rect 86654 47846 86666 47898
rect 86718 47846 86730 47898
rect 86782 47846 88596 47898
rect 85284 47824 88596 47846
rect 85814 47548 85820 47600
rect 85872 47588 85878 47600
rect 87957 47591 88015 47597
rect 87957 47588 87969 47591
rect 85872 47560 87969 47588
rect 85872 47548 85878 47560
rect 87957 47557 87969 47560
rect 88003 47557 88015 47591
rect 87957 47551 88015 47557
rect 88206 47461 88212 47464
rect 88163 47455 88212 47461
rect 88163 47421 88175 47455
rect 88209 47421 88212 47455
rect 88163 47415 88212 47421
rect 88206 47412 88212 47415
rect 88264 47412 88270 47464
rect 4876 47354 7912 47376
rect 4876 47302 6618 47354
rect 6670 47302 6682 47354
rect 6734 47302 6746 47354
rect 6798 47302 6810 47354
rect 6862 47302 6874 47354
rect 6926 47302 7912 47354
rect 4876 47280 7912 47302
rect 85284 47354 88596 47376
rect 85284 47302 87210 47354
rect 87262 47302 87274 47354
rect 87326 47302 87338 47354
rect 87390 47302 87402 47354
rect 87454 47302 87466 47354
rect 87518 47302 88596 47354
rect 85284 47280 88596 47302
rect 88206 46868 88212 46920
rect 88264 46868 88270 46920
rect 4876 46810 7912 46832
rect 4876 46758 5882 46810
rect 5934 46758 5946 46810
rect 5998 46758 6010 46810
rect 6062 46758 6074 46810
rect 6126 46758 6138 46810
rect 6190 46758 7912 46810
rect 4876 46736 7912 46758
rect 85284 46810 88596 46832
rect 85284 46758 86474 46810
rect 86526 46758 86538 46810
rect 86590 46758 86602 46810
rect 86654 46758 86666 46810
rect 86718 46758 86730 46810
rect 86782 46758 88596 46810
rect 85284 46736 88596 46758
rect 4876 46266 7912 46288
rect 4876 46214 6618 46266
rect 6670 46214 6682 46266
rect 6734 46214 6746 46266
rect 6798 46214 6810 46266
rect 6862 46214 6874 46266
rect 6926 46214 7912 46266
rect 4876 46192 7912 46214
rect 85284 46266 88596 46288
rect 85284 46214 87210 46266
rect 87262 46214 87274 46266
rect 87326 46214 87338 46266
rect 87390 46214 87402 46266
rect 87454 46214 87466 46266
rect 87518 46214 88596 46266
rect 85284 46192 88596 46214
rect 46990 45984 46996 46036
rect 47048 46024 47054 46036
rect 47048 45996 48554 46024
rect 47048 45984 47054 45996
rect 48526 45956 48554 45996
rect 50164 45956 50170 45968
rect 48526 45928 50170 45956
rect 50164 45916 50170 45928
rect 50222 45956 50228 45968
rect 51130 45956 51136 45968
rect 50222 45928 51136 45956
rect 50222 45916 50228 45928
rect 51130 45916 51136 45928
rect 51188 45916 51194 45968
rect 10558 45888 10564 45900
rect 9932 45860 10564 45888
rect 4876 45722 7912 45744
rect 4876 45670 5882 45722
rect 5934 45670 5946 45722
rect 5998 45670 6010 45722
rect 6062 45670 6074 45722
rect 6126 45670 6138 45722
rect 6190 45670 7912 45722
rect 4876 45648 7912 45670
rect 7338 45508 7344 45560
rect 7396 45548 7402 45560
rect 9932 45548 9960 45860
rect 10558 45848 10564 45860
rect 10616 45848 10622 45900
rect 46438 45848 46444 45900
rect 46496 45888 46502 45900
rect 51268 45888 51274 45900
rect 46496 45860 51274 45888
rect 46496 45848 46502 45860
rect 51268 45848 51274 45860
rect 51326 45888 51332 45900
rect 85814 45888 85820 45900
rect 51326 45860 85820 45888
rect 51326 45848 51332 45860
rect 85814 45848 85820 45860
rect 85872 45848 85878 45900
rect 85284 45722 88596 45744
rect 85284 45670 86474 45722
rect 86526 45670 86538 45722
rect 86590 45670 86602 45722
rect 86654 45670 86666 45722
rect 86718 45670 86730 45722
rect 86782 45670 88596 45722
rect 85284 45648 88596 45670
rect 7396 45520 9960 45548
rect 7396 45508 7402 45520
rect 85814 45508 85820 45560
rect 85872 45508 85878 45560
rect 7157 45483 7215 45489
rect 7157 45449 7169 45483
rect 7203 45480 7215 45483
rect 8994 45480 9000 45492
rect 7203 45452 9000 45480
rect 7203 45449 7215 45452
rect 7157 45443 7215 45449
rect 8994 45440 9000 45452
rect 9052 45440 9058 45492
rect 4302 45372 4308 45424
rect 4360 45412 4366 45424
rect 5161 45415 5219 45421
rect 5161 45412 5173 45415
rect 4360 45384 5173 45412
rect 4360 45372 4366 45384
rect 5161 45381 5173 45384
rect 5207 45412 5219 45415
rect 5501 45415 5559 45421
rect 5501 45412 5513 45415
rect 5207 45384 5513 45412
rect 5207 45381 5219 45384
rect 5161 45375 5219 45381
rect 5501 45381 5513 45384
rect 5547 45381 5559 45415
rect 5501 45375 5559 45381
rect 85998 45372 86004 45424
rect 86056 45372 86062 45424
rect 88206 45372 88212 45424
rect 88264 45372 88270 45424
rect 5363 45347 5421 45353
rect 5363 45313 5375 45347
rect 5409 45344 5421 45347
rect 5682 45344 5688 45356
rect 5409 45316 5688 45344
rect 5409 45313 5421 45316
rect 5363 45307 5421 45313
rect 5682 45304 5688 45316
rect 5740 45304 5746 45356
rect 85630 45236 85636 45288
rect 85688 45236 85694 45288
rect 86182 45236 86188 45288
rect 86240 45236 86246 45288
rect 4876 45178 7912 45200
rect 4876 45126 6618 45178
rect 6670 45126 6682 45178
rect 6734 45126 6746 45178
rect 6798 45126 6810 45178
rect 6862 45126 6874 45178
rect 6926 45126 7912 45178
rect 4876 45104 7912 45126
rect 85284 45178 88596 45200
rect 85284 45126 87210 45178
rect 87262 45126 87274 45178
rect 87326 45126 87338 45178
rect 87390 45126 87402 45178
rect 87454 45126 87466 45178
rect 87518 45126 88596 45178
rect 85284 45104 88596 45126
rect 7525 45007 7583 45013
rect 7525 44973 7537 45007
rect 7571 45004 7583 45007
rect 7614 45004 7620 45016
rect 7571 44976 7620 45004
rect 7571 44973 7583 44976
rect 7525 44967 7583 44973
rect 7614 44964 7620 44976
rect 7672 44964 7678 45016
rect 5409 44939 5467 44945
rect 5409 44905 5421 44939
rect 5455 44936 5467 44939
rect 8534 44936 8540 44948
rect 5455 44908 8540 44936
rect 5455 44905 5467 44908
rect 5409 44899 5467 44905
rect 8534 44896 8540 44908
rect 8592 44896 8598 44948
rect 4210 44692 4216 44744
rect 4268 44732 4274 44744
rect 5245 44735 5303 44741
rect 5245 44732 5257 44735
rect 4268 44704 5257 44732
rect 4268 44692 4274 44704
rect 5245 44701 5257 44704
rect 5291 44701 5303 44735
rect 5245 44695 5303 44701
rect 88206 44692 88212 44744
rect 88264 44692 88270 44744
rect 4876 44634 7912 44656
rect 4876 44582 5882 44634
rect 5934 44582 5946 44634
rect 5998 44582 6010 44634
rect 6062 44582 6074 44634
rect 6126 44582 6138 44634
rect 6190 44582 7912 44634
rect 4876 44560 7912 44582
rect 85284 44634 88596 44656
rect 85284 44582 86474 44634
rect 86526 44582 86538 44634
rect 86590 44582 86602 44634
rect 86654 44582 86666 44634
rect 86718 44582 86730 44634
rect 86782 44582 88596 44634
rect 85284 44560 88596 44582
rect 83606 44352 83612 44404
rect 83664 44392 83670 44404
rect 88049 44395 88107 44401
rect 88049 44392 88061 44395
rect 83664 44364 88061 44392
rect 83664 44352 83670 44364
rect 88049 44361 88061 44364
rect 88095 44361 88107 44395
rect 88049 44355 88107 44361
rect 87749 44327 87807 44333
rect 87749 44293 87761 44327
rect 87795 44324 87807 44327
rect 88206 44324 88212 44336
rect 87795 44296 88212 44324
rect 87795 44293 87807 44296
rect 87749 44287 87807 44293
rect 88206 44284 88212 44296
rect 88264 44284 88270 44336
rect 4876 44090 7912 44112
rect 4876 44038 6618 44090
rect 6670 44038 6682 44090
rect 6734 44038 6746 44090
rect 6798 44038 6810 44090
rect 6862 44038 6874 44090
rect 6926 44038 7912 44090
rect 4876 44016 7912 44038
rect 85284 44090 88596 44112
rect 85284 44038 87210 44090
rect 87262 44038 87274 44090
rect 87326 44038 87338 44090
rect 87390 44038 87402 44090
rect 87454 44038 87466 44090
rect 87518 44038 88596 44090
rect 85284 44016 88596 44038
rect 4876 43546 7912 43568
rect 4876 43494 5882 43546
rect 5934 43494 5946 43546
rect 5998 43494 6010 43546
rect 6062 43494 6074 43546
rect 6126 43494 6138 43546
rect 6190 43494 7912 43546
rect 4876 43472 7912 43494
rect 85284 43546 88596 43568
rect 85284 43494 86474 43546
rect 86526 43494 86538 43546
rect 86590 43494 86602 43546
rect 86654 43494 86666 43546
rect 86718 43494 86730 43546
rect 86782 43494 88596 43546
rect 85284 43472 88596 43494
rect 85814 43332 85820 43384
rect 85872 43372 85878 43384
rect 88049 43375 88107 43381
rect 88049 43372 88061 43375
rect 85872 43344 88061 43372
rect 85872 43332 85878 43344
rect 88049 43341 88061 43344
rect 88095 43341 88107 43375
rect 88049 43335 88107 43341
rect 4118 43196 4124 43248
rect 4176 43236 4182 43248
rect 5245 43239 5303 43245
rect 5245 43236 5257 43239
rect 4176 43208 5257 43236
rect 4176 43196 4182 43208
rect 5245 43205 5257 43208
rect 5291 43205 5303 43239
rect 5245 43199 5303 43205
rect 5409 43239 5467 43245
rect 5409 43205 5421 43239
rect 5455 43236 5467 43239
rect 8534 43236 8540 43248
rect 5455 43208 8540 43236
rect 5455 43205 5467 43208
rect 5409 43199 5467 43205
rect 8534 43196 8540 43208
rect 8592 43196 8598 43248
rect 87749 43239 87807 43245
rect 87749 43205 87761 43239
rect 87795 43236 87807 43239
rect 88206 43236 88212 43248
rect 87795 43208 88212 43236
rect 87795 43205 87807 43208
rect 87749 43199 87807 43205
rect 88206 43196 88212 43208
rect 88264 43196 88270 43248
rect 4876 43002 7912 43024
rect 4876 42950 6618 43002
rect 6670 42950 6682 43002
rect 6734 42950 6746 43002
rect 6798 42950 6810 43002
rect 6862 42950 6874 43002
rect 6926 42950 7912 43002
rect 4876 42928 7912 42950
rect 85284 43002 88596 43024
rect 85284 42950 87210 43002
rect 87262 42950 87274 43002
rect 87326 42950 87338 43002
rect 87390 42950 87402 43002
rect 87454 42950 87466 43002
rect 87518 42950 88596 43002
rect 85284 42928 88596 42950
rect 5409 42763 5467 42769
rect 5409 42729 5421 42763
rect 5455 42760 5467 42763
rect 8534 42760 8540 42772
rect 5455 42732 8540 42760
rect 5455 42729 5467 42732
rect 5409 42723 5467 42729
rect 8534 42720 8540 42732
rect 8592 42720 8598 42772
rect 87933 42763 87991 42769
rect 87933 42729 87945 42763
rect 87979 42760 87991 42763
rect 88206 42760 88212 42772
rect 87979 42732 88212 42760
rect 87979 42729 87991 42732
rect 87933 42723 87991 42729
rect 88206 42720 88212 42732
rect 88264 42720 88270 42772
rect 85814 42584 85820 42636
rect 85872 42624 85878 42636
rect 88049 42627 88107 42633
rect 88049 42624 88061 42627
rect 85872 42596 88061 42624
rect 85872 42584 85878 42596
rect 88049 42593 88061 42596
rect 88095 42593 88107 42627
rect 88049 42587 88107 42593
rect 4118 42516 4124 42568
rect 4176 42556 4182 42568
rect 5245 42559 5303 42565
rect 5245 42556 5257 42559
rect 4176 42528 5257 42556
rect 4176 42516 4182 42528
rect 5245 42525 5257 42528
rect 5291 42525 5303 42559
rect 5245 42519 5303 42525
rect 4876 42458 7912 42480
rect 4876 42406 5882 42458
rect 5934 42406 5946 42458
rect 5998 42406 6010 42458
rect 6062 42406 6074 42458
rect 6126 42406 6138 42458
rect 6190 42406 7912 42458
rect 4876 42384 7912 42406
rect 85284 42458 88596 42480
rect 85284 42406 86474 42458
rect 86526 42406 86538 42458
rect 86590 42406 86602 42458
rect 86654 42406 86666 42458
rect 86718 42406 86730 42458
rect 86782 42406 88596 42458
rect 85284 42384 88596 42406
rect 4876 41914 7912 41936
rect 4876 41862 6618 41914
rect 6670 41862 6682 41914
rect 6734 41862 6746 41914
rect 6798 41862 6810 41914
rect 6862 41862 6874 41914
rect 6926 41862 7912 41914
rect 4876 41840 7912 41862
rect 85284 41914 88596 41936
rect 85284 41862 87210 41914
rect 87262 41862 87274 41914
rect 87326 41862 87338 41914
rect 87390 41862 87402 41914
rect 87454 41862 87466 41914
rect 87518 41862 88596 41914
rect 85284 41840 88596 41862
rect 4118 41632 4124 41684
rect 4176 41672 4182 41684
rect 5245 41675 5303 41681
rect 5245 41672 5257 41675
rect 4176 41644 5257 41672
rect 4176 41632 4182 41644
rect 5245 41641 5257 41644
rect 5291 41641 5303 41675
rect 5245 41635 5303 41641
rect 5406 41632 5412 41684
rect 5464 41632 5470 41684
rect 87562 41632 87568 41684
rect 87620 41672 87626 41684
rect 88049 41675 88107 41681
rect 88049 41672 88061 41675
rect 87620 41644 88061 41672
rect 87620 41632 87626 41644
rect 88049 41641 88061 41644
rect 88095 41641 88107 41675
rect 88049 41635 88107 41641
rect 88206 41632 88212 41684
rect 88264 41632 88270 41684
rect 87933 41607 87991 41613
rect 87933 41573 87945 41607
rect 87979 41604 87991 41607
rect 88224 41604 88252 41632
rect 87979 41576 88252 41604
rect 87979 41573 87991 41576
rect 87933 41567 87991 41573
rect 4876 41370 7912 41392
rect 4876 41318 5882 41370
rect 5934 41318 5946 41370
rect 5998 41318 6010 41370
rect 6062 41318 6074 41370
rect 6126 41318 6138 41370
rect 6190 41318 7912 41370
rect 4876 41296 7912 41318
rect 85284 41370 88596 41392
rect 85284 41318 86474 41370
rect 86526 41318 86538 41370
rect 86590 41318 86602 41370
rect 86654 41318 86666 41370
rect 86718 41318 86730 41370
rect 86782 41318 88596 41370
rect 85284 41296 88596 41318
rect 4876 40826 7912 40848
rect 4876 40774 6618 40826
rect 6670 40774 6682 40826
rect 6734 40774 6746 40826
rect 6798 40774 6810 40826
rect 6862 40774 6874 40826
rect 6926 40774 7912 40826
rect 4876 40752 7912 40774
rect 85284 40826 88596 40848
rect 85284 40774 87210 40826
rect 87262 40774 87274 40826
rect 87326 40774 87338 40826
rect 87390 40774 87402 40826
rect 87454 40774 87466 40826
rect 87518 40774 88596 40826
rect 85284 40752 88596 40774
rect 5409 40587 5467 40593
rect 5409 40553 5421 40587
rect 5455 40584 5467 40587
rect 8534 40584 8540 40596
rect 5455 40556 8540 40584
rect 5455 40553 5467 40556
rect 5409 40547 5467 40553
rect 8534 40544 8540 40556
rect 8592 40544 8598 40596
rect 87930 40476 87936 40528
rect 87988 40476 87994 40528
rect 88206 40476 88212 40528
rect 88264 40476 88270 40528
rect 3934 40408 3940 40460
rect 3992 40448 3998 40460
rect 5245 40451 5303 40457
rect 5245 40448 5257 40451
rect 3992 40420 5257 40448
rect 3992 40408 3998 40420
rect 5245 40417 5257 40420
rect 5291 40417 5303 40451
rect 5245 40411 5303 40417
rect 4876 40282 7912 40304
rect 4876 40230 5882 40282
rect 5934 40230 5946 40282
rect 5998 40230 6010 40282
rect 6062 40230 6074 40282
rect 6126 40230 6138 40282
rect 6190 40230 7912 40282
rect 4876 40208 7912 40230
rect 85284 40282 88596 40304
rect 85284 40230 86474 40282
rect 86526 40230 86538 40282
rect 86590 40230 86602 40282
rect 86654 40230 86666 40282
rect 86718 40230 86730 40282
rect 86782 40230 88596 40282
rect 85284 40208 88596 40230
rect 88206 40068 88212 40120
rect 88264 40068 88270 40120
rect 4876 39738 7912 39760
rect 4876 39686 6618 39738
rect 6670 39686 6682 39738
rect 6734 39686 6746 39738
rect 6798 39686 6810 39738
rect 6862 39686 6874 39738
rect 6926 39686 7912 39738
rect 4876 39664 7912 39686
rect 85284 39738 88596 39760
rect 85284 39686 87210 39738
rect 87262 39686 87274 39738
rect 87326 39686 87338 39738
rect 87390 39686 87402 39738
rect 87454 39686 87466 39738
rect 87518 39686 88596 39738
rect 85284 39664 88596 39686
rect 5409 39499 5467 39505
rect 5409 39465 5421 39499
rect 5455 39496 5467 39499
rect 8534 39496 8540 39508
rect 5455 39468 8540 39496
rect 5455 39465 5467 39468
rect 5409 39459 5467 39465
rect 8534 39456 8540 39468
rect 8592 39456 8598 39508
rect 87841 39499 87899 39505
rect 87841 39465 87853 39499
rect 87887 39496 87899 39499
rect 88206 39496 88212 39508
rect 87887 39468 88212 39496
rect 87887 39465 87899 39468
rect 87841 39459 87899 39465
rect 88206 39456 88212 39468
rect 88264 39456 88270 39508
rect 87562 39320 87568 39372
rect 87620 39360 87626 39372
rect 88045 39363 88103 39369
rect 88045 39360 88057 39363
rect 87620 39332 88057 39360
rect 87620 39320 87626 39332
rect 88045 39329 88057 39332
rect 88091 39329 88103 39363
rect 88045 39323 88103 39329
rect 4210 39252 4216 39304
rect 4268 39292 4274 39304
rect 5245 39295 5303 39301
rect 5245 39292 5257 39295
rect 4268 39264 5257 39292
rect 4268 39252 4274 39264
rect 5245 39261 5257 39264
rect 5291 39261 5303 39295
rect 5245 39255 5303 39261
rect 4876 39194 7912 39216
rect 4876 39142 5882 39194
rect 5934 39142 5946 39194
rect 5998 39142 6010 39194
rect 6062 39142 6074 39194
rect 6126 39142 6138 39194
rect 6190 39142 7912 39194
rect 4876 39120 7912 39142
rect 85284 39194 88596 39216
rect 85284 39142 86474 39194
rect 86526 39142 86538 39194
rect 86590 39142 86602 39194
rect 86654 39142 86666 39194
rect 86718 39142 86730 39194
rect 86782 39142 88596 39194
rect 85284 39120 88596 39142
rect 4876 38650 7912 38672
rect 4876 38598 6618 38650
rect 6670 38598 6682 38650
rect 6734 38598 6746 38650
rect 6798 38598 6810 38650
rect 6862 38598 6874 38650
rect 6926 38598 7912 38650
rect 4876 38576 7912 38598
rect 85284 38650 88596 38672
rect 85284 38598 87210 38650
rect 87262 38598 87274 38650
rect 87326 38598 87338 38650
rect 87390 38598 87402 38650
rect 87454 38598 87466 38650
rect 87518 38598 88596 38650
rect 85284 38576 88596 38598
rect 4876 38106 7912 38128
rect 4876 38054 5882 38106
rect 5934 38054 5946 38106
rect 5998 38054 6010 38106
rect 6062 38054 6074 38106
rect 6126 38054 6138 38106
rect 6190 38054 7912 38106
rect 4876 38032 7912 38054
rect 85284 38106 88596 38128
rect 85284 38054 86474 38106
rect 86526 38054 86538 38106
rect 86590 38054 86602 38106
rect 86654 38054 86666 38106
rect 86718 38054 86730 38106
rect 86782 38054 88596 38106
rect 85284 38032 88596 38054
rect 85814 37892 85820 37944
rect 85872 37932 85878 37944
rect 88045 37935 88103 37941
rect 88045 37932 88057 37935
rect 85872 37904 88057 37932
rect 85872 37892 85878 37904
rect 88045 37901 88057 37904
rect 88091 37901 88103 37935
rect 88045 37895 88103 37901
rect 4210 37756 4216 37808
rect 4268 37796 4274 37808
rect 5245 37799 5303 37805
rect 5245 37796 5257 37799
rect 4268 37768 5257 37796
rect 4268 37756 4274 37768
rect 5245 37765 5257 37768
rect 5291 37765 5303 37799
rect 5245 37759 5303 37765
rect 5409 37799 5467 37805
rect 5409 37765 5421 37799
rect 5455 37796 5467 37799
rect 8534 37796 8540 37808
rect 5455 37768 8540 37796
rect 5455 37765 5467 37768
rect 5409 37759 5467 37765
rect 8534 37756 8540 37768
rect 8592 37756 8598 37808
rect 87749 37799 87807 37805
rect 87749 37765 87761 37799
rect 87795 37796 87807 37799
rect 88206 37796 88212 37808
rect 87795 37768 88212 37796
rect 87795 37765 87807 37768
rect 87749 37759 87807 37765
rect 88206 37756 88212 37768
rect 88264 37756 88270 37808
rect 4876 37562 7912 37584
rect 4876 37510 6618 37562
rect 6670 37510 6682 37562
rect 6734 37510 6746 37562
rect 6798 37510 6810 37562
rect 6862 37510 6874 37562
rect 6926 37510 7912 37562
rect 4876 37488 7912 37510
rect 85284 37562 88596 37584
rect 85284 37510 87210 37562
rect 87262 37510 87274 37562
rect 87326 37510 87338 37562
rect 87390 37510 87402 37562
rect 87454 37510 87466 37562
rect 87518 37510 88596 37562
rect 85284 37488 88596 37510
rect 5409 37323 5467 37329
rect 5409 37289 5421 37323
rect 5455 37320 5467 37323
rect 8534 37320 8540 37332
rect 5455 37292 8540 37320
rect 5455 37289 5467 37292
rect 5409 37283 5467 37289
rect 8534 37280 8540 37292
rect 8592 37280 8598 37332
rect 87933 37323 87991 37329
rect 87933 37289 87945 37323
rect 87979 37320 87991 37323
rect 88206 37320 88212 37332
rect 87979 37292 88212 37320
rect 87979 37289 87991 37292
rect 87933 37283 87991 37289
rect 88206 37280 88212 37292
rect 88264 37280 88270 37332
rect 85814 37144 85820 37196
rect 85872 37184 85878 37196
rect 88050 37187 88108 37193
rect 88050 37184 88062 37187
rect 85872 37156 88062 37184
rect 85872 37144 85878 37156
rect 88050 37153 88062 37156
rect 88096 37153 88108 37187
rect 88050 37147 88108 37153
rect 4118 37076 4124 37128
rect 4176 37116 4182 37128
rect 5245 37119 5303 37125
rect 5245 37116 5257 37119
rect 4176 37088 5257 37116
rect 4176 37076 4182 37088
rect 5245 37085 5257 37088
rect 5291 37085 5303 37119
rect 5245 37079 5303 37085
rect 4876 37018 7912 37040
rect 4876 36966 5882 37018
rect 5934 36966 5946 37018
rect 5998 36966 6010 37018
rect 6062 36966 6074 37018
rect 6126 36966 6138 37018
rect 6190 36966 7912 37018
rect 4876 36944 7912 36966
rect 85284 37018 88596 37040
rect 85284 36966 86474 37018
rect 86526 36966 86538 37018
rect 86590 36966 86602 37018
rect 86654 36966 86666 37018
rect 86718 36966 86730 37018
rect 86782 36966 88596 37018
rect 85284 36944 88596 36966
rect 4876 36474 7912 36496
rect 4876 36422 6618 36474
rect 6670 36422 6682 36474
rect 6734 36422 6746 36474
rect 6798 36422 6810 36474
rect 6862 36422 6874 36474
rect 6926 36422 7912 36474
rect 4876 36400 7912 36422
rect 85284 36474 88596 36496
rect 85284 36422 87210 36474
rect 87262 36422 87274 36474
rect 87326 36422 87338 36474
rect 87390 36422 87402 36474
rect 87454 36422 87466 36474
rect 87518 36422 88596 36474
rect 85284 36400 88596 36422
rect 5406 36192 5412 36244
rect 5464 36192 5470 36244
rect 87933 36235 87991 36241
rect 87933 36201 87945 36235
rect 87979 36232 87991 36235
rect 88209 36235 88267 36241
rect 88209 36232 88221 36235
rect 87979 36204 88221 36232
rect 87979 36201 87991 36204
rect 87933 36195 87991 36201
rect 88209 36201 88221 36204
rect 88255 36232 88267 36235
rect 88574 36232 88580 36244
rect 88255 36204 88580 36232
rect 88255 36201 88267 36204
rect 88209 36195 88267 36201
rect 88574 36192 88580 36204
rect 88632 36192 88638 36244
rect 4118 36124 4124 36176
rect 4176 36164 4182 36176
rect 5245 36167 5303 36173
rect 5245 36164 5257 36167
rect 4176 36136 5257 36164
rect 4176 36124 4182 36136
rect 5245 36133 5257 36136
rect 5291 36133 5303 36167
rect 5245 36127 5303 36133
rect 84802 36124 84808 36176
rect 84860 36164 84866 36176
rect 88050 36167 88108 36173
rect 88050 36164 88062 36167
rect 84860 36136 88062 36164
rect 84860 36124 84866 36136
rect 88050 36133 88062 36136
rect 88096 36133 88108 36167
rect 88050 36127 88108 36133
rect 4876 35930 7912 35952
rect 4876 35878 5882 35930
rect 5934 35878 5946 35930
rect 5998 35878 6010 35930
rect 6062 35878 6074 35930
rect 6126 35878 6138 35930
rect 6190 35878 7912 35930
rect 4876 35856 7912 35878
rect 85284 35930 88596 35952
rect 85284 35878 86474 35930
rect 86526 35878 86538 35930
rect 86590 35878 86602 35930
rect 86654 35878 86666 35930
rect 86718 35878 86730 35930
rect 86782 35878 88596 35930
rect 85284 35856 88596 35878
rect 4876 35386 7912 35408
rect 4876 35334 6618 35386
rect 6670 35334 6682 35386
rect 6734 35334 6746 35386
rect 6798 35334 6810 35386
rect 6862 35334 6874 35386
rect 6926 35334 7912 35386
rect 4876 35312 7912 35334
rect 85284 35386 88596 35408
rect 85284 35334 87210 35386
rect 87262 35334 87274 35386
rect 87326 35334 87338 35386
rect 87390 35334 87402 35386
rect 87454 35334 87466 35386
rect 87518 35334 88596 35386
rect 85284 35312 88596 35334
rect 5409 35147 5467 35153
rect 5409 35113 5421 35147
rect 5455 35144 5467 35147
rect 8534 35144 8540 35156
rect 5455 35116 8540 35144
rect 5455 35113 5467 35116
rect 5409 35107 5467 35113
rect 8534 35104 8540 35116
rect 8592 35104 8598 35156
rect 87933 35147 87991 35153
rect 87933 35113 87945 35147
rect 87979 35144 87991 35147
rect 88206 35144 88212 35156
rect 87979 35116 88212 35144
rect 87979 35113 87991 35116
rect 87933 35107 87991 35113
rect 88206 35104 88212 35116
rect 88264 35104 88270 35156
rect 4210 35036 4216 35088
rect 4268 35076 4274 35088
rect 5245 35079 5303 35085
rect 5245 35076 5257 35079
rect 4268 35048 5257 35076
rect 4268 35036 4274 35048
rect 5245 35045 5257 35048
rect 5291 35045 5303 35079
rect 5245 35039 5303 35045
rect 85814 34968 85820 35020
rect 85872 35008 85878 35020
rect 88050 35011 88108 35017
rect 88050 35008 88062 35011
rect 85872 34980 88062 35008
rect 85872 34968 85878 34980
rect 88050 34977 88062 34980
rect 88096 34977 88108 35011
rect 88050 34971 88108 34977
rect 4876 34842 7912 34864
rect 4876 34790 5882 34842
rect 5934 34790 5946 34842
rect 5998 34790 6010 34842
rect 6062 34790 6074 34842
rect 6126 34790 6138 34842
rect 6190 34790 7912 34842
rect 4876 34768 7912 34790
rect 85284 34842 88596 34864
rect 85284 34790 86474 34842
rect 86526 34790 86538 34842
rect 86590 34790 86602 34842
rect 86654 34790 86666 34842
rect 86718 34790 86730 34842
rect 86782 34790 88596 34842
rect 85284 34768 88596 34790
rect 4876 34298 7912 34320
rect 4876 34246 6618 34298
rect 6670 34246 6682 34298
rect 6734 34246 6746 34298
rect 6798 34246 6810 34298
rect 6862 34246 6874 34298
rect 6926 34246 7912 34298
rect 4876 34224 7912 34246
rect 85284 34298 88596 34320
rect 85284 34246 87210 34298
rect 87262 34246 87274 34298
rect 87326 34246 87338 34298
rect 87390 34246 87402 34298
rect 87454 34246 87466 34298
rect 87518 34246 88596 34298
rect 85284 34224 88596 34246
rect 5409 34059 5467 34065
rect 5409 34025 5421 34059
rect 5455 34056 5467 34059
rect 8534 34056 8540 34068
rect 5455 34028 8540 34056
rect 5455 34025 5467 34028
rect 5409 34019 5467 34025
rect 8534 34016 8540 34028
rect 8592 34016 8598 34068
rect 87933 34059 87991 34065
rect 87933 34025 87945 34059
rect 87979 34056 87991 34059
rect 88206 34056 88212 34068
rect 87979 34028 88212 34056
rect 87979 34025 87991 34028
rect 87933 34019 87991 34025
rect 88206 34016 88212 34028
rect 88264 34016 88270 34068
rect 85814 33880 85820 33932
rect 85872 33920 85878 33932
rect 88049 33923 88107 33929
rect 88049 33920 88061 33923
rect 85872 33892 88061 33920
rect 85872 33880 85878 33892
rect 88049 33889 88061 33892
rect 88095 33889 88107 33923
rect 88049 33883 88107 33889
rect 4210 33812 4216 33864
rect 4268 33852 4274 33864
rect 5245 33855 5303 33861
rect 5245 33852 5257 33855
rect 4268 33824 5257 33852
rect 4268 33812 4274 33824
rect 5245 33821 5257 33824
rect 5291 33821 5303 33855
rect 5245 33815 5303 33821
rect 4876 33754 7912 33776
rect 4876 33702 5882 33754
rect 5934 33702 5946 33754
rect 5998 33702 6010 33754
rect 6062 33702 6074 33754
rect 6126 33702 6138 33754
rect 6190 33702 7912 33754
rect 4876 33680 7912 33702
rect 85284 33754 88596 33776
rect 85284 33702 86474 33754
rect 86526 33702 86538 33754
rect 86590 33702 86602 33754
rect 86654 33702 86666 33754
rect 86718 33702 86730 33754
rect 86782 33702 88596 33754
rect 85284 33680 88596 33702
rect 4876 33210 7912 33232
rect 4876 33158 6618 33210
rect 6670 33158 6682 33210
rect 6734 33158 6746 33210
rect 6798 33158 6810 33210
rect 6862 33158 6874 33210
rect 6926 33158 7912 33210
rect 4876 33136 7912 33158
rect 85284 33210 88596 33232
rect 85284 33158 87210 33210
rect 87262 33158 87274 33210
rect 87326 33158 87338 33210
rect 87390 33158 87402 33210
rect 87454 33158 87466 33210
rect 87518 33158 88596 33210
rect 85284 33136 88596 33158
rect 4876 32666 7912 32688
rect 4876 32614 5882 32666
rect 5934 32614 5946 32666
rect 5998 32614 6010 32666
rect 6062 32614 6074 32666
rect 6126 32614 6138 32666
rect 6190 32614 7912 32666
rect 4876 32592 7912 32614
rect 85284 32666 88596 32688
rect 85284 32614 86474 32666
rect 86526 32614 86538 32666
rect 86590 32614 86602 32666
rect 86654 32614 86666 32666
rect 86718 32614 86730 32666
rect 86782 32614 88596 32666
rect 85284 32592 88596 32614
rect 85814 32452 85820 32504
rect 85872 32492 85878 32504
rect 88050 32495 88108 32501
rect 88050 32492 88062 32495
rect 85872 32464 88062 32492
rect 85872 32452 85878 32464
rect 88050 32461 88062 32464
rect 88096 32461 88108 32495
rect 88050 32455 88108 32461
rect 4210 32316 4216 32368
rect 4268 32356 4274 32368
rect 5245 32359 5303 32365
rect 5245 32356 5257 32359
rect 4268 32328 5257 32356
rect 4268 32316 4274 32328
rect 5245 32325 5257 32328
rect 5291 32325 5303 32359
rect 5245 32319 5303 32325
rect 5409 32359 5467 32365
rect 5409 32325 5421 32359
rect 5455 32356 5467 32359
rect 8534 32356 8540 32368
rect 5455 32328 8540 32356
rect 5455 32325 5467 32328
rect 5409 32319 5467 32325
rect 8534 32316 8540 32328
rect 8592 32316 8598 32368
rect 87749 32359 87807 32365
rect 87749 32325 87761 32359
rect 87795 32356 87807 32359
rect 88206 32356 88212 32368
rect 87795 32328 88212 32356
rect 87795 32325 87807 32328
rect 87749 32319 87807 32325
rect 88206 32316 88212 32328
rect 88264 32316 88270 32368
rect 4876 32122 7912 32144
rect 4876 32070 6618 32122
rect 6670 32070 6682 32122
rect 6734 32070 6746 32122
rect 6798 32070 6810 32122
rect 6862 32070 6874 32122
rect 6926 32070 7912 32122
rect 4876 32048 7912 32070
rect 85284 32122 88596 32144
rect 85284 32070 87210 32122
rect 87262 32070 87274 32122
rect 87326 32070 87338 32122
rect 87390 32070 87402 32122
rect 87454 32070 87466 32122
rect 87518 32070 88596 32122
rect 85284 32048 88596 32070
rect 5409 31883 5467 31889
rect 5409 31849 5421 31883
rect 5455 31880 5467 31883
rect 8534 31880 8540 31892
rect 5455 31852 8540 31880
rect 5455 31849 5467 31852
rect 5409 31843 5467 31849
rect 8534 31840 8540 31852
rect 8592 31840 8598 31892
rect 87933 31883 87991 31889
rect 87933 31849 87945 31883
rect 87979 31880 87991 31883
rect 88206 31880 88212 31892
rect 87979 31852 88212 31880
rect 87979 31849 87991 31852
rect 87933 31843 87991 31849
rect 88206 31840 88212 31852
rect 88264 31840 88270 31892
rect 85814 31704 85820 31756
rect 85872 31744 85878 31756
rect 88049 31747 88107 31753
rect 88049 31744 88061 31747
rect 85872 31716 88061 31744
rect 85872 31704 85878 31716
rect 88049 31713 88061 31716
rect 88095 31713 88107 31747
rect 88049 31707 88107 31713
rect 4118 31636 4124 31688
rect 4176 31676 4182 31688
rect 5245 31679 5303 31685
rect 5245 31676 5257 31679
rect 4176 31648 5257 31676
rect 4176 31636 4182 31648
rect 5245 31645 5257 31648
rect 5291 31645 5303 31679
rect 5245 31639 5303 31645
rect 4876 31578 7912 31600
rect 4876 31526 5882 31578
rect 5934 31526 5946 31578
rect 5998 31526 6010 31578
rect 6062 31526 6074 31578
rect 6126 31526 6138 31578
rect 6190 31526 7912 31578
rect 4876 31504 7912 31526
rect 85284 31578 88596 31600
rect 85284 31526 86474 31578
rect 86526 31526 86538 31578
rect 86590 31526 86602 31578
rect 86654 31526 86666 31578
rect 86718 31526 86730 31578
rect 86782 31526 88596 31578
rect 85284 31504 88596 31526
rect 4876 31034 7912 31056
rect 4876 30982 6618 31034
rect 6670 30982 6682 31034
rect 6734 30982 6746 31034
rect 6798 30982 6810 31034
rect 6862 30982 6874 31034
rect 6926 30982 7912 31034
rect 4876 30960 7912 30982
rect 85284 31034 88596 31056
rect 85284 30982 87210 31034
rect 87262 30982 87274 31034
rect 87326 30982 87338 31034
rect 87390 30982 87402 31034
rect 87454 30982 87466 31034
rect 87518 30982 88596 31034
rect 85284 30960 88596 30982
rect 5406 30752 5412 30804
rect 5464 30752 5470 30804
rect 87933 30795 87991 30801
rect 87933 30761 87945 30795
rect 87979 30792 87991 30795
rect 88209 30795 88267 30801
rect 88209 30792 88221 30795
rect 87979 30764 88221 30792
rect 87979 30761 87991 30764
rect 87933 30755 87991 30761
rect 88209 30761 88221 30764
rect 88255 30792 88267 30795
rect 88574 30792 88580 30804
rect 88255 30764 88580 30792
rect 88255 30761 88267 30764
rect 88209 30755 88267 30761
rect 88574 30752 88580 30764
rect 88632 30752 88638 30804
rect 4118 30616 4124 30668
rect 4176 30656 4182 30668
rect 5245 30659 5303 30665
rect 5245 30656 5257 30659
rect 4176 30628 5257 30656
rect 4176 30616 4182 30628
rect 5245 30625 5257 30628
rect 5291 30625 5303 30659
rect 5245 30619 5303 30625
rect 84802 30616 84808 30668
rect 84860 30656 84866 30668
rect 88050 30659 88108 30665
rect 88050 30656 88062 30659
rect 84860 30628 88062 30656
rect 84860 30616 84866 30628
rect 88050 30625 88062 30628
rect 88096 30625 88108 30659
rect 88050 30619 88108 30625
rect 4876 30490 7912 30512
rect 4876 30438 5882 30490
rect 5934 30438 5946 30490
rect 5998 30438 6010 30490
rect 6062 30438 6074 30490
rect 6126 30438 6138 30490
rect 6190 30438 7912 30490
rect 4876 30416 7912 30438
rect 85284 30490 88596 30512
rect 85284 30438 86474 30490
rect 86526 30438 86538 30490
rect 86590 30438 86602 30490
rect 86654 30438 86666 30490
rect 86718 30438 86730 30490
rect 86782 30438 88596 30490
rect 85284 30416 88596 30438
rect 4876 29946 7912 29968
rect 4876 29894 6618 29946
rect 6670 29894 6682 29946
rect 6734 29894 6746 29946
rect 6798 29894 6810 29946
rect 6862 29894 6874 29946
rect 6926 29894 7912 29946
rect 4876 29872 7912 29894
rect 85284 29946 88596 29968
rect 85284 29894 87210 29946
rect 87262 29894 87274 29946
rect 87326 29894 87338 29946
rect 87390 29894 87402 29946
rect 87454 29894 87466 29946
rect 87518 29894 88596 29946
rect 85284 29872 88596 29894
rect 4302 29664 4308 29716
rect 4360 29704 4366 29716
rect 5161 29707 5219 29713
rect 5161 29704 5173 29707
rect 4360 29676 5173 29704
rect 4360 29664 4366 29676
rect 5161 29673 5173 29676
rect 5207 29704 5219 29707
rect 5501 29707 5559 29713
rect 5501 29704 5513 29707
rect 5207 29676 5513 29704
rect 5207 29673 5219 29676
rect 5161 29667 5219 29673
rect 5501 29673 5513 29676
rect 5547 29673 5559 29707
rect 5501 29667 5559 29673
rect 85814 29664 85820 29716
rect 85872 29704 85878 29716
rect 87957 29707 88015 29713
rect 87957 29704 87969 29707
rect 85872 29676 87969 29704
rect 85872 29664 85878 29676
rect 87957 29673 87969 29676
rect 88003 29673 88015 29707
rect 87957 29667 88015 29673
rect 5363 29571 5421 29577
rect 5363 29537 5375 29571
rect 5409 29568 5421 29571
rect 8534 29568 8540 29580
rect 5409 29540 8540 29568
rect 5409 29537 5421 29540
rect 5363 29531 5421 29537
rect 8534 29528 8540 29540
rect 8592 29528 8598 29580
rect 88163 29503 88221 29509
rect 88163 29469 88175 29503
rect 88209 29500 88221 29503
rect 88390 29500 88396 29512
rect 88209 29472 88396 29500
rect 88209 29469 88221 29472
rect 88163 29463 88221 29469
rect 88390 29460 88396 29472
rect 88448 29460 88454 29512
rect 4876 29402 7912 29424
rect 4876 29350 5882 29402
rect 5934 29350 5946 29402
rect 5998 29350 6010 29402
rect 6062 29350 6074 29402
rect 6126 29350 6138 29402
rect 6190 29350 7912 29402
rect 4876 29328 7912 29350
rect 85284 29402 88596 29424
rect 85284 29350 86474 29402
rect 86526 29350 86538 29402
rect 86590 29350 86602 29402
rect 86654 29350 86666 29402
rect 86718 29350 86730 29402
rect 86782 29350 88596 29402
rect 85284 29328 88596 29350
rect 4876 28858 7912 28880
rect 4876 28806 6618 28858
rect 6670 28806 6682 28858
rect 6734 28806 6746 28858
rect 6798 28806 6810 28858
rect 6862 28806 6874 28858
rect 6926 28806 7912 28858
rect 4876 28784 7912 28806
rect 85284 28858 88596 28880
rect 85284 28806 87210 28858
rect 87262 28806 87274 28858
rect 87326 28806 87338 28858
rect 87390 28806 87402 28858
rect 87454 28806 87466 28858
rect 87518 28806 88596 28858
rect 85284 28784 88596 28806
rect 4302 28576 4308 28628
rect 4360 28616 4366 28628
rect 5161 28619 5219 28625
rect 5161 28616 5173 28619
rect 4360 28588 5173 28616
rect 4360 28576 4366 28588
rect 5161 28585 5173 28588
rect 5207 28616 5219 28619
rect 5501 28619 5559 28625
rect 5501 28616 5513 28619
rect 5207 28588 5513 28616
rect 5207 28585 5219 28588
rect 5161 28579 5219 28585
rect 5501 28585 5513 28588
rect 5547 28585 5559 28619
rect 5501 28579 5559 28585
rect 85814 28576 85820 28628
rect 85872 28616 85878 28628
rect 87957 28619 88015 28625
rect 87957 28616 87969 28619
rect 85872 28588 87969 28616
rect 85872 28576 85878 28588
rect 87957 28585 87969 28588
rect 88003 28585 88015 28619
rect 87957 28579 88015 28585
rect 5363 28483 5421 28489
rect 5363 28449 5375 28483
rect 5409 28480 5421 28483
rect 8534 28480 8540 28492
rect 5409 28452 8540 28480
rect 5409 28449 5421 28452
rect 5363 28443 5421 28449
rect 8534 28440 8540 28452
rect 8592 28440 8598 28492
rect 88206 28421 88212 28424
rect 88163 28415 88212 28421
rect 88163 28381 88175 28415
rect 88209 28381 88212 28415
rect 88163 28375 88212 28381
rect 88206 28372 88212 28375
rect 88264 28372 88270 28424
rect 4876 28314 7912 28336
rect 4876 28262 5882 28314
rect 5934 28262 5946 28314
rect 5998 28262 6010 28314
rect 6062 28262 6074 28314
rect 6126 28262 6138 28314
rect 6190 28262 7912 28314
rect 4876 28240 7912 28262
rect 85284 28314 88596 28336
rect 85284 28262 86474 28314
rect 86526 28262 86538 28314
rect 86590 28262 86602 28314
rect 86654 28262 86666 28314
rect 86718 28262 86730 28314
rect 86782 28262 88596 28314
rect 85284 28240 88596 28262
rect 4876 27770 7912 27792
rect 4876 27718 6618 27770
rect 6670 27718 6682 27770
rect 6734 27718 6746 27770
rect 6798 27718 6810 27770
rect 6862 27718 6874 27770
rect 6926 27718 7912 27770
rect 4876 27696 7912 27718
rect 85284 27770 88596 27792
rect 85284 27718 87210 27770
rect 87262 27718 87274 27770
rect 87326 27718 87338 27770
rect 87390 27718 87402 27770
rect 87454 27718 87466 27770
rect 87518 27718 88596 27770
rect 85284 27696 88596 27718
rect 4876 27226 7912 27248
rect 4876 27174 5882 27226
rect 5934 27174 5946 27226
rect 5998 27174 6010 27226
rect 6062 27174 6074 27226
rect 6126 27174 6138 27226
rect 6190 27174 7912 27226
rect 4876 27152 7912 27174
rect 85284 27226 88596 27248
rect 85284 27174 86474 27226
rect 86526 27174 86538 27226
rect 86590 27174 86602 27226
rect 86654 27174 86666 27226
rect 86718 27174 86730 27226
rect 86782 27174 88596 27226
rect 85284 27152 88596 27174
rect 5363 27055 5421 27061
rect 5363 27021 5375 27055
rect 5409 27052 5421 27055
rect 8534 27052 8540 27064
rect 5409 27024 8540 27052
rect 5409 27021 5421 27024
rect 5363 27015 5421 27021
rect 8534 27012 8540 27024
rect 8592 27012 8598 27064
rect 4302 26876 4308 26928
rect 4360 26916 4366 26928
rect 5161 26919 5219 26925
rect 5161 26916 5173 26919
rect 4360 26888 5173 26916
rect 4360 26876 4366 26888
rect 5161 26885 5173 26888
rect 5207 26916 5219 26919
rect 5501 26919 5559 26925
rect 5501 26916 5513 26919
rect 5207 26888 5513 26916
rect 5207 26885 5219 26888
rect 5161 26879 5219 26885
rect 5501 26885 5513 26888
rect 5547 26885 5559 26919
rect 5501 26879 5559 26885
rect 85814 26876 85820 26928
rect 85872 26916 85878 26928
rect 87957 26919 88015 26925
rect 87957 26916 87969 26919
rect 85872 26888 87969 26916
rect 85872 26876 85878 26888
rect 87957 26885 87969 26888
rect 88003 26885 88015 26919
rect 87957 26879 88015 26885
rect 88163 26783 88221 26789
rect 88163 26749 88175 26783
rect 88209 26780 88221 26783
rect 88390 26780 88396 26792
rect 88209 26752 88396 26780
rect 88209 26749 88221 26752
rect 88163 26743 88221 26749
rect 88390 26740 88396 26752
rect 88448 26740 88454 26792
rect 4876 26682 7912 26704
rect 4876 26630 6618 26682
rect 6670 26630 6682 26682
rect 6734 26630 6746 26682
rect 6798 26630 6810 26682
rect 6862 26630 6874 26682
rect 6926 26630 7912 26682
rect 4876 26608 7912 26630
rect 85284 26682 88596 26704
rect 85284 26630 87210 26682
rect 87262 26630 87274 26682
rect 87326 26630 87338 26682
rect 87390 26630 87402 26682
rect 87454 26630 87466 26682
rect 87518 26630 88596 26682
rect 85284 26608 88596 26630
rect 4302 26400 4308 26452
rect 4360 26440 4366 26452
rect 5161 26443 5219 26449
rect 5161 26440 5173 26443
rect 4360 26412 5173 26440
rect 4360 26400 4366 26412
rect 5161 26409 5173 26412
rect 5207 26440 5219 26443
rect 5501 26443 5559 26449
rect 5501 26440 5513 26443
rect 5207 26412 5513 26440
rect 5207 26409 5219 26412
rect 5161 26403 5219 26409
rect 5501 26409 5513 26412
rect 5547 26409 5559 26443
rect 5501 26403 5559 26409
rect 87562 26400 87568 26452
rect 87620 26440 87626 26452
rect 87957 26443 88015 26449
rect 87957 26440 87969 26443
rect 87620 26412 87969 26440
rect 87620 26400 87626 26412
rect 87957 26409 87969 26412
rect 88003 26409 88015 26443
rect 87957 26403 88015 26409
rect 5363 26307 5421 26313
rect 5363 26273 5375 26307
rect 5409 26304 5421 26307
rect 8534 26304 8540 26316
rect 5409 26276 8540 26304
rect 5409 26273 5421 26276
rect 5363 26267 5421 26273
rect 8534 26264 8540 26276
rect 8592 26264 8598 26316
rect 88206 26245 88212 26248
rect 88163 26239 88212 26245
rect 88163 26205 88175 26239
rect 88209 26205 88212 26239
rect 88163 26199 88212 26205
rect 88206 26196 88212 26199
rect 88264 26196 88270 26248
rect 4876 26138 7912 26160
rect 4876 26086 5882 26138
rect 5934 26086 5946 26138
rect 5998 26086 6010 26138
rect 6062 26086 6074 26138
rect 6126 26086 6138 26138
rect 6190 26086 7912 26138
rect 4876 26064 7912 26086
rect 85284 26138 88596 26160
rect 85284 26086 86474 26138
rect 86526 26086 86538 26138
rect 86590 26086 86602 26138
rect 86654 26086 86666 26138
rect 86718 26086 86730 26138
rect 86782 26086 88596 26138
rect 85284 26064 88596 26086
rect 4876 25594 7912 25616
rect 4876 25542 6618 25594
rect 6670 25542 6682 25594
rect 6734 25542 6746 25594
rect 6798 25542 6810 25594
rect 6862 25542 6874 25594
rect 6926 25542 7912 25594
rect 4876 25520 7912 25542
rect 85284 25594 88596 25616
rect 85284 25542 87210 25594
rect 87262 25542 87274 25594
rect 87326 25542 87338 25594
rect 87390 25542 87402 25594
rect 87454 25542 87466 25594
rect 87518 25542 88596 25594
rect 85284 25520 88596 25542
rect 4302 25312 4308 25364
rect 4360 25352 4366 25364
rect 5161 25355 5219 25361
rect 5161 25352 5173 25355
rect 4360 25324 5173 25352
rect 4360 25312 4366 25324
rect 5161 25321 5173 25324
rect 5207 25352 5219 25355
rect 5501 25355 5559 25361
rect 5501 25352 5513 25355
rect 5207 25324 5513 25352
rect 5207 25321 5219 25324
rect 5161 25315 5219 25321
rect 5501 25321 5513 25324
rect 5547 25321 5559 25355
rect 5501 25315 5559 25321
rect 84802 25312 84808 25364
rect 84860 25352 84866 25364
rect 87957 25355 88015 25361
rect 87957 25352 87969 25355
rect 84860 25324 87969 25352
rect 84860 25312 84866 25324
rect 87957 25321 87969 25324
rect 88003 25321 88015 25355
rect 87957 25315 88015 25321
rect 5406 25157 5412 25160
rect 5363 25151 5412 25157
rect 5363 25117 5375 25151
rect 5409 25117 5412 25151
rect 5363 25111 5412 25117
rect 5406 25108 5412 25111
rect 5464 25108 5470 25160
rect 88163 25151 88221 25157
rect 88163 25117 88175 25151
rect 88209 25148 88221 25151
rect 88574 25148 88580 25160
rect 88209 25120 88580 25148
rect 88209 25117 88221 25120
rect 88163 25111 88221 25117
rect 88574 25108 88580 25120
rect 88632 25108 88638 25160
rect 4876 25050 7912 25072
rect 4876 24998 5882 25050
rect 5934 24998 5946 25050
rect 5998 24998 6010 25050
rect 6062 24998 6074 25050
rect 6126 24998 6138 25050
rect 6190 24998 7912 25050
rect 4876 24976 7912 24998
rect 85284 25050 88596 25072
rect 85284 24998 86474 25050
rect 86526 24998 86538 25050
rect 86590 24998 86602 25050
rect 86654 24998 86666 25050
rect 86718 24998 86730 25050
rect 86782 24998 88596 25050
rect 85284 24976 88596 24998
rect 4876 24506 7912 24528
rect 4876 24454 6618 24506
rect 6670 24454 6682 24506
rect 6734 24454 6746 24506
rect 6798 24454 6810 24506
rect 6862 24454 6874 24506
rect 6926 24454 7912 24506
rect 4876 24432 7912 24454
rect 85284 24506 88596 24528
rect 85284 24454 87210 24506
rect 87262 24454 87274 24506
rect 87326 24454 87338 24506
rect 87390 24454 87402 24506
rect 87454 24454 87466 24506
rect 87518 24454 88596 24506
rect 85284 24432 88596 24454
rect 4302 24224 4308 24276
rect 4360 24264 4366 24276
rect 5161 24267 5219 24273
rect 5161 24264 5173 24267
rect 4360 24236 5173 24264
rect 4360 24224 4366 24236
rect 5161 24233 5173 24236
rect 5207 24264 5219 24267
rect 5501 24267 5559 24273
rect 5501 24264 5513 24267
rect 5207 24236 5513 24264
rect 5207 24233 5219 24236
rect 5161 24227 5219 24233
rect 5501 24233 5513 24236
rect 5547 24233 5559 24267
rect 5501 24227 5559 24233
rect 87562 24224 87568 24276
rect 87620 24264 87626 24276
rect 87957 24267 88015 24273
rect 87957 24264 87969 24267
rect 87620 24236 87969 24264
rect 87620 24224 87626 24236
rect 87957 24233 87969 24236
rect 88003 24233 88015 24267
rect 87957 24227 88015 24233
rect 5363 24131 5421 24137
rect 5363 24097 5375 24131
rect 5409 24128 5421 24131
rect 8534 24128 8540 24140
rect 5409 24100 8540 24128
rect 5409 24097 5421 24100
rect 5363 24091 5421 24097
rect 8534 24088 8540 24100
rect 8592 24088 8598 24140
rect 88163 24131 88221 24137
rect 88163 24097 88175 24131
rect 88209 24128 88221 24131
rect 88482 24128 88488 24140
rect 88209 24100 88488 24128
rect 88209 24097 88221 24100
rect 88163 24091 88221 24097
rect 88482 24088 88488 24100
rect 88540 24088 88546 24140
rect 4876 23962 7912 23984
rect 4876 23910 5882 23962
rect 5934 23910 5946 23962
rect 5998 23910 6010 23962
rect 6062 23910 6074 23962
rect 6126 23910 6138 23962
rect 6190 23910 7912 23962
rect 4876 23888 7912 23910
rect 85284 23962 88596 23984
rect 85284 23910 86474 23962
rect 86526 23910 86538 23962
rect 86590 23910 86602 23962
rect 86654 23910 86666 23962
rect 86718 23910 86730 23962
rect 86782 23910 88596 23962
rect 85284 23888 88596 23910
rect 4876 23418 7912 23440
rect 4876 23366 6618 23418
rect 6670 23366 6682 23418
rect 6734 23366 6746 23418
rect 6798 23366 6810 23418
rect 6862 23366 6874 23418
rect 6926 23366 7912 23418
rect 4876 23344 7912 23366
rect 85284 23418 88596 23440
rect 85284 23366 87210 23418
rect 87262 23366 87274 23418
rect 87326 23366 87338 23418
rect 87390 23366 87402 23418
rect 87454 23366 87466 23418
rect 87518 23366 88596 23418
rect 85284 23344 88596 23366
rect 4302 23136 4308 23188
rect 4360 23176 4366 23188
rect 5161 23179 5219 23185
rect 5161 23176 5173 23179
rect 4360 23148 5173 23176
rect 4360 23136 4366 23148
rect 5161 23145 5173 23148
rect 5207 23176 5219 23179
rect 5501 23179 5559 23185
rect 5501 23176 5513 23179
rect 5207 23148 5513 23176
rect 5207 23145 5219 23148
rect 5161 23139 5219 23145
rect 5501 23145 5513 23148
rect 5547 23145 5559 23179
rect 5501 23139 5559 23145
rect 85814 23136 85820 23188
rect 85872 23176 85878 23188
rect 87957 23179 88015 23185
rect 87957 23176 87969 23179
rect 85872 23148 87969 23176
rect 85872 23136 85878 23148
rect 87957 23145 87969 23148
rect 88003 23145 88015 23179
rect 87957 23139 88015 23145
rect 5363 23043 5421 23049
rect 5363 23009 5375 23043
rect 5409 23040 5421 23043
rect 8534 23040 8540 23052
rect 5409 23012 8540 23040
rect 5409 23009 5421 23012
rect 5363 23003 5421 23009
rect 8534 23000 8540 23012
rect 8592 23000 8598 23052
rect 88206 22981 88212 22984
rect 88163 22975 88212 22981
rect 88163 22941 88175 22975
rect 88209 22941 88212 22975
rect 88163 22935 88212 22941
rect 88206 22932 88212 22935
rect 88264 22932 88270 22984
rect 4876 22874 7912 22896
rect 4876 22822 5882 22874
rect 5934 22822 5946 22874
rect 5998 22822 6010 22874
rect 6062 22822 6074 22874
rect 6126 22822 6138 22874
rect 6190 22822 7912 22874
rect 4876 22800 7912 22822
rect 85284 22874 88596 22896
rect 85284 22822 86474 22874
rect 86526 22822 86538 22874
rect 86590 22822 86602 22874
rect 86654 22822 86666 22874
rect 86718 22822 86730 22874
rect 86782 22822 88596 22874
rect 85284 22800 88596 22822
rect 4876 22330 7912 22352
rect 4876 22278 6618 22330
rect 6670 22278 6682 22330
rect 6734 22278 6746 22330
rect 6798 22278 6810 22330
rect 6862 22278 6874 22330
rect 6926 22278 7912 22330
rect 4876 22256 7912 22278
rect 85284 22330 88596 22352
rect 85284 22278 87210 22330
rect 87262 22278 87274 22330
rect 87326 22278 87338 22330
rect 87390 22278 87402 22330
rect 87454 22278 87466 22330
rect 87518 22278 88596 22330
rect 85284 22256 88596 22278
rect 4876 21786 7912 21808
rect 4876 21734 5882 21786
rect 5934 21734 5946 21786
rect 5998 21734 6010 21786
rect 6062 21734 6074 21786
rect 6126 21734 6138 21786
rect 6190 21734 7912 21786
rect 4876 21712 7912 21734
rect 85284 21786 88596 21808
rect 85284 21734 86474 21786
rect 86526 21734 86538 21786
rect 86590 21734 86602 21786
rect 86654 21734 86666 21786
rect 86718 21734 86730 21786
rect 86782 21734 88596 21786
rect 85284 21712 88596 21734
rect 5363 21615 5421 21621
rect 5363 21581 5375 21615
rect 5409 21612 5421 21615
rect 8534 21612 8540 21624
rect 5409 21584 8540 21612
rect 5409 21581 5421 21584
rect 5363 21575 5421 21581
rect 8534 21572 8540 21584
rect 8592 21572 8598 21624
rect 4302 21436 4308 21488
rect 4360 21476 4366 21488
rect 5161 21479 5219 21485
rect 5161 21476 5173 21479
rect 4360 21448 5173 21476
rect 4360 21436 4366 21448
rect 5161 21445 5173 21448
rect 5207 21476 5219 21479
rect 5501 21479 5559 21485
rect 5501 21476 5513 21479
rect 5207 21448 5513 21476
rect 5207 21445 5219 21448
rect 5161 21439 5219 21445
rect 5501 21445 5513 21448
rect 5547 21445 5559 21479
rect 5501 21439 5559 21445
rect 85814 21436 85820 21488
rect 85872 21476 85878 21488
rect 87957 21479 88015 21485
rect 87957 21476 87969 21479
rect 85872 21448 87969 21476
rect 85872 21436 85878 21448
rect 87957 21445 87969 21448
rect 88003 21445 88015 21479
rect 87957 21439 88015 21445
rect 88163 21343 88221 21349
rect 88163 21309 88175 21343
rect 88209 21340 88221 21343
rect 88390 21340 88396 21352
rect 88209 21312 88396 21340
rect 88209 21309 88221 21312
rect 88163 21303 88221 21309
rect 88390 21300 88396 21312
rect 88448 21300 88454 21352
rect 4876 21242 7912 21264
rect 4876 21190 6618 21242
rect 6670 21190 6682 21242
rect 6734 21190 6746 21242
rect 6798 21190 6810 21242
rect 6862 21190 6874 21242
rect 6926 21190 7912 21242
rect 4876 21168 7912 21190
rect 85284 21242 88596 21264
rect 85284 21190 87210 21242
rect 87262 21190 87274 21242
rect 87326 21190 87338 21242
rect 87390 21190 87402 21242
rect 87454 21190 87466 21242
rect 87518 21190 88596 21242
rect 85284 21168 88596 21190
rect 5363 21071 5421 21077
rect 5363 21037 5375 21071
rect 5409 21068 5421 21071
rect 5682 21068 5688 21080
rect 5409 21040 5688 21068
rect 5409 21037 5421 21040
rect 5363 21031 5421 21037
rect 5682 21028 5688 21040
rect 5740 21028 5746 21080
rect 88163 21071 88221 21077
rect 88163 21037 88175 21071
rect 88209 21068 88221 21071
rect 88574 21068 88580 21080
rect 88209 21040 88580 21068
rect 88209 21037 88221 21040
rect 88163 21031 88221 21037
rect 88574 21028 88580 21040
rect 88632 21028 88638 21080
rect 4302 20960 4308 21012
rect 4360 21000 4366 21012
rect 5161 21003 5219 21009
rect 5161 21000 5173 21003
rect 4360 20972 5173 21000
rect 4360 20960 4366 20972
rect 5161 20969 5173 20972
rect 5207 21000 5219 21003
rect 5501 21003 5559 21009
rect 5501 21000 5513 21003
rect 5207 20972 5513 21000
rect 5207 20969 5219 20972
rect 5161 20963 5219 20969
rect 5501 20969 5513 20972
rect 5547 20969 5559 21003
rect 5501 20963 5559 20969
rect 84802 20960 84808 21012
rect 84860 21000 84866 21012
rect 87957 21003 88015 21009
rect 87957 21000 87969 21003
rect 84860 20972 87969 21000
rect 84860 20960 84866 20972
rect 87957 20969 87969 20972
rect 88003 20969 88015 21003
rect 87957 20963 88015 20969
rect 4876 20698 7912 20720
rect 4876 20646 5882 20698
rect 5934 20646 5946 20698
rect 5998 20646 6010 20698
rect 6062 20646 6074 20698
rect 6126 20646 6138 20698
rect 6190 20646 7912 20698
rect 4876 20624 7912 20646
rect 85284 20698 88596 20720
rect 85284 20646 86474 20698
rect 86526 20646 86538 20698
rect 86590 20646 86602 20698
rect 86654 20646 86666 20698
rect 86718 20646 86730 20698
rect 86782 20646 88596 20698
rect 85284 20624 88596 20646
rect 4876 20154 7912 20176
rect 4876 20102 6618 20154
rect 6670 20102 6682 20154
rect 6734 20102 6746 20154
rect 6798 20102 6810 20154
rect 6862 20102 6874 20154
rect 6926 20102 7912 20154
rect 4876 20080 7912 20102
rect 85284 20154 88596 20176
rect 85284 20102 87210 20154
rect 87262 20102 87274 20154
rect 87326 20102 87338 20154
rect 87390 20102 87402 20154
rect 87454 20102 87466 20154
rect 87518 20102 88596 20154
rect 85284 20080 88596 20102
rect 4302 19872 4308 19924
rect 4360 19912 4366 19924
rect 5161 19915 5219 19921
rect 5161 19912 5173 19915
rect 4360 19884 5173 19912
rect 4360 19872 4366 19884
rect 5161 19881 5173 19884
rect 5207 19912 5219 19915
rect 5501 19915 5559 19921
rect 5501 19912 5513 19915
rect 5207 19884 5513 19912
rect 5207 19881 5219 19884
rect 5161 19875 5219 19881
rect 5501 19881 5513 19884
rect 5547 19881 5559 19915
rect 5501 19875 5559 19881
rect 87562 19872 87568 19924
rect 87620 19912 87626 19924
rect 87957 19915 88015 19921
rect 87957 19912 87969 19915
rect 87620 19884 87969 19912
rect 87620 19872 87626 19884
rect 87957 19881 87969 19884
rect 88003 19881 88015 19915
rect 87957 19875 88015 19881
rect 5363 19779 5421 19785
rect 5363 19745 5375 19779
rect 5409 19776 5421 19779
rect 8534 19776 8540 19788
rect 5409 19748 8540 19776
rect 5409 19745 5421 19748
rect 5363 19739 5421 19745
rect 8534 19736 8540 19748
rect 8592 19736 8598 19788
rect 88163 19711 88221 19717
rect 88163 19677 88175 19711
rect 88209 19708 88221 19711
rect 88666 19708 88672 19720
rect 88209 19680 88672 19708
rect 88209 19677 88221 19680
rect 88163 19671 88221 19677
rect 88666 19668 88672 19680
rect 88724 19668 88730 19720
rect 4876 19610 7912 19632
rect 4876 19558 5882 19610
rect 5934 19558 5946 19610
rect 5998 19558 6010 19610
rect 6062 19558 6074 19610
rect 6126 19558 6138 19610
rect 6190 19558 7912 19610
rect 4876 19536 7912 19558
rect 85284 19610 88596 19632
rect 85284 19558 86474 19610
rect 86526 19558 86538 19610
rect 86590 19558 86602 19610
rect 86654 19558 86666 19610
rect 86718 19558 86730 19610
rect 86782 19558 88596 19610
rect 85284 19536 88596 19558
rect 4876 19066 7912 19088
rect 4876 19014 6618 19066
rect 6670 19014 6682 19066
rect 6734 19014 6746 19066
rect 6798 19014 6810 19066
rect 6862 19014 6874 19066
rect 6926 19014 7912 19066
rect 4876 18992 7912 19014
rect 85284 19066 88596 19088
rect 85284 19014 87210 19066
rect 87262 19014 87274 19066
rect 87326 19014 87338 19066
rect 87390 19014 87402 19066
rect 87454 19014 87466 19066
rect 87518 19014 88596 19066
rect 85284 18992 88596 19014
rect 4302 18784 4308 18836
rect 4360 18824 4366 18836
rect 5161 18827 5219 18833
rect 5161 18824 5173 18827
rect 4360 18796 5173 18824
rect 4360 18784 4366 18796
rect 5161 18793 5173 18796
rect 5207 18824 5219 18827
rect 5501 18827 5559 18833
rect 5501 18824 5513 18827
rect 5207 18796 5513 18824
rect 5207 18793 5219 18796
rect 5161 18787 5219 18793
rect 5501 18793 5513 18796
rect 5547 18793 5559 18827
rect 5501 18787 5559 18793
rect 87286 18784 87292 18836
rect 87344 18824 87350 18836
rect 87957 18827 88015 18833
rect 87957 18824 87969 18827
rect 87344 18796 87969 18824
rect 87344 18784 87350 18796
rect 87957 18793 87969 18796
rect 88003 18793 88015 18827
rect 87957 18787 88015 18793
rect 5363 18691 5421 18697
rect 5363 18657 5375 18691
rect 5409 18688 5421 18691
rect 8534 18688 8540 18700
rect 5409 18660 8540 18688
rect 5409 18657 5421 18660
rect 5363 18651 5421 18657
rect 8534 18648 8540 18660
rect 8592 18648 8598 18700
rect 88206 18697 88212 18700
rect 88163 18691 88212 18697
rect 88163 18657 88175 18691
rect 88209 18657 88212 18691
rect 88163 18651 88212 18657
rect 88206 18648 88212 18651
rect 88264 18648 88270 18700
rect 4876 18522 7912 18544
rect 4876 18470 5882 18522
rect 5934 18470 5946 18522
rect 5998 18470 6010 18522
rect 6062 18470 6074 18522
rect 6126 18470 6138 18522
rect 6190 18470 7912 18522
rect 4876 18448 7912 18470
rect 85284 18522 88596 18544
rect 85284 18470 86474 18522
rect 86526 18470 86538 18522
rect 86590 18470 86602 18522
rect 86654 18470 86666 18522
rect 86718 18470 86730 18522
rect 86782 18470 88596 18522
rect 85284 18448 88596 18470
rect 4876 17978 7912 18000
rect 4876 17926 6618 17978
rect 6670 17926 6682 17978
rect 6734 17926 6746 17978
rect 6798 17926 6810 17978
rect 6862 17926 6874 17978
rect 6926 17926 7912 17978
rect 4876 17904 7912 17926
rect 85284 17978 88596 18000
rect 85284 17926 87210 17978
rect 87262 17926 87274 17978
rect 87326 17926 87338 17978
rect 87390 17926 87402 17978
rect 87454 17926 87466 17978
rect 87518 17926 88596 17978
rect 85284 17904 88596 17926
rect 4302 17696 4308 17748
rect 4360 17736 4366 17748
rect 5161 17739 5219 17745
rect 5161 17736 5173 17739
rect 4360 17708 5173 17736
rect 4360 17696 4366 17708
rect 5161 17705 5173 17708
rect 5207 17736 5219 17739
rect 5501 17739 5559 17745
rect 5501 17736 5513 17739
rect 5207 17708 5513 17736
rect 5207 17705 5219 17708
rect 5161 17699 5219 17705
rect 5501 17705 5513 17708
rect 5547 17705 5559 17739
rect 5501 17699 5559 17705
rect 85814 17696 85820 17748
rect 85872 17736 85878 17748
rect 87957 17739 88015 17745
rect 87957 17736 87969 17739
rect 85872 17708 87969 17736
rect 85872 17696 85878 17708
rect 87957 17705 87969 17708
rect 88003 17705 88015 17739
rect 87957 17699 88015 17705
rect 5363 17603 5421 17609
rect 5363 17569 5375 17603
rect 5409 17600 5421 17603
rect 8534 17600 8540 17612
rect 5409 17572 8540 17600
rect 5409 17569 5421 17572
rect 5363 17563 5421 17569
rect 8534 17560 8540 17572
rect 8592 17560 8598 17612
rect 88206 17541 88212 17544
rect 88163 17535 88212 17541
rect 88163 17501 88175 17535
rect 88209 17501 88212 17535
rect 88163 17495 88212 17501
rect 88206 17492 88212 17495
rect 88264 17492 88270 17544
rect 4876 17434 7912 17456
rect 4876 17382 5882 17434
rect 5934 17382 5946 17434
rect 5998 17382 6010 17434
rect 6062 17382 6074 17434
rect 6126 17382 6138 17434
rect 6190 17382 7912 17434
rect 4876 17360 7912 17382
rect 85284 17434 88596 17456
rect 85284 17382 86474 17434
rect 86526 17382 86538 17434
rect 86590 17382 86602 17434
rect 86654 17382 86666 17434
rect 86718 17382 86730 17434
rect 86782 17382 88596 17434
rect 85284 17360 88596 17382
rect 4876 16890 7912 16912
rect 4876 16838 6618 16890
rect 6670 16838 6682 16890
rect 6734 16838 6746 16890
rect 6798 16838 6810 16890
rect 6862 16838 6874 16890
rect 6926 16838 7912 16890
rect 4876 16816 7912 16838
rect 85284 16890 88596 16912
rect 85284 16838 87210 16890
rect 87262 16838 87274 16890
rect 87326 16838 87338 16890
rect 87390 16838 87402 16890
rect 87454 16838 87466 16890
rect 87518 16838 88596 16890
rect 85284 16816 88596 16838
rect 4876 16346 7912 16368
rect 4876 16294 5882 16346
rect 5934 16294 5946 16346
rect 5998 16294 6010 16346
rect 6062 16294 6074 16346
rect 6126 16294 6138 16346
rect 6190 16294 7912 16346
rect 4876 16272 7912 16294
rect 85284 16346 88596 16368
rect 85284 16294 86474 16346
rect 86526 16294 86538 16346
rect 86590 16294 86602 16346
rect 86654 16294 86666 16346
rect 86718 16294 86730 16346
rect 86782 16294 88596 16346
rect 85284 16272 88596 16294
rect 5363 16175 5421 16181
rect 5363 16141 5375 16175
rect 5409 16172 5421 16175
rect 8534 16172 8540 16184
rect 5409 16144 8540 16172
rect 5409 16141 5421 16144
rect 5363 16135 5421 16141
rect 8534 16132 8540 16144
rect 8592 16132 8598 16184
rect 4302 15996 4308 16048
rect 4360 16036 4366 16048
rect 5161 16039 5219 16045
rect 5161 16036 5173 16039
rect 4360 16008 5173 16036
rect 4360 15996 4366 16008
rect 5161 16005 5173 16008
rect 5207 16036 5219 16039
rect 5501 16039 5559 16045
rect 5501 16036 5513 16039
rect 5207 16008 5513 16036
rect 5207 16005 5219 16008
rect 5161 15999 5219 16005
rect 5501 16005 5513 16008
rect 5547 16005 5559 16039
rect 5501 15999 5559 16005
rect 85814 15996 85820 16048
rect 85872 16036 85878 16048
rect 87957 16039 88015 16045
rect 87957 16036 87969 16039
rect 85872 16008 87969 16036
rect 85872 15996 85878 16008
rect 87957 16005 87969 16008
rect 88003 16005 88015 16039
rect 87957 15999 88015 16005
rect 88206 15909 88212 15912
rect 88163 15903 88212 15909
rect 88163 15869 88175 15903
rect 88209 15869 88212 15903
rect 88163 15863 88212 15869
rect 88206 15860 88212 15863
rect 88264 15860 88270 15912
rect 4876 15802 7912 15824
rect 4876 15750 6618 15802
rect 6670 15750 6682 15802
rect 6734 15750 6746 15802
rect 6798 15750 6810 15802
rect 6862 15750 6874 15802
rect 6926 15750 7912 15802
rect 4876 15728 7912 15750
rect 85284 15802 88596 15824
rect 85284 15750 87210 15802
rect 87262 15750 87274 15802
rect 87326 15750 87338 15802
rect 87390 15750 87402 15802
rect 87454 15750 87466 15802
rect 87518 15750 88596 15802
rect 85284 15728 88596 15750
rect 5363 15631 5421 15637
rect 5363 15597 5375 15631
rect 5409 15628 5421 15631
rect 5682 15628 5688 15640
rect 5409 15600 5688 15628
rect 5409 15597 5421 15600
rect 5363 15591 5421 15597
rect 5682 15588 5688 15600
rect 5740 15588 5746 15640
rect 88163 15631 88221 15637
rect 88163 15597 88175 15631
rect 88209 15628 88221 15631
rect 88574 15628 88580 15640
rect 88209 15600 88580 15628
rect 88209 15597 88221 15600
rect 88163 15591 88221 15597
rect 88574 15588 88580 15600
rect 88632 15588 88638 15640
rect 4302 15520 4308 15572
rect 4360 15560 4366 15572
rect 5161 15563 5219 15569
rect 5161 15560 5173 15563
rect 4360 15532 5173 15560
rect 4360 15520 4366 15532
rect 5161 15529 5173 15532
rect 5207 15560 5219 15563
rect 5501 15563 5559 15569
rect 5501 15560 5513 15563
rect 5207 15532 5513 15560
rect 5207 15529 5219 15532
rect 5161 15523 5219 15529
rect 5501 15529 5513 15532
rect 5547 15529 5559 15563
rect 5501 15523 5559 15529
rect 84802 15520 84808 15572
rect 84860 15560 84866 15572
rect 87957 15563 88015 15569
rect 87957 15560 87969 15563
rect 84860 15532 87969 15560
rect 84860 15520 84866 15532
rect 87957 15529 87969 15532
rect 88003 15529 88015 15563
rect 87957 15523 88015 15529
rect 4876 15258 7912 15280
rect 4876 15206 5882 15258
rect 5934 15206 5946 15258
rect 5998 15206 6010 15258
rect 6062 15206 6074 15258
rect 6126 15206 6138 15258
rect 6190 15206 7912 15258
rect 4876 15184 7912 15206
rect 85284 15258 88596 15280
rect 85284 15206 86474 15258
rect 86526 15206 86538 15258
rect 86590 15206 86602 15258
rect 86654 15206 86666 15258
rect 86718 15206 86730 15258
rect 86782 15206 88596 15258
rect 85284 15184 88596 15206
rect 85446 14976 85452 15028
rect 85504 15016 85510 15028
rect 85630 15016 85636 15028
rect 85504 14988 85636 15016
rect 85504 14976 85510 14988
rect 85630 14976 85636 14988
rect 85688 15016 85694 15028
rect 87473 15019 87531 15025
rect 87473 15016 87485 15019
rect 85688 14988 87485 15016
rect 85688 14976 85694 14988
rect 87473 14985 87485 14988
rect 87519 15016 87531 15019
rect 88209 15019 88267 15025
rect 88209 15016 88221 15019
rect 87519 14988 88221 15016
rect 87519 14985 87531 14988
rect 87473 14979 87531 14985
rect 88209 14985 88221 14988
rect 88255 14985 88267 15019
rect 88209 14979 88267 14985
rect 87796 14951 87854 14957
rect 87796 14917 87808 14951
rect 87842 14948 87854 14951
rect 87842 14920 88068 14948
rect 87842 14917 87854 14920
rect 87796 14911 87854 14917
rect 88040 14824 88068 14920
rect 88022 14772 88028 14824
rect 88080 14772 88086 14824
rect 4876 14714 7912 14736
rect 4876 14662 6618 14714
rect 6670 14662 6682 14714
rect 6734 14662 6746 14714
rect 6798 14662 6810 14714
rect 6862 14662 6874 14714
rect 6926 14662 7912 14714
rect 4876 14640 7912 14662
rect 85284 14714 88596 14736
rect 85284 14662 87210 14714
rect 87262 14662 87274 14714
rect 87326 14662 87338 14714
rect 87390 14662 87402 14714
rect 87454 14662 87466 14714
rect 87518 14662 88596 14714
rect 85284 14640 88596 14662
rect 83422 14228 83428 14280
rect 83480 14268 83486 14280
rect 85630 14268 85636 14280
rect 83480 14240 85636 14268
rect 83480 14228 83486 14240
rect 85630 14228 85636 14240
rect 85688 14228 85694 14280
rect 4876 14170 7912 14192
rect 4876 14118 5882 14170
rect 5934 14118 5946 14170
rect 5998 14118 6010 14170
rect 6062 14118 6074 14170
rect 6126 14118 6138 14170
rect 6190 14118 7912 14170
rect 4876 14096 7912 14118
rect 85284 14170 88596 14192
rect 85284 14118 86474 14170
rect 86526 14118 86538 14170
rect 86590 14118 86602 14170
rect 86654 14118 86666 14170
rect 86718 14118 86730 14170
rect 86782 14118 88596 14170
rect 85284 14096 88596 14118
rect 4876 13626 7912 13648
rect 4876 13574 6618 13626
rect 6670 13574 6682 13626
rect 6734 13574 6746 13626
rect 6798 13574 6810 13626
rect 6862 13574 6874 13626
rect 6926 13574 7912 13626
rect 4876 13552 7912 13574
rect 85284 13626 88596 13648
rect 85284 13574 87210 13626
rect 87262 13574 87274 13626
rect 87326 13574 87338 13626
rect 87390 13574 87402 13626
rect 87454 13574 87466 13626
rect 87518 13574 88596 13626
rect 85284 13552 88596 13574
rect 83606 13412 83612 13464
rect 83664 13452 83670 13464
rect 85538 13452 85544 13464
rect 83664 13424 85544 13452
rect 83664 13412 83670 13424
rect 85538 13412 85544 13424
rect 85596 13452 85602 13464
rect 85633 13455 85691 13461
rect 85633 13452 85645 13455
rect 85596 13424 85645 13452
rect 85596 13412 85602 13424
rect 85633 13421 85645 13424
rect 85679 13452 85691 13455
rect 87657 13455 87715 13461
rect 85679 13424 87194 13452
rect 85679 13421 85691 13424
rect 85633 13415 85691 13421
rect 87166 13316 87194 13424
rect 87657 13421 87669 13455
rect 87703 13452 87715 13455
rect 87703 13424 88252 13452
rect 87703 13421 87715 13424
rect 87657 13415 87715 13421
rect 88224 13396 88252 13424
rect 88206 13344 88212 13396
rect 88264 13384 88270 13396
rect 88264 13344 88272 13384
rect 88214 13338 88272 13344
rect 87930 13316 87936 13328
rect 87166 13288 87936 13316
rect 87930 13276 87936 13288
rect 87988 13276 87994 13328
rect 4876 13082 7912 13104
rect 4876 13030 5882 13082
rect 5934 13030 5946 13082
rect 5998 13030 6010 13082
rect 6062 13030 6074 13082
rect 6126 13030 6138 13082
rect 6190 13030 7912 13082
rect 4876 13008 7912 13030
rect 85284 13082 88596 13104
rect 85284 13030 86474 13082
rect 86526 13030 86538 13082
rect 86590 13030 86602 13082
rect 86654 13030 86666 13082
rect 86718 13030 86730 13082
rect 86782 13030 88596 13082
rect 85284 13008 88596 13030
rect 87930 12868 87936 12920
rect 87988 12908 87994 12920
rect 88209 12911 88267 12917
rect 88209 12908 88221 12911
rect 87988 12880 88221 12908
rect 87988 12868 87994 12880
rect 88209 12877 88221 12880
rect 88255 12877 88267 12911
rect 88209 12871 88267 12877
rect 87796 12775 87854 12781
rect 87796 12741 87808 12775
rect 87842 12772 87854 12775
rect 87842 12744 88068 12772
rect 87842 12741 87854 12744
rect 87796 12735 87854 12741
rect 87473 12707 87531 12713
rect 87473 12704 87485 12707
rect 87166 12676 87485 12704
rect 85354 12596 85360 12648
rect 85412 12636 85418 12648
rect 87166 12636 87194 12676
rect 87473 12673 87485 12676
rect 87519 12704 87531 12707
rect 87562 12704 87568 12716
rect 87519 12676 87568 12704
rect 87519 12673 87531 12676
rect 87473 12667 87531 12673
rect 87562 12664 87568 12676
rect 87620 12664 87626 12716
rect 88040 12713 88068 12744
rect 88025 12707 88083 12713
rect 88025 12673 88037 12707
rect 88071 12704 88083 12707
rect 88574 12704 88580 12716
rect 88071 12676 88580 12704
rect 88071 12673 88083 12676
rect 88025 12667 88083 12673
rect 88574 12664 88580 12676
rect 88632 12664 88638 12716
rect 85412 12608 87194 12636
rect 85412 12596 85418 12608
rect 4876 12538 7912 12560
rect 4876 12486 6618 12538
rect 6670 12486 6682 12538
rect 6734 12486 6746 12538
rect 6798 12486 6810 12538
rect 6862 12486 6874 12538
rect 6926 12486 7912 12538
rect 4876 12464 7912 12486
rect 85284 12538 88596 12560
rect 85284 12486 87210 12538
rect 87262 12486 87274 12538
rect 87326 12486 87338 12538
rect 87390 12486 87402 12538
rect 87454 12486 87466 12538
rect 87518 12486 88596 12538
rect 85284 12464 88596 12486
rect 83606 12324 83612 12376
rect 83664 12364 83670 12376
rect 85354 12364 85360 12376
rect 83664 12336 85360 12364
rect 83664 12324 83670 12336
rect 85354 12324 85360 12336
rect 85412 12364 85418 12376
rect 85633 12367 85691 12373
rect 85633 12364 85645 12367
rect 85412 12336 85645 12364
rect 85412 12324 85418 12336
rect 85633 12333 85645 12336
rect 85679 12333 85691 12367
rect 85633 12327 85691 12333
rect 87562 12324 87568 12376
rect 87620 12364 87626 12376
rect 88117 12367 88175 12373
rect 88117 12364 88129 12367
rect 87620 12336 88129 12364
rect 87620 12324 87626 12336
rect 88117 12333 88129 12336
rect 88163 12333 88175 12367
rect 88117 12327 88175 12333
rect 4876 11994 7912 12016
rect 4876 11942 5882 11994
rect 5934 11942 5946 11994
rect 5998 11942 6010 11994
rect 6062 11942 6074 11994
rect 6126 11942 6138 11994
rect 6190 11942 7912 11994
rect 4876 11920 7912 11942
rect 85284 11994 88596 12016
rect 85284 11942 86474 11994
rect 86526 11942 86538 11994
rect 86590 11942 86602 11994
rect 86654 11942 86666 11994
rect 86718 11942 86730 11994
rect 86782 11942 88596 11994
rect 85284 11920 88596 11942
rect 4876 11450 7912 11472
rect 4876 11398 6618 11450
rect 6670 11398 6682 11450
rect 6734 11398 6746 11450
rect 6798 11398 6810 11450
rect 6862 11398 6874 11450
rect 6926 11398 7912 11450
rect 4876 11376 7912 11398
rect 85284 11450 88596 11472
rect 85284 11398 87210 11450
rect 87262 11398 87274 11450
rect 87326 11398 87338 11450
rect 87390 11398 87402 11450
rect 87454 11398 87466 11450
rect 87518 11398 88596 11450
rect 85284 11376 88596 11398
rect 83238 11236 83244 11288
rect 83296 11276 83302 11288
rect 85633 11279 85691 11285
rect 85633 11276 85645 11279
rect 83296 11248 85645 11276
rect 83296 11236 83302 11248
rect 85633 11245 85645 11248
rect 85679 11245 85691 11279
rect 85633 11239 85691 11245
rect 4876 10906 7912 10928
rect 4876 10854 5882 10906
rect 5934 10854 5946 10906
rect 5998 10854 6010 10906
rect 6062 10854 6074 10906
rect 6126 10854 6138 10906
rect 6190 10854 7912 10906
rect 4876 10832 7912 10854
rect 85284 10906 88596 10928
rect 85284 10854 86474 10906
rect 86526 10854 86538 10906
rect 86590 10854 86602 10906
rect 86654 10854 86666 10906
rect 86718 10854 86730 10906
rect 86782 10854 88596 10906
rect 85284 10832 88596 10854
rect 87749 10599 87807 10605
rect 87749 10565 87761 10599
rect 87795 10596 87807 10599
rect 88206 10596 88212 10608
rect 87795 10568 88212 10596
rect 87795 10565 87807 10568
rect 87749 10559 87807 10565
rect 88206 10556 88212 10568
rect 88264 10556 88270 10608
rect 88049 10531 88107 10537
rect 88049 10528 88061 10531
rect 84728 10500 88061 10528
rect 84728 10392 84756 10500
rect 88049 10497 88061 10500
rect 88095 10497 88107 10531
rect 88049 10491 88107 10497
rect 4876 10362 7912 10384
rect 4876 10310 6618 10362
rect 6670 10310 6682 10362
rect 6734 10310 6746 10362
rect 6798 10310 6810 10362
rect 6862 10310 6874 10362
rect 6926 10310 7912 10362
rect 4876 10288 7912 10310
rect 82520 10364 84756 10392
rect 82520 10200 82548 10364
rect 85284 10362 88596 10384
rect 85284 10310 87210 10362
rect 87262 10310 87274 10362
rect 87326 10310 87338 10362
rect 87390 10310 87402 10362
rect 87454 10310 87466 10362
rect 87518 10310 88596 10362
rect 85284 10288 88596 10310
rect 45702 10148 45708 10200
rect 45760 10188 45766 10200
rect 46070 10188 46076 10200
rect 45760 10160 46076 10188
rect 45760 10148 45766 10160
rect 46070 10148 46076 10160
rect 46128 10148 46134 10200
rect 82502 10148 82508 10200
rect 82560 10148 82566 10200
rect 4876 9818 7912 9840
rect 4876 9766 5882 9818
rect 5934 9766 5946 9818
rect 5998 9766 6010 9818
rect 6062 9766 6074 9818
rect 6126 9766 6138 9818
rect 6190 9766 7912 9818
rect 4876 9744 7912 9766
rect 85284 9818 88596 9840
rect 85284 9766 86474 9818
rect 86526 9766 86538 9818
rect 86590 9766 86602 9818
rect 86654 9766 86666 9818
rect 86718 9766 86730 9818
rect 86782 9766 88596 9818
rect 85284 9744 88596 9766
rect 4876 9274 7912 9296
rect 4876 9222 6618 9274
rect 6670 9222 6682 9274
rect 6734 9222 6746 9274
rect 6798 9222 6810 9274
rect 6862 9222 6874 9274
rect 6926 9222 7912 9274
rect 4876 9200 7912 9222
rect 85284 9274 88596 9296
rect 85284 9222 87210 9274
rect 87262 9222 87274 9274
rect 87326 9222 87338 9274
rect 87390 9222 87402 9274
rect 87454 9222 87466 9274
rect 87518 9222 88596 9274
rect 85284 9200 88596 9222
rect 4876 8730 7912 8752
rect 4876 8678 5882 8730
rect 5934 8678 5946 8730
rect 5998 8678 6010 8730
rect 6062 8678 6074 8730
rect 6126 8678 6138 8730
rect 6190 8678 7912 8730
rect 4876 8656 7912 8678
rect 85284 8730 88596 8752
rect 85284 8678 86474 8730
rect 86526 8678 86538 8730
rect 86590 8678 86602 8730
rect 86654 8678 86666 8730
rect 86718 8678 86730 8730
rect 86782 8678 88596 8730
rect 85284 8656 88596 8678
rect 4876 8186 7912 8208
rect 4876 8134 6618 8186
rect 6670 8134 6682 8186
rect 6734 8134 6746 8186
rect 6798 8134 6810 8186
rect 6862 8134 6874 8186
rect 6926 8134 7912 8186
rect 4876 8112 7912 8134
rect 85284 8186 88596 8208
rect 85284 8134 87210 8186
rect 87262 8134 87274 8186
rect 87326 8134 87338 8186
rect 87390 8134 87402 8186
rect 87454 8134 87466 8186
rect 87518 8134 88596 8186
rect 85284 8112 88596 8134
rect 4876 7642 88596 7664
rect 4876 7590 5882 7642
rect 5934 7590 5946 7642
rect 5998 7590 6010 7642
rect 6062 7590 6074 7642
rect 6126 7590 6138 7642
rect 6190 7590 17722 7642
rect 17774 7590 17786 7642
rect 17838 7590 17850 7642
rect 17902 7590 17914 7642
rect 17966 7590 17978 7642
rect 18030 7590 36122 7642
rect 36174 7590 36186 7642
rect 36238 7590 36250 7642
rect 36302 7590 36314 7642
rect 36366 7590 36378 7642
rect 36430 7590 54522 7642
rect 54574 7590 54586 7642
rect 54638 7590 54650 7642
rect 54702 7590 54714 7642
rect 54766 7590 54778 7642
rect 54830 7590 72922 7642
rect 72974 7590 72986 7642
rect 73038 7590 73050 7642
rect 73102 7590 73114 7642
rect 73166 7590 73178 7642
rect 73230 7590 86474 7642
rect 86526 7590 86538 7642
rect 86590 7590 86602 7642
rect 86654 7590 86666 7642
rect 86718 7590 86730 7642
rect 86782 7590 88596 7642
rect 4876 7568 88596 7590
rect 45426 7428 45432 7480
rect 45484 7428 45490 7480
rect 45613 7471 45671 7477
rect 45613 7437 45625 7471
rect 45659 7468 45671 7471
rect 45702 7468 45708 7480
rect 45659 7440 45708 7468
rect 45659 7437 45671 7440
rect 45613 7431 45671 7437
rect 45702 7428 45708 7440
rect 45760 7428 45766 7480
rect 45797 7471 45855 7477
rect 45797 7437 45809 7471
rect 45843 7468 45855 7471
rect 45886 7468 45892 7480
rect 45843 7440 45892 7468
rect 45843 7437 45855 7440
rect 45797 7431 45855 7437
rect 45886 7428 45892 7440
rect 45944 7428 45950 7480
rect 45978 7428 45984 7480
rect 46036 7428 46042 7480
rect 45904 7332 45932 7428
rect 83514 7332 83520 7344
rect 45904 7304 83520 7332
rect 83514 7292 83520 7304
rect 83572 7292 83578 7344
rect 45978 7224 45984 7276
rect 46036 7264 46042 7276
rect 83330 7264 83336 7276
rect 46036 7236 83336 7264
rect 46036 7224 46042 7236
rect 83330 7224 83336 7236
rect 83388 7224 83394 7276
rect 45702 7156 45708 7208
rect 45760 7196 45766 7208
rect 83606 7196 83612 7208
rect 45760 7168 83612 7196
rect 45760 7156 45766 7168
rect 83606 7156 83612 7168
rect 83664 7156 83670 7208
rect 4876 7098 88596 7120
rect 4876 7046 6618 7098
rect 6670 7046 6682 7098
rect 6734 7046 6746 7098
rect 6798 7046 6810 7098
rect 6862 7046 6874 7098
rect 6926 7046 18382 7098
rect 18434 7046 18446 7098
rect 18498 7046 18510 7098
rect 18562 7046 18574 7098
rect 18626 7046 18638 7098
rect 18690 7046 36782 7098
rect 36834 7046 36846 7098
rect 36898 7046 36910 7098
rect 36962 7046 36974 7098
rect 37026 7046 37038 7098
rect 37090 7046 55182 7098
rect 55234 7046 55246 7098
rect 55298 7046 55310 7098
rect 55362 7046 55374 7098
rect 55426 7046 55438 7098
rect 55490 7046 73582 7098
rect 73634 7046 73646 7098
rect 73698 7046 73710 7098
rect 73762 7046 73774 7098
rect 73826 7046 73838 7098
rect 73890 7046 87210 7098
rect 87262 7046 87274 7098
rect 87326 7046 87338 7098
rect 87390 7046 87402 7098
rect 87454 7046 87466 7098
rect 87518 7046 88596 7098
rect 4876 7024 88596 7046
rect 4876 6554 88596 6576
rect 4876 6502 17722 6554
rect 17774 6502 17786 6554
rect 17838 6502 17850 6554
rect 17902 6502 17914 6554
rect 17966 6502 17978 6554
rect 18030 6502 36122 6554
rect 36174 6502 36186 6554
rect 36238 6502 36250 6554
rect 36302 6502 36314 6554
rect 36366 6502 36378 6554
rect 36430 6502 54522 6554
rect 54574 6502 54586 6554
rect 54638 6502 54650 6554
rect 54702 6502 54714 6554
rect 54766 6502 54778 6554
rect 54830 6502 72922 6554
rect 72974 6502 72986 6554
rect 73038 6502 73050 6554
rect 73102 6502 73114 6554
rect 73166 6502 73178 6554
rect 73230 6502 88596 6554
rect 4876 6480 88596 6502
rect 4876 6010 88596 6032
rect 4876 5958 18382 6010
rect 18434 5958 18446 6010
rect 18498 5958 18510 6010
rect 18562 5958 18574 6010
rect 18626 5958 18638 6010
rect 18690 5958 36782 6010
rect 36834 5958 36846 6010
rect 36898 5958 36910 6010
rect 36962 5958 36974 6010
rect 37026 5958 37038 6010
rect 37090 5958 55182 6010
rect 55234 5958 55246 6010
rect 55298 5958 55310 6010
rect 55362 5958 55374 6010
rect 55426 5958 55438 6010
rect 55490 5958 73582 6010
rect 73634 5958 73646 6010
rect 73698 5958 73710 6010
rect 73762 5958 73774 6010
rect 73826 5958 73838 6010
rect 73890 5958 88596 6010
rect 4876 5936 88596 5958
rect 4876 5466 88596 5488
rect 4876 5414 17722 5466
rect 17774 5414 17786 5466
rect 17838 5414 17850 5466
rect 17902 5414 17914 5466
rect 17966 5414 17978 5466
rect 18030 5414 36122 5466
rect 36174 5414 36186 5466
rect 36238 5414 36250 5466
rect 36302 5414 36314 5466
rect 36366 5414 36378 5466
rect 36430 5414 54522 5466
rect 54574 5414 54586 5466
rect 54638 5414 54650 5466
rect 54702 5414 54714 5466
rect 54766 5414 54778 5466
rect 54830 5414 72922 5466
rect 72974 5414 72986 5466
rect 73038 5414 73050 5466
rect 73102 5414 73114 5466
rect 73166 5414 73178 5466
rect 73230 5414 88596 5466
rect 4876 5392 88596 5414
rect 30430 5252 30436 5304
rect 30488 5292 30494 5304
rect 30733 5295 30791 5301
rect 30733 5292 30745 5295
rect 30488 5264 30745 5292
rect 30488 5252 30494 5264
rect 30733 5261 30745 5264
rect 30779 5261 30791 5295
rect 30733 5255 30791 5261
rect 31534 5252 31540 5304
rect 31592 5301 31598 5304
rect 31592 5295 31641 5301
rect 31592 5261 31595 5295
rect 31629 5261 31641 5295
rect 31592 5255 31641 5261
rect 31592 5252 31598 5255
rect 32638 5252 32644 5304
rect 32696 5301 32702 5304
rect 32696 5295 32724 5301
rect 32712 5261 32724 5295
rect 32696 5255 32724 5261
rect 32696 5252 32702 5255
rect 33742 5252 33748 5304
rect 33800 5292 33806 5304
rect 34846 5301 34852 5304
rect 33954 5295 34012 5301
rect 33954 5292 33966 5295
rect 33800 5264 33966 5292
rect 33800 5252 33806 5264
rect 33954 5261 33966 5264
rect 34000 5261 34012 5295
rect 33954 5255 34012 5261
rect 34803 5295 34852 5301
rect 34803 5261 34815 5295
rect 34849 5261 34852 5295
rect 34803 5255 34852 5261
rect 34846 5252 34852 5255
rect 34904 5252 34910 5304
rect 35950 5301 35956 5304
rect 35895 5295 35956 5301
rect 35895 5261 35907 5295
rect 35941 5261 35956 5295
rect 35895 5255 35956 5261
rect 35950 5252 35956 5255
rect 36008 5252 36014 5304
rect 37146 5252 37152 5304
rect 37204 5301 37210 5304
rect 37204 5295 37232 5301
rect 37220 5261 37232 5295
rect 37204 5255 37232 5261
rect 37204 5252 37210 5255
rect 38158 5252 38164 5304
rect 38216 5292 38222 5304
rect 38462 5295 38520 5301
rect 38462 5292 38474 5295
rect 38216 5264 38474 5292
rect 38216 5252 38222 5264
rect 38462 5261 38474 5264
rect 38508 5261 38520 5295
rect 38462 5255 38520 5261
rect 39262 5252 39268 5304
rect 39320 5301 39326 5304
rect 39320 5295 39369 5301
rect 39320 5261 39323 5295
rect 39357 5261 39369 5295
rect 39320 5255 39369 5261
rect 39320 5252 39326 5255
rect 40366 5252 40372 5304
rect 40424 5301 40430 5304
rect 40424 5295 40452 5301
rect 40440 5261 40452 5295
rect 40424 5255 40452 5261
rect 40424 5252 40430 5255
rect 41470 5252 41476 5304
rect 41528 5292 41534 5304
rect 42574 5301 42580 5304
rect 41681 5295 41739 5301
rect 41681 5292 41693 5295
rect 41528 5264 41693 5292
rect 41528 5252 41534 5264
rect 41681 5261 41693 5264
rect 41727 5261 41739 5295
rect 41681 5255 41739 5261
rect 42531 5295 42580 5301
rect 42531 5261 42543 5295
rect 42577 5261 42580 5295
rect 42531 5255 42580 5261
rect 42574 5252 42580 5255
rect 42632 5252 42638 5304
rect 43678 5301 43684 5304
rect 43623 5295 43684 5301
rect 43623 5261 43635 5295
rect 43669 5261 43684 5295
rect 43623 5255 43684 5261
rect 43678 5252 43684 5255
rect 43736 5252 43742 5304
rect 44782 5252 44788 5304
rect 44840 5292 44846 5304
rect 44901 5295 44959 5301
rect 44901 5292 44913 5295
rect 44840 5264 44913 5292
rect 44840 5252 44846 5264
rect 44901 5261 44913 5264
rect 44947 5261 44959 5295
rect 44901 5255 44959 5261
rect 68058 5252 68064 5304
rect 68116 5301 68122 5304
rect 68978 5301 68984 5304
rect 68116 5295 68143 5301
rect 68131 5261 68143 5295
rect 68116 5255 68143 5261
rect 68935 5295 68984 5301
rect 68935 5261 68947 5295
rect 68981 5261 68984 5295
rect 68935 5255 68984 5261
rect 68116 5252 68122 5255
rect 68978 5252 68984 5255
rect 69036 5252 69042 5304
rect 69990 5252 69996 5304
rect 70048 5301 70054 5304
rect 70048 5295 70076 5301
rect 70064 5261 70076 5295
rect 70048 5255 70076 5261
rect 70048 5252 70054 5255
rect 71278 5252 71284 5304
rect 71336 5301 71342 5304
rect 71336 5295 71364 5301
rect 71352 5261 71364 5295
rect 71336 5255 71364 5261
rect 71336 5252 71342 5255
rect 72566 5252 72572 5304
rect 72624 5301 72630 5304
rect 72624 5295 72652 5301
rect 72640 5261 72652 5295
rect 72624 5255 72652 5261
rect 72624 5252 72630 5255
rect 73394 5252 73400 5304
rect 73452 5301 73458 5304
rect 73452 5295 73501 5301
rect 73452 5261 73455 5295
rect 73489 5261 73501 5295
rect 73452 5255 73501 5261
rect 73452 5252 73458 5255
rect 74498 5252 74504 5304
rect 74556 5301 74562 5304
rect 74556 5295 74584 5301
rect 74572 5261 74584 5295
rect 74556 5255 74584 5261
rect 74556 5252 74562 5255
rect 75786 5252 75792 5304
rect 75844 5301 75850 5304
rect 76706 5301 76712 5304
rect 75844 5295 75872 5301
rect 75860 5261 75872 5295
rect 75844 5255 75872 5261
rect 76663 5295 76712 5301
rect 76663 5261 76675 5295
rect 76709 5261 76712 5295
rect 76663 5255 76712 5261
rect 75844 5252 75850 5255
rect 76706 5252 76712 5255
rect 76764 5252 76770 5304
rect 77718 5252 77724 5304
rect 77776 5301 77782 5304
rect 77776 5295 77804 5301
rect 77792 5261 77804 5295
rect 77776 5255 77804 5261
rect 77776 5252 77782 5255
rect 79006 5252 79012 5304
rect 79064 5301 79070 5304
rect 79064 5295 79091 5301
rect 79079 5261 79091 5295
rect 79064 5255 79091 5261
rect 79064 5252 79070 5255
rect 80110 5252 80116 5304
rect 80168 5292 80174 5304
rect 80321 5295 80379 5301
rect 80321 5292 80333 5295
rect 80168 5264 80333 5292
rect 80168 5252 80174 5264
rect 80321 5261 80333 5264
rect 80367 5261 80379 5295
rect 80321 5255 80379 5261
rect 81122 5252 81128 5304
rect 81180 5301 81186 5304
rect 81180 5295 81229 5301
rect 81180 5261 81183 5295
rect 81217 5261 81229 5295
rect 81180 5255 81229 5261
rect 81180 5252 81186 5255
rect 14974 5116 14980 5168
rect 15032 5156 15038 5168
rect 15277 5159 15335 5165
rect 15277 5156 15289 5159
rect 15032 5128 15289 5156
rect 15032 5116 15038 5128
rect 15277 5125 15289 5128
rect 15323 5125 15335 5159
rect 15277 5119 15335 5125
rect 16170 5116 16176 5168
rect 16228 5116 16234 5168
rect 17182 5116 17188 5168
rect 17240 5165 17246 5168
rect 17240 5159 17267 5165
rect 17255 5125 17267 5159
rect 17240 5119 17267 5125
rect 17240 5116 17246 5119
rect 18286 5116 18292 5168
rect 18344 5156 18350 5168
rect 18497 5159 18555 5165
rect 18497 5156 18509 5159
rect 18344 5128 18509 5156
rect 18344 5116 18350 5128
rect 18497 5125 18509 5128
rect 18543 5125 18555 5159
rect 18497 5119 18555 5125
rect 19390 5116 19396 5168
rect 19448 5116 19454 5168
rect 20494 5165 20500 5168
rect 20466 5159 20500 5165
rect 20466 5125 20478 5159
rect 20466 5119 20500 5125
rect 20494 5116 20500 5119
rect 20552 5116 20558 5168
rect 21598 5116 21604 5168
rect 21656 5156 21662 5168
rect 21717 5159 21775 5165
rect 21717 5156 21729 5159
rect 21656 5128 21729 5156
rect 21656 5116 21662 5128
rect 21717 5125 21729 5128
rect 21763 5125 21775 5159
rect 21717 5119 21775 5125
rect 22702 5116 22708 5168
rect 22760 5156 22766 5168
rect 23005 5159 23063 5165
rect 23005 5156 23017 5159
rect 22760 5128 23017 5156
rect 22760 5116 22766 5128
rect 23005 5125 23017 5128
rect 23051 5125 23063 5159
rect 23005 5119 23063 5125
rect 23898 5116 23904 5168
rect 23956 5116 23962 5168
rect 24910 5116 24916 5168
rect 24968 5165 24974 5168
rect 24968 5159 24995 5165
rect 24983 5125 24995 5159
rect 24968 5119 24995 5125
rect 24968 5116 24974 5119
rect 26014 5116 26020 5168
rect 26072 5156 26078 5168
rect 26225 5159 26283 5165
rect 26225 5156 26237 5159
rect 26072 5128 26237 5156
rect 26072 5116 26078 5128
rect 26225 5125 26237 5128
rect 26271 5125 26283 5159
rect 26225 5119 26283 5125
rect 27118 5116 27124 5168
rect 27176 5116 27182 5168
rect 28222 5165 28228 5168
rect 28194 5159 28228 5165
rect 28194 5125 28206 5159
rect 28194 5119 28228 5125
rect 28222 5116 28228 5119
rect 28280 5116 28286 5168
rect 29326 5116 29332 5168
rect 29384 5156 29390 5168
rect 29445 5159 29503 5165
rect 29445 5156 29457 5159
rect 29384 5128 29457 5156
rect 29384 5116 29390 5128
rect 29445 5125 29457 5128
rect 29491 5125 29503 5159
rect 29445 5119 29503 5125
rect 30706 5116 30712 5168
rect 30764 5156 30770 5168
rect 30893 5159 30951 5165
rect 30893 5156 30905 5159
rect 30764 5128 30905 5156
rect 30764 5116 30770 5128
rect 30893 5125 30905 5128
rect 30939 5156 30951 5159
rect 31077 5159 31135 5165
rect 31077 5156 31089 5159
rect 30939 5128 31089 5156
rect 30939 5125 30951 5128
rect 30893 5119 30951 5125
rect 31077 5125 31089 5128
rect 31123 5125 31135 5159
rect 31077 5119 31135 5125
rect 31350 5116 31356 5168
rect 31408 5165 31414 5168
rect 31408 5159 31439 5165
rect 31427 5156 31439 5159
rect 31721 5159 31779 5165
rect 31721 5156 31733 5159
rect 31427 5128 31733 5156
rect 31427 5125 31439 5128
rect 31408 5119 31439 5125
rect 31721 5125 31733 5128
rect 31767 5125 31779 5159
rect 31721 5119 31779 5125
rect 31408 5116 31414 5119
rect 32638 5116 32644 5168
rect 32696 5156 32702 5168
rect 32825 5159 32883 5165
rect 32825 5156 32837 5159
rect 32696 5128 32837 5156
rect 32696 5116 32702 5128
rect 32825 5125 32837 5128
rect 32871 5156 32883 5159
rect 33009 5159 33067 5165
rect 33009 5156 33021 5159
rect 32871 5128 33021 5156
rect 32871 5125 32883 5128
rect 32825 5119 32883 5125
rect 33009 5125 33021 5128
rect 33055 5125 33067 5159
rect 33009 5119 33067 5125
rect 33926 5116 33932 5168
rect 33984 5156 33990 5168
rect 34113 5159 34171 5165
rect 34113 5156 34125 5159
rect 33984 5128 34125 5156
rect 33984 5116 33990 5128
rect 34113 5125 34125 5128
rect 34159 5156 34171 5159
rect 34297 5159 34355 5165
rect 34297 5156 34309 5159
rect 34159 5128 34309 5156
rect 34159 5125 34171 5128
rect 34113 5119 34171 5125
rect 34297 5125 34309 5128
rect 34343 5125 34355 5159
rect 34297 5119 34355 5125
rect 34570 5116 34576 5168
rect 34628 5165 34634 5168
rect 34628 5159 34659 5165
rect 34647 5156 34659 5159
rect 34941 5159 34999 5165
rect 34941 5156 34953 5159
rect 34647 5128 34953 5156
rect 34647 5125 34659 5128
rect 34628 5119 34659 5125
rect 34941 5125 34953 5128
rect 34987 5125 34999 5159
rect 34941 5119 34999 5125
rect 34628 5116 34634 5119
rect 35858 5116 35864 5168
rect 35916 5156 35922 5168
rect 36045 5159 36103 5165
rect 36045 5156 36057 5159
rect 35916 5128 36057 5156
rect 35916 5116 35922 5128
rect 36045 5125 36057 5128
rect 36091 5156 36103 5159
rect 36229 5159 36287 5165
rect 36229 5156 36241 5159
rect 36091 5128 36241 5156
rect 36091 5125 36103 5128
rect 36045 5119 36103 5125
rect 36229 5125 36241 5128
rect 36275 5125 36287 5159
rect 36229 5119 36287 5125
rect 37146 5116 37152 5168
rect 37204 5156 37210 5168
rect 37333 5159 37391 5165
rect 37333 5156 37345 5159
rect 37204 5128 37345 5156
rect 37204 5116 37210 5128
rect 37333 5125 37345 5128
rect 37379 5156 37391 5159
rect 37517 5159 37575 5165
rect 37517 5156 37529 5159
rect 37379 5128 37529 5156
rect 37379 5125 37391 5128
rect 37333 5119 37391 5125
rect 37517 5125 37529 5128
rect 37563 5125 37575 5159
rect 37517 5119 37575 5125
rect 38434 5116 38440 5168
rect 38492 5156 38498 5168
rect 38621 5159 38679 5165
rect 38621 5156 38633 5159
rect 38492 5128 38633 5156
rect 38492 5116 38498 5128
rect 38621 5125 38633 5128
rect 38667 5156 38679 5159
rect 38805 5159 38863 5165
rect 38805 5156 38817 5159
rect 38667 5128 38817 5156
rect 38667 5125 38679 5128
rect 38621 5119 38679 5125
rect 38805 5125 38817 5128
rect 38851 5125 38863 5159
rect 38805 5119 38863 5125
rect 39078 5116 39084 5168
rect 39136 5165 39142 5168
rect 39136 5159 39167 5165
rect 39155 5156 39167 5159
rect 39449 5159 39507 5165
rect 39449 5156 39461 5159
rect 39155 5128 39461 5156
rect 39155 5125 39167 5128
rect 39136 5119 39167 5125
rect 39449 5125 39461 5128
rect 39495 5125 39507 5159
rect 39449 5119 39507 5125
rect 39136 5116 39142 5119
rect 40366 5116 40372 5168
rect 40424 5156 40430 5168
rect 40553 5159 40611 5165
rect 40553 5156 40565 5159
rect 40424 5128 40565 5156
rect 40424 5116 40430 5128
rect 40553 5125 40565 5128
rect 40599 5156 40611 5159
rect 40737 5159 40795 5165
rect 40737 5156 40749 5159
rect 40599 5128 40749 5156
rect 40599 5125 40611 5128
rect 40553 5119 40611 5125
rect 40737 5125 40749 5128
rect 40783 5125 40795 5159
rect 40737 5119 40795 5125
rect 41654 5116 41660 5168
rect 41712 5156 41718 5168
rect 41841 5159 41899 5165
rect 41841 5156 41853 5159
rect 41712 5128 41853 5156
rect 41712 5116 41718 5128
rect 41841 5125 41853 5128
rect 41887 5156 41899 5159
rect 42025 5159 42083 5165
rect 42025 5156 42037 5159
rect 41887 5128 42037 5156
rect 41887 5125 41899 5128
rect 41841 5119 41899 5125
rect 42025 5125 42037 5128
rect 42071 5125 42083 5159
rect 42025 5119 42083 5125
rect 42298 5116 42304 5168
rect 42356 5165 42362 5168
rect 42356 5159 42387 5165
rect 42375 5156 42387 5159
rect 42669 5159 42727 5165
rect 42669 5156 42681 5159
rect 42375 5128 42681 5156
rect 42375 5125 42387 5128
rect 42356 5119 42387 5125
rect 42669 5125 42681 5128
rect 42715 5125 42727 5159
rect 42669 5119 42727 5125
rect 42356 5116 42362 5119
rect 43586 5116 43592 5168
rect 43644 5156 43650 5168
rect 43773 5159 43831 5165
rect 43773 5156 43785 5159
rect 43644 5128 43785 5156
rect 43644 5116 43650 5128
rect 43773 5125 43785 5128
rect 43819 5156 43831 5159
rect 43957 5159 44015 5165
rect 43957 5156 43969 5159
rect 43819 5128 43969 5156
rect 43819 5125 43831 5128
rect 43773 5119 43831 5125
rect 43957 5125 43969 5128
rect 44003 5125 44015 5159
rect 43957 5119 44015 5125
rect 44874 5116 44880 5168
rect 44932 5156 44938 5168
rect 45061 5159 45119 5165
rect 45061 5156 45073 5159
rect 44932 5128 45073 5156
rect 44932 5116 44938 5128
rect 45061 5125 45073 5128
rect 45107 5156 45119 5159
rect 45245 5159 45303 5165
rect 45245 5156 45257 5159
rect 45107 5128 45257 5156
rect 45107 5125 45119 5128
rect 45061 5119 45119 5125
rect 45245 5125 45257 5128
rect 45291 5125 45303 5159
rect 45245 5119 45303 5125
rect 52602 5116 52608 5168
rect 52660 5165 52666 5168
rect 52660 5159 52687 5165
rect 52675 5125 52687 5159
rect 52660 5119 52687 5125
rect 52660 5116 52666 5119
rect 53522 5116 53528 5168
rect 53580 5116 53586 5168
rect 54442 5116 54448 5168
rect 54500 5156 54506 5168
rect 54561 5159 54619 5165
rect 54561 5156 54573 5159
rect 54500 5128 54573 5156
rect 54500 5116 54506 5128
rect 54561 5125 54573 5128
rect 54607 5125 54619 5159
rect 54561 5119 54619 5125
rect 55822 5116 55828 5168
rect 55880 5165 55886 5168
rect 55880 5159 55907 5165
rect 55895 5125 55907 5159
rect 55880 5119 55907 5125
rect 55880 5116 55886 5119
rect 57018 5116 57024 5168
rect 57076 5156 57082 5168
rect 57137 5159 57195 5165
rect 57137 5156 57149 5159
rect 57076 5128 57149 5156
rect 57076 5116 57082 5128
rect 57137 5125 57149 5128
rect 57183 5125 57195 5159
rect 57137 5119 57195 5125
rect 58030 5116 58036 5168
rect 58088 5116 58094 5168
rect 59042 5116 59048 5168
rect 59100 5165 59106 5168
rect 59100 5159 59127 5165
rect 59115 5125 59127 5159
rect 59100 5119 59127 5125
rect 59100 5116 59106 5119
rect 60330 5116 60336 5168
rect 60388 5165 60394 5168
rect 60388 5159 60415 5165
rect 60403 5125 60415 5159
rect 60388 5119 60415 5125
rect 60388 5116 60394 5119
rect 61250 5116 61256 5168
rect 61308 5116 61314 5168
rect 62354 5165 62360 5168
rect 62326 5159 62360 5165
rect 62326 5125 62338 5159
rect 62326 5119 62360 5125
rect 62354 5116 62360 5119
rect 62412 5116 62418 5168
rect 63550 5116 63556 5168
rect 63608 5165 63614 5168
rect 63608 5159 63635 5165
rect 63623 5125 63635 5159
rect 63608 5119 63635 5125
rect 63608 5116 63614 5119
rect 64746 5116 64752 5168
rect 64804 5156 64810 5168
rect 64865 5159 64923 5165
rect 64865 5156 64877 5159
rect 64804 5128 64877 5156
rect 64804 5116 64810 5128
rect 64865 5125 64877 5128
rect 64911 5125 64923 5159
rect 64865 5119 64923 5125
rect 65758 5116 65764 5168
rect 65816 5116 65822 5168
rect 66770 5116 66776 5168
rect 66828 5165 66834 5168
rect 66828 5159 66855 5165
rect 66843 5125 66855 5159
rect 66828 5119 66855 5125
rect 66828 5116 66834 5119
rect 68058 5116 68064 5168
rect 68116 5156 68122 5168
rect 68245 5159 68303 5165
rect 68245 5156 68257 5159
rect 68116 5128 68257 5156
rect 68116 5116 68122 5128
rect 68245 5125 68257 5128
rect 68291 5156 68303 5159
rect 68429 5159 68487 5165
rect 68429 5156 68441 5159
rect 68291 5128 68441 5156
rect 68291 5125 68303 5128
rect 68245 5119 68303 5125
rect 68429 5125 68441 5128
rect 68475 5125 68487 5159
rect 68429 5119 68487 5125
rect 68702 5116 68708 5168
rect 68760 5165 68766 5168
rect 68760 5159 68791 5165
rect 68779 5156 68791 5159
rect 69073 5159 69131 5165
rect 69073 5156 69085 5159
rect 68779 5128 69085 5156
rect 68779 5125 68791 5128
rect 68760 5119 68791 5125
rect 69073 5125 69085 5128
rect 69119 5125 69131 5159
rect 69073 5119 69131 5125
rect 68760 5116 68766 5119
rect 69990 5116 69996 5168
rect 70048 5156 70054 5168
rect 70177 5159 70235 5165
rect 70177 5156 70189 5159
rect 70048 5128 70189 5156
rect 70048 5116 70054 5128
rect 70177 5125 70189 5128
rect 70223 5156 70235 5159
rect 70361 5159 70419 5165
rect 70361 5156 70373 5159
rect 70223 5128 70373 5156
rect 70223 5125 70235 5128
rect 70177 5119 70235 5125
rect 70361 5125 70373 5128
rect 70407 5125 70419 5159
rect 70361 5119 70419 5125
rect 71278 5116 71284 5168
rect 71336 5156 71342 5168
rect 71465 5159 71523 5165
rect 71465 5156 71477 5159
rect 71336 5128 71477 5156
rect 71336 5116 71342 5128
rect 71465 5125 71477 5128
rect 71511 5156 71523 5159
rect 71649 5159 71707 5165
rect 71649 5156 71661 5159
rect 71511 5128 71661 5156
rect 71511 5125 71523 5128
rect 71465 5119 71523 5125
rect 71649 5125 71661 5128
rect 71695 5125 71707 5159
rect 71649 5119 71707 5125
rect 72566 5116 72572 5168
rect 72624 5156 72630 5168
rect 72753 5159 72811 5165
rect 72753 5156 72765 5159
rect 72624 5128 72765 5156
rect 72624 5116 72630 5128
rect 72753 5125 72765 5128
rect 72799 5156 72811 5159
rect 72937 5159 72995 5165
rect 72937 5156 72949 5159
rect 72799 5128 72949 5156
rect 72799 5125 72811 5128
rect 72753 5119 72811 5125
rect 72937 5125 72949 5128
rect 72983 5125 72995 5159
rect 72937 5119 72995 5125
rect 73210 5116 73216 5168
rect 73268 5165 73274 5168
rect 73268 5159 73299 5165
rect 73287 5156 73299 5159
rect 73581 5159 73639 5165
rect 73581 5156 73593 5159
rect 73287 5128 73593 5156
rect 73287 5125 73299 5128
rect 73268 5119 73299 5125
rect 73581 5125 73593 5128
rect 73627 5125 73639 5159
rect 73581 5119 73639 5125
rect 73268 5116 73274 5119
rect 74498 5116 74504 5168
rect 74556 5156 74562 5168
rect 74685 5159 74743 5165
rect 74685 5156 74697 5159
rect 74556 5128 74697 5156
rect 74556 5116 74562 5128
rect 74685 5125 74697 5128
rect 74731 5156 74743 5159
rect 74869 5159 74927 5165
rect 74869 5156 74881 5159
rect 74731 5128 74881 5156
rect 74731 5125 74743 5128
rect 74685 5119 74743 5125
rect 74869 5125 74881 5128
rect 74915 5125 74927 5159
rect 74869 5119 74927 5125
rect 75786 5116 75792 5168
rect 75844 5156 75850 5168
rect 75973 5159 76031 5165
rect 75973 5156 75985 5159
rect 75844 5128 75985 5156
rect 75844 5116 75850 5128
rect 75973 5125 75985 5128
rect 76019 5156 76031 5159
rect 76157 5159 76215 5165
rect 76157 5156 76169 5159
rect 76019 5128 76169 5156
rect 76019 5125 76031 5128
rect 75973 5119 76031 5125
rect 76157 5125 76169 5128
rect 76203 5125 76215 5159
rect 76157 5119 76215 5125
rect 76430 5116 76436 5168
rect 76488 5165 76494 5168
rect 76488 5159 76519 5165
rect 76507 5156 76519 5159
rect 76801 5159 76859 5165
rect 76801 5156 76813 5159
rect 76507 5128 76813 5156
rect 76507 5125 76519 5128
rect 76488 5119 76519 5125
rect 76801 5125 76813 5128
rect 76847 5125 76859 5159
rect 76801 5119 76859 5125
rect 76488 5116 76494 5119
rect 77718 5116 77724 5168
rect 77776 5156 77782 5168
rect 77905 5159 77963 5165
rect 77905 5156 77917 5159
rect 77776 5128 77917 5156
rect 77776 5116 77782 5128
rect 77905 5125 77917 5128
rect 77951 5156 77963 5159
rect 78089 5159 78147 5165
rect 78089 5156 78101 5159
rect 77951 5128 78101 5156
rect 77951 5125 77963 5128
rect 77905 5119 77963 5125
rect 78089 5125 78101 5128
rect 78135 5125 78147 5159
rect 78089 5119 78147 5125
rect 79006 5116 79012 5168
rect 79064 5156 79070 5168
rect 79193 5159 79251 5165
rect 79193 5156 79205 5159
rect 79064 5128 79205 5156
rect 79064 5116 79070 5128
rect 79193 5125 79205 5128
rect 79239 5156 79251 5159
rect 79377 5159 79435 5165
rect 79377 5156 79389 5159
rect 79239 5128 79389 5156
rect 79239 5125 79251 5128
rect 79193 5119 79251 5125
rect 79377 5125 79389 5128
rect 79423 5125 79435 5159
rect 79377 5119 79435 5125
rect 80294 5116 80300 5168
rect 80352 5156 80358 5168
rect 80481 5159 80539 5165
rect 80481 5156 80493 5159
rect 80352 5128 80493 5156
rect 80352 5116 80358 5128
rect 80481 5125 80493 5128
rect 80527 5156 80539 5159
rect 80665 5159 80723 5165
rect 80665 5156 80677 5159
rect 80527 5128 80677 5156
rect 80527 5125 80539 5128
rect 80481 5119 80539 5125
rect 80665 5125 80677 5128
rect 80711 5125 80723 5159
rect 80665 5119 80723 5125
rect 80938 5116 80944 5168
rect 80996 5165 81002 5168
rect 80996 5159 81027 5165
rect 81015 5156 81027 5159
rect 81309 5159 81367 5165
rect 81309 5156 81321 5159
rect 81015 5128 81321 5156
rect 81015 5125 81027 5128
rect 80996 5119 81027 5125
rect 81309 5125 81321 5128
rect 81355 5125 81367 5159
rect 81309 5119 81367 5125
rect 80996 5116 81002 5119
rect 15250 4980 15256 5032
rect 15308 5020 15314 5032
rect 15483 5023 15541 5029
rect 15483 5020 15495 5023
rect 15308 4992 15495 5020
rect 15308 4980 15314 4992
rect 15483 4989 15495 4992
rect 15529 4989 15541 5023
rect 15483 4983 15541 4989
rect 15894 4980 15900 5032
rect 15952 5020 15958 5032
rect 16009 5023 16067 5029
rect 16009 5020 16021 5023
rect 15952 4992 16021 5020
rect 15952 4980 15958 4992
rect 16009 4989 16021 4992
rect 16055 4989 16067 5023
rect 16009 4983 16067 4989
rect 17182 4980 17188 5032
rect 17240 5020 17246 5032
rect 18746 5029 18752 5032
rect 17415 5023 17473 5029
rect 17415 5020 17427 5023
rect 17240 4992 17427 5020
rect 17240 4980 17246 4992
rect 17415 4989 17427 4992
rect 17461 4989 17473 5023
rect 17415 4983 17473 4989
rect 18703 5023 18752 5029
rect 18703 4989 18715 5023
rect 18749 4989 18752 5023
rect 18703 4983 18752 4989
rect 18746 4980 18752 4983
rect 18804 4980 18810 5032
rect 19114 4980 19120 5032
rect 19172 5020 19178 5032
rect 19229 5023 19287 5029
rect 19229 5020 19241 5023
rect 19172 4992 19241 5020
rect 19172 4980 19178 4992
rect 19229 4989 19241 4992
rect 19275 4989 19287 5023
rect 19229 4983 19287 4989
rect 20402 4980 20408 5032
rect 20460 5020 20466 5032
rect 20635 5023 20693 5029
rect 20635 5020 20647 5023
rect 20460 4992 20647 5020
rect 20460 4980 20466 4992
rect 20635 4989 20647 4992
rect 20681 4989 20693 5023
rect 20635 4983 20693 4989
rect 21690 4980 21696 5032
rect 21748 5020 21754 5032
rect 21923 5023 21981 5029
rect 21923 5020 21935 5023
rect 21748 4992 21935 5020
rect 21748 4980 21754 4992
rect 21923 4989 21935 4992
rect 21969 4989 21981 5023
rect 21923 4983 21981 4989
rect 22978 4980 22984 5032
rect 23036 5020 23042 5032
rect 23211 5023 23269 5029
rect 23211 5020 23223 5023
rect 23036 4992 23223 5020
rect 23036 4980 23042 4992
rect 23211 4989 23223 4992
rect 23257 4989 23269 5023
rect 23211 4983 23269 4989
rect 23622 4980 23628 5032
rect 23680 5020 23686 5032
rect 23737 5023 23795 5029
rect 23737 5020 23749 5023
rect 23680 4992 23749 5020
rect 23680 4980 23686 4992
rect 23737 4989 23749 4992
rect 23783 4989 23795 5023
rect 23737 4983 23795 4989
rect 24910 4980 24916 5032
rect 24968 5020 24974 5032
rect 25143 5023 25201 5029
rect 25143 5020 25155 5023
rect 24968 4992 25155 5020
rect 24968 4980 24974 4992
rect 25143 4989 25155 4992
rect 25189 4989 25201 5023
rect 25143 4983 25201 4989
rect 26198 4980 26204 5032
rect 26256 5020 26262 5032
rect 26431 5023 26489 5029
rect 26431 5020 26443 5023
rect 26256 4992 26443 5020
rect 26256 4980 26262 4992
rect 26431 4989 26443 4992
rect 26477 4989 26489 5023
rect 26431 4983 26489 4989
rect 26842 4980 26848 5032
rect 26900 5020 26906 5032
rect 26957 5023 27015 5029
rect 26957 5020 26969 5023
rect 26900 4992 26969 5020
rect 26900 4980 26906 4992
rect 26957 4989 26969 4992
rect 27003 4989 27015 5023
rect 26957 4983 27015 4989
rect 28130 4980 28136 5032
rect 28188 5020 28194 5032
rect 28363 5023 28421 5029
rect 28363 5020 28375 5023
rect 28188 4992 28375 5020
rect 28188 4980 28194 4992
rect 28363 4989 28375 4992
rect 28409 4989 28421 5023
rect 28363 4983 28421 4989
rect 29418 4980 29424 5032
rect 29476 5020 29482 5032
rect 29651 5023 29709 5029
rect 29651 5020 29663 5023
rect 29476 4992 29663 5020
rect 29476 4980 29482 4992
rect 29651 4989 29663 4992
rect 29697 4989 29709 5023
rect 29651 4983 29709 4989
rect 52602 4980 52608 5032
rect 52660 5020 52666 5032
rect 52835 5023 52893 5029
rect 52835 5020 52847 5023
rect 52660 4992 52847 5020
rect 52660 4980 52666 4992
rect 52835 4989 52847 4992
rect 52881 4989 52893 5023
rect 52835 4983 52893 4989
rect 53246 4980 53252 5032
rect 53304 5020 53310 5032
rect 53361 5023 53419 5029
rect 53361 5020 53373 5023
rect 53304 4992 53373 5020
rect 53304 4980 53310 4992
rect 53361 4989 53373 4992
rect 53407 4989 53419 5023
rect 53361 4983 53419 4989
rect 54534 4980 54540 5032
rect 54592 5020 54598 5032
rect 54767 5023 54825 5029
rect 54767 5020 54779 5023
rect 54592 4992 54779 5020
rect 54592 4980 54598 4992
rect 54767 4989 54779 4992
rect 54813 4989 54825 5023
rect 54767 4983 54825 4989
rect 55822 4980 55828 5032
rect 55880 5020 55886 5032
rect 56055 5023 56113 5029
rect 56055 5020 56067 5023
rect 55880 4992 56067 5020
rect 55880 4980 55886 4992
rect 56055 4989 56067 4992
rect 56101 4989 56113 5023
rect 56055 4983 56113 4989
rect 57110 4980 57116 5032
rect 57168 5020 57174 5032
rect 57343 5023 57401 5029
rect 57343 5020 57355 5023
rect 57168 4992 57355 5020
rect 57168 4980 57174 4992
rect 57343 4989 57355 4992
rect 57389 4989 57401 5023
rect 57343 4983 57401 4989
rect 57754 4980 57760 5032
rect 57812 5020 57818 5032
rect 57869 5023 57927 5029
rect 57869 5020 57881 5023
rect 57812 4992 57881 5020
rect 57812 4980 57818 4992
rect 57869 4989 57881 4992
rect 57915 4989 57927 5023
rect 57869 4983 57927 4989
rect 59042 4980 59048 5032
rect 59100 5020 59106 5032
rect 59275 5023 59333 5029
rect 59275 5020 59287 5023
rect 59100 4992 59287 5020
rect 59100 4980 59106 4992
rect 59275 4989 59287 4992
rect 59321 4989 59333 5023
rect 59275 4983 59333 4989
rect 60330 4980 60336 5032
rect 60388 5020 60394 5032
rect 60563 5023 60621 5029
rect 60563 5020 60575 5023
rect 60388 4992 60575 5020
rect 60388 4980 60394 4992
rect 60563 4989 60575 4992
rect 60609 4989 60621 5023
rect 60563 4983 60621 4989
rect 60974 4980 60980 5032
rect 61032 5020 61038 5032
rect 61089 5023 61147 5029
rect 61089 5020 61101 5023
rect 61032 4992 61101 5020
rect 61032 4980 61038 4992
rect 61089 4989 61101 4992
rect 61135 4989 61147 5023
rect 61089 4983 61147 4989
rect 62262 4980 62268 5032
rect 62320 5020 62326 5032
rect 62495 5023 62553 5029
rect 62495 5020 62507 5023
rect 62320 4992 62507 5020
rect 62320 4980 62326 4992
rect 62495 4989 62507 4992
rect 62541 4989 62553 5023
rect 62495 4983 62553 4989
rect 63550 4980 63556 5032
rect 63608 5020 63614 5032
rect 63783 5023 63841 5029
rect 63783 5020 63795 5023
rect 63608 4992 63795 5020
rect 63608 4980 63614 4992
rect 63783 4989 63795 4992
rect 63829 4989 63841 5023
rect 63783 4983 63841 4989
rect 64838 4980 64844 5032
rect 64896 5020 64902 5032
rect 65071 5023 65129 5029
rect 65071 5020 65083 5023
rect 64896 4992 65083 5020
rect 64896 4980 64902 4992
rect 65071 4989 65083 4992
rect 65117 4989 65129 5023
rect 65071 4983 65129 4989
rect 65482 4980 65488 5032
rect 65540 5020 65546 5032
rect 65597 5023 65655 5029
rect 65597 5020 65609 5023
rect 65540 4992 65609 5020
rect 65540 4980 65546 4992
rect 65597 4989 65609 4992
rect 65643 4989 65655 5023
rect 65597 4983 65655 4989
rect 66770 4980 66776 5032
rect 66828 5020 66834 5032
rect 67003 5023 67061 5029
rect 67003 5020 67015 5023
rect 66828 4992 67015 5020
rect 66828 4980 66834 4992
rect 67003 4989 67015 4992
rect 67049 4989 67061 5023
rect 67003 4983 67061 4989
rect 4876 4922 88596 4944
rect 4876 4870 18382 4922
rect 18434 4870 18446 4922
rect 18498 4870 18510 4922
rect 18562 4870 18574 4922
rect 18626 4870 18638 4922
rect 18690 4870 36782 4922
rect 36834 4870 36846 4922
rect 36898 4870 36910 4922
rect 36962 4870 36974 4922
rect 37026 4870 37038 4922
rect 37090 4870 55182 4922
rect 55234 4870 55246 4922
rect 55298 4870 55310 4922
rect 55362 4870 55374 4922
rect 55426 4870 55438 4922
rect 55490 4870 73582 4922
rect 73634 4870 73646 4922
rect 73698 4870 73710 4922
rect 73762 4870 73774 4922
rect 73826 4870 73838 4922
rect 73890 4870 88596 4922
rect 4876 4848 88596 4870
<< via1 >>
rect 36508 87668 36560 87720
rect 37520 87668 37572 87720
rect 18382 87558 18434 87610
rect 18446 87558 18498 87610
rect 18510 87558 18562 87610
rect 18574 87558 18626 87610
rect 18638 87558 18690 87610
rect 36782 87558 36834 87610
rect 36846 87558 36898 87610
rect 36910 87558 36962 87610
rect 36974 87558 37026 87610
rect 37038 87558 37090 87610
rect 55182 87558 55234 87610
rect 55246 87558 55298 87610
rect 55310 87558 55362 87610
rect 55374 87558 55426 87610
rect 55438 87558 55490 87610
rect 73582 87558 73634 87610
rect 73646 87558 73698 87610
rect 73710 87558 73762 87610
rect 73774 87558 73826 87610
rect 73838 87558 73890 87610
rect 15256 87371 15308 87380
rect 15256 87337 15289 87371
rect 15289 87337 15308 87371
rect 34576 87396 34628 87448
rect 37152 87396 37204 87448
rect 39084 87396 39136 87448
rect 41016 87396 41068 87448
rect 42304 87396 42356 87448
rect 44236 87396 44288 87448
rect 15256 87328 15308 87337
rect 15900 87328 15952 87380
rect 17188 87328 17240 87380
rect 18752 87328 18804 87380
rect 19120 87371 19172 87380
rect 19120 87337 19157 87371
rect 19157 87337 19172 87371
rect 19120 87328 19172 87337
rect 20408 87328 20460 87380
rect 21696 87328 21748 87380
rect 22984 87328 23036 87380
rect 23628 87371 23680 87380
rect 23628 87337 23665 87371
rect 23665 87337 23680 87371
rect 23628 87328 23680 87337
rect 24916 87328 24968 87380
rect 26204 87328 26256 87380
rect 26848 87371 26900 87380
rect 26848 87337 26885 87371
rect 26885 87337 26900 87371
rect 26848 87328 26900 87337
rect 28136 87328 28188 87380
rect 29424 87328 29476 87380
rect 30620 87328 30672 87380
rect 31540 87328 31592 87380
rect 32644 87371 32696 87380
rect 32644 87337 32677 87371
rect 32677 87337 32696 87371
rect 32644 87328 32696 87337
rect 33748 87328 33800 87380
rect 34852 87371 34904 87380
rect 34852 87337 34861 87371
rect 34861 87337 34895 87371
rect 34895 87337 34904 87371
rect 34852 87328 34904 87337
rect 35956 87371 36008 87380
rect 35956 87337 35968 87371
rect 35968 87337 36008 87371
rect 35956 87328 36008 87337
rect 37428 87371 37480 87380
rect 37428 87337 37456 87371
rect 37456 87337 37480 87371
rect 37428 87328 37480 87337
rect 37612 87371 37664 87380
rect 37612 87337 37624 87371
rect 37624 87337 37664 87371
rect 37612 87328 37664 87337
rect 38164 87328 38216 87380
rect 38440 87371 38492 87380
rect 38440 87337 38473 87371
rect 38473 87337 38492 87371
rect 38440 87328 38492 87337
rect 39268 87328 39320 87380
rect 40372 87371 40424 87380
rect 40372 87337 40405 87371
rect 40405 87337 40424 87371
rect 40372 87328 40424 87337
rect 41476 87328 41528 87380
rect 41660 87328 41712 87380
rect 42580 87371 42632 87380
rect 42580 87337 42589 87371
rect 42589 87337 42623 87371
rect 42623 87337 42632 87371
rect 42580 87328 42632 87337
rect 42948 87328 43000 87380
rect 43684 87371 43736 87380
rect 43684 87337 43696 87371
rect 43696 87337 43736 87371
rect 43684 87328 43736 87337
rect 44788 87328 44840 87380
rect 44880 87328 44932 87380
rect 45524 87328 45576 87380
rect 46168 87328 46220 87380
rect 46812 87328 46864 87380
rect 47456 87328 47508 87380
rect 48100 87328 48152 87380
rect 48744 87328 48796 87380
rect 49388 87328 49440 87380
rect 50032 87328 50084 87380
rect 52608 87371 52660 87380
rect 52608 87337 52641 87371
rect 52641 87337 52660 87371
rect 68708 87396 68760 87448
rect 76436 87396 76488 87448
rect 52608 87328 52660 87337
rect 53252 87328 53304 87380
rect 54540 87328 54592 87380
rect 55828 87328 55880 87380
rect 57116 87328 57168 87380
rect 57760 87371 57812 87380
rect 57760 87337 57797 87371
rect 57797 87337 57812 87371
rect 57760 87328 57812 87337
rect 59048 87328 59100 87380
rect 60336 87328 60388 87380
rect 60980 87371 61032 87380
rect 60980 87337 61017 87371
rect 61017 87337 61032 87371
rect 60980 87328 61032 87337
rect 62268 87328 62320 87380
rect 63556 87328 63608 87380
rect 64844 87328 64896 87380
rect 65488 87371 65540 87380
rect 65488 87337 65525 87371
rect 65525 87337 65540 87371
rect 65488 87328 65540 87337
rect 66776 87328 66828 87380
rect 67880 87328 67932 87380
rect 68984 87371 69036 87380
rect 68984 87337 68993 87371
rect 68993 87337 69027 87371
rect 69027 87337 69036 87371
rect 68984 87328 69036 87337
rect 69996 87371 70048 87380
rect 69996 87337 70029 87371
rect 70029 87337 70048 87371
rect 69996 87328 70048 87337
rect 71192 87328 71244 87380
rect 72296 87328 72348 87380
rect 73400 87328 73452 87380
rect 74504 87371 74556 87380
rect 74504 87337 74537 87371
rect 74537 87337 74556 87371
rect 74504 87328 74556 87337
rect 75608 87328 75660 87380
rect 76712 87371 76764 87380
rect 76712 87337 76721 87371
rect 76721 87337 76755 87371
rect 76755 87337 76764 87371
rect 76712 87328 76764 87337
rect 77724 87371 77776 87380
rect 77724 87337 77757 87371
rect 77757 87337 77776 87371
rect 77724 87328 77776 87337
rect 78920 87328 78972 87380
rect 80392 87371 80444 87380
rect 80392 87337 80404 87371
rect 80404 87337 80444 87371
rect 80392 87328 80444 87337
rect 81128 87328 81180 87380
rect 82232 87371 82284 87380
rect 82232 87337 82265 87371
rect 82265 87337 82284 87371
rect 82232 87328 82284 87337
rect 36600 87303 36652 87312
rect 36600 87269 36609 87303
rect 36609 87269 36643 87303
rect 36643 87269 36652 87303
rect 36600 87260 36652 87269
rect 39084 87260 39136 87312
rect 15532 87235 15584 87244
rect 15532 87201 15541 87235
rect 15541 87201 15575 87235
rect 15575 87201 15584 87235
rect 15532 87192 15584 87201
rect 16084 87192 16136 87244
rect 17188 87235 17240 87244
rect 17188 87201 17222 87235
rect 17222 87201 17240 87235
rect 17188 87192 17240 87201
rect 18292 87192 18344 87244
rect 19396 87192 19448 87244
rect 20408 87235 20460 87244
rect 20408 87201 20442 87235
rect 20442 87201 20460 87235
rect 20408 87192 20460 87201
rect 21604 87192 21656 87244
rect 22708 87192 22760 87244
rect 23812 87192 23864 87244
rect 24916 87235 24968 87244
rect 24916 87201 24950 87235
rect 24950 87201 24968 87235
rect 24916 87192 24968 87201
rect 26020 87192 26072 87244
rect 27124 87192 27176 87244
rect 28136 87235 28188 87244
rect 28136 87201 28169 87235
rect 28169 87201 28188 87235
rect 28136 87192 28188 87201
rect 29332 87192 29384 87244
rect 30712 87192 30764 87244
rect 31356 87192 31408 87244
rect 32736 87192 32788 87244
rect 33932 87192 33984 87244
rect 35864 87192 35916 87244
rect 38348 87192 38400 87244
rect 40464 87192 40516 87244
rect 43592 87192 43644 87244
rect 52884 87235 52936 87244
rect 52884 87201 52893 87235
rect 52893 87201 52927 87235
rect 52927 87201 52936 87235
rect 52884 87192 52936 87201
rect 53528 87235 53580 87244
rect 53528 87201 53562 87235
rect 53562 87201 53580 87235
rect 53528 87192 53580 87201
rect 54448 87192 54500 87244
rect 55736 87192 55788 87244
rect 56840 87192 56892 87244
rect 57944 87192 57996 87244
rect 59048 87235 59100 87244
rect 59048 87201 59082 87235
rect 59082 87201 59100 87235
rect 59048 87192 59100 87201
rect 60152 87192 60204 87244
rect 61164 87192 61216 87244
rect 62452 87192 62504 87244
rect 63464 87192 63516 87244
rect 64568 87192 64620 87244
rect 65672 87192 65724 87244
rect 66776 87235 66828 87244
rect 66776 87201 66810 87235
rect 66810 87201 66828 87235
rect 66776 87192 66828 87201
rect 68064 87192 68116 87244
rect 70088 87192 70140 87244
rect 71284 87192 71336 87244
rect 72572 87192 72624 87244
rect 73216 87192 73268 87244
rect 74596 87192 74648 87244
rect 75792 87192 75844 87244
rect 77816 87192 77868 87244
rect 79012 87192 79064 87244
rect 80300 87192 80352 87244
rect 80944 87192 80996 87244
rect 82324 87192 82376 87244
rect 17722 87014 17774 87066
rect 17786 87014 17838 87066
rect 17850 87014 17902 87066
rect 17914 87014 17966 87066
rect 17978 87014 18030 87066
rect 36122 87014 36174 87066
rect 36186 87014 36238 87066
rect 36250 87014 36302 87066
rect 36314 87014 36366 87066
rect 36378 87014 36430 87066
rect 54522 87014 54574 87066
rect 54586 87014 54638 87066
rect 54650 87014 54702 87066
rect 54714 87014 54766 87066
rect 54778 87014 54830 87066
rect 72922 87014 72974 87066
rect 72986 87014 73038 87066
rect 73050 87014 73102 87066
rect 73114 87014 73166 87066
rect 73178 87014 73230 87066
rect 37520 86852 37572 86904
rect 37796 86852 37848 86904
rect 38440 86852 38492 86904
rect 36600 86580 36652 86632
rect 46996 86580 47048 86632
rect 50308 86580 50360 86632
rect 18382 86470 18434 86522
rect 18446 86470 18498 86522
rect 18510 86470 18562 86522
rect 18574 86470 18626 86522
rect 18638 86470 18690 86522
rect 36782 86470 36834 86522
rect 36846 86470 36898 86522
rect 36910 86470 36962 86522
rect 36974 86470 37026 86522
rect 37038 86470 37090 86522
rect 55182 86470 55234 86522
rect 55246 86470 55298 86522
rect 55310 86470 55362 86522
rect 55374 86470 55426 86522
rect 55438 86470 55490 86522
rect 73582 86470 73634 86522
rect 73646 86470 73698 86522
rect 73710 86470 73762 86522
rect 73774 86470 73826 86522
rect 73838 86470 73890 86522
rect 17722 85926 17774 85978
rect 17786 85926 17838 85978
rect 17850 85926 17902 85978
rect 17914 85926 17966 85978
rect 17978 85926 18030 85978
rect 36122 85926 36174 85978
rect 36186 85926 36238 85978
rect 36250 85926 36302 85978
rect 36314 85926 36366 85978
rect 36378 85926 36430 85978
rect 54522 85926 54574 85978
rect 54586 85926 54638 85978
rect 54650 85926 54702 85978
rect 54714 85926 54766 85978
rect 54778 85926 54830 85978
rect 72922 85926 72974 85978
rect 72986 85926 73038 85978
rect 73050 85926 73102 85978
rect 73114 85926 73166 85978
rect 73178 85926 73230 85978
rect 18382 85382 18434 85434
rect 18446 85382 18498 85434
rect 18510 85382 18562 85434
rect 18574 85382 18626 85434
rect 18638 85382 18690 85434
rect 36782 85382 36834 85434
rect 36846 85382 36898 85434
rect 36910 85382 36962 85434
rect 36974 85382 37026 85434
rect 37038 85382 37090 85434
rect 55182 85382 55234 85434
rect 55246 85382 55298 85434
rect 55310 85382 55362 85434
rect 55374 85382 55426 85434
rect 55438 85382 55490 85434
rect 73582 85382 73634 85434
rect 73646 85382 73698 85434
rect 73710 85382 73762 85434
rect 73774 85382 73826 85434
rect 73838 85382 73890 85434
rect 5882 84838 5934 84890
rect 5946 84838 5998 84890
rect 6010 84838 6062 84890
rect 6074 84838 6126 84890
rect 6138 84838 6190 84890
rect 17722 84838 17774 84890
rect 17786 84838 17838 84890
rect 17850 84838 17902 84890
rect 17914 84838 17966 84890
rect 17978 84838 18030 84890
rect 36122 84838 36174 84890
rect 36186 84838 36238 84890
rect 36250 84838 36302 84890
rect 36314 84838 36366 84890
rect 36378 84838 36430 84890
rect 54522 84838 54574 84890
rect 54586 84838 54638 84890
rect 54650 84838 54702 84890
rect 54714 84838 54766 84890
rect 54778 84838 54830 84890
rect 72922 84838 72974 84890
rect 72986 84838 73038 84890
rect 73050 84838 73102 84890
rect 73114 84838 73166 84890
rect 73178 84838 73230 84890
rect 86474 84838 86526 84890
rect 86538 84838 86590 84890
rect 86602 84838 86654 84890
rect 86666 84838 86718 84890
rect 86730 84838 86782 84890
rect 46168 84676 46220 84728
rect 12772 84608 12824 84660
rect 36600 84608 36652 84660
rect 11668 84540 11720 84592
rect 39084 84608 39136 84660
rect 49112 84608 49164 84660
rect 50308 84719 50360 84728
rect 50308 84685 50317 84719
rect 50317 84685 50351 84719
rect 50351 84685 50360 84719
rect 50308 84676 50360 84685
rect 51320 84608 51372 84660
rect 46076 84540 46128 84592
rect 7528 84472 7580 84524
rect 10564 84404 10616 84456
rect 13876 84404 13928 84456
rect 39728 84472 39780 84524
rect 45892 84404 45944 84456
rect 45984 84447 46036 84456
rect 45984 84413 45993 84447
rect 45993 84413 46027 84447
rect 46027 84413 46036 84447
rect 45984 84404 46036 84413
rect 48008 84404 48060 84456
rect 49112 84404 49164 84456
rect 51320 84404 51372 84456
rect 6618 84294 6670 84346
rect 6682 84294 6734 84346
rect 6746 84294 6798 84346
rect 6810 84294 6862 84346
rect 6874 84294 6926 84346
rect 18382 84294 18434 84346
rect 18446 84294 18498 84346
rect 18510 84294 18562 84346
rect 18574 84294 18626 84346
rect 18638 84294 18690 84346
rect 36782 84294 36834 84346
rect 36846 84294 36898 84346
rect 36910 84294 36962 84346
rect 36974 84294 37026 84346
rect 37038 84294 37090 84346
rect 55182 84294 55234 84346
rect 55246 84294 55298 84346
rect 55310 84294 55362 84346
rect 55374 84294 55426 84346
rect 55438 84294 55490 84346
rect 73582 84294 73634 84346
rect 73646 84294 73698 84346
rect 73710 84294 73762 84346
rect 73774 84294 73826 84346
rect 73838 84294 73890 84346
rect 87210 84294 87262 84346
rect 87274 84294 87326 84346
rect 87338 84294 87390 84346
rect 87402 84294 87454 84346
rect 87466 84294 87518 84346
rect 5882 83750 5934 83802
rect 5946 83750 5998 83802
rect 6010 83750 6062 83802
rect 6074 83750 6126 83802
rect 6138 83750 6190 83802
rect 86474 83750 86526 83802
rect 86538 83750 86590 83802
rect 86602 83750 86654 83802
rect 86666 83750 86718 83802
rect 86730 83750 86782 83802
rect 6618 83206 6670 83258
rect 6682 83206 6734 83258
rect 6746 83206 6798 83258
rect 6810 83206 6862 83258
rect 6874 83206 6926 83258
rect 87210 83206 87262 83258
rect 87274 83206 87326 83258
rect 87338 83206 87390 83258
rect 87402 83206 87454 83258
rect 87466 83206 87518 83258
rect 13876 83112 13928 83164
rect 83244 83112 83296 83164
rect 9828 83044 9880 83096
rect 12772 83044 12824 83096
rect 14980 82976 15032 83028
rect 15532 82976 15584 83028
rect 37060 82976 37112 83028
rect 37612 82976 37664 83028
rect 5882 82662 5934 82714
rect 5946 82662 5998 82714
rect 6010 82662 6062 82714
rect 6074 82662 6126 82714
rect 6138 82662 6190 82714
rect 86474 82662 86526 82714
rect 86538 82662 86590 82714
rect 86602 82662 86654 82714
rect 86666 82662 86718 82714
rect 86730 82662 86782 82714
rect 7620 82364 7672 82416
rect 11668 82364 11720 82416
rect 7804 82296 7856 82348
rect 10564 82296 10616 82348
rect 52378 82296 52430 82348
rect 52884 82296 52936 82348
rect 79978 82296 80030 82348
rect 80392 82296 80444 82348
rect 6618 82118 6670 82170
rect 6682 82118 6734 82170
rect 6746 82118 6798 82170
rect 6810 82118 6862 82170
rect 6874 82118 6926 82170
rect 87210 82118 87262 82170
rect 87274 82118 87326 82170
rect 87338 82118 87390 82170
rect 87402 82118 87454 82170
rect 87466 82118 87518 82170
rect 5882 81574 5934 81626
rect 5946 81574 5998 81626
rect 6010 81574 6062 81626
rect 6074 81574 6126 81626
rect 6138 81574 6190 81626
rect 86474 81574 86526 81626
rect 86538 81574 86590 81626
rect 86602 81574 86654 81626
rect 86666 81574 86718 81626
rect 86730 81574 86782 81626
rect 4124 81276 4176 81328
rect 8540 81276 8592 81328
rect 88212 81319 88264 81328
rect 88212 81285 88221 81319
rect 88221 81285 88255 81319
rect 88255 81285 88264 81319
rect 88212 81276 88264 81285
rect 84348 81208 84400 81260
rect 6618 81030 6670 81082
rect 6682 81030 6734 81082
rect 6746 81030 6798 81082
rect 6810 81030 6862 81082
rect 6874 81030 6926 81082
rect 87210 81030 87262 81082
rect 87274 81030 87326 81082
rect 87338 81030 87390 81082
rect 87402 81030 87454 81082
rect 87466 81030 87518 81082
rect 5882 80486 5934 80538
rect 5946 80486 5998 80538
rect 6010 80486 6062 80538
rect 6074 80486 6126 80538
rect 6138 80486 6190 80538
rect 86474 80486 86526 80538
rect 86538 80486 86590 80538
rect 86602 80486 86654 80538
rect 86666 80486 86718 80538
rect 86730 80486 86782 80538
rect 8540 80188 8592 80240
rect 88212 80231 88264 80240
rect 88212 80197 88221 80231
rect 88221 80197 88255 80231
rect 88255 80197 88264 80231
rect 88212 80188 88264 80197
rect 85820 80120 85872 80172
rect 4124 80052 4176 80104
rect 6618 79942 6670 79994
rect 6682 79942 6734 79994
rect 6746 79942 6798 79994
rect 6810 79942 6862 79994
rect 6874 79942 6926 79994
rect 87210 79942 87262 79994
rect 87274 79942 87326 79994
rect 87338 79942 87390 79994
rect 87402 79942 87454 79994
rect 87466 79942 87518 79994
rect 5882 79398 5934 79450
rect 5946 79398 5998 79450
rect 6010 79398 6062 79450
rect 6074 79398 6126 79450
rect 6138 79398 6190 79450
rect 86474 79398 86526 79450
rect 86538 79398 86590 79450
rect 86602 79398 86654 79450
rect 86666 79398 86718 79450
rect 86730 79398 86782 79450
rect 6618 78854 6670 78906
rect 6682 78854 6734 78906
rect 6746 78854 6798 78906
rect 6810 78854 6862 78906
rect 6874 78854 6926 78906
rect 87210 78854 87262 78906
rect 87274 78854 87326 78906
rect 87338 78854 87390 78906
rect 87402 78854 87454 78906
rect 87466 78854 87518 78906
rect 85820 78692 85872 78744
rect 8540 78624 8592 78676
rect 88212 78667 88264 78676
rect 88212 78633 88221 78667
rect 88221 78633 88255 78667
rect 88255 78633 88264 78667
rect 88212 78624 88264 78633
rect 4124 78488 4176 78540
rect 5882 78310 5934 78362
rect 5946 78310 5998 78362
rect 6010 78310 6062 78362
rect 6074 78310 6126 78362
rect 6138 78310 6190 78362
rect 86474 78310 86526 78362
rect 86538 78310 86590 78362
rect 86602 78310 86654 78362
rect 86666 78310 86718 78362
rect 86730 78310 86782 78362
rect 8540 78012 8592 78064
rect 88212 78055 88264 78064
rect 88212 78021 88221 78055
rect 88221 78021 88255 78055
rect 88255 78021 88264 78055
rect 88212 78012 88264 78021
rect 85820 77944 85872 77996
rect 4124 77876 4176 77928
rect 6618 77766 6670 77818
rect 6682 77766 6734 77818
rect 6746 77766 6798 77818
rect 6810 77766 6862 77818
rect 6874 77766 6926 77818
rect 87210 77766 87262 77818
rect 87274 77766 87326 77818
rect 87338 77766 87390 77818
rect 87402 77766 87454 77818
rect 87466 77766 87518 77818
rect 5882 77222 5934 77274
rect 5946 77222 5998 77274
rect 6010 77222 6062 77274
rect 6074 77222 6126 77274
rect 6138 77222 6190 77274
rect 86474 77222 86526 77274
rect 86538 77222 86590 77274
rect 86602 77222 86654 77274
rect 86666 77222 86718 77274
rect 86730 77222 86782 77274
rect 8540 76924 8592 76976
rect 4216 76788 4268 76840
rect 85820 76788 85872 76840
rect 88028 76831 88080 76840
rect 88028 76797 88037 76831
rect 88037 76797 88071 76831
rect 88071 76797 88080 76831
rect 88028 76788 88080 76797
rect 6618 76678 6670 76730
rect 6682 76678 6734 76730
rect 6746 76678 6798 76730
rect 6810 76678 6862 76730
rect 6874 76678 6926 76730
rect 87210 76678 87262 76730
rect 87274 76678 87326 76730
rect 87338 76678 87390 76730
rect 87402 76678 87454 76730
rect 87466 76678 87518 76730
rect 5882 76134 5934 76186
rect 5946 76134 5998 76186
rect 6010 76134 6062 76186
rect 6074 76134 6126 76186
rect 6138 76134 6190 76186
rect 86474 76134 86526 76186
rect 86538 76134 86590 76186
rect 86602 76134 86654 76186
rect 86666 76134 86718 76186
rect 86730 76134 86782 76186
rect 8540 75836 8592 75888
rect 88212 75879 88264 75888
rect 88212 75845 88221 75879
rect 88221 75845 88255 75879
rect 88255 75845 88264 75879
rect 88212 75836 88264 75845
rect 4124 75768 4176 75820
rect 85820 75768 85872 75820
rect 6618 75590 6670 75642
rect 6682 75590 6734 75642
rect 6746 75590 6798 75642
rect 6810 75590 6862 75642
rect 6874 75590 6926 75642
rect 87210 75590 87262 75642
rect 87274 75590 87326 75642
rect 87338 75590 87390 75642
rect 87402 75590 87454 75642
rect 87466 75590 87518 75642
rect 5882 75046 5934 75098
rect 5946 75046 5998 75098
rect 6010 75046 6062 75098
rect 6074 75046 6126 75098
rect 6138 75046 6190 75098
rect 86474 75046 86526 75098
rect 86538 75046 86590 75098
rect 86602 75046 86654 75098
rect 86666 75046 86718 75098
rect 86730 75046 86782 75098
rect 4124 74748 4176 74800
rect 5412 74791 5464 74800
rect 5412 74757 5421 74791
rect 5421 74757 5455 74791
rect 5455 74757 5464 74791
rect 5412 74748 5464 74757
rect 84532 74748 84584 74800
rect 88580 74748 88632 74800
rect 6618 74502 6670 74554
rect 6682 74502 6734 74554
rect 6746 74502 6798 74554
rect 6810 74502 6862 74554
rect 6874 74502 6926 74554
rect 87210 74502 87262 74554
rect 87274 74502 87326 74554
rect 87338 74502 87390 74554
rect 87402 74502 87454 74554
rect 87466 74502 87518 74554
rect 5882 73958 5934 74010
rect 5946 73958 5998 74010
rect 6010 73958 6062 74010
rect 6074 73958 6126 74010
rect 6138 73958 6190 74010
rect 86474 73958 86526 74010
rect 86538 73958 86590 74010
rect 86602 73958 86654 74010
rect 86666 73958 86718 74010
rect 86730 73958 86782 74010
rect 6618 73414 6670 73466
rect 6682 73414 6734 73466
rect 6746 73414 6798 73466
rect 6810 73414 6862 73466
rect 6874 73414 6926 73466
rect 87210 73414 87262 73466
rect 87274 73414 87326 73466
rect 87338 73414 87390 73466
rect 87402 73414 87454 73466
rect 87466 73414 87518 73466
rect 84808 73252 84860 73304
rect 5412 73227 5464 73236
rect 5412 73193 5421 73227
rect 5421 73193 5455 73227
rect 5455 73193 5464 73227
rect 5412 73184 5464 73193
rect 88212 73227 88264 73236
rect 88212 73193 88221 73227
rect 88221 73193 88255 73227
rect 88255 73193 88264 73227
rect 88212 73184 88264 73193
rect 4124 73048 4176 73100
rect 5882 72870 5934 72922
rect 5946 72870 5998 72922
rect 6010 72870 6062 72922
rect 6074 72870 6126 72922
rect 6138 72870 6190 72922
rect 86474 72870 86526 72922
rect 86538 72870 86590 72922
rect 86602 72870 86654 72922
rect 86666 72870 86718 72922
rect 86730 72870 86782 72922
rect 8540 72572 8592 72624
rect 88212 72615 88264 72624
rect 88212 72581 88221 72615
rect 88221 72581 88255 72615
rect 88255 72581 88264 72615
rect 88212 72572 88264 72581
rect 4124 72436 4176 72488
rect 87844 72436 87896 72488
rect 6618 72326 6670 72378
rect 6682 72326 6734 72378
rect 6746 72326 6798 72378
rect 6810 72326 6862 72378
rect 6874 72326 6926 72378
rect 87210 72326 87262 72378
rect 87274 72326 87326 72378
rect 87338 72326 87390 72378
rect 87402 72326 87454 72378
rect 87466 72326 87518 72378
rect 5882 71782 5934 71834
rect 5946 71782 5998 71834
rect 6010 71782 6062 71834
rect 6074 71782 6126 71834
rect 6138 71782 6190 71834
rect 86474 71782 86526 71834
rect 86538 71782 86590 71834
rect 86602 71782 86654 71834
rect 86666 71782 86718 71834
rect 86730 71782 86782 71834
rect 8540 71484 8592 71536
rect 88212 71527 88264 71536
rect 88212 71493 88221 71527
rect 88221 71493 88255 71527
rect 88255 71493 88264 71527
rect 88212 71484 88264 71493
rect 85820 71416 85872 71468
rect 4216 71348 4268 71400
rect 6618 71238 6670 71290
rect 6682 71238 6734 71290
rect 6746 71238 6798 71290
rect 6810 71238 6862 71290
rect 6874 71238 6926 71290
rect 87210 71238 87262 71290
rect 87274 71238 87326 71290
rect 87338 71238 87390 71290
rect 87402 71238 87454 71290
rect 87466 71238 87518 71290
rect 5882 70694 5934 70746
rect 5946 70694 5998 70746
rect 6010 70694 6062 70746
rect 6074 70694 6126 70746
rect 6138 70694 6190 70746
rect 86474 70694 86526 70746
rect 86538 70694 86590 70746
rect 86602 70694 86654 70746
rect 86666 70694 86718 70746
rect 86730 70694 86782 70746
rect 8540 70396 8592 70448
rect 88212 70439 88264 70448
rect 88212 70405 88221 70439
rect 88221 70405 88255 70439
rect 88255 70405 88264 70439
rect 88212 70396 88264 70405
rect 4124 70328 4176 70380
rect 85820 70328 85872 70380
rect 6618 70150 6670 70202
rect 6682 70150 6734 70202
rect 6746 70150 6798 70202
rect 6810 70150 6862 70202
rect 6874 70150 6926 70202
rect 87210 70150 87262 70202
rect 87274 70150 87326 70202
rect 87338 70150 87390 70202
rect 87402 70150 87454 70202
rect 87466 70150 87518 70202
rect 5882 69606 5934 69658
rect 5946 69606 5998 69658
rect 6010 69606 6062 69658
rect 6074 69606 6126 69658
rect 6138 69606 6190 69658
rect 86474 69606 86526 69658
rect 86538 69606 86590 69658
rect 86602 69606 86654 69658
rect 86666 69606 86718 69658
rect 86730 69606 86782 69658
rect 5412 69351 5464 69360
rect 5412 69317 5421 69351
rect 5421 69317 5455 69351
rect 5455 69317 5464 69351
rect 5412 69308 5464 69317
rect 88580 69308 88632 69360
rect 4124 69240 4176 69292
rect 84808 69240 84860 69292
rect 6618 69062 6670 69114
rect 6682 69062 6734 69114
rect 6746 69062 6798 69114
rect 6810 69062 6862 69114
rect 6874 69062 6926 69114
rect 87210 69062 87262 69114
rect 87274 69062 87326 69114
rect 87338 69062 87390 69114
rect 87402 69062 87454 69114
rect 87466 69062 87518 69114
rect 5882 68518 5934 68570
rect 5946 68518 5998 68570
rect 6010 68518 6062 68570
rect 6074 68518 6126 68570
rect 6138 68518 6190 68570
rect 86474 68518 86526 68570
rect 86538 68518 86590 68570
rect 86602 68518 86654 68570
rect 86666 68518 86718 68570
rect 86730 68518 86782 68570
rect 6618 67974 6670 68026
rect 6682 67974 6734 68026
rect 6746 67974 6798 68026
rect 6810 67974 6862 68026
rect 6874 67974 6926 68026
rect 87210 67974 87262 68026
rect 87274 67974 87326 68026
rect 87338 67974 87390 68026
rect 87402 67974 87454 68026
rect 87466 67974 87518 68026
rect 85268 67812 85320 67864
rect 5412 67787 5464 67796
rect 5412 67753 5421 67787
rect 5421 67753 5455 67787
rect 5455 67753 5464 67787
rect 5412 67744 5464 67753
rect 88212 67787 88264 67796
rect 88212 67753 88221 67787
rect 88221 67753 88255 67787
rect 88255 67753 88264 67787
rect 88212 67744 88264 67753
rect 4032 67608 4084 67660
rect 5882 67430 5934 67482
rect 5946 67430 5998 67482
rect 6010 67430 6062 67482
rect 6074 67430 6126 67482
rect 6138 67430 6190 67482
rect 86474 67430 86526 67482
rect 86538 67430 86590 67482
rect 86602 67430 86654 67482
rect 86666 67430 86718 67482
rect 86730 67430 86782 67482
rect 8540 67132 8592 67184
rect 88212 67175 88264 67184
rect 88212 67141 88221 67175
rect 88221 67141 88255 67175
rect 88255 67141 88264 67175
rect 88212 67132 88264 67141
rect 85820 67064 85872 67116
rect 4124 66996 4176 67048
rect 6618 66886 6670 66938
rect 6682 66886 6734 66938
rect 6746 66886 6798 66938
rect 6810 66886 6862 66938
rect 6874 66886 6926 66938
rect 87210 66886 87262 66938
rect 87274 66886 87326 66938
rect 87338 66886 87390 66938
rect 87402 66886 87454 66938
rect 87466 66886 87518 66938
rect 5882 66342 5934 66394
rect 5946 66342 5998 66394
rect 6010 66342 6062 66394
rect 6074 66342 6126 66394
rect 6138 66342 6190 66394
rect 86474 66342 86526 66394
rect 86538 66342 86590 66394
rect 86602 66342 86654 66394
rect 86666 66342 86718 66394
rect 86730 66342 86782 66394
rect 8540 66112 8592 66164
rect 4308 66044 4360 66096
rect 85820 66044 85872 66096
rect 88212 65908 88264 65960
rect 6618 65798 6670 65850
rect 6682 65798 6734 65850
rect 6746 65798 6798 65850
rect 6810 65798 6862 65850
rect 6874 65798 6926 65850
rect 87210 65798 87262 65850
rect 87274 65798 87326 65850
rect 87338 65798 87390 65850
rect 87402 65798 87454 65850
rect 87466 65798 87518 65850
rect 5882 65254 5934 65306
rect 5946 65254 5998 65306
rect 6010 65254 6062 65306
rect 6074 65254 6126 65306
rect 6138 65254 6190 65306
rect 86474 65254 86526 65306
rect 86538 65254 86590 65306
rect 86602 65254 86654 65306
rect 86666 65254 86718 65306
rect 86730 65254 86782 65306
rect 8540 65024 8592 65076
rect 4308 64956 4360 65008
rect 85820 64956 85872 65008
rect 88396 64820 88448 64872
rect 6618 64710 6670 64762
rect 6682 64710 6734 64762
rect 6746 64710 6798 64762
rect 6810 64710 6862 64762
rect 6874 64710 6926 64762
rect 87210 64710 87262 64762
rect 87274 64710 87326 64762
rect 87338 64710 87390 64762
rect 87402 64710 87454 64762
rect 87466 64710 87518 64762
rect 7528 64591 7580 64600
rect 7528 64557 7537 64591
rect 7537 64557 7571 64591
rect 7571 64557 7580 64591
rect 7528 64548 7580 64557
rect 5882 64166 5934 64218
rect 5946 64166 5998 64218
rect 6010 64166 6062 64218
rect 6074 64166 6126 64218
rect 6138 64166 6190 64218
rect 86474 64166 86526 64218
rect 86538 64166 86590 64218
rect 86602 64166 86654 64218
rect 86666 64166 86718 64218
rect 86730 64166 86782 64218
rect 4308 63868 4360 63920
rect 7528 63868 7580 63920
rect 84532 63868 84584 63920
rect 5688 63732 5740 63784
rect 7804 63732 7856 63784
rect 88580 63732 88632 63784
rect 6618 63622 6670 63674
rect 6682 63622 6734 63674
rect 6746 63622 6798 63674
rect 6810 63622 6862 63674
rect 6874 63622 6926 63674
rect 87210 63622 87262 63674
rect 87274 63622 87326 63674
rect 87338 63622 87390 63674
rect 87402 63622 87454 63674
rect 87466 63622 87518 63674
rect 7344 63460 7396 63512
rect 7804 63460 7856 63512
rect 5882 63078 5934 63130
rect 5946 63078 5998 63130
rect 6010 63078 6062 63130
rect 6074 63078 6126 63130
rect 6138 63078 6190 63130
rect 86474 63078 86526 63130
rect 86538 63078 86590 63130
rect 86602 63078 86654 63130
rect 86666 63078 86718 63130
rect 86730 63078 86782 63130
rect 6618 62534 6670 62586
rect 6682 62534 6734 62586
rect 6746 62534 6798 62586
rect 6810 62534 6862 62586
rect 6874 62534 6926 62586
rect 87210 62534 87262 62586
rect 87274 62534 87326 62586
rect 87338 62534 87390 62586
rect 87402 62534 87454 62586
rect 87466 62534 87518 62586
rect 4308 62304 4360 62356
rect 84808 62304 84860 62356
rect 5688 62168 5740 62220
rect 88396 62100 88448 62152
rect 5882 61990 5934 62042
rect 5946 61990 5998 62042
rect 6010 61990 6062 62042
rect 6074 61990 6126 62042
rect 6138 61990 6190 62042
rect 86474 61990 86526 62042
rect 86538 61990 86590 62042
rect 86602 61990 86654 62042
rect 86666 61990 86718 62042
rect 86730 61990 86782 62042
rect 4308 61692 4360 61744
rect 85820 61692 85872 61744
rect 8540 61624 8592 61676
rect 88212 61556 88264 61608
rect 6618 61446 6670 61498
rect 6682 61446 6734 61498
rect 6746 61446 6798 61498
rect 6810 61446 6862 61498
rect 6874 61446 6926 61498
rect 87210 61446 87262 61498
rect 87274 61446 87326 61498
rect 87338 61446 87390 61498
rect 87402 61446 87454 61498
rect 87466 61446 87518 61498
rect 5882 60902 5934 60954
rect 5946 60902 5998 60954
rect 6010 60902 6062 60954
rect 6074 60902 6126 60954
rect 6138 60902 6190 60954
rect 86474 60902 86526 60954
rect 86538 60902 86590 60954
rect 86602 60902 86654 60954
rect 86666 60902 86718 60954
rect 86730 60902 86782 60954
rect 4308 60604 4360 60656
rect 85820 60604 85872 60656
rect 8540 60536 8592 60588
rect 88212 60468 88264 60520
rect 6618 60358 6670 60410
rect 6682 60358 6734 60410
rect 6746 60358 6798 60410
rect 6810 60358 6862 60410
rect 6874 60358 6926 60410
rect 87210 60358 87262 60410
rect 87274 60358 87326 60410
rect 87338 60358 87390 60410
rect 87402 60358 87454 60410
rect 87466 60358 87518 60410
rect 5882 59814 5934 59866
rect 5946 59814 5998 59866
rect 6010 59814 6062 59866
rect 6074 59814 6126 59866
rect 6138 59814 6190 59866
rect 86474 59814 86526 59866
rect 86538 59814 86590 59866
rect 86602 59814 86654 59866
rect 86666 59814 86718 59866
rect 86730 59814 86782 59866
rect 4308 59516 4360 59568
rect 87476 59516 87528 59568
rect 8540 59448 8592 59500
rect 88212 59380 88264 59432
rect 6618 59270 6670 59322
rect 6682 59270 6734 59322
rect 6746 59270 6798 59322
rect 6810 59270 6862 59322
rect 6874 59270 6926 59322
rect 87210 59270 87262 59322
rect 87274 59270 87326 59322
rect 87338 59270 87390 59322
rect 87402 59270 87454 59322
rect 87466 59270 87518 59322
rect 5882 58726 5934 58778
rect 5946 58726 5998 58778
rect 6010 58726 6062 58778
rect 6074 58726 6126 58778
rect 6138 58726 6190 58778
rect 86474 58726 86526 58778
rect 86538 58726 86590 58778
rect 86602 58726 86654 58778
rect 86666 58726 86718 58778
rect 86730 58726 86782 58778
rect 4308 58428 4360 58480
rect 85084 58428 85136 58480
rect 5412 58292 5464 58344
rect 88580 58292 88632 58344
rect 6618 58182 6670 58234
rect 6682 58182 6734 58234
rect 6746 58182 6798 58234
rect 6810 58182 6862 58234
rect 6874 58182 6926 58234
rect 87210 58182 87262 58234
rect 87274 58182 87326 58234
rect 87338 58182 87390 58234
rect 87402 58182 87454 58234
rect 87466 58182 87518 58234
rect 5882 57638 5934 57690
rect 5946 57638 5998 57690
rect 6010 57638 6062 57690
rect 6074 57638 6126 57690
rect 6138 57638 6190 57690
rect 86474 57638 86526 57690
rect 86538 57638 86590 57690
rect 86602 57638 86654 57690
rect 86666 57638 86718 57690
rect 86730 57638 86782 57690
rect 6618 57094 6670 57146
rect 6682 57094 6734 57146
rect 6746 57094 6798 57146
rect 6810 57094 6862 57146
rect 6874 57094 6926 57146
rect 87210 57094 87262 57146
rect 87274 57094 87326 57146
rect 87338 57094 87390 57146
rect 87402 57094 87454 57146
rect 87466 57094 87518 57146
rect 9920 56932 9972 56984
rect 88580 56932 88632 56984
rect 4308 56864 4360 56916
rect 87568 56864 87620 56916
rect 5882 56550 5934 56602
rect 5946 56550 5998 56602
rect 6010 56550 6062 56602
rect 6074 56550 6126 56602
rect 6138 56550 6190 56602
rect 86474 56550 86526 56602
rect 86538 56550 86590 56602
rect 86602 56550 86654 56602
rect 86666 56550 86718 56602
rect 86730 56550 86782 56602
rect 9920 56320 9972 56372
rect 4308 56252 4360 56304
rect 85820 56252 85872 56304
rect 88212 56116 88264 56168
rect 6618 56006 6670 56058
rect 6682 56006 6734 56058
rect 6746 56006 6798 56058
rect 6810 56006 6862 56058
rect 6874 56006 6926 56058
rect 87210 56006 87262 56058
rect 87274 56006 87326 56058
rect 87338 56006 87390 56058
rect 87402 56006 87454 56058
rect 87466 56006 87518 56058
rect 5882 55462 5934 55514
rect 5946 55462 5998 55514
rect 6010 55462 6062 55514
rect 6074 55462 6126 55514
rect 6138 55462 6190 55514
rect 86474 55462 86526 55514
rect 86538 55462 86590 55514
rect 86602 55462 86654 55514
rect 86666 55462 86718 55514
rect 86730 55462 86782 55514
rect 8540 55232 8592 55284
rect 4308 55164 4360 55216
rect 85820 55164 85872 55216
rect 88212 55028 88264 55080
rect 6618 54918 6670 54970
rect 6682 54918 6734 54970
rect 6746 54918 6798 54970
rect 6810 54918 6862 54970
rect 6874 54918 6926 54970
rect 87210 54918 87262 54970
rect 87274 54918 87326 54970
rect 87338 54918 87390 54970
rect 87402 54918 87454 54970
rect 87466 54918 87518 54970
rect 5882 54374 5934 54426
rect 5946 54374 5998 54426
rect 6010 54374 6062 54426
rect 6074 54374 6126 54426
rect 6138 54374 6190 54426
rect 86474 54374 86526 54426
rect 86538 54374 86590 54426
rect 86602 54374 86654 54426
rect 86666 54374 86718 54426
rect 86730 54374 86782 54426
rect 5688 54144 5740 54196
rect 4308 54076 4360 54128
rect 84532 54076 84584 54128
rect 88212 54076 88264 54128
rect 6618 53830 6670 53882
rect 6682 53830 6734 53882
rect 6746 53830 6798 53882
rect 6810 53830 6862 53882
rect 6874 53830 6926 53882
rect 87210 53830 87262 53882
rect 87274 53830 87326 53882
rect 87338 53830 87390 53882
rect 87402 53830 87454 53882
rect 87466 53830 87518 53882
rect 5882 53286 5934 53338
rect 5946 53286 5998 53338
rect 6010 53286 6062 53338
rect 6074 53286 6126 53338
rect 6138 53286 6190 53338
rect 86474 53286 86526 53338
rect 86538 53286 86590 53338
rect 86602 53286 86654 53338
rect 86666 53286 86718 53338
rect 86730 53286 86782 53338
rect 8540 53056 8592 53108
rect 4308 52988 4360 53040
rect 87568 52988 87620 53040
rect 88212 52852 88264 52904
rect 6618 52742 6670 52794
rect 6682 52742 6734 52794
rect 6746 52742 6798 52794
rect 6810 52742 6862 52794
rect 6874 52742 6926 52794
rect 87210 52742 87262 52794
rect 87274 52742 87326 52794
rect 87338 52742 87390 52794
rect 87402 52742 87454 52794
rect 87466 52742 87518 52794
rect 5882 52198 5934 52250
rect 5946 52198 5998 52250
rect 6010 52198 6062 52250
rect 6074 52198 6126 52250
rect 6138 52198 6190 52250
rect 86474 52198 86526 52250
rect 86538 52198 86590 52250
rect 86602 52198 86654 52250
rect 86666 52198 86718 52250
rect 86730 52198 86782 52250
rect 6618 51654 6670 51706
rect 6682 51654 6734 51706
rect 6746 51654 6798 51706
rect 6810 51654 6862 51706
rect 6874 51654 6926 51706
rect 87210 51654 87262 51706
rect 87274 51654 87326 51706
rect 87338 51654 87390 51706
rect 87402 51654 87454 51706
rect 87466 51654 87518 51706
rect 8540 51492 8592 51544
rect 4308 51424 4360 51476
rect 87568 51424 87620 51476
rect 88212 51288 88264 51340
rect 5882 51110 5934 51162
rect 5946 51110 5998 51162
rect 6010 51110 6062 51162
rect 6074 51110 6126 51162
rect 6138 51110 6190 51162
rect 86474 51110 86526 51162
rect 86538 51110 86590 51162
rect 86602 51110 86654 51162
rect 86666 51110 86718 51162
rect 86730 51110 86782 51162
rect 85636 50719 85688 50728
rect 85636 50685 85645 50719
rect 85645 50685 85679 50719
rect 85679 50685 85688 50719
rect 85636 50676 85688 50685
rect 6618 50566 6670 50618
rect 6682 50566 6734 50618
rect 6746 50566 6798 50618
rect 6810 50566 6862 50618
rect 6874 50566 6926 50618
rect 87210 50566 87262 50618
rect 87274 50566 87326 50618
rect 87338 50566 87390 50618
rect 87402 50566 87454 50618
rect 87466 50566 87518 50618
rect 5882 50022 5934 50074
rect 5946 50022 5998 50074
rect 6010 50022 6062 50074
rect 6074 50022 6126 50074
rect 6138 50022 6190 50074
rect 86474 50022 86526 50074
rect 86538 50022 86590 50074
rect 86602 50022 86654 50074
rect 86666 50022 86718 50074
rect 86730 50022 86782 50074
rect 85636 49631 85688 49640
rect 85636 49597 85645 49631
rect 85645 49597 85679 49631
rect 85679 49597 85688 49631
rect 85636 49588 85688 49597
rect 6618 49478 6670 49530
rect 6682 49478 6734 49530
rect 6746 49478 6798 49530
rect 6810 49478 6862 49530
rect 6874 49478 6926 49530
rect 87210 49478 87262 49530
rect 87274 49478 87326 49530
rect 87338 49478 87390 49530
rect 87402 49478 87454 49530
rect 87466 49478 87518 49530
rect 5882 48934 5934 48986
rect 5946 48934 5998 48986
rect 6010 48934 6062 48986
rect 6074 48934 6126 48986
rect 6138 48934 6190 48986
rect 86474 48934 86526 48986
rect 86538 48934 86590 48986
rect 86602 48934 86654 48986
rect 86666 48934 86718 48986
rect 86730 48934 86782 48986
rect 88212 48679 88264 48688
rect 88212 48645 88221 48679
rect 88221 48645 88255 48679
rect 88255 48645 88264 48679
rect 88212 48636 88264 48645
rect 85360 48568 85412 48620
rect 6618 48390 6670 48442
rect 6682 48390 6734 48442
rect 6746 48390 6798 48442
rect 6810 48390 6862 48442
rect 6874 48390 6926 48442
rect 87210 48390 87262 48442
rect 87274 48390 87326 48442
rect 87338 48390 87390 48442
rect 87402 48390 87454 48442
rect 87466 48390 87518 48442
rect 88212 47999 88264 48008
rect 88212 47965 88221 47999
rect 88221 47965 88255 47999
rect 88255 47965 88264 47999
rect 88212 47956 88264 47965
rect 5882 47846 5934 47898
rect 5946 47846 5998 47898
rect 6010 47846 6062 47898
rect 6074 47846 6126 47898
rect 6138 47846 6190 47898
rect 86474 47846 86526 47898
rect 86538 47846 86590 47898
rect 86602 47846 86654 47898
rect 86666 47846 86718 47898
rect 86730 47846 86782 47898
rect 85820 47548 85872 47600
rect 88212 47412 88264 47464
rect 6618 47302 6670 47354
rect 6682 47302 6734 47354
rect 6746 47302 6798 47354
rect 6810 47302 6862 47354
rect 6874 47302 6926 47354
rect 87210 47302 87262 47354
rect 87274 47302 87326 47354
rect 87338 47302 87390 47354
rect 87402 47302 87454 47354
rect 87466 47302 87518 47354
rect 88212 46911 88264 46920
rect 88212 46877 88221 46911
rect 88221 46877 88255 46911
rect 88255 46877 88264 46911
rect 88212 46868 88264 46877
rect 5882 46758 5934 46810
rect 5946 46758 5998 46810
rect 6010 46758 6062 46810
rect 6074 46758 6126 46810
rect 6138 46758 6190 46810
rect 86474 46758 86526 46810
rect 86538 46758 86590 46810
rect 86602 46758 86654 46810
rect 86666 46758 86718 46810
rect 86730 46758 86782 46810
rect 6618 46214 6670 46266
rect 6682 46214 6734 46266
rect 6746 46214 6798 46266
rect 6810 46214 6862 46266
rect 6874 46214 6926 46266
rect 87210 46214 87262 46266
rect 87274 46214 87326 46266
rect 87338 46214 87390 46266
rect 87402 46214 87454 46266
rect 87466 46214 87518 46266
rect 46996 45984 47048 46036
rect 50170 45916 50222 45968
rect 51136 45916 51188 45968
rect 5882 45670 5934 45722
rect 5946 45670 5998 45722
rect 6010 45670 6062 45722
rect 6074 45670 6126 45722
rect 6138 45670 6190 45722
rect 7344 45551 7396 45560
rect 7344 45517 7353 45551
rect 7353 45517 7387 45551
rect 7387 45517 7396 45551
rect 10564 45848 10616 45900
rect 46444 45848 46496 45900
rect 51274 45848 51326 45900
rect 85820 45848 85872 45900
rect 86474 45670 86526 45722
rect 86538 45670 86590 45722
rect 86602 45670 86654 45722
rect 86666 45670 86718 45722
rect 86730 45670 86782 45722
rect 7344 45508 7396 45517
rect 85820 45551 85872 45560
rect 85820 45517 85829 45551
rect 85829 45517 85863 45551
rect 85863 45517 85872 45551
rect 85820 45508 85872 45517
rect 9000 45440 9052 45492
rect 4308 45372 4360 45424
rect 86004 45415 86056 45424
rect 86004 45381 86013 45415
rect 86013 45381 86047 45415
rect 86047 45381 86056 45415
rect 86004 45372 86056 45381
rect 88212 45415 88264 45424
rect 88212 45381 88221 45415
rect 88221 45381 88255 45415
rect 88255 45381 88264 45415
rect 88212 45372 88264 45381
rect 5688 45304 5740 45356
rect 85636 45279 85688 45288
rect 85636 45245 85645 45279
rect 85645 45245 85679 45279
rect 85679 45245 85688 45279
rect 85636 45236 85688 45245
rect 86188 45279 86240 45288
rect 86188 45245 86197 45279
rect 86197 45245 86231 45279
rect 86231 45245 86240 45279
rect 86188 45236 86240 45245
rect 6618 45126 6670 45178
rect 6682 45126 6734 45178
rect 6746 45126 6798 45178
rect 6810 45126 6862 45178
rect 6874 45126 6926 45178
rect 87210 45126 87262 45178
rect 87274 45126 87326 45178
rect 87338 45126 87390 45178
rect 87402 45126 87454 45178
rect 87466 45126 87518 45178
rect 7620 44964 7672 45016
rect 8540 44896 8592 44948
rect 4216 44692 4268 44744
rect 88212 44735 88264 44744
rect 88212 44701 88221 44735
rect 88221 44701 88255 44735
rect 88255 44701 88264 44735
rect 88212 44692 88264 44701
rect 5882 44582 5934 44634
rect 5946 44582 5998 44634
rect 6010 44582 6062 44634
rect 6074 44582 6126 44634
rect 6138 44582 6190 44634
rect 86474 44582 86526 44634
rect 86538 44582 86590 44634
rect 86602 44582 86654 44634
rect 86666 44582 86718 44634
rect 86730 44582 86782 44634
rect 83612 44352 83664 44404
rect 88212 44327 88264 44336
rect 88212 44293 88221 44327
rect 88221 44293 88255 44327
rect 88255 44293 88264 44327
rect 88212 44284 88264 44293
rect 6618 44038 6670 44090
rect 6682 44038 6734 44090
rect 6746 44038 6798 44090
rect 6810 44038 6862 44090
rect 6874 44038 6926 44090
rect 87210 44038 87262 44090
rect 87274 44038 87326 44090
rect 87338 44038 87390 44090
rect 87402 44038 87454 44090
rect 87466 44038 87518 44090
rect 5882 43494 5934 43546
rect 5946 43494 5998 43546
rect 6010 43494 6062 43546
rect 6074 43494 6126 43546
rect 6138 43494 6190 43546
rect 86474 43494 86526 43546
rect 86538 43494 86590 43546
rect 86602 43494 86654 43546
rect 86666 43494 86718 43546
rect 86730 43494 86782 43546
rect 85820 43332 85872 43384
rect 4124 43196 4176 43248
rect 8540 43196 8592 43248
rect 88212 43239 88264 43248
rect 88212 43205 88221 43239
rect 88221 43205 88255 43239
rect 88255 43205 88264 43239
rect 88212 43196 88264 43205
rect 6618 42950 6670 43002
rect 6682 42950 6734 43002
rect 6746 42950 6798 43002
rect 6810 42950 6862 43002
rect 6874 42950 6926 43002
rect 87210 42950 87262 43002
rect 87274 42950 87326 43002
rect 87338 42950 87390 43002
rect 87402 42950 87454 43002
rect 87466 42950 87518 43002
rect 8540 42720 8592 42772
rect 88212 42763 88264 42772
rect 88212 42729 88221 42763
rect 88221 42729 88255 42763
rect 88255 42729 88264 42763
rect 88212 42720 88264 42729
rect 85820 42584 85872 42636
rect 4124 42516 4176 42568
rect 5882 42406 5934 42458
rect 5946 42406 5998 42458
rect 6010 42406 6062 42458
rect 6074 42406 6126 42458
rect 6138 42406 6190 42458
rect 86474 42406 86526 42458
rect 86538 42406 86590 42458
rect 86602 42406 86654 42458
rect 86666 42406 86718 42458
rect 86730 42406 86782 42458
rect 6618 41862 6670 41914
rect 6682 41862 6734 41914
rect 6746 41862 6798 41914
rect 6810 41862 6862 41914
rect 6874 41862 6926 41914
rect 87210 41862 87262 41914
rect 87274 41862 87326 41914
rect 87338 41862 87390 41914
rect 87402 41862 87454 41914
rect 87466 41862 87518 41914
rect 4124 41632 4176 41684
rect 5412 41675 5464 41684
rect 5412 41641 5421 41675
rect 5421 41641 5455 41675
rect 5455 41641 5464 41675
rect 5412 41632 5464 41641
rect 87568 41632 87620 41684
rect 88212 41675 88264 41684
rect 88212 41641 88221 41675
rect 88221 41641 88255 41675
rect 88255 41641 88264 41675
rect 88212 41632 88264 41641
rect 5882 41318 5934 41370
rect 5946 41318 5998 41370
rect 6010 41318 6062 41370
rect 6074 41318 6126 41370
rect 6138 41318 6190 41370
rect 86474 41318 86526 41370
rect 86538 41318 86590 41370
rect 86602 41318 86654 41370
rect 86666 41318 86718 41370
rect 86730 41318 86782 41370
rect 6618 40774 6670 40826
rect 6682 40774 6734 40826
rect 6746 40774 6798 40826
rect 6810 40774 6862 40826
rect 6874 40774 6926 40826
rect 87210 40774 87262 40826
rect 87274 40774 87326 40826
rect 87338 40774 87390 40826
rect 87402 40774 87454 40826
rect 87466 40774 87518 40826
rect 8540 40544 8592 40596
rect 87936 40519 87988 40528
rect 87936 40485 87945 40519
rect 87945 40485 87979 40519
rect 87979 40485 87988 40519
rect 87936 40476 87988 40485
rect 88212 40519 88264 40528
rect 88212 40485 88221 40519
rect 88221 40485 88255 40519
rect 88255 40485 88264 40519
rect 88212 40476 88264 40485
rect 3940 40408 3992 40460
rect 5882 40230 5934 40282
rect 5946 40230 5998 40282
rect 6010 40230 6062 40282
rect 6074 40230 6126 40282
rect 6138 40230 6190 40282
rect 86474 40230 86526 40282
rect 86538 40230 86590 40282
rect 86602 40230 86654 40282
rect 86666 40230 86718 40282
rect 86730 40230 86782 40282
rect 88212 40111 88264 40120
rect 88212 40077 88221 40111
rect 88221 40077 88255 40111
rect 88255 40077 88264 40111
rect 88212 40068 88264 40077
rect 6618 39686 6670 39738
rect 6682 39686 6734 39738
rect 6746 39686 6798 39738
rect 6810 39686 6862 39738
rect 6874 39686 6926 39738
rect 87210 39686 87262 39738
rect 87274 39686 87326 39738
rect 87338 39686 87390 39738
rect 87402 39686 87454 39738
rect 87466 39686 87518 39738
rect 8540 39456 8592 39508
rect 88212 39499 88264 39508
rect 88212 39465 88221 39499
rect 88221 39465 88255 39499
rect 88255 39465 88264 39499
rect 88212 39456 88264 39465
rect 87568 39320 87620 39372
rect 4216 39252 4268 39304
rect 5882 39142 5934 39194
rect 5946 39142 5998 39194
rect 6010 39142 6062 39194
rect 6074 39142 6126 39194
rect 6138 39142 6190 39194
rect 86474 39142 86526 39194
rect 86538 39142 86590 39194
rect 86602 39142 86654 39194
rect 86666 39142 86718 39194
rect 86730 39142 86782 39194
rect 6618 38598 6670 38650
rect 6682 38598 6734 38650
rect 6746 38598 6798 38650
rect 6810 38598 6862 38650
rect 6874 38598 6926 38650
rect 87210 38598 87262 38650
rect 87274 38598 87326 38650
rect 87338 38598 87390 38650
rect 87402 38598 87454 38650
rect 87466 38598 87518 38650
rect 5882 38054 5934 38106
rect 5946 38054 5998 38106
rect 6010 38054 6062 38106
rect 6074 38054 6126 38106
rect 6138 38054 6190 38106
rect 86474 38054 86526 38106
rect 86538 38054 86590 38106
rect 86602 38054 86654 38106
rect 86666 38054 86718 38106
rect 86730 38054 86782 38106
rect 85820 37892 85872 37944
rect 4216 37756 4268 37808
rect 8540 37756 8592 37808
rect 88212 37799 88264 37808
rect 88212 37765 88221 37799
rect 88221 37765 88255 37799
rect 88255 37765 88264 37799
rect 88212 37756 88264 37765
rect 6618 37510 6670 37562
rect 6682 37510 6734 37562
rect 6746 37510 6798 37562
rect 6810 37510 6862 37562
rect 6874 37510 6926 37562
rect 87210 37510 87262 37562
rect 87274 37510 87326 37562
rect 87338 37510 87390 37562
rect 87402 37510 87454 37562
rect 87466 37510 87518 37562
rect 8540 37280 8592 37332
rect 88212 37323 88264 37332
rect 88212 37289 88221 37323
rect 88221 37289 88255 37323
rect 88255 37289 88264 37323
rect 88212 37280 88264 37289
rect 85820 37144 85872 37196
rect 4124 37076 4176 37128
rect 5882 36966 5934 37018
rect 5946 36966 5998 37018
rect 6010 36966 6062 37018
rect 6074 36966 6126 37018
rect 6138 36966 6190 37018
rect 86474 36966 86526 37018
rect 86538 36966 86590 37018
rect 86602 36966 86654 37018
rect 86666 36966 86718 37018
rect 86730 36966 86782 37018
rect 6618 36422 6670 36474
rect 6682 36422 6734 36474
rect 6746 36422 6798 36474
rect 6810 36422 6862 36474
rect 6874 36422 6926 36474
rect 87210 36422 87262 36474
rect 87274 36422 87326 36474
rect 87338 36422 87390 36474
rect 87402 36422 87454 36474
rect 87466 36422 87518 36474
rect 5412 36235 5464 36244
rect 5412 36201 5421 36235
rect 5421 36201 5455 36235
rect 5455 36201 5464 36235
rect 5412 36192 5464 36201
rect 88580 36192 88632 36244
rect 4124 36124 4176 36176
rect 84808 36124 84860 36176
rect 5882 35878 5934 35930
rect 5946 35878 5998 35930
rect 6010 35878 6062 35930
rect 6074 35878 6126 35930
rect 6138 35878 6190 35930
rect 86474 35878 86526 35930
rect 86538 35878 86590 35930
rect 86602 35878 86654 35930
rect 86666 35878 86718 35930
rect 86730 35878 86782 35930
rect 6618 35334 6670 35386
rect 6682 35334 6734 35386
rect 6746 35334 6798 35386
rect 6810 35334 6862 35386
rect 6874 35334 6926 35386
rect 87210 35334 87262 35386
rect 87274 35334 87326 35386
rect 87338 35334 87390 35386
rect 87402 35334 87454 35386
rect 87466 35334 87518 35386
rect 8540 35104 8592 35156
rect 88212 35147 88264 35156
rect 88212 35113 88221 35147
rect 88221 35113 88255 35147
rect 88255 35113 88264 35147
rect 88212 35104 88264 35113
rect 4216 35036 4268 35088
rect 85820 34968 85872 35020
rect 5882 34790 5934 34842
rect 5946 34790 5998 34842
rect 6010 34790 6062 34842
rect 6074 34790 6126 34842
rect 6138 34790 6190 34842
rect 86474 34790 86526 34842
rect 86538 34790 86590 34842
rect 86602 34790 86654 34842
rect 86666 34790 86718 34842
rect 86730 34790 86782 34842
rect 6618 34246 6670 34298
rect 6682 34246 6734 34298
rect 6746 34246 6798 34298
rect 6810 34246 6862 34298
rect 6874 34246 6926 34298
rect 87210 34246 87262 34298
rect 87274 34246 87326 34298
rect 87338 34246 87390 34298
rect 87402 34246 87454 34298
rect 87466 34246 87518 34298
rect 8540 34016 8592 34068
rect 88212 34059 88264 34068
rect 88212 34025 88221 34059
rect 88221 34025 88255 34059
rect 88255 34025 88264 34059
rect 88212 34016 88264 34025
rect 85820 33880 85872 33932
rect 4216 33812 4268 33864
rect 5882 33702 5934 33754
rect 5946 33702 5998 33754
rect 6010 33702 6062 33754
rect 6074 33702 6126 33754
rect 6138 33702 6190 33754
rect 86474 33702 86526 33754
rect 86538 33702 86590 33754
rect 86602 33702 86654 33754
rect 86666 33702 86718 33754
rect 86730 33702 86782 33754
rect 6618 33158 6670 33210
rect 6682 33158 6734 33210
rect 6746 33158 6798 33210
rect 6810 33158 6862 33210
rect 6874 33158 6926 33210
rect 87210 33158 87262 33210
rect 87274 33158 87326 33210
rect 87338 33158 87390 33210
rect 87402 33158 87454 33210
rect 87466 33158 87518 33210
rect 5882 32614 5934 32666
rect 5946 32614 5998 32666
rect 6010 32614 6062 32666
rect 6074 32614 6126 32666
rect 6138 32614 6190 32666
rect 86474 32614 86526 32666
rect 86538 32614 86590 32666
rect 86602 32614 86654 32666
rect 86666 32614 86718 32666
rect 86730 32614 86782 32666
rect 85820 32452 85872 32504
rect 4216 32316 4268 32368
rect 8540 32316 8592 32368
rect 88212 32359 88264 32368
rect 88212 32325 88221 32359
rect 88221 32325 88255 32359
rect 88255 32325 88264 32359
rect 88212 32316 88264 32325
rect 6618 32070 6670 32122
rect 6682 32070 6734 32122
rect 6746 32070 6798 32122
rect 6810 32070 6862 32122
rect 6874 32070 6926 32122
rect 87210 32070 87262 32122
rect 87274 32070 87326 32122
rect 87338 32070 87390 32122
rect 87402 32070 87454 32122
rect 87466 32070 87518 32122
rect 8540 31840 8592 31892
rect 88212 31883 88264 31892
rect 88212 31849 88221 31883
rect 88221 31849 88255 31883
rect 88255 31849 88264 31883
rect 88212 31840 88264 31849
rect 85820 31704 85872 31756
rect 4124 31636 4176 31688
rect 5882 31526 5934 31578
rect 5946 31526 5998 31578
rect 6010 31526 6062 31578
rect 6074 31526 6126 31578
rect 6138 31526 6190 31578
rect 86474 31526 86526 31578
rect 86538 31526 86590 31578
rect 86602 31526 86654 31578
rect 86666 31526 86718 31578
rect 86730 31526 86782 31578
rect 6618 30982 6670 31034
rect 6682 30982 6734 31034
rect 6746 30982 6798 31034
rect 6810 30982 6862 31034
rect 6874 30982 6926 31034
rect 87210 30982 87262 31034
rect 87274 30982 87326 31034
rect 87338 30982 87390 31034
rect 87402 30982 87454 31034
rect 87466 30982 87518 31034
rect 5412 30795 5464 30804
rect 5412 30761 5421 30795
rect 5421 30761 5455 30795
rect 5455 30761 5464 30795
rect 5412 30752 5464 30761
rect 88580 30752 88632 30804
rect 4124 30616 4176 30668
rect 84808 30616 84860 30668
rect 5882 30438 5934 30490
rect 5946 30438 5998 30490
rect 6010 30438 6062 30490
rect 6074 30438 6126 30490
rect 6138 30438 6190 30490
rect 86474 30438 86526 30490
rect 86538 30438 86590 30490
rect 86602 30438 86654 30490
rect 86666 30438 86718 30490
rect 86730 30438 86782 30490
rect 6618 29894 6670 29946
rect 6682 29894 6734 29946
rect 6746 29894 6798 29946
rect 6810 29894 6862 29946
rect 6874 29894 6926 29946
rect 87210 29894 87262 29946
rect 87274 29894 87326 29946
rect 87338 29894 87390 29946
rect 87402 29894 87454 29946
rect 87466 29894 87518 29946
rect 4308 29664 4360 29716
rect 85820 29664 85872 29716
rect 8540 29528 8592 29580
rect 88396 29460 88448 29512
rect 5882 29350 5934 29402
rect 5946 29350 5998 29402
rect 6010 29350 6062 29402
rect 6074 29350 6126 29402
rect 6138 29350 6190 29402
rect 86474 29350 86526 29402
rect 86538 29350 86590 29402
rect 86602 29350 86654 29402
rect 86666 29350 86718 29402
rect 86730 29350 86782 29402
rect 6618 28806 6670 28858
rect 6682 28806 6734 28858
rect 6746 28806 6798 28858
rect 6810 28806 6862 28858
rect 6874 28806 6926 28858
rect 87210 28806 87262 28858
rect 87274 28806 87326 28858
rect 87338 28806 87390 28858
rect 87402 28806 87454 28858
rect 87466 28806 87518 28858
rect 4308 28576 4360 28628
rect 85820 28576 85872 28628
rect 8540 28440 8592 28492
rect 88212 28372 88264 28424
rect 5882 28262 5934 28314
rect 5946 28262 5998 28314
rect 6010 28262 6062 28314
rect 6074 28262 6126 28314
rect 6138 28262 6190 28314
rect 86474 28262 86526 28314
rect 86538 28262 86590 28314
rect 86602 28262 86654 28314
rect 86666 28262 86718 28314
rect 86730 28262 86782 28314
rect 6618 27718 6670 27770
rect 6682 27718 6734 27770
rect 6746 27718 6798 27770
rect 6810 27718 6862 27770
rect 6874 27718 6926 27770
rect 87210 27718 87262 27770
rect 87274 27718 87326 27770
rect 87338 27718 87390 27770
rect 87402 27718 87454 27770
rect 87466 27718 87518 27770
rect 5882 27174 5934 27226
rect 5946 27174 5998 27226
rect 6010 27174 6062 27226
rect 6074 27174 6126 27226
rect 6138 27174 6190 27226
rect 86474 27174 86526 27226
rect 86538 27174 86590 27226
rect 86602 27174 86654 27226
rect 86666 27174 86718 27226
rect 86730 27174 86782 27226
rect 8540 27012 8592 27064
rect 4308 26876 4360 26928
rect 85820 26876 85872 26928
rect 88396 26740 88448 26792
rect 6618 26630 6670 26682
rect 6682 26630 6734 26682
rect 6746 26630 6798 26682
rect 6810 26630 6862 26682
rect 6874 26630 6926 26682
rect 87210 26630 87262 26682
rect 87274 26630 87326 26682
rect 87338 26630 87390 26682
rect 87402 26630 87454 26682
rect 87466 26630 87518 26682
rect 4308 26400 4360 26452
rect 87568 26400 87620 26452
rect 8540 26264 8592 26316
rect 88212 26196 88264 26248
rect 5882 26086 5934 26138
rect 5946 26086 5998 26138
rect 6010 26086 6062 26138
rect 6074 26086 6126 26138
rect 6138 26086 6190 26138
rect 86474 26086 86526 26138
rect 86538 26086 86590 26138
rect 86602 26086 86654 26138
rect 86666 26086 86718 26138
rect 86730 26086 86782 26138
rect 6618 25542 6670 25594
rect 6682 25542 6734 25594
rect 6746 25542 6798 25594
rect 6810 25542 6862 25594
rect 6874 25542 6926 25594
rect 87210 25542 87262 25594
rect 87274 25542 87326 25594
rect 87338 25542 87390 25594
rect 87402 25542 87454 25594
rect 87466 25542 87518 25594
rect 4308 25312 4360 25364
rect 84808 25312 84860 25364
rect 5412 25108 5464 25160
rect 88580 25108 88632 25160
rect 5882 24998 5934 25050
rect 5946 24998 5998 25050
rect 6010 24998 6062 25050
rect 6074 24998 6126 25050
rect 6138 24998 6190 25050
rect 86474 24998 86526 25050
rect 86538 24998 86590 25050
rect 86602 24998 86654 25050
rect 86666 24998 86718 25050
rect 86730 24998 86782 25050
rect 6618 24454 6670 24506
rect 6682 24454 6734 24506
rect 6746 24454 6798 24506
rect 6810 24454 6862 24506
rect 6874 24454 6926 24506
rect 87210 24454 87262 24506
rect 87274 24454 87326 24506
rect 87338 24454 87390 24506
rect 87402 24454 87454 24506
rect 87466 24454 87518 24506
rect 4308 24224 4360 24276
rect 87568 24224 87620 24276
rect 8540 24088 8592 24140
rect 88488 24088 88540 24140
rect 5882 23910 5934 23962
rect 5946 23910 5998 23962
rect 6010 23910 6062 23962
rect 6074 23910 6126 23962
rect 6138 23910 6190 23962
rect 86474 23910 86526 23962
rect 86538 23910 86590 23962
rect 86602 23910 86654 23962
rect 86666 23910 86718 23962
rect 86730 23910 86782 23962
rect 6618 23366 6670 23418
rect 6682 23366 6734 23418
rect 6746 23366 6798 23418
rect 6810 23366 6862 23418
rect 6874 23366 6926 23418
rect 87210 23366 87262 23418
rect 87274 23366 87326 23418
rect 87338 23366 87390 23418
rect 87402 23366 87454 23418
rect 87466 23366 87518 23418
rect 4308 23136 4360 23188
rect 85820 23136 85872 23188
rect 8540 23000 8592 23052
rect 88212 22932 88264 22984
rect 5882 22822 5934 22874
rect 5946 22822 5998 22874
rect 6010 22822 6062 22874
rect 6074 22822 6126 22874
rect 6138 22822 6190 22874
rect 86474 22822 86526 22874
rect 86538 22822 86590 22874
rect 86602 22822 86654 22874
rect 86666 22822 86718 22874
rect 86730 22822 86782 22874
rect 6618 22278 6670 22330
rect 6682 22278 6734 22330
rect 6746 22278 6798 22330
rect 6810 22278 6862 22330
rect 6874 22278 6926 22330
rect 87210 22278 87262 22330
rect 87274 22278 87326 22330
rect 87338 22278 87390 22330
rect 87402 22278 87454 22330
rect 87466 22278 87518 22330
rect 5882 21734 5934 21786
rect 5946 21734 5998 21786
rect 6010 21734 6062 21786
rect 6074 21734 6126 21786
rect 6138 21734 6190 21786
rect 86474 21734 86526 21786
rect 86538 21734 86590 21786
rect 86602 21734 86654 21786
rect 86666 21734 86718 21786
rect 86730 21734 86782 21786
rect 8540 21572 8592 21624
rect 4308 21436 4360 21488
rect 85820 21436 85872 21488
rect 88396 21300 88448 21352
rect 6618 21190 6670 21242
rect 6682 21190 6734 21242
rect 6746 21190 6798 21242
rect 6810 21190 6862 21242
rect 6874 21190 6926 21242
rect 87210 21190 87262 21242
rect 87274 21190 87326 21242
rect 87338 21190 87390 21242
rect 87402 21190 87454 21242
rect 87466 21190 87518 21242
rect 5688 21028 5740 21080
rect 88580 21028 88632 21080
rect 4308 20960 4360 21012
rect 84808 20960 84860 21012
rect 5882 20646 5934 20698
rect 5946 20646 5998 20698
rect 6010 20646 6062 20698
rect 6074 20646 6126 20698
rect 6138 20646 6190 20698
rect 86474 20646 86526 20698
rect 86538 20646 86590 20698
rect 86602 20646 86654 20698
rect 86666 20646 86718 20698
rect 86730 20646 86782 20698
rect 6618 20102 6670 20154
rect 6682 20102 6734 20154
rect 6746 20102 6798 20154
rect 6810 20102 6862 20154
rect 6874 20102 6926 20154
rect 87210 20102 87262 20154
rect 87274 20102 87326 20154
rect 87338 20102 87390 20154
rect 87402 20102 87454 20154
rect 87466 20102 87518 20154
rect 4308 19872 4360 19924
rect 87568 19872 87620 19924
rect 8540 19736 8592 19788
rect 88672 19668 88724 19720
rect 5882 19558 5934 19610
rect 5946 19558 5998 19610
rect 6010 19558 6062 19610
rect 6074 19558 6126 19610
rect 6138 19558 6190 19610
rect 86474 19558 86526 19610
rect 86538 19558 86590 19610
rect 86602 19558 86654 19610
rect 86666 19558 86718 19610
rect 86730 19558 86782 19610
rect 6618 19014 6670 19066
rect 6682 19014 6734 19066
rect 6746 19014 6798 19066
rect 6810 19014 6862 19066
rect 6874 19014 6926 19066
rect 87210 19014 87262 19066
rect 87274 19014 87326 19066
rect 87338 19014 87390 19066
rect 87402 19014 87454 19066
rect 87466 19014 87518 19066
rect 4308 18784 4360 18836
rect 87292 18784 87344 18836
rect 8540 18648 8592 18700
rect 88212 18648 88264 18700
rect 5882 18470 5934 18522
rect 5946 18470 5998 18522
rect 6010 18470 6062 18522
rect 6074 18470 6126 18522
rect 6138 18470 6190 18522
rect 86474 18470 86526 18522
rect 86538 18470 86590 18522
rect 86602 18470 86654 18522
rect 86666 18470 86718 18522
rect 86730 18470 86782 18522
rect 6618 17926 6670 17978
rect 6682 17926 6734 17978
rect 6746 17926 6798 17978
rect 6810 17926 6862 17978
rect 6874 17926 6926 17978
rect 87210 17926 87262 17978
rect 87274 17926 87326 17978
rect 87338 17926 87390 17978
rect 87402 17926 87454 17978
rect 87466 17926 87518 17978
rect 4308 17696 4360 17748
rect 85820 17696 85872 17748
rect 8540 17560 8592 17612
rect 88212 17492 88264 17544
rect 5882 17382 5934 17434
rect 5946 17382 5998 17434
rect 6010 17382 6062 17434
rect 6074 17382 6126 17434
rect 6138 17382 6190 17434
rect 86474 17382 86526 17434
rect 86538 17382 86590 17434
rect 86602 17382 86654 17434
rect 86666 17382 86718 17434
rect 86730 17382 86782 17434
rect 6618 16838 6670 16890
rect 6682 16838 6734 16890
rect 6746 16838 6798 16890
rect 6810 16838 6862 16890
rect 6874 16838 6926 16890
rect 87210 16838 87262 16890
rect 87274 16838 87326 16890
rect 87338 16838 87390 16890
rect 87402 16838 87454 16890
rect 87466 16838 87518 16890
rect 5882 16294 5934 16346
rect 5946 16294 5998 16346
rect 6010 16294 6062 16346
rect 6074 16294 6126 16346
rect 6138 16294 6190 16346
rect 86474 16294 86526 16346
rect 86538 16294 86590 16346
rect 86602 16294 86654 16346
rect 86666 16294 86718 16346
rect 86730 16294 86782 16346
rect 8540 16132 8592 16184
rect 4308 15996 4360 16048
rect 85820 15996 85872 16048
rect 88212 15860 88264 15912
rect 6618 15750 6670 15802
rect 6682 15750 6734 15802
rect 6746 15750 6798 15802
rect 6810 15750 6862 15802
rect 6874 15750 6926 15802
rect 87210 15750 87262 15802
rect 87274 15750 87326 15802
rect 87338 15750 87390 15802
rect 87402 15750 87454 15802
rect 87466 15750 87518 15802
rect 5688 15588 5740 15640
rect 88580 15588 88632 15640
rect 4308 15520 4360 15572
rect 84808 15520 84860 15572
rect 5882 15206 5934 15258
rect 5946 15206 5998 15258
rect 6010 15206 6062 15258
rect 6074 15206 6126 15258
rect 6138 15206 6190 15258
rect 86474 15206 86526 15258
rect 86538 15206 86590 15258
rect 86602 15206 86654 15258
rect 86666 15206 86718 15258
rect 86730 15206 86782 15258
rect 85452 14976 85504 15028
rect 85636 14976 85688 15028
rect 88028 14815 88080 14824
rect 88028 14781 88037 14815
rect 88037 14781 88071 14815
rect 88071 14781 88080 14815
rect 88028 14772 88080 14781
rect 6618 14662 6670 14714
rect 6682 14662 6734 14714
rect 6746 14662 6798 14714
rect 6810 14662 6862 14714
rect 6874 14662 6926 14714
rect 87210 14662 87262 14714
rect 87274 14662 87326 14714
rect 87338 14662 87390 14714
rect 87402 14662 87454 14714
rect 87466 14662 87518 14714
rect 83428 14228 83480 14280
rect 85636 14271 85688 14280
rect 85636 14237 85645 14271
rect 85645 14237 85679 14271
rect 85679 14237 85688 14271
rect 85636 14228 85688 14237
rect 5882 14118 5934 14170
rect 5946 14118 5998 14170
rect 6010 14118 6062 14170
rect 6074 14118 6126 14170
rect 6138 14118 6190 14170
rect 86474 14118 86526 14170
rect 86538 14118 86590 14170
rect 86602 14118 86654 14170
rect 86666 14118 86718 14170
rect 86730 14118 86782 14170
rect 6618 13574 6670 13626
rect 6682 13574 6734 13626
rect 6746 13574 6798 13626
rect 6810 13574 6862 13626
rect 6874 13574 6926 13626
rect 87210 13574 87262 13626
rect 87274 13574 87326 13626
rect 87338 13574 87390 13626
rect 87402 13574 87454 13626
rect 87466 13574 87518 13626
rect 83612 13412 83664 13464
rect 85544 13412 85596 13464
rect 88212 13378 88264 13396
rect 88212 13344 88226 13378
rect 88226 13344 88260 13378
rect 88260 13344 88264 13378
rect 87936 13319 87988 13328
rect 87936 13285 87945 13319
rect 87945 13285 87979 13319
rect 87979 13285 87988 13319
rect 87936 13276 87988 13285
rect 5882 13030 5934 13082
rect 5946 13030 5998 13082
rect 6010 13030 6062 13082
rect 6074 13030 6126 13082
rect 6138 13030 6190 13082
rect 86474 13030 86526 13082
rect 86538 13030 86590 13082
rect 86602 13030 86654 13082
rect 86666 13030 86718 13082
rect 86730 13030 86782 13082
rect 87936 12868 87988 12920
rect 85360 12596 85412 12648
rect 87568 12664 87620 12716
rect 88580 12664 88632 12716
rect 6618 12486 6670 12538
rect 6682 12486 6734 12538
rect 6746 12486 6798 12538
rect 6810 12486 6862 12538
rect 6874 12486 6926 12538
rect 87210 12486 87262 12538
rect 87274 12486 87326 12538
rect 87338 12486 87390 12538
rect 87402 12486 87454 12538
rect 87466 12486 87518 12538
rect 83612 12324 83664 12376
rect 85360 12324 85412 12376
rect 87568 12324 87620 12376
rect 5882 11942 5934 11994
rect 5946 11942 5998 11994
rect 6010 11942 6062 11994
rect 6074 11942 6126 11994
rect 6138 11942 6190 11994
rect 86474 11942 86526 11994
rect 86538 11942 86590 11994
rect 86602 11942 86654 11994
rect 86666 11942 86718 11994
rect 86730 11942 86782 11994
rect 6618 11398 6670 11450
rect 6682 11398 6734 11450
rect 6746 11398 6798 11450
rect 6810 11398 6862 11450
rect 6874 11398 6926 11450
rect 87210 11398 87262 11450
rect 87274 11398 87326 11450
rect 87338 11398 87390 11450
rect 87402 11398 87454 11450
rect 87466 11398 87518 11450
rect 83244 11236 83296 11288
rect 5882 10854 5934 10906
rect 5946 10854 5998 10906
rect 6010 10854 6062 10906
rect 6074 10854 6126 10906
rect 6138 10854 6190 10906
rect 86474 10854 86526 10906
rect 86538 10854 86590 10906
rect 86602 10854 86654 10906
rect 86666 10854 86718 10906
rect 86730 10854 86782 10906
rect 88212 10599 88264 10608
rect 88212 10565 88221 10599
rect 88221 10565 88255 10599
rect 88255 10565 88264 10599
rect 88212 10556 88264 10565
rect 6618 10310 6670 10362
rect 6682 10310 6734 10362
rect 6746 10310 6798 10362
rect 6810 10310 6862 10362
rect 6874 10310 6926 10362
rect 87210 10310 87262 10362
rect 87274 10310 87326 10362
rect 87338 10310 87390 10362
rect 87402 10310 87454 10362
rect 87466 10310 87518 10362
rect 45708 10148 45760 10200
rect 46076 10148 46128 10200
rect 82508 10148 82560 10200
rect 5882 9766 5934 9818
rect 5946 9766 5998 9818
rect 6010 9766 6062 9818
rect 6074 9766 6126 9818
rect 6138 9766 6190 9818
rect 86474 9766 86526 9818
rect 86538 9766 86590 9818
rect 86602 9766 86654 9818
rect 86666 9766 86718 9818
rect 86730 9766 86782 9818
rect 6618 9222 6670 9274
rect 6682 9222 6734 9274
rect 6746 9222 6798 9274
rect 6810 9222 6862 9274
rect 6874 9222 6926 9274
rect 87210 9222 87262 9274
rect 87274 9222 87326 9274
rect 87338 9222 87390 9274
rect 87402 9222 87454 9274
rect 87466 9222 87518 9274
rect 5882 8678 5934 8730
rect 5946 8678 5998 8730
rect 6010 8678 6062 8730
rect 6074 8678 6126 8730
rect 6138 8678 6190 8730
rect 86474 8678 86526 8730
rect 86538 8678 86590 8730
rect 86602 8678 86654 8730
rect 86666 8678 86718 8730
rect 86730 8678 86782 8730
rect 6618 8134 6670 8186
rect 6682 8134 6734 8186
rect 6746 8134 6798 8186
rect 6810 8134 6862 8186
rect 6874 8134 6926 8186
rect 87210 8134 87262 8186
rect 87274 8134 87326 8186
rect 87338 8134 87390 8186
rect 87402 8134 87454 8186
rect 87466 8134 87518 8186
rect 5882 7590 5934 7642
rect 5946 7590 5998 7642
rect 6010 7590 6062 7642
rect 6074 7590 6126 7642
rect 6138 7590 6190 7642
rect 17722 7590 17774 7642
rect 17786 7590 17838 7642
rect 17850 7590 17902 7642
rect 17914 7590 17966 7642
rect 17978 7590 18030 7642
rect 36122 7590 36174 7642
rect 36186 7590 36238 7642
rect 36250 7590 36302 7642
rect 36314 7590 36366 7642
rect 36378 7590 36430 7642
rect 54522 7590 54574 7642
rect 54586 7590 54638 7642
rect 54650 7590 54702 7642
rect 54714 7590 54766 7642
rect 54778 7590 54830 7642
rect 72922 7590 72974 7642
rect 72986 7590 73038 7642
rect 73050 7590 73102 7642
rect 73114 7590 73166 7642
rect 73178 7590 73230 7642
rect 86474 7590 86526 7642
rect 86538 7590 86590 7642
rect 86602 7590 86654 7642
rect 86666 7590 86718 7642
rect 86730 7590 86782 7642
rect 45432 7471 45484 7480
rect 45432 7437 45441 7471
rect 45441 7437 45475 7471
rect 45475 7437 45484 7471
rect 45432 7428 45484 7437
rect 45708 7428 45760 7480
rect 45892 7428 45944 7480
rect 45984 7471 46036 7480
rect 45984 7437 45993 7471
rect 45993 7437 46027 7471
rect 46027 7437 46036 7471
rect 45984 7428 46036 7437
rect 83520 7292 83572 7344
rect 45984 7224 46036 7276
rect 83336 7224 83388 7276
rect 45708 7156 45760 7208
rect 83612 7156 83664 7208
rect 6618 7046 6670 7098
rect 6682 7046 6734 7098
rect 6746 7046 6798 7098
rect 6810 7046 6862 7098
rect 6874 7046 6926 7098
rect 18382 7046 18434 7098
rect 18446 7046 18498 7098
rect 18510 7046 18562 7098
rect 18574 7046 18626 7098
rect 18638 7046 18690 7098
rect 36782 7046 36834 7098
rect 36846 7046 36898 7098
rect 36910 7046 36962 7098
rect 36974 7046 37026 7098
rect 37038 7046 37090 7098
rect 55182 7046 55234 7098
rect 55246 7046 55298 7098
rect 55310 7046 55362 7098
rect 55374 7046 55426 7098
rect 55438 7046 55490 7098
rect 73582 7046 73634 7098
rect 73646 7046 73698 7098
rect 73710 7046 73762 7098
rect 73774 7046 73826 7098
rect 73838 7046 73890 7098
rect 87210 7046 87262 7098
rect 87274 7046 87326 7098
rect 87338 7046 87390 7098
rect 87402 7046 87454 7098
rect 87466 7046 87518 7098
rect 17722 6502 17774 6554
rect 17786 6502 17838 6554
rect 17850 6502 17902 6554
rect 17914 6502 17966 6554
rect 17978 6502 18030 6554
rect 36122 6502 36174 6554
rect 36186 6502 36238 6554
rect 36250 6502 36302 6554
rect 36314 6502 36366 6554
rect 36378 6502 36430 6554
rect 54522 6502 54574 6554
rect 54586 6502 54638 6554
rect 54650 6502 54702 6554
rect 54714 6502 54766 6554
rect 54778 6502 54830 6554
rect 72922 6502 72974 6554
rect 72986 6502 73038 6554
rect 73050 6502 73102 6554
rect 73114 6502 73166 6554
rect 73178 6502 73230 6554
rect 18382 5958 18434 6010
rect 18446 5958 18498 6010
rect 18510 5958 18562 6010
rect 18574 5958 18626 6010
rect 18638 5958 18690 6010
rect 36782 5958 36834 6010
rect 36846 5958 36898 6010
rect 36910 5958 36962 6010
rect 36974 5958 37026 6010
rect 37038 5958 37090 6010
rect 55182 5958 55234 6010
rect 55246 5958 55298 6010
rect 55310 5958 55362 6010
rect 55374 5958 55426 6010
rect 55438 5958 55490 6010
rect 73582 5958 73634 6010
rect 73646 5958 73698 6010
rect 73710 5958 73762 6010
rect 73774 5958 73826 6010
rect 73838 5958 73890 6010
rect 17722 5414 17774 5466
rect 17786 5414 17838 5466
rect 17850 5414 17902 5466
rect 17914 5414 17966 5466
rect 17978 5414 18030 5466
rect 36122 5414 36174 5466
rect 36186 5414 36238 5466
rect 36250 5414 36302 5466
rect 36314 5414 36366 5466
rect 36378 5414 36430 5466
rect 54522 5414 54574 5466
rect 54586 5414 54638 5466
rect 54650 5414 54702 5466
rect 54714 5414 54766 5466
rect 54778 5414 54830 5466
rect 72922 5414 72974 5466
rect 72986 5414 73038 5466
rect 73050 5414 73102 5466
rect 73114 5414 73166 5466
rect 73178 5414 73230 5466
rect 30436 5252 30488 5304
rect 31540 5252 31592 5304
rect 32644 5295 32696 5304
rect 32644 5261 32678 5295
rect 32678 5261 32696 5295
rect 32644 5252 32696 5261
rect 33748 5252 33800 5304
rect 34852 5252 34904 5304
rect 35956 5252 36008 5304
rect 37152 5295 37204 5304
rect 37152 5261 37186 5295
rect 37186 5261 37204 5295
rect 37152 5252 37204 5261
rect 38164 5252 38216 5304
rect 39268 5252 39320 5304
rect 40372 5295 40424 5304
rect 40372 5261 40406 5295
rect 40406 5261 40424 5295
rect 40372 5252 40424 5261
rect 41476 5252 41528 5304
rect 42580 5252 42632 5304
rect 43684 5252 43736 5304
rect 44788 5252 44840 5304
rect 68064 5295 68116 5304
rect 68064 5261 68097 5295
rect 68097 5261 68116 5295
rect 68064 5252 68116 5261
rect 68984 5252 69036 5304
rect 69996 5295 70048 5304
rect 69996 5261 70030 5295
rect 70030 5261 70048 5295
rect 69996 5252 70048 5261
rect 71284 5295 71336 5304
rect 71284 5261 71318 5295
rect 71318 5261 71336 5295
rect 71284 5252 71336 5261
rect 72572 5295 72624 5304
rect 72572 5261 72606 5295
rect 72606 5261 72624 5295
rect 72572 5252 72624 5261
rect 73400 5252 73452 5304
rect 74504 5295 74556 5304
rect 74504 5261 74538 5295
rect 74538 5261 74556 5295
rect 74504 5252 74556 5261
rect 75792 5295 75844 5304
rect 75792 5261 75826 5295
rect 75826 5261 75844 5295
rect 75792 5252 75844 5261
rect 76712 5252 76764 5304
rect 77724 5295 77776 5304
rect 77724 5261 77758 5295
rect 77758 5261 77776 5295
rect 77724 5252 77776 5261
rect 79012 5295 79064 5304
rect 79012 5261 79045 5295
rect 79045 5261 79064 5295
rect 79012 5252 79064 5261
rect 80116 5252 80168 5304
rect 81128 5252 81180 5304
rect 14980 5116 15032 5168
rect 16176 5159 16228 5168
rect 16176 5125 16185 5159
rect 16185 5125 16219 5159
rect 16219 5125 16228 5159
rect 16176 5116 16228 5125
rect 17188 5159 17240 5168
rect 17188 5125 17221 5159
rect 17221 5125 17240 5159
rect 17188 5116 17240 5125
rect 18292 5116 18344 5168
rect 19396 5159 19448 5168
rect 19396 5125 19405 5159
rect 19405 5125 19439 5159
rect 19439 5125 19448 5159
rect 19396 5116 19448 5125
rect 20500 5159 20552 5168
rect 20500 5125 20512 5159
rect 20512 5125 20552 5159
rect 20500 5116 20552 5125
rect 21604 5116 21656 5168
rect 22708 5116 22760 5168
rect 23904 5159 23956 5168
rect 23904 5125 23913 5159
rect 23913 5125 23947 5159
rect 23947 5125 23956 5159
rect 23904 5116 23956 5125
rect 24916 5159 24968 5168
rect 24916 5125 24949 5159
rect 24949 5125 24968 5159
rect 24916 5116 24968 5125
rect 26020 5116 26072 5168
rect 27124 5159 27176 5168
rect 27124 5125 27133 5159
rect 27133 5125 27167 5159
rect 27167 5125 27176 5159
rect 27124 5116 27176 5125
rect 28228 5159 28280 5168
rect 28228 5125 28240 5159
rect 28240 5125 28280 5159
rect 28228 5116 28280 5125
rect 29332 5116 29384 5168
rect 30712 5116 30764 5168
rect 31356 5159 31408 5168
rect 31356 5125 31393 5159
rect 31393 5125 31408 5159
rect 31356 5116 31408 5125
rect 32644 5116 32696 5168
rect 33932 5116 33984 5168
rect 34576 5159 34628 5168
rect 34576 5125 34613 5159
rect 34613 5125 34628 5159
rect 34576 5116 34628 5125
rect 35864 5116 35916 5168
rect 37152 5116 37204 5168
rect 38440 5116 38492 5168
rect 39084 5159 39136 5168
rect 39084 5125 39121 5159
rect 39121 5125 39136 5159
rect 39084 5116 39136 5125
rect 40372 5116 40424 5168
rect 41660 5116 41712 5168
rect 42304 5159 42356 5168
rect 42304 5125 42341 5159
rect 42341 5125 42356 5159
rect 42304 5116 42356 5125
rect 43592 5116 43644 5168
rect 44880 5116 44932 5168
rect 52608 5159 52660 5168
rect 52608 5125 52641 5159
rect 52641 5125 52660 5159
rect 52608 5116 52660 5125
rect 53528 5159 53580 5168
rect 53528 5125 53537 5159
rect 53537 5125 53571 5159
rect 53571 5125 53580 5159
rect 53528 5116 53580 5125
rect 54448 5116 54500 5168
rect 55828 5159 55880 5168
rect 55828 5125 55861 5159
rect 55861 5125 55880 5159
rect 55828 5116 55880 5125
rect 57024 5116 57076 5168
rect 58036 5159 58088 5168
rect 58036 5125 58045 5159
rect 58045 5125 58079 5159
rect 58079 5125 58088 5159
rect 58036 5116 58088 5125
rect 59048 5159 59100 5168
rect 59048 5125 59081 5159
rect 59081 5125 59100 5159
rect 59048 5116 59100 5125
rect 60336 5159 60388 5168
rect 60336 5125 60369 5159
rect 60369 5125 60388 5159
rect 60336 5116 60388 5125
rect 61256 5159 61308 5168
rect 61256 5125 61265 5159
rect 61265 5125 61299 5159
rect 61299 5125 61308 5159
rect 61256 5116 61308 5125
rect 62360 5159 62412 5168
rect 62360 5125 62372 5159
rect 62372 5125 62412 5159
rect 62360 5116 62412 5125
rect 63556 5159 63608 5168
rect 63556 5125 63589 5159
rect 63589 5125 63608 5159
rect 63556 5116 63608 5125
rect 64752 5116 64804 5168
rect 65764 5159 65816 5168
rect 65764 5125 65773 5159
rect 65773 5125 65807 5159
rect 65807 5125 65816 5159
rect 65764 5116 65816 5125
rect 66776 5159 66828 5168
rect 66776 5125 66809 5159
rect 66809 5125 66828 5159
rect 66776 5116 66828 5125
rect 68064 5116 68116 5168
rect 68708 5159 68760 5168
rect 68708 5125 68745 5159
rect 68745 5125 68760 5159
rect 68708 5116 68760 5125
rect 69996 5116 70048 5168
rect 71284 5116 71336 5168
rect 72572 5116 72624 5168
rect 73216 5159 73268 5168
rect 73216 5125 73253 5159
rect 73253 5125 73268 5159
rect 73216 5116 73268 5125
rect 74504 5116 74556 5168
rect 75792 5116 75844 5168
rect 76436 5159 76488 5168
rect 76436 5125 76473 5159
rect 76473 5125 76488 5159
rect 76436 5116 76488 5125
rect 77724 5116 77776 5168
rect 79012 5116 79064 5168
rect 80300 5116 80352 5168
rect 80944 5159 80996 5168
rect 80944 5125 80981 5159
rect 80981 5125 80996 5159
rect 80944 5116 80996 5125
rect 15256 4980 15308 5032
rect 15900 4980 15952 5032
rect 17188 4980 17240 5032
rect 18752 4980 18804 5032
rect 19120 4980 19172 5032
rect 20408 4980 20460 5032
rect 21696 4980 21748 5032
rect 22984 4980 23036 5032
rect 23628 4980 23680 5032
rect 24916 4980 24968 5032
rect 26204 4980 26256 5032
rect 26848 4980 26900 5032
rect 28136 4980 28188 5032
rect 29424 4980 29476 5032
rect 52608 4980 52660 5032
rect 53252 4980 53304 5032
rect 54540 4980 54592 5032
rect 55828 4980 55880 5032
rect 57116 4980 57168 5032
rect 57760 4980 57812 5032
rect 59048 4980 59100 5032
rect 60336 4980 60388 5032
rect 60980 4980 61032 5032
rect 62268 4980 62320 5032
rect 63556 4980 63608 5032
rect 64844 4980 64896 5032
rect 65488 4980 65540 5032
rect 66776 4980 66828 5032
rect 18382 4870 18434 4922
rect 18446 4870 18498 4922
rect 18510 4870 18562 4922
rect 18574 4870 18626 4922
rect 18638 4870 18690 4922
rect 36782 4870 36834 4922
rect 36846 4870 36898 4922
rect 36910 4870 36962 4922
rect 36974 4870 37026 4922
rect 37038 4870 37090 4922
rect 55182 4870 55234 4922
rect 55246 4870 55298 4922
rect 55310 4870 55362 4922
rect 55374 4870 55426 4922
rect 55438 4870 55490 4922
rect 73582 4870 73634 4922
rect 73646 4870 73698 4922
rect 73710 4870 73762 4922
rect 73774 4870 73826 4922
rect 73838 4870 73890 4922
<< metal2 >>
rect 15254 88000 15310 88800
rect 15898 88000 15954 88800
rect 17186 88000 17242 88800
rect 18474 88000 18530 88800
rect 18580 88054 18792 88082
rect 15268 87386 15296 88000
rect 15912 87386 15940 88000
rect 17200 87386 17228 88000
rect 18488 87946 18516 88000
rect 18580 87946 18608 88054
rect 18488 87918 18608 87946
rect 18382 87612 18690 87621
rect 18382 87610 18388 87612
rect 18444 87610 18468 87612
rect 18524 87610 18548 87612
rect 18604 87610 18628 87612
rect 18684 87610 18690 87612
rect 18444 87558 18446 87610
rect 18626 87558 18628 87610
rect 18382 87556 18388 87558
rect 18444 87556 18468 87558
rect 18524 87556 18548 87558
rect 18604 87556 18628 87558
rect 18684 87556 18690 87558
rect 18382 87547 18690 87556
rect 18764 87386 18792 88054
rect 19118 88000 19174 88800
rect 20406 88000 20462 88800
rect 21694 88000 21750 88800
rect 22982 88000 23038 88800
rect 23626 88000 23682 88800
rect 24914 88000 24970 88800
rect 26202 88000 26258 88800
rect 26846 88000 26902 88800
rect 28134 88000 28190 88800
rect 29422 88000 29478 88800
rect 30710 88000 30766 88800
rect 31354 88000 31410 88800
rect 32642 88000 32698 88800
rect 33930 88000 33986 88800
rect 34574 88000 34630 88800
rect 35862 88000 35918 88800
rect 36506 88000 36562 88800
rect 37150 88000 37206 88800
rect 37794 88000 37850 88800
rect 38438 88000 38494 88800
rect 39082 88000 39138 88800
rect 39726 88000 39782 88800
rect 40370 88000 40426 88800
rect 41014 88000 41070 88800
rect 41658 88000 41714 88800
rect 42302 88000 42358 88800
rect 42946 88000 43002 88800
rect 43590 88000 43646 88800
rect 44234 88000 44290 88800
rect 44878 88000 44934 88800
rect 45522 88000 45578 88800
rect 46166 88000 46222 88800
rect 46810 88000 46866 88800
rect 47454 88000 47510 88800
rect 48098 88000 48154 88800
rect 48742 88000 48798 88800
rect 49386 88000 49442 88800
rect 50030 88000 50086 88800
rect 52606 88000 52662 88800
rect 53250 88000 53306 88800
rect 54538 88000 54594 88800
rect 55826 88000 55882 88800
rect 57114 88000 57170 88800
rect 57758 88000 57814 88800
rect 59046 88000 59102 88800
rect 60334 88000 60390 88800
rect 60978 88000 61034 88800
rect 62266 88000 62322 88800
rect 63554 88000 63610 88800
rect 64842 88000 64898 88800
rect 65486 88000 65542 88800
rect 66774 88000 66830 88800
rect 68062 88000 68118 88800
rect 68706 88000 68762 88800
rect 69994 88000 70050 88800
rect 71282 88000 71338 88800
rect 72570 88000 72626 88800
rect 73214 88000 73270 88800
rect 74502 88000 74558 88800
rect 75790 88000 75846 88800
rect 76434 88000 76490 88800
rect 77722 88000 77778 88800
rect 79010 88000 79066 88800
rect 80298 88000 80354 88800
rect 80942 88000 80998 88800
rect 82230 88000 82286 88800
rect 19132 87386 19160 88000
rect 20420 87386 20448 88000
rect 21708 87386 21736 88000
rect 22996 87386 23024 88000
rect 23640 87386 23668 88000
rect 24928 87386 24956 88000
rect 26216 87386 26244 88000
rect 26860 87386 26888 88000
rect 28148 87386 28176 88000
rect 29436 87386 29464 88000
rect 15256 87380 15308 87386
rect 15256 87322 15308 87328
rect 15900 87380 15952 87386
rect 15900 87322 15952 87328
rect 17188 87380 17240 87386
rect 17188 87322 17240 87328
rect 18752 87380 18804 87386
rect 18752 87322 18804 87328
rect 19120 87380 19172 87386
rect 19120 87322 19172 87328
rect 20408 87380 20460 87386
rect 20408 87322 20460 87328
rect 21696 87380 21748 87386
rect 21696 87322 21748 87328
rect 22984 87380 23036 87386
rect 22984 87322 23036 87328
rect 23628 87380 23680 87386
rect 23628 87322 23680 87328
rect 24916 87380 24968 87386
rect 24916 87322 24968 87328
rect 26204 87380 26256 87386
rect 26204 87322 26256 87328
rect 26848 87380 26900 87386
rect 26848 87322 26900 87328
rect 28136 87380 28188 87386
rect 28136 87322 28188 87328
rect 29424 87380 29476 87386
rect 29424 87322 29476 87328
rect 30620 87380 30672 87386
rect 30620 87322 30672 87328
rect 15532 87244 15584 87250
rect 15532 87186 15584 87192
rect 16084 87244 16136 87250
rect 16084 87186 16136 87192
rect 17188 87244 17240 87250
rect 17188 87186 17240 87192
rect 18292 87244 18344 87250
rect 18292 87186 18344 87192
rect 19396 87244 19448 87250
rect 19396 87186 19448 87192
rect 20408 87244 20460 87250
rect 21604 87244 21656 87250
rect 20460 87192 20540 87194
rect 20408 87186 20540 87192
rect 21604 87186 21656 87192
rect 22708 87244 22760 87250
rect 22708 87186 22760 87192
rect 23812 87244 23864 87250
rect 23812 87186 23864 87192
rect 24916 87244 24968 87250
rect 24916 87186 24968 87192
rect 26020 87244 26072 87250
rect 26020 87186 26072 87192
rect 27124 87244 27176 87250
rect 27124 87186 27176 87192
rect 28136 87244 28188 87250
rect 29332 87244 29384 87250
rect 28188 87192 28268 87194
rect 28136 87186 28268 87192
rect 29332 87186 29384 87192
rect 5882 84892 6190 84901
rect 5882 84890 5888 84892
rect 5944 84890 5968 84892
rect 6024 84890 6048 84892
rect 6104 84890 6128 84892
rect 6184 84890 6190 84892
rect 5944 84838 5946 84890
rect 6126 84838 6128 84890
rect 5882 84836 5888 84838
rect 5944 84836 5968 84838
rect 6024 84836 6048 84838
rect 6104 84836 6128 84838
rect 6184 84836 6190 84838
rect 5882 84827 6190 84836
rect 12772 84660 12824 84666
rect 12772 84602 12824 84608
rect 11668 84592 11720 84598
rect 11668 84534 11720 84540
rect 7528 84524 7580 84530
rect 7528 84466 7580 84472
rect 6618 84348 6926 84357
rect 6618 84346 6624 84348
rect 6680 84346 6704 84348
rect 6760 84346 6784 84348
rect 6840 84346 6864 84348
rect 6920 84346 6926 84348
rect 6680 84294 6682 84346
rect 6862 84294 6864 84346
rect 6618 84292 6624 84294
rect 6680 84292 6704 84294
rect 6760 84292 6784 84294
rect 6840 84292 6864 84294
rect 6920 84292 6926 84294
rect 6618 84283 6926 84292
rect 5882 83804 6190 83813
rect 5882 83802 5888 83804
rect 5944 83802 5968 83804
rect 6024 83802 6048 83804
rect 6104 83802 6128 83804
rect 6184 83802 6190 83804
rect 5944 83750 5946 83802
rect 6126 83750 6128 83802
rect 5882 83748 5888 83750
rect 5944 83748 5968 83750
rect 6024 83748 6048 83750
rect 6104 83748 6128 83750
rect 6184 83748 6190 83750
rect 5882 83739 6190 83748
rect 6618 83260 6926 83269
rect 6618 83258 6624 83260
rect 6680 83258 6704 83260
rect 6760 83258 6784 83260
rect 6840 83258 6864 83260
rect 6920 83258 6926 83260
rect 6680 83206 6682 83258
rect 6862 83206 6864 83258
rect 6618 83204 6624 83206
rect 6680 83204 6704 83206
rect 6760 83204 6784 83206
rect 6840 83204 6864 83206
rect 6920 83204 6926 83206
rect 6618 83195 6926 83204
rect 5882 82716 6190 82725
rect 5882 82714 5888 82716
rect 5944 82714 5968 82716
rect 6024 82714 6048 82716
rect 6104 82714 6128 82716
rect 6184 82714 6190 82716
rect 5944 82662 5946 82714
rect 6126 82662 6128 82714
rect 5882 82660 5888 82662
rect 5944 82660 5968 82662
rect 6024 82660 6048 82662
rect 6104 82660 6128 82662
rect 6184 82660 6190 82662
rect 5882 82651 6190 82660
rect 6618 82172 6926 82181
rect 6618 82170 6624 82172
rect 6680 82170 6704 82172
rect 6760 82170 6784 82172
rect 6840 82170 6864 82172
rect 6920 82170 6926 82172
rect 6680 82118 6682 82170
rect 6862 82118 6864 82170
rect 6618 82116 6624 82118
rect 6680 82116 6704 82118
rect 6760 82116 6784 82118
rect 6840 82116 6864 82118
rect 6920 82116 6926 82118
rect 6618 82107 6926 82116
rect 5882 81628 6190 81637
rect 5882 81626 5888 81628
rect 5944 81626 5968 81628
rect 6024 81626 6048 81628
rect 6104 81626 6128 81628
rect 6184 81626 6190 81628
rect 5944 81574 5946 81626
rect 6126 81574 6128 81626
rect 5882 81572 5888 81574
rect 5944 81572 5968 81574
rect 6024 81572 6048 81574
rect 6104 81572 6128 81574
rect 6184 81572 6190 81574
rect 5882 81563 6190 81572
rect 4124 81328 4176 81334
rect 4122 81296 4124 81305
rect 4176 81296 4178 81305
rect 4122 81231 4178 81240
rect 6618 81084 6926 81093
rect 6618 81082 6624 81084
rect 6680 81082 6704 81084
rect 6760 81082 6784 81084
rect 6840 81082 6864 81084
rect 6920 81082 6926 81084
rect 6680 81030 6682 81082
rect 6862 81030 6864 81082
rect 6618 81028 6624 81030
rect 6680 81028 6704 81030
rect 6760 81028 6784 81030
rect 6840 81028 6864 81030
rect 6920 81028 6926 81030
rect 6618 81019 6926 81028
rect 5882 80540 6190 80549
rect 5882 80538 5888 80540
rect 5944 80538 5968 80540
rect 6024 80538 6048 80540
rect 6104 80538 6128 80540
rect 6184 80538 6190 80540
rect 5944 80486 5946 80538
rect 6126 80486 6128 80538
rect 5882 80484 5888 80486
rect 5944 80484 5968 80486
rect 6024 80484 6048 80486
rect 6104 80484 6128 80486
rect 6184 80484 6190 80486
rect 5882 80475 6190 80484
rect 4124 80104 4176 80110
rect 4124 80046 4176 80052
rect 4136 79945 4164 80046
rect 6618 79996 6926 80005
rect 6618 79994 6624 79996
rect 6680 79994 6704 79996
rect 6760 79994 6784 79996
rect 6840 79994 6864 79996
rect 6920 79994 6926 79996
rect 4122 79936 4178 79945
rect 6680 79942 6682 79994
rect 6862 79942 6864 79994
rect 6618 79940 6624 79942
rect 6680 79940 6704 79942
rect 6760 79940 6784 79942
rect 6840 79940 6864 79942
rect 6920 79940 6926 79942
rect 6618 79931 6926 79940
rect 4122 79871 4178 79880
rect 5882 79452 6190 79461
rect 5882 79450 5888 79452
rect 5944 79450 5968 79452
rect 6024 79450 6048 79452
rect 6104 79450 6128 79452
rect 6184 79450 6190 79452
rect 5944 79398 5946 79450
rect 6126 79398 6128 79450
rect 5882 79396 5888 79398
rect 5944 79396 5968 79398
rect 6024 79396 6048 79398
rect 6104 79396 6128 79398
rect 6184 79396 6190 79398
rect 5882 79387 6190 79396
rect 6618 78908 6926 78917
rect 6618 78906 6624 78908
rect 6680 78906 6704 78908
rect 6760 78906 6784 78908
rect 6840 78906 6864 78908
rect 6920 78906 6926 78908
rect 6680 78854 6682 78906
rect 6862 78854 6864 78906
rect 6618 78852 6624 78854
rect 6680 78852 6704 78854
rect 6760 78852 6784 78854
rect 6840 78852 6864 78854
rect 6920 78852 6926 78854
rect 6618 78843 6926 78852
rect 4122 78576 4178 78585
rect 4122 78511 4124 78520
rect 4176 78511 4178 78520
rect 4124 78482 4176 78488
rect 5882 78364 6190 78373
rect 5882 78362 5888 78364
rect 5944 78362 5968 78364
rect 6024 78362 6048 78364
rect 6104 78362 6128 78364
rect 6184 78362 6190 78364
rect 5944 78310 5946 78362
rect 6126 78310 6128 78362
rect 5882 78308 5888 78310
rect 5944 78308 5968 78310
rect 6024 78308 6048 78310
rect 6104 78308 6128 78310
rect 6184 78308 6190 78310
rect 5882 78299 6190 78308
rect 4124 77928 4176 77934
rect 4122 77896 4124 77905
rect 4176 77896 4178 77905
rect 4122 77831 4178 77840
rect 6618 77820 6926 77829
rect 6618 77818 6624 77820
rect 6680 77818 6704 77820
rect 6760 77818 6784 77820
rect 6840 77818 6864 77820
rect 6920 77818 6926 77820
rect 6680 77766 6682 77818
rect 6862 77766 6864 77818
rect 6618 77764 6624 77766
rect 6680 77764 6704 77766
rect 6760 77764 6784 77766
rect 6840 77764 6864 77766
rect 6920 77764 6926 77766
rect 6618 77755 6926 77764
rect 5882 77276 6190 77285
rect 5882 77274 5888 77276
rect 5944 77274 5968 77276
rect 6024 77274 6048 77276
rect 6104 77274 6128 77276
rect 6184 77274 6190 77276
rect 5944 77222 5946 77274
rect 6126 77222 6128 77274
rect 5882 77220 5888 77222
rect 5944 77220 5968 77222
rect 6024 77220 6048 77222
rect 6104 77220 6128 77222
rect 6184 77220 6190 77222
rect 5882 77211 6190 77220
rect 4216 76840 4268 76846
rect 4216 76782 4268 76788
rect 4228 76545 4256 76782
rect 6618 76732 6926 76741
rect 6618 76730 6624 76732
rect 6680 76730 6704 76732
rect 6760 76730 6784 76732
rect 6840 76730 6864 76732
rect 6920 76730 6926 76732
rect 6680 76678 6682 76730
rect 6862 76678 6864 76730
rect 6618 76676 6624 76678
rect 6680 76676 6704 76678
rect 6760 76676 6784 76678
rect 6840 76676 6864 76678
rect 6920 76676 6926 76678
rect 6618 76667 6926 76676
rect 4214 76536 4270 76545
rect 4214 76471 4270 76480
rect 5882 76188 6190 76197
rect 5882 76186 5888 76188
rect 5944 76186 5968 76188
rect 6024 76186 6048 76188
rect 6104 76186 6128 76188
rect 6184 76186 6190 76188
rect 5944 76134 5946 76186
rect 6126 76134 6128 76186
rect 5882 76132 5888 76134
rect 5944 76132 5968 76134
rect 6024 76132 6048 76134
rect 6104 76132 6128 76134
rect 6184 76132 6190 76134
rect 5882 76123 6190 76132
rect 4122 75856 4178 75865
rect 4122 75791 4124 75800
rect 4176 75791 4178 75800
rect 4124 75762 4176 75768
rect 6618 75644 6926 75653
rect 6618 75642 6624 75644
rect 6680 75642 6704 75644
rect 6760 75642 6784 75644
rect 6840 75642 6864 75644
rect 6920 75642 6926 75644
rect 6680 75590 6682 75642
rect 6862 75590 6864 75642
rect 6618 75588 6624 75590
rect 6680 75588 6704 75590
rect 6760 75588 6784 75590
rect 6840 75588 6864 75590
rect 6920 75588 6926 75590
rect 6618 75579 6926 75588
rect 5882 75100 6190 75109
rect 5882 75098 5888 75100
rect 5944 75098 5968 75100
rect 6024 75098 6048 75100
rect 6104 75098 6128 75100
rect 6184 75098 6190 75100
rect 5944 75046 5946 75098
rect 6126 75046 6128 75098
rect 5882 75044 5888 75046
rect 5944 75044 5968 75046
rect 6024 75044 6048 75046
rect 6104 75044 6128 75046
rect 6184 75044 6190 75046
rect 5882 75035 6190 75044
rect 4124 74800 4176 74806
rect 5412 74800 5464 74806
rect 4124 74742 4176 74748
rect 5410 74768 5412 74777
rect 5464 74768 5466 74777
rect 4136 74505 4164 74742
rect 5410 74703 5466 74712
rect 6618 74556 6926 74565
rect 6618 74554 6624 74556
rect 6680 74554 6704 74556
rect 6760 74554 6784 74556
rect 6840 74554 6864 74556
rect 6920 74554 6926 74556
rect 4122 74496 4178 74505
rect 6680 74502 6682 74554
rect 6862 74502 6864 74554
rect 6618 74500 6624 74502
rect 6680 74500 6704 74502
rect 6760 74500 6784 74502
rect 6840 74500 6864 74502
rect 6920 74500 6926 74502
rect 6618 74491 6926 74500
rect 4122 74431 4178 74440
rect 5882 74012 6190 74021
rect 5882 74010 5888 74012
rect 5944 74010 5968 74012
rect 6024 74010 6048 74012
rect 6104 74010 6128 74012
rect 6184 74010 6190 74012
rect 5944 73958 5946 74010
rect 6126 73958 6128 74010
rect 5882 73956 5888 73958
rect 5944 73956 5968 73958
rect 6024 73956 6048 73958
rect 6104 73956 6128 73958
rect 6184 73956 6190 73958
rect 5882 73947 6190 73956
rect 5410 73680 5466 73689
rect 5410 73615 5466 73624
rect 5424 73242 5452 73615
rect 6618 73468 6926 73477
rect 6618 73466 6624 73468
rect 6680 73466 6704 73468
rect 6760 73466 6784 73468
rect 6840 73466 6864 73468
rect 6920 73466 6926 73468
rect 6680 73414 6682 73466
rect 6862 73414 6864 73466
rect 6618 73412 6624 73414
rect 6680 73412 6704 73414
rect 6760 73412 6784 73414
rect 6840 73412 6864 73414
rect 6920 73412 6926 73414
rect 6618 73403 6926 73412
rect 5412 73236 5464 73242
rect 5412 73178 5464 73184
rect 4122 73136 4178 73145
rect 4122 73071 4124 73080
rect 4176 73071 4178 73080
rect 4124 73042 4176 73048
rect 5882 72924 6190 72933
rect 5882 72922 5888 72924
rect 5944 72922 5968 72924
rect 6024 72922 6048 72924
rect 6104 72922 6128 72924
rect 6184 72922 6190 72924
rect 5944 72870 5946 72922
rect 6126 72870 6128 72922
rect 5882 72868 5888 72870
rect 5944 72868 5968 72870
rect 6024 72868 6048 72870
rect 6104 72868 6128 72870
rect 6184 72868 6190 72870
rect 5882 72859 6190 72868
rect 4124 72488 4176 72494
rect 4122 72456 4124 72465
rect 4176 72456 4178 72465
rect 4122 72391 4178 72400
rect 6618 72380 6926 72389
rect 6618 72378 6624 72380
rect 6680 72378 6704 72380
rect 6760 72378 6784 72380
rect 6840 72378 6864 72380
rect 6920 72378 6926 72380
rect 6680 72326 6682 72378
rect 6862 72326 6864 72378
rect 6618 72324 6624 72326
rect 6680 72324 6704 72326
rect 6760 72324 6784 72326
rect 6840 72324 6864 72326
rect 6920 72324 6926 72326
rect 6618 72315 6926 72324
rect 5882 71836 6190 71845
rect 5882 71834 5888 71836
rect 5944 71834 5968 71836
rect 6024 71834 6048 71836
rect 6104 71834 6128 71836
rect 6184 71834 6190 71836
rect 5944 71782 5946 71834
rect 6126 71782 6128 71834
rect 5882 71780 5888 71782
rect 5944 71780 5968 71782
rect 6024 71780 6048 71782
rect 6104 71780 6128 71782
rect 6184 71780 6190 71782
rect 5882 71771 6190 71780
rect 4216 71400 4268 71406
rect 4216 71342 4268 71348
rect 4228 71105 4256 71342
rect 6618 71292 6926 71301
rect 6618 71290 6624 71292
rect 6680 71290 6704 71292
rect 6760 71290 6784 71292
rect 6840 71290 6864 71292
rect 6920 71290 6926 71292
rect 6680 71238 6682 71290
rect 6862 71238 6864 71290
rect 6618 71236 6624 71238
rect 6680 71236 6704 71238
rect 6760 71236 6784 71238
rect 6840 71236 6864 71238
rect 6920 71236 6926 71238
rect 6618 71227 6926 71236
rect 4214 71096 4270 71105
rect 4214 71031 4270 71040
rect 5882 70748 6190 70757
rect 5882 70746 5888 70748
rect 5944 70746 5968 70748
rect 6024 70746 6048 70748
rect 6104 70746 6128 70748
rect 6184 70746 6190 70748
rect 5944 70694 5946 70746
rect 6126 70694 6128 70746
rect 5882 70692 5888 70694
rect 5944 70692 5968 70694
rect 6024 70692 6048 70694
rect 6104 70692 6128 70694
rect 6184 70692 6190 70694
rect 5882 70683 6190 70692
rect 4122 70416 4178 70425
rect 4122 70351 4124 70360
rect 4176 70351 4178 70360
rect 4124 70322 4176 70328
rect 6618 70204 6926 70213
rect 6618 70202 6624 70204
rect 6680 70202 6704 70204
rect 6760 70202 6784 70204
rect 6840 70202 6864 70204
rect 6920 70202 6926 70204
rect 6680 70150 6682 70202
rect 6862 70150 6864 70202
rect 6618 70148 6624 70150
rect 6680 70148 6704 70150
rect 6760 70148 6784 70150
rect 6840 70148 6864 70150
rect 6920 70148 6926 70150
rect 6618 70139 6926 70148
rect 5882 69660 6190 69669
rect 5882 69658 5888 69660
rect 5944 69658 5968 69660
rect 6024 69658 6048 69660
rect 6104 69658 6128 69660
rect 6184 69658 6190 69660
rect 5944 69606 5946 69658
rect 6126 69606 6128 69658
rect 5882 69604 5888 69606
rect 5944 69604 5968 69606
rect 6024 69604 6048 69606
rect 6104 69604 6128 69606
rect 6184 69604 6190 69606
rect 5882 69595 6190 69604
rect 5412 69360 5464 69366
rect 5412 69302 5464 69308
rect 4124 69292 4176 69298
rect 4124 69234 4176 69240
rect 4136 69065 4164 69234
rect 4122 69056 4178 69065
rect 4122 68991 4178 69000
rect 5424 68929 5452 69302
rect 6618 69116 6926 69125
rect 6618 69114 6624 69116
rect 6680 69114 6704 69116
rect 6760 69114 6784 69116
rect 6840 69114 6864 69116
rect 6920 69114 6926 69116
rect 6680 69062 6682 69114
rect 6862 69062 6864 69114
rect 6618 69060 6624 69062
rect 6680 69060 6704 69062
rect 6760 69060 6784 69062
rect 6840 69060 6864 69062
rect 6920 69060 6926 69062
rect 6618 69051 6926 69060
rect 5410 68920 5466 68929
rect 5410 68855 5466 68864
rect 5882 68572 6190 68581
rect 5882 68570 5888 68572
rect 5944 68570 5968 68572
rect 6024 68570 6048 68572
rect 6104 68570 6128 68572
rect 6184 68570 6190 68572
rect 5944 68518 5946 68570
rect 6126 68518 6128 68570
rect 5882 68516 5888 68518
rect 5944 68516 5968 68518
rect 6024 68516 6048 68518
rect 6104 68516 6128 68518
rect 6184 68516 6190 68518
rect 5882 68507 6190 68516
rect 5410 68240 5466 68249
rect 5410 68175 5466 68184
rect 5424 67802 5452 68175
rect 6618 68028 6926 68037
rect 6618 68026 6624 68028
rect 6680 68026 6704 68028
rect 6760 68026 6784 68028
rect 6840 68026 6864 68028
rect 6920 68026 6926 68028
rect 6680 67974 6682 68026
rect 6862 67974 6864 68026
rect 6618 67972 6624 67974
rect 6680 67972 6704 67974
rect 6760 67972 6784 67974
rect 6840 67972 6864 67974
rect 6920 67972 6926 67974
rect 6618 67963 6926 67972
rect 5412 67796 5464 67802
rect 5412 67738 5464 67744
rect 4030 67696 4086 67705
rect 4030 67631 4032 67640
rect 4084 67631 4086 67640
rect 4032 67602 4084 67608
rect 5882 67484 6190 67493
rect 5882 67482 5888 67484
rect 5944 67482 5968 67484
rect 6024 67482 6048 67484
rect 6104 67482 6128 67484
rect 6184 67482 6190 67484
rect 5944 67430 5946 67482
rect 6126 67430 6128 67482
rect 5882 67428 5888 67430
rect 5944 67428 5968 67430
rect 6024 67428 6048 67430
rect 6104 67428 6128 67430
rect 6184 67428 6190 67430
rect 5882 67419 6190 67428
rect 4124 67048 4176 67054
rect 4122 67016 4124 67025
rect 4176 67016 4178 67025
rect 4122 66951 4178 66960
rect 6618 66940 6926 66949
rect 6618 66938 6624 66940
rect 6680 66938 6704 66940
rect 6760 66938 6784 66940
rect 6840 66938 6864 66940
rect 6920 66938 6926 66940
rect 6680 66886 6682 66938
rect 6862 66886 6864 66938
rect 6618 66884 6624 66886
rect 6680 66884 6704 66886
rect 6760 66884 6784 66886
rect 6840 66884 6864 66886
rect 6920 66884 6926 66886
rect 6618 66875 6926 66884
rect 5882 66396 6190 66405
rect 5882 66394 5888 66396
rect 5944 66394 5968 66396
rect 6024 66394 6048 66396
rect 6104 66394 6128 66396
rect 6184 66394 6190 66396
rect 5944 66342 5946 66394
rect 6126 66342 6128 66394
rect 5882 66340 5888 66342
rect 5944 66340 5968 66342
rect 6024 66340 6048 66342
rect 6104 66340 6128 66342
rect 6184 66340 6190 66342
rect 5882 66331 6190 66340
rect 4308 66096 4360 66102
rect 4308 66038 4360 66044
rect 4320 65665 4348 66038
rect 6618 65852 6926 65861
rect 6618 65850 6624 65852
rect 6680 65850 6704 65852
rect 6760 65850 6784 65852
rect 6840 65850 6864 65852
rect 6920 65850 6926 65852
rect 6680 65798 6682 65850
rect 6862 65798 6864 65850
rect 6618 65796 6624 65798
rect 6680 65796 6704 65798
rect 6760 65796 6784 65798
rect 6840 65796 6864 65798
rect 6920 65796 6926 65798
rect 6618 65787 6926 65796
rect 4306 65656 4362 65665
rect 4306 65591 4362 65600
rect 5882 65308 6190 65317
rect 5882 65306 5888 65308
rect 5944 65306 5968 65308
rect 6024 65306 6048 65308
rect 6104 65306 6128 65308
rect 6184 65306 6190 65308
rect 5944 65254 5946 65306
rect 6126 65254 6128 65306
rect 5882 65252 5888 65254
rect 5944 65252 5968 65254
rect 6024 65252 6048 65254
rect 6104 65252 6128 65254
rect 6184 65252 6190 65254
rect 5882 65243 6190 65252
rect 4308 65008 4360 65014
rect 4306 64976 4308 64985
rect 4360 64976 4362 64985
rect 4306 64911 4362 64920
rect 6618 64764 6926 64773
rect 6618 64762 6624 64764
rect 6680 64762 6704 64764
rect 6760 64762 6784 64764
rect 6840 64762 6864 64764
rect 6920 64762 6926 64764
rect 6680 64710 6682 64762
rect 6862 64710 6864 64762
rect 6618 64708 6624 64710
rect 6680 64708 6704 64710
rect 6760 64708 6784 64710
rect 6840 64708 6864 64710
rect 6920 64708 6926 64710
rect 6618 64699 6926 64708
rect 7540 64606 7568 84466
rect 10564 84456 10616 84462
rect 10564 84398 10616 84404
rect 9828 83096 9880 83102
rect 9828 83038 9880 83044
rect 7620 82416 7672 82422
rect 7620 82358 7672 82364
rect 7528 64600 7580 64606
rect 7528 64542 7580 64548
rect 5882 64220 6190 64229
rect 5882 64218 5888 64220
rect 5944 64218 5968 64220
rect 6024 64218 6048 64220
rect 6104 64218 6128 64220
rect 6184 64218 6190 64220
rect 5944 64166 5946 64218
rect 6126 64166 6128 64218
rect 5882 64164 5888 64166
rect 5944 64164 5968 64166
rect 6024 64164 6048 64166
rect 6104 64164 6128 64166
rect 6184 64164 6190 64166
rect 5882 64155 6190 64164
rect 7540 63926 7568 64542
rect 4308 63920 4360 63926
rect 4308 63862 4360 63868
rect 7528 63920 7580 63926
rect 7528 63862 7580 63868
rect 4320 63625 4348 63862
rect 5688 63784 5740 63790
rect 5688 63726 5740 63732
rect 4306 63616 4362 63625
rect 4306 63551 4362 63560
rect 5700 63489 5728 63726
rect 6618 63676 6926 63685
rect 6618 63674 6624 63676
rect 6680 63674 6704 63676
rect 6760 63674 6784 63676
rect 6840 63674 6864 63676
rect 6920 63674 6926 63676
rect 6680 63622 6682 63674
rect 6862 63622 6864 63674
rect 6618 63620 6624 63622
rect 6680 63620 6704 63622
rect 6760 63620 6784 63622
rect 6840 63620 6864 63622
rect 6920 63620 6926 63622
rect 6618 63611 6926 63620
rect 7344 63512 7396 63518
rect 5686 63480 5742 63489
rect 7344 63454 7396 63460
rect 5686 63415 5742 63424
rect 5882 63132 6190 63141
rect 5882 63130 5888 63132
rect 5944 63130 5968 63132
rect 6024 63130 6048 63132
rect 6104 63130 6128 63132
rect 6184 63130 6190 63132
rect 5944 63078 5946 63130
rect 6126 63078 6128 63130
rect 5882 63076 5888 63078
rect 5944 63076 5968 63078
rect 6024 63076 6048 63078
rect 6104 63076 6128 63078
rect 6184 63076 6190 63078
rect 5882 63067 6190 63076
rect 6618 62588 6926 62597
rect 6618 62586 6624 62588
rect 6680 62586 6704 62588
rect 6760 62586 6784 62588
rect 6840 62586 6864 62588
rect 6920 62586 6926 62588
rect 6680 62534 6682 62586
rect 6862 62534 6864 62586
rect 6618 62532 6624 62534
rect 6680 62532 6704 62534
rect 6760 62532 6784 62534
rect 6840 62532 6864 62534
rect 6920 62532 6926 62534
rect 6618 62523 6926 62532
rect 5686 62392 5742 62401
rect 4308 62356 4360 62362
rect 5686 62327 5742 62336
rect 4308 62298 4360 62304
rect 4320 62265 4348 62298
rect 4306 62256 4362 62265
rect 5700 62226 5728 62327
rect 4306 62191 4362 62200
rect 5688 62220 5740 62226
rect 5688 62162 5740 62168
rect 5882 62044 6190 62053
rect 5882 62042 5888 62044
rect 5944 62042 5968 62044
rect 6024 62042 6048 62044
rect 6104 62042 6128 62044
rect 6184 62042 6190 62044
rect 5944 61990 5946 62042
rect 6126 61990 6128 62042
rect 5882 61988 5888 61990
rect 5944 61988 5968 61990
rect 6024 61988 6048 61990
rect 6104 61988 6128 61990
rect 6184 61988 6190 61990
rect 5882 61979 6190 61988
rect 4308 61744 4360 61750
rect 4308 61686 4360 61692
rect 4320 61585 4348 61686
rect 4306 61576 4362 61585
rect 4306 61511 4362 61520
rect 6618 61500 6926 61509
rect 6618 61498 6624 61500
rect 6680 61498 6704 61500
rect 6760 61498 6784 61500
rect 6840 61498 6864 61500
rect 6920 61498 6926 61500
rect 6680 61446 6682 61498
rect 6862 61446 6864 61498
rect 6618 61444 6624 61446
rect 6680 61444 6704 61446
rect 6760 61444 6784 61446
rect 6840 61444 6864 61446
rect 6920 61444 6926 61446
rect 6618 61435 6926 61444
rect 5882 60956 6190 60965
rect 5882 60954 5888 60956
rect 5944 60954 5968 60956
rect 6024 60954 6048 60956
rect 6104 60954 6128 60956
rect 6184 60954 6190 60956
rect 5944 60902 5946 60954
rect 6126 60902 6128 60954
rect 5882 60900 5888 60902
rect 5944 60900 5968 60902
rect 6024 60900 6048 60902
rect 6104 60900 6128 60902
rect 6184 60900 6190 60902
rect 5882 60891 6190 60900
rect 4308 60656 4360 60662
rect 4308 60598 4360 60604
rect 4320 60225 4348 60598
rect 6618 60412 6926 60421
rect 6618 60410 6624 60412
rect 6680 60410 6704 60412
rect 6760 60410 6784 60412
rect 6840 60410 6864 60412
rect 6920 60410 6926 60412
rect 6680 60358 6682 60410
rect 6862 60358 6864 60410
rect 6618 60356 6624 60358
rect 6680 60356 6704 60358
rect 6760 60356 6784 60358
rect 6840 60356 6864 60358
rect 6920 60356 6926 60358
rect 6618 60347 6926 60356
rect 4306 60216 4362 60225
rect 4306 60151 4362 60160
rect 5882 59868 6190 59877
rect 5882 59866 5888 59868
rect 5944 59866 5968 59868
rect 6024 59866 6048 59868
rect 6104 59866 6128 59868
rect 6184 59866 6190 59868
rect 5944 59814 5946 59866
rect 6126 59814 6128 59866
rect 5882 59812 5888 59814
rect 5944 59812 5968 59814
rect 6024 59812 6048 59814
rect 6104 59812 6128 59814
rect 6184 59812 6190 59814
rect 5882 59803 6190 59812
rect 4308 59568 4360 59574
rect 4306 59536 4308 59545
rect 4360 59536 4362 59545
rect 4306 59471 4362 59480
rect 6618 59324 6926 59333
rect 6618 59322 6624 59324
rect 6680 59322 6704 59324
rect 6760 59322 6784 59324
rect 6840 59322 6864 59324
rect 6920 59322 6926 59324
rect 6680 59270 6682 59322
rect 6862 59270 6864 59322
rect 6618 59268 6624 59270
rect 6680 59268 6704 59270
rect 6760 59268 6784 59270
rect 6840 59268 6864 59270
rect 6920 59268 6926 59270
rect 6618 59259 6926 59268
rect 5882 58780 6190 58789
rect 5882 58778 5888 58780
rect 5944 58778 5968 58780
rect 6024 58778 6048 58780
rect 6104 58778 6128 58780
rect 6184 58778 6190 58780
rect 5944 58726 5946 58778
rect 6126 58726 6128 58778
rect 5882 58724 5888 58726
rect 5944 58724 5968 58726
rect 6024 58724 6048 58726
rect 6104 58724 6128 58726
rect 6184 58724 6190 58726
rect 5882 58715 6190 58724
rect 4308 58480 4360 58486
rect 4308 58422 4360 58428
rect 4320 58185 4348 58422
rect 5412 58344 5464 58350
rect 5412 58286 5464 58292
rect 4306 58176 4362 58185
rect 4306 58111 4362 58120
rect 5424 58049 5452 58286
rect 6618 58236 6926 58245
rect 6618 58234 6624 58236
rect 6680 58234 6704 58236
rect 6760 58234 6784 58236
rect 6840 58234 6864 58236
rect 6920 58234 6926 58236
rect 6680 58182 6682 58234
rect 6862 58182 6864 58234
rect 6618 58180 6624 58182
rect 6680 58180 6704 58182
rect 6760 58180 6784 58182
rect 6840 58180 6864 58182
rect 6920 58180 6926 58182
rect 6618 58171 6926 58180
rect 5410 58040 5466 58049
rect 5410 57975 5466 57984
rect 5882 57692 6190 57701
rect 5882 57690 5888 57692
rect 5944 57690 5968 57692
rect 6024 57690 6048 57692
rect 6104 57690 6128 57692
rect 6184 57690 6190 57692
rect 5944 57638 5946 57690
rect 6126 57638 6128 57690
rect 5882 57636 5888 57638
rect 5944 57636 5968 57638
rect 6024 57636 6048 57638
rect 6104 57636 6128 57638
rect 6184 57636 6190 57638
rect 5882 57627 6190 57636
rect 6618 57148 6926 57157
rect 6618 57146 6624 57148
rect 6680 57146 6704 57148
rect 6760 57146 6784 57148
rect 6840 57146 6864 57148
rect 6920 57146 6926 57148
rect 6680 57094 6682 57146
rect 6862 57094 6864 57146
rect 6618 57092 6624 57094
rect 6680 57092 6704 57094
rect 6760 57092 6784 57094
rect 6840 57092 6864 57094
rect 6920 57092 6926 57094
rect 6618 57083 6926 57092
rect 4308 56916 4360 56922
rect 4308 56858 4360 56864
rect 4320 56825 4348 56858
rect 4306 56816 4362 56825
rect 4306 56751 4362 56760
rect 5882 56604 6190 56613
rect 5882 56602 5888 56604
rect 5944 56602 5968 56604
rect 6024 56602 6048 56604
rect 6104 56602 6128 56604
rect 6184 56602 6190 56604
rect 5944 56550 5946 56602
rect 6126 56550 6128 56602
rect 5882 56548 5888 56550
rect 5944 56548 5968 56550
rect 6024 56548 6048 56550
rect 6104 56548 6128 56550
rect 6184 56548 6190 56550
rect 5882 56539 6190 56548
rect 4308 56304 4360 56310
rect 4308 56246 4360 56252
rect 4320 56145 4348 56246
rect 4306 56136 4362 56145
rect 4306 56071 4362 56080
rect 6618 56060 6926 56069
rect 6618 56058 6624 56060
rect 6680 56058 6704 56060
rect 6760 56058 6784 56060
rect 6840 56058 6864 56060
rect 6920 56058 6926 56060
rect 6680 56006 6682 56058
rect 6862 56006 6864 56058
rect 6618 56004 6624 56006
rect 6680 56004 6704 56006
rect 6760 56004 6784 56006
rect 6840 56004 6864 56006
rect 6920 56004 6926 56006
rect 6618 55995 6926 56004
rect 5882 55516 6190 55525
rect 5882 55514 5888 55516
rect 5944 55514 5968 55516
rect 6024 55514 6048 55516
rect 6104 55514 6128 55516
rect 6184 55514 6190 55516
rect 5944 55462 5946 55514
rect 6126 55462 6128 55514
rect 5882 55460 5888 55462
rect 5944 55460 5968 55462
rect 6024 55460 6048 55462
rect 6104 55460 6128 55462
rect 6184 55460 6190 55462
rect 5882 55451 6190 55460
rect 4308 55216 4360 55222
rect 4308 55158 4360 55164
rect 4320 54785 4348 55158
rect 6618 54972 6926 54981
rect 6618 54970 6624 54972
rect 6680 54970 6704 54972
rect 6760 54970 6784 54972
rect 6840 54970 6864 54972
rect 6920 54970 6926 54972
rect 6680 54918 6682 54970
rect 6862 54918 6864 54970
rect 6618 54916 6624 54918
rect 6680 54916 6704 54918
rect 6760 54916 6784 54918
rect 6840 54916 6864 54918
rect 6920 54916 6926 54918
rect 6618 54907 6926 54916
rect 4306 54776 4362 54785
rect 4306 54711 4362 54720
rect 5882 54428 6190 54437
rect 5882 54426 5888 54428
rect 5944 54426 5968 54428
rect 6024 54426 6048 54428
rect 6104 54426 6128 54428
rect 6184 54426 6190 54428
rect 5944 54374 5946 54426
rect 6126 54374 6128 54426
rect 5882 54372 5888 54374
rect 5944 54372 5968 54374
rect 6024 54372 6048 54374
rect 6104 54372 6128 54374
rect 6184 54372 6190 54374
rect 5882 54363 6190 54372
rect 5688 54196 5740 54202
rect 5688 54138 5740 54144
rect 4308 54128 4360 54134
rect 4306 54096 4308 54105
rect 4360 54096 4362 54105
rect 4306 54031 4362 54040
rect 5700 53697 5728 54138
rect 6618 53884 6926 53893
rect 6618 53882 6624 53884
rect 6680 53882 6704 53884
rect 6760 53882 6784 53884
rect 6840 53882 6864 53884
rect 6920 53882 6926 53884
rect 6680 53830 6682 53882
rect 6862 53830 6864 53882
rect 6618 53828 6624 53830
rect 6680 53828 6704 53830
rect 6760 53828 6784 53830
rect 6840 53828 6864 53830
rect 6920 53828 6926 53830
rect 6618 53819 6926 53828
rect 5686 53688 5742 53697
rect 5686 53623 5742 53632
rect 5882 53340 6190 53349
rect 5882 53338 5888 53340
rect 5944 53338 5968 53340
rect 6024 53338 6048 53340
rect 6104 53338 6128 53340
rect 6184 53338 6190 53340
rect 5944 53286 5946 53338
rect 6126 53286 6128 53338
rect 5882 53284 5888 53286
rect 5944 53284 5968 53286
rect 6024 53284 6048 53286
rect 6104 53284 6128 53286
rect 6184 53284 6190 53286
rect 5882 53275 6190 53284
rect 4308 53040 4360 53046
rect 4308 52982 4360 52988
rect 4320 52745 4348 52982
rect 6618 52796 6926 52805
rect 6618 52794 6624 52796
rect 6680 52794 6704 52796
rect 6760 52794 6784 52796
rect 6840 52794 6864 52796
rect 6920 52794 6926 52796
rect 4306 52736 4362 52745
rect 6680 52742 6682 52794
rect 6862 52742 6864 52794
rect 6618 52740 6624 52742
rect 6680 52740 6704 52742
rect 6760 52740 6784 52742
rect 6840 52740 6864 52742
rect 6920 52740 6926 52742
rect 6618 52731 6926 52740
rect 4306 52671 4362 52680
rect 5882 52252 6190 52261
rect 5882 52250 5888 52252
rect 5944 52250 5968 52252
rect 6024 52250 6048 52252
rect 6104 52250 6128 52252
rect 6184 52250 6190 52252
rect 5944 52198 5946 52250
rect 6126 52198 6128 52250
rect 5882 52196 5888 52198
rect 5944 52196 5968 52198
rect 6024 52196 6048 52198
rect 6104 52196 6128 52198
rect 6184 52196 6190 52198
rect 5882 52187 6190 52196
rect 6618 51708 6926 51717
rect 6618 51706 6624 51708
rect 6680 51706 6704 51708
rect 6760 51706 6784 51708
rect 6840 51706 6864 51708
rect 6920 51706 6926 51708
rect 6680 51654 6682 51706
rect 6862 51654 6864 51706
rect 6618 51652 6624 51654
rect 6680 51652 6704 51654
rect 6760 51652 6784 51654
rect 6840 51652 6864 51654
rect 6920 51652 6926 51654
rect 6618 51643 6926 51652
rect 4308 51476 4360 51482
rect 4308 51418 4360 51424
rect 4320 51385 4348 51418
rect 4306 51376 4362 51385
rect 4306 51311 4362 51320
rect 5882 51164 6190 51173
rect 5882 51162 5888 51164
rect 5944 51162 5968 51164
rect 6024 51162 6048 51164
rect 6104 51162 6128 51164
rect 6184 51162 6190 51164
rect 5944 51110 5946 51162
rect 6126 51110 6128 51162
rect 5882 51108 5888 51110
rect 5944 51108 5968 51110
rect 6024 51108 6048 51110
rect 6104 51108 6128 51110
rect 6184 51108 6190 51110
rect 5882 51099 6190 51108
rect 6618 50620 6926 50629
rect 6618 50618 6624 50620
rect 6680 50618 6704 50620
rect 6760 50618 6784 50620
rect 6840 50618 6864 50620
rect 6920 50618 6926 50620
rect 6680 50566 6682 50618
rect 6862 50566 6864 50618
rect 6618 50564 6624 50566
rect 6680 50564 6704 50566
rect 6760 50564 6784 50566
rect 6840 50564 6864 50566
rect 6920 50564 6926 50566
rect 6618 50555 6926 50564
rect 5882 50076 6190 50085
rect 5882 50074 5888 50076
rect 5944 50074 5968 50076
rect 6024 50074 6048 50076
rect 6104 50074 6128 50076
rect 6184 50074 6190 50076
rect 5944 50022 5946 50074
rect 6126 50022 6128 50074
rect 5882 50020 5888 50022
rect 5944 50020 5968 50022
rect 6024 50020 6048 50022
rect 6104 50020 6128 50022
rect 6184 50020 6190 50022
rect 5882 50011 6190 50020
rect 6618 49532 6926 49541
rect 6618 49530 6624 49532
rect 6680 49530 6704 49532
rect 6760 49530 6784 49532
rect 6840 49530 6864 49532
rect 6920 49530 6926 49532
rect 6680 49478 6682 49530
rect 6862 49478 6864 49530
rect 6618 49476 6624 49478
rect 6680 49476 6704 49478
rect 6760 49476 6784 49478
rect 6840 49476 6864 49478
rect 6920 49476 6926 49478
rect 6618 49467 6926 49476
rect 5882 48988 6190 48997
rect 5882 48986 5888 48988
rect 5944 48986 5968 48988
rect 6024 48986 6048 48988
rect 6104 48986 6128 48988
rect 6184 48986 6190 48988
rect 5944 48934 5946 48986
rect 6126 48934 6128 48986
rect 5882 48932 5888 48934
rect 5944 48932 5968 48934
rect 6024 48932 6048 48934
rect 6104 48932 6128 48934
rect 6184 48932 6190 48934
rect 5882 48923 6190 48932
rect 6618 48444 6926 48453
rect 6618 48442 6624 48444
rect 6680 48442 6704 48444
rect 6760 48442 6784 48444
rect 6840 48442 6864 48444
rect 6920 48442 6926 48444
rect 6680 48390 6682 48442
rect 6862 48390 6864 48442
rect 6618 48388 6624 48390
rect 6680 48388 6704 48390
rect 6760 48388 6784 48390
rect 6840 48388 6864 48390
rect 6920 48388 6926 48390
rect 6618 48379 6926 48388
rect 5882 47900 6190 47909
rect 5882 47898 5888 47900
rect 5944 47898 5968 47900
rect 6024 47898 6048 47900
rect 6104 47898 6128 47900
rect 6184 47898 6190 47900
rect 5944 47846 5946 47898
rect 6126 47846 6128 47898
rect 5882 47844 5888 47846
rect 5944 47844 5968 47846
rect 6024 47844 6048 47846
rect 6104 47844 6128 47846
rect 6184 47844 6190 47846
rect 5882 47835 6190 47844
rect 6618 47356 6926 47365
rect 6618 47354 6624 47356
rect 6680 47354 6704 47356
rect 6760 47354 6784 47356
rect 6840 47354 6864 47356
rect 6920 47354 6926 47356
rect 6680 47302 6682 47354
rect 6862 47302 6864 47354
rect 6618 47300 6624 47302
rect 6680 47300 6704 47302
rect 6760 47300 6784 47302
rect 6840 47300 6864 47302
rect 6920 47300 6926 47302
rect 6618 47291 6926 47300
rect 5882 46812 6190 46821
rect 5882 46810 5888 46812
rect 5944 46810 5968 46812
rect 6024 46810 6048 46812
rect 6104 46810 6128 46812
rect 6184 46810 6190 46812
rect 5944 46758 5946 46810
rect 6126 46758 6128 46810
rect 5882 46756 5888 46758
rect 5944 46756 5968 46758
rect 6024 46756 6048 46758
rect 6104 46756 6128 46758
rect 6184 46756 6190 46758
rect 5882 46747 6190 46756
rect 6618 46268 6926 46277
rect 6618 46266 6624 46268
rect 6680 46266 6704 46268
rect 6760 46266 6784 46268
rect 6840 46266 6864 46268
rect 6920 46266 6926 46268
rect 6680 46214 6682 46266
rect 6862 46214 6864 46266
rect 6618 46212 6624 46214
rect 6680 46212 6704 46214
rect 6760 46212 6784 46214
rect 6840 46212 6864 46214
rect 6920 46212 6926 46214
rect 6618 46203 6926 46212
rect 5882 45724 6190 45733
rect 5882 45722 5888 45724
rect 5944 45722 5968 45724
rect 6024 45722 6048 45724
rect 6104 45722 6128 45724
rect 6184 45722 6190 45724
rect 5944 45670 5946 45722
rect 6126 45670 6128 45722
rect 5882 45668 5888 45670
rect 5944 45668 5968 45670
rect 6024 45668 6048 45670
rect 6104 45668 6128 45670
rect 6184 45668 6190 45670
rect 5882 45659 6190 45668
rect 7356 45566 7384 63454
rect 7632 45809 7660 82358
rect 7804 82348 7856 82354
rect 7804 82290 7856 82296
rect 7816 63790 7844 82290
rect 8540 81328 8592 81334
rect 8540 81270 8592 81276
rect 8552 81033 8580 81270
rect 8538 81024 8594 81033
rect 8538 80959 8594 80968
rect 8540 80240 8592 80246
rect 8540 80182 8592 80188
rect 8552 79945 8580 80182
rect 8538 79936 8594 79945
rect 8538 79871 8594 79880
rect 8538 78848 8594 78857
rect 8538 78783 8594 78792
rect 8552 78682 8580 78783
rect 8540 78676 8592 78682
rect 8540 78618 8592 78624
rect 8540 78064 8592 78070
rect 8540 78006 8592 78012
rect 8552 77769 8580 78006
rect 8538 77760 8594 77769
rect 8538 77695 8594 77704
rect 8540 76976 8592 76982
rect 8540 76918 8592 76924
rect 8552 76681 8580 76918
rect 8538 76672 8594 76681
rect 8538 76607 8594 76616
rect 8540 75888 8592 75894
rect 8540 75830 8592 75836
rect 8552 75593 8580 75830
rect 8538 75584 8594 75593
rect 8538 75519 8594 75528
rect 8540 72624 8592 72630
rect 8540 72566 8592 72572
rect 8552 72329 8580 72566
rect 8538 72320 8594 72329
rect 8538 72255 8594 72264
rect 8540 71536 8592 71542
rect 8540 71478 8592 71484
rect 8552 71241 8580 71478
rect 8538 71232 8594 71241
rect 8538 71167 8594 71176
rect 8540 70448 8592 70454
rect 8540 70390 8592 70396
rect 8552 70153 8580 70390
rect 8538 70144 8594 70153
rect 8538 70079 8594 70088
rect 8540 67184 8592 67190
rect 8540 67126 8592 67132
rect 8552 66889 8580 67126
rect 8538 66880 8594 66889
rect 8538 66815 8594 66824
rect 8540 66164 8592 66170
rect 8540 66106 8592 66112
rect 8552 65801 8580 66106
rect 8538 65792 8594 65801
rect 8538 65727 8594 65736
rect 8540 65076 8592 65082
rect 8540 65018 8592 65024
rect 8552 64713 8580 65018
rect 8538 64704 8594 64713
rect 8538 64639 8594 64648
rect 7804 63784 7856 63790
rect 7804 63726 7856 63732
rect 7816 63518 7844 63726
rect 7804 63512 7856 63518
rect 7804 63454 7856 63460
rect 8540 61676 8592 61682
rect 8540 61618 8592 61624
rect 8552 61449 8580 61618
rect 8538 61440 8594 61449
rect 8538 61375 8594 61384
rect 8540 60588 8592 60594
rect 8540 60530 8592 60536
rect 8552 60361 8580 60530
rect 8538 60352 8594 60361
rect 8538 60287 8594 60296
rect 8540 59500 8592 59506
rect 8540 59442 8592 59448
rect 8552 59273 8580 59442
rect 8538 59264 8594 59273
rect 8538 59199 8594 59208
rect 8540 55284 8592 55290
rect 8540 55226 8592 55232
rect 8552 54921 8580 55226
rect 8538 54912 8594 54921
rect 8538 54847 8594 54856
rect 8540 53108 8592 53114
rect 8540 53050 8592 53056
rect 8552 52745 8580 53050
rect 8538 52736 8594 52745
rect 8538 52671 8594 52680
rect 8538 51648 8594 51657
rect 8538 51583 8594 51592
rect 8552 51550 8580 51583
rect 8540 51544 8592 51550
rect 8540 51486 8592 51492
rect 7618 45800 7674 45809
rect 7618 45735 7674 45744
rect 7344 45560 7396 45566
rect 7344 45502 7396 45508
rect 4308 45424 4360 45430
rect 4308 45366 4360 45372
rect 5686 45392 5742 45401
rect 4320 45265 4348 45366
rect 5686 45327 5688 45336
rect 5740 45327 5742 45336
rect 5688 45298 5740 45304
rect 4306 45256 4362 45265
rect 4306 45191 4362 45200
rect 6618 45180 6926 45189
rect 6618 45178 6624 45180
rect 6680 45178 6704 45180
rect 6760 45178 6784 45180
rect 6840 45178 6864 45180
rect 6920 45178 6926 45180
rect 6680 45126 6682 45178
rect 6862 45126 6864 45178
rect 6618 45124 6624 45126
rect 6680 45124 6704 45126
rect 6760 45124 6784 45126
rect 6840 45124 6864 45126
rect 6920 45124 6926 45126
rect 6618 45115 6926 45124
rect 7632 45022 7660 45735
rect 9840 45537 9868 83038
rect 10576 82354 10604 84398
rect 11680 82422 11708 84534
rect 12784 83102 12812 84602
rect 13876 84456 13928 84462
rect 13876 84398 13928 84404
rect 13888 83170 13916 84398
rect 13876 83164 13928 83170
rect 13876 83106 13928 83112
rect 12772 83096 12824 83102
rect 12772 83038 12824 83044
rect 11668 82416 11720 82422
rect 11668 82358 11720 82364
rect 10564 82348 10616 82354
rect 10564 82290 10616 82296
rect 10576 82084 10604 82290
rect 11680 82084 11708 82358
rect 12784 82084 12812 83038
rect 13888 82084 13916 83106
rect 15544 83034 15572 87186
rect 14980 83028 15032 83034
rect 14980 82970 15032 82976
rect 15532 83028 15584 83034
rect 15532 82970 15584 82976
rect 14992 82084 15020 82970
rect 16096 82084 16124 87186
rect 17200 82084 17228 87186
rect 17722 87068 18030 87077
rect 17722 87066 17728 87068
rect 17784 87066 17808 87068
rect 17864 87066 17888 87068
rect 17944 87066 17968 87068
rect 18024 87066 18030 87068
rect 17784 87014 17786 87066
rect 17966 87014 17968 87066
rect 17722 87012 17728 87014
rect 17784 87012 17808 87014
rect 17864 87012 17888 87014
rect 17944 87012 17968 87014
rect 18024 87012 18030 87014
rect 17722 87003 18030 87012
rect 17722 85980 18030 85989
rect 17722 85978 17728 85980
rect 17784 85978 17808 85980
rect 17864 85978 17888 85980
rect 17944 85978 17968 85980
rect 18024 85978 18030 85980
rect 17784 85926 17786 85978
rect 17966 85926 17968 85978
rect 17722 85924 17728 85926
rect 17784 85924 17808 85926
rect 17864 85924 17888 85926
rect 17944 85924 17968 85926
rect 18024 85924 18030 85926
rect 17722 85915 18030 85924
rect 17722 84892 18030 84901
rect 17722 84890 17728 84892
rect 17784 84890 17808 84892
rect 17864 84890 17888 84892
rect 17944 84890 17968 84892
rect 18024 84890 18030 84892
rect 17784 84838 17786 84890
rect 17966 84838 17968 84890
rect 17722 84836 17728 84838
rect 17784 84836 17808 84838
rect 17864 84836 17888 84838
rect 17944 84836 17968 84838
rect 18024 84836 18030 84838
rect 17722 84827 18030 84836
rect 18304 82084 18332 87186
rect 18382 86524 18690 86533
rect 18382 86522 18388 86524
rect 18444 86522 18468 86524
rect 18524 86522 18548 86524
rect 18604 86522 18628 86524
rect 18684 86522 18690 86524
rect 18444 86470 18446 86522
rect 18626 86470 18628 86522
rect 18382 86468 18388 86470
rect 18444 86468 18468 86470
rect 18524 86468 18548 86470
rect 18604 86468 18628 86470
rect 18684 86468 18690 86470
rect 18382 86459 18690 86468
rect 18382 85436 18690 85445
rect 18382 85434 18388 85436
rect 18444 85434 18468 85436
rect 18524 85434 18548 85436
rect 18604 85434 18628 85436
rect 18684 85434 18690 85436
rect 18444 85382 18446 85434
rect 18626 85382 18628 85434
rect 18382 85380 18388 85382
rect 18444 85380 18468 85382
rect 18524 85380 18548 85382
rect 18604 85380 18628 85382
rect 18684 85380 18690 85382
rect 18382 85371 18690 85380
rect 18382 84348 18690 84357
rect 18382 84346 18388 84348
rect 18444 84346 18468 84348
rect 18524 84346 18548 84348
rect 18604 84346 18628 84348
rect 18684 84346 18690 84348
rect 18444 84294 18446 84346
rect 18626 84294 18628 84346
rect 18382 84292 18388 84294
rect 18444 84292 18468 84294
rect 18524 84292 18548 84294
rect 18604 84292 18628 84294
rect 18684 84292 18690 84294
rect 18382 84283 18690 84292
rect 19408 82084 19436 87186
rect 20420 87166 20540 87186
rect 20512 82084 20540 87166
rect 21616 82084 21644 87186
rect 22720 82084 22748 87186
rect 23824 82084 23852 87186
rect 24928 82084 24956 87186
rect 26032 82084 26060 87186
rect 27136 82084 27164 87186
rect 28148 87166 28268 87186
rect 28240 82084 28268 87166
rect 29344 82084 29372 87186
rect 30632 83050 30660 87322
rect 30724 87250 30752 88000
rect 31368 87250 31396 88000
rect 32656 87538 32684 88000
rect 32656 87510 32776 87538
rect 31540 87380 31592 87386
rect 31540 87322 31592 87328
rect 32644 87380 32696 87386
rect 32644 87322 32696 87328
rect 30712 87244 30764 87250
rect 30712 87186 30764 87192
rect 31356 87244 31408 87250
rect 31356 87186 31408 87192
rect 30448 83022 30660 83050
rect 30448 82084 30476 83022
rect 31552 82084 31580 87322
rect 32656 82084 32684 87322
rect 32748 87250 32776 87510
rect 33748 87380 33800 87386
rect 33748 87322 33800 87328
rect 32736 87244 32788 87250
rect 32736 87186 32788 87192
rect 33760 82084 33788 87322
rect 33944 87250 33972 88000
rect 34588 87454 34616 88000
rect 34576 87448 34628 87454
rect 34576 87390 34628 87396
rect 34852 87380 34904 87386
rect 34852 87322 34904 87328
rect 33932 87244 33984 87250
rect 33932 87186 33984 87192
rect 34864 82084 34892 87322
rect 35876 87250 35904 88000
rect 36520 87726 36548 88000
rect 36508 87720 36560 87726
rect 36508 87662 36560 87668
rect 36782 87612 37090 87621
rect 36782 87610 36788 87612
rect 36844 87610 36868 87612
rect 36924 87610 36948 87612
rect 37004 87610 37028 87612
rect 37084 87610 37090 87612
rect 36844 87558 36846 87610
rect 37026 87558 37028 87610
rect 36782 87556 36788 87558
rect 36844 87556 36868 87558
rect 36924 87556 36948 87558
rect 37004 87556 37028 87558
rect 37084 87556 37090 87558
rect 36782 87547 37090 87556
rect 37164 87454 37192 88000
rect 37520 87720 37572 87726
rect 37520 87662 37572 87668
rect 37152 87448 37204 87454
rect 37152 87390 37204 87396
rect 35956 87380 36008 87386
rect 35956 87322 36008 87328
rect 37428 87380 37480 87386
rect 37532 87368 37560 87662
rect 37480 87340 37560 87368
rect 37428 87322 37480 87328
rect 35864 87244 35916 87250
rect 35864 87186 35916 87192
rect 35968 82084 35996 87322
rect 36600 87312 36652 87318
rect 36600 87254 36652 87260
rect 36122 87068 36430 87077
rect 36122 87066 36128 87068
rect 36184 87066 36208 87068
rect 36264 87066 36288 87068
rect 36344 87066 36368 87068
rect 36424 87066 36430 87068
rect 36184 87014 36186 87066
rect 36366 87014 36368 87066
rect 36122 87012 36128 87014
rect 36184 87012 36208 87014
rect 36264 87012 36288 87014
rect 36344 87012 36368 87014
rect 36424 87012 36430 87014
rect 36122 87003 36430 87012
rect 36612 86638 36640 87254
rect 37532 86910 37560 87340
rect 37612 87380 37664 87386
rect 37612 87322 37664 87328
rect 37520 86904 37572 86910
rect 37520 86846 37572 86852
rect 36600 86632 36652 86638
rect 36600 86574 36652 86580
rect 36122 85980 36430 85989
rect 36122 85978 36128 85980
rect 36184 85978 36208 85980
rect 36264 85978 36288 85980
rect 36344 85978 36368 85980
rect 36424 85978 36430 85980
rect 36184 85926 36186 85978
rect 36366 85926 36368 85978
rect 36122 85924 36128 85926
rect 36184 85924 36208 85926
rect 36264 85924 36288 85926
rect 36344 85924 36368 85926
rect 36424 85924 36430 85926
rect 36122 85915 36430 85924
rect 36122 84892 36430 84901
rect 36122 84890 36128 84892
rect 36184 84890 36208 84892
rect 36264 84890 36288 84892
rect 36344 84890 36368 84892
rect 36424 84890 36430 84892
rect 36184 84838 36186 84890
rect 36366 84838 36368 84890
rect 36122 84836 36128 84838
rect 36184 84836 36208 84838
rect 36264 84836 36288 84838
rect 36344 84836 36368 84838
rect 36424 84836 36430 84838
rect 36122 84827 36430 84836
rect 36612 84666 36640 86574
rect 36782 86524 37090 86533
rect 36782 86522 36788 86524
rect 36844 86522 36868 86524
rect 36924 86522 36948 86524
rect 37004 86522 37028 86524
rect 37084 86522 37090 86524
rect 36844 86470 36846 86522
rect 37026 86470 37028 86522
rect 36782 86468 36788 86470
rect 36844 86468 36868 86470
rect 36924 86468 36948 86470
rect 37004 86468 37028 86470
rect 37084 86468 37090 86470
rect 36782 86459 37090 86468
rect 36782 85436 37090 85445
rect 36782 85434 36788 85436
rect 36844 85434 36868 85436
rect 36924 85434 36948 85436
rect 37004 85434 37028 85436
rect 37084 85434 37090 85436
rect 36844 85382 36846 85434
rect 37026 85382 37028 85434
rect 36782 85380 36788 85382
rect 36844 85380 36868 85382
rect 36924 85380 36948 85382
rect 37004 85380 37028 85382
rect 37084 85380 37090 85382
rect 36782 85371 37090 85380
rect 36600 84660 36652 84666
rect 36600 84602 36652 84608
rect 36782 84348 37090 84357
rect 36782 84346 36788 84348
rect 36844 84346 36868 84348
rect 36924 84346 36948 84348
rect 37004 84346 37028 84348
rect 37084 84346 37090 84348
rect 36844 84294 36846 84346
rect 37026 84294 37028 84346
rect 36782 84292 36788 84294
rect 36844 84292 36868 84294
rect 36924 84292 36948 84294
rect 37004 84292 37028 84294
rect 37084 84292 37090 84294
rect 36782 84283 37090 84292
rect 37624 83034 37652 87322
rect 37808 86910 37836 88000
rect 38452 87538 38480 88000
rect 38360 87510 38480 87538
rect 38164 87380 38216 87386
rect 38164 87322 38216 87328
rect 37796 86904 37848 86910
rect 37796 86846 37848 86852
rect 37060 83028 37112 83034
rect 37060 82970 37112 82976
rect 37612 83028 37664 83034
rect 37612 82970 37664 82976
rect 37072 82084 37100 82970
rect 38176 82084 38204 87322
rect 38360 87250 38388 87510
rect 39096 87454 39124 88000
rect 39084 87448 39136 87454
rect 39084 87390 39136 87396
rect 38440 87380 38492 87386
rect 38440 87322 38492 87328
rect 39268 87380 39320 87386
rect 39268 87322 39320 87328
rect 38348 87244 38400 87250
rect 38348 87186 38400 87192
rect 38452 86910 38480 87322
rect 39084 87312 39136 87318
rect 39084 87254 39136 87260
rect 38440 86904 38492 86910
rect 38440 86846 38492 86852
rect 39096 84666 39124 87254
rect 39084 84660 39136 84666
rect 39084 84602 39136 84608
rect 39280 82084 39308 87322
rect 39740 84530 39768 88000
rect 40384 87538 40412 88000
rect 40384 87510 40504 87538
rect 40372 87380 40424 87386
rect 40372 87322 40424 87328
rect 39728 84524 39780 84530
rect 39728 84466 39780 84472
rect 40384 82084 40412 87322
rect 40476 87250 40504 87510
rect 41028 87454 41056 88000
rect 41016 87448 41068 87454
rect 41016 87390 41068 87396
rect 41672 87386 41700 88000
rect 42316 87454 42344 88000
rect 42304 87448 42356 87454
rect 42304 87390 42356 87396
rect 42960 87386 42988 88000
rect 41476 87380 41528 87386
rect 41476 87322 41528 87328
rect 41660 87380 41712 87386
rect 41660 87322 41712 87328
rect 42580 87380 42632 87386
rect 42580 87322 42632 87328
rect 42948 87380 43000 87386
rect 42948 87322 43000 87328
rect 40464 87244 40516 87250
rect 40464 87186 40516 87192
rect 41488 82084 41516 87322
rect 42592 82084 42620 87322
rect 43604 87250 43632 88000
rect 44248 87454 44276 88000
rect 44236 87448 44288 87454
rect 44236 87390 44288 87396
rect 44892 87386 44920 88000
rect 45536 87386 45564 88000
rect 46180 87386 46208 88000
rect 46824 87386 46852 88000
rect 47468 87386 47496 88000
rect 48112 87386 48140 88000
rect 48756 87386 48784 88000
rect 49400 87386 49428 88000
rect 50044 87386 50072 88000
rect 52620 87386 52648 88000
rect 53264 87386 53292 88000
rect 54552 87386 54580 88000
rect 55182 87612 55490 87621
rect 55182 87610 55188 87612
rect 55244 87610 55268 87612
rect 55324 87610 55348 87612
rect 55404 87610 55428 87612
rect 55484 87610 55490 87612
rect 55244 87558 55246 87610
rect 55426 87558 55428 87610
rect 55182 87556 55188 87558
rect 55244 87556 55268 87558
rect 55324 87556 55348 87558
rect 55404 87556 55428 87558
rect 55484 87556 55490 87558
rect 55182 87547 55490 87556
rect 55840 87386 55868 88000
rect 57128 87386 57156 88000
rect 57772 87386 57800 88000
rect 59060 87386 59088 88000
rect 60348 87386 60376 88000
rect 60992 87386 61020 88000
rect 62280 87386 62308 88000
rect 63568 87386 63596 88000
rect 64856 87386 64884 88000
rect 65500 87386 65528 88000
rect 66788 87386 66816 88000
rect 43684 87380 43736 87386
rect 43684 87322 43736 87328
rect 44788 87380 44840 87386
rect 44788 87322 44840 87328
rect 44880 87380 44932 87386
rect 44880 87322 44932 87328
rect 45524 87380 45576 87386
rect 45524 87322 45576 87328
rect 46168 87380 46220 87386
rect 46168 87322 46220 87328
rect 46812 87380 46864 87386
rect 46812 87322 46864 87328
rect 47456 87380 47508 87386
rect 47456 87322 47508 87328
rect 48100 87380 48152 87386
rect 48100 87322 48152 87328
rect 48744 87380 48796 87386
rect 48744 87322 48796 87328
rect 49388 87380 49440 87386
rect 49388 87322 49440 87328
rect 50032 87380 50084 87386
rect 50032 87322 50084 87328
rect 52608 87380 52660 87386
rect 52608 87322 52660 87328
rect 53252 87380 53304 87386
rect 53252 87322 53304 87328
rect 54540 87380 54592 87386
rect 54540 87322 54592 87328
rect 55828 87380 55880 87386
rect 55828 87322 55880 87328
rect 57116 87380 57168 87386
rect 57116 87322 57168 87328
rect 57760 87380 57812 87386
rect 57760 87322 57812 87328
rect 59048 87380 59100 87386
rect 59048 87322 59100 87328
rect 60336 87380 60388 87386
rect 60336 87322 60388 87328
rect 60980 87380 61032 87386
rect 60980 87322 61032 87328
rect 62268 87380 62320 87386
rect 62268 87322 62320 87328
rect 63556 87380 63608 87386
rect 63556 87322 63608 87328
rect 64844 87380 64896 87386
rect 64844 87322 64896 87328
rect 65488 87380 65540 87386
rect 65488 87322 65540 87328
rect 66776 87380 66828 87386
rect 66776 87322 66828 87328
rect 67880 87380 67932 87386
rect 67880 87322 67932 87328
rect 43592 87244 43644 87250
rect 43592 87186 43644 87192
rect 43696 82084 43724 87322
rect 44800 82084 44828 87322
rect 52884 87244 52936 87250
rect 52884 87186 52936 87192
rect 53528 87244 53580 87250
rect 53528 87186 53580 87192
rect 54448 87244 54500 87250
rect 54448 87186 54500 87192
rect 55736 87244 55788 87250
rect 55736 87186 55788 87192
rect 56840 87244 56892 87250
rect 56840 87186 56892 87192
rect 57944 87244 57996 87250
rect 57944 87186 57996 87192
rect 59048 87244 59100 87250
rect 59048 87186 59100 87192
rect 60152 87244 60204 87250
rect 60152 87186 60204 87192
rect 61164 87244 61216 87250
rect 62452 87244 62504 87250
rect 61164 87186 61216 87192
rect 62372 87192 62452 87194
rect 62372 87186 62504 87192
rect 63464 87244 63516 87250
rect 63464 87186 63516 87192
rect 64568 87244 64620 87250
rect 64568 87186 64620 87192
rect 65672 87244 65724 87250
rect 65672 87186 65724 87192
rect 66776 87244 66828 87250
rect 66776 87186 66828 87192
rect 46996 86632 47048 86638
rect 46996 86574 47048 86580
rect 50308 86632 50360 86638
rect 50308 86574 50360 86580
rect 46168 84728 46220 84734
rect 46168 84670 46220 84676
rect 46076 84592 46128 84598
rect 46076 84534 46128 84540
rect 45892 84456 45944 84462
rect 45892 84398 45944 84404
rect 45984 84456 46036 84462
rect 45984 84398 46036 84404
rect 9920 56984 9972 56990
rect 9918 56952 9920 56961
rect 9972 56952 9974 56961
rect 9918 56887 9974 56896
rect 9920 56372 9972 56378
rect 9920 56314 9972 56320
rect 9932 56281 9960 56314
rect 9918 56272 9974 56281
rect 9918 56207 9974 56216
rect 45904 49481 45932 84398
rect 45996 50569 46024 84398
rect 45982 50560 46038 50569
rect 45982 50495 46038 50504
rect 45890 49472 45946 49481
rect 45890 49407 45946 49416
rect 11666 45936 11722 45945
rect 10564 45900 10616 45906
rect 11666 45871 11722 45880
rect 12770 45936 12826 45945
rect 12770 45871 12826 45880
rect 13874 45936 13930 45945
rect 13874 45871 13930 45880
rect 10564 45842 10616 45848
rect 10576 45772 10604 45842
rect 11680 45772 11708 45871
rect 12784 45772 12812 45871
rect 13888 45772 13916 45871
rect 14992 45772 15020 46452
rect 16096 45772 16124 46452
rect 17200 45772 17228 46452
rect 18304 45772 18332 46452
rect 19408 45772 19436 46452
rect 20512 45772 20540 46452
rect 21616 45772 21644 46452
rect 22720 45772 22748 46452
rect 23824 45772 23852 46452
rect 24928 45772 24956 46452
rect 26032 45772 26060 46452
rect 27136 45772 27164 46452
rect 28240 45772 28268 46452
rect 29344 45772 29372 46452
rect 30448 45772 30476 46452
rect 31552 45772 31580 46452
rect 32656 45772 32684 46452
rect 33760 45772 33788 46452
rect 34864 45772 34892 46452
rect 35968 45772 35996 46452
rect 37072 45772 37100 46452
rect 38176 45772 38204 46452
rect 39280 45772 39308 46452
rect 40384 45772 40412 46452
rect 41488 45772 41516 46452
rect 42592 45772 42620 46452
rect 43696 45772 43724 46452
rect 44800 45772 44828 46452
rect 8998 45528 9054 45537
rect 8998 45463 9000 45472
rect 9052 45463 9054 45472
rect 9826 45528 9882 45537
rect 9826 45463 9882 45472
rect 9000 45434 9052 45440
rect 7620 45016 7672 45022
rect 7620 44958 7672 44964
rect 8540 44948 8592 44954
rect 8540 44890 8592 44896
rect 4216 44744 4268 44750
rect 8552 44721 8580 44890
rect 4216 44686 4268 44692
rect 8538 44712 8594 44721
rect 4228 44585 4256 44686
rect 8538 44647 8594 44656
rect 5882 44636 6190 44645
rect 5882 44634 5888 44636
rect 5944 44634 5968 44636
rect 6024 44634 6048 44636
rect 6104 44634 6128 44636
rect 6184 44634 6190 44636
rect 4214 44576 4270 44585
rect 5944 44582 5946 44634
rect 6126 44582 6128 44634
rect 5882 44580 5888 44582
rect 5944 44580 5968 44582
rect 6024 44580 6048 44582
rect 6104 44580 6128 44582
rect 6184 44580 6190 44582
rect 5882 44571 6190 44580
rect 4214 44511 4270 44520
rect 6618 44092 6926 44101
rect 6618 44090 6624 44092
rect 6680 44090 6704 44092
rect 6760 44090 6784 44092
rect 6840 44090 6864 44092
rect 6920 44090 6926 44092
rect 6680 44038 6682 44090
rect 6862 44038 6864 44090
rect 6618 44036 6624 44038
rect 6680 44036 6704 44038
rect 6760 44036 6784 44038
rect 6840 44036 6864 44038
rect 6920 44036 6926 44038
rect 6618 44027 6926 44036
rect 5882 43548 6190 43557
rect 5882 43546 5888 43548
rect 5944 43546 5968 43548
rect 6024 43546 6048 43548
rect 6104 43546 6128 43548
rect 6184 43546 6190 43548
rect 5944 43494 5946 43546
rect 6126 43494 6128 43546
rect 5882 43492 5888 43494
rect 5944 43492 5968 43494
rect 6024 43492 6048 43494
rect 6104 43492 6128 43494
rect 6184 43492 6190 43494
rect 5882 43483 6190 43492
rect 8538 43488 8594 43497
rect 8538 43423 8594 43432
rect 8552 43254 8580 43423
rect 4124 43248 4176 43254
rect 4122 43216 4124 43225
rect 8540 43248 8592 43254
rect 4176 43216 4178 43225
rect 8540 43190 8592 43196
rect 4122 43151 4178 43160
rect 6618 43004 6926 43013
rect 6618 43002 6624 43004
rect 6680 43002 6704 43004
rect 6760 43002 6784 43004
rect 6840 43002 6864 43004
rect 6920 43002 6926 43004
rect 6680 42950 6682 43002
rect 6862 42950 6864 43002
rect 6618 42948 6624 42950
rect 6680 42948 6704 42950
rect 6760 42948 6784 42950
rect 6840 42948 6864 42950
rect 6920 42948 6926 42950
rect 6618 42939 6926 42948
rect 8540 42772 8592 42778
rect 8540 42714 8592 42720
rect 4124 42568 4176 42574
rect 4122 42536 4124 42545
rect 8552 42545 8580 42714
rect 4176 42536 4178 42545
rect 4122 42471 4178 42480
rect 8538 42536 8594 42545
rect 8538 42471 8594 42480
rect 5882 42460 6190 42469
rect 5882 42458 5888 42460
rect 5944 42458 5968 42460
rect 6024 42458 6048 42460
rect 6104 42458 6128 42460
rect 6184 42458 6190 42460
rect 5944 42406 5946 42458
rect 6126 42406 6128 42458
rect 5882 42404 5888 42406
rect 5944 42404 5968 42406
rect 6024 42404 6048 42406
rect 6104 42404 6128 42406
rect 6184 42404 6190 42406
rect 5882 42395 6190 42404
rect 6618 41916 6926 41925
rect 6618 41914 6624 41916
rect 6680 41914 6704 41916
rect 6760 41914 6784 41916
rect 6840 41914 6864 41916
rect 6920 41914 6926 41916
rect 6680 41862 6682 41914
rect 6862 41862 6864 41914
rect 6618 41860 6624 41862
rect 6680 41860 6704 41862
rect 6760 41860 6784 41862
rect 6840 41860 6864 41862
rect 6920 41860 6926 41862
rect 6618 41851 6926 41860
rect 4124 41684 4176 41690
rect 4124 41626 4176 41632
rect 5412 41684 5464 41690
rect 5412 41626 5464 41632
rect 4136 41185 4164 41626
rect 5424 41593 5452 41626
rect 5410 41584 5466 41593
rect 5410 41519 5466 41528
rect 5882 41372 6190 41381
rect 5882 41370 5888 41372
rect 5944 41370 5968 41372
rect 6024 41370 6048 41372
rect 6104 41370 6128 41372
rect 6184 41370 6190 41372
rect 5944 41318 5946 41370
rect 6126 41318 6128 41370
rect 5882 41316 5888 41318
rect 5944 41316 5968 41318
rect 6024 41316 6048 41318
rect 6104 41316 6128 41318
rect 6184 41316 6190 41318
rect 5882 41307 6190 41316
rect 4122 41176 4178 41185
rect 4122 41111 4178 41120
rect 6618 40828 6926 40837
rect 6618 40826 6624 40828
rect 6680 40826 6704 40828
rect 6760 40826 6784 40828
rect 6840 40826 6864 40828
rect 6920 40826 6926 40828
rect 6680 40774 6682 40826
rect 6862 40774 6864 40826
rect 6618 40772 6624 40774
rect 6680 40772 6704 40774
rect 6760 40772 6784 40774
rect 6840 40772 6864 40774
rect 6920 40772 6926 40774
rect 6618 40763 6926 40772
rect 8540 40596 8592 40602
rect 8540 40538 8592 40544
rect 3938 40496 3994 40505
rect 3938 40431 3940 40440
rect 3992 40431 3994 40440
rect 3940 40402 3992 40408
rect 8552 40369 8580 40538
rect 8538 40360 8594 40369
rect 8538 40295 8594 40304
rect 5882 40284 6190 40293
rect 5882 40282 5888 40284
rect 5944 40282 5968 40284
rect 6024 40282 6048 40284
rect 6104 40282 6128 40284
rect 6184 40282 6190 40284
rect 5944 40230 5946 40282
rect 6126 40230 6128 40282
rect 5882 40228 5888 40230
rect 5944 40228 5968 40230
rect 6024 40228 6048 40230
rect 6104 40228 6128 40230
rect 6184 40228 6190 40230
rect 5882 40219 6190 40228
rect 6618 39740 6926 39749
rect 6618 39738 6624 39740
rect 6680 39738 6704 39740
rect 6760 39738 6784 39740
rect 6840 39738 6864 39740
rect 6920 39738 6926 39740
rect 6680 39686 6682 39738
rect 6862 39686 6864 39738
rect 6618 39684 6624 39686
rect 6680 39684 6704 39686
rect 6760 39684 6784 39686
rect 6840 39684 6864 39686
rect 6920 39684 6926 39686
rect 6618 39675 6926 39684
rect 8540 39508 8592 39514
rect 8540 39450 8592 39456
rect 4216 39304 4268 39310
rect 8552 39281 8580 39450
rect 4216 39246 4268 39252
rect 8538 39272 8594 39281
rect 4228 39145 4256 39246
rect 8538 39207 8594 39216
rect 5882 39196 6190 39205
rect 5882 39194 5888 39196
rect 5944 39194 5968 39196
rect 6024 39194 6048 39196
rect 6104 39194 6128 39196
rect 6184 39194 6190 39196
rect 4214 39136 4270 39145
rect 5944 39142 5946 39194
rect 6126 39142 6128 39194
rect 5882 39140 5888 39142
rect 5944 39140 5968 39142
rect 6024 39140 6048 39142
rect 6104 39140 6128 39142
rect 6184 39140 6190 39142
rect 5882 39131 6190 39140
rect 4214 39071 4270 39080
rect 6618 38652 6926 38661
rect 6618 38650 6624 38652
rect 6680 38650 6704 38652
rect 6760 38650 6784 38652
rect 6840 38650 6864 38652
rect 6920 38650 6926 38652
rect 6680 38598 6682 38650
rect 6862 38598 6864 38650
rect 6618 38596 6624 38598
rect 6680 38596 6704 38598
rect 6760 38596 6784 38598
rect 6840 38596 6864 38598
rect 6920 38596 6926 38598
rect 6618 38587 6926 38596
rect 5882 38108 6190 38117
rect 5882 38106 5888 38108
rect 5944 38106 5968 38108
rect 6024 38106 6048 38108
rect 6104 38106 6128 38108
rect 6184 38106 6190 38108
rect 5944 38054 5946 38106
rect 6126 38054 6128 38106
rect 5882 38052 5888 38054
rect 5944 38052 5968 38054
rect 6024 38052 6048 38054
rect 6104 38052 6128 38054
rect 6184 38052 6190 38054
rect 5882 38043 6190 38052
rect 8538 38048 8594 38057
rect 8538 37983 8594 37992
rect 8552 37814 8580 37983
rect 4216 37808 4268 37814
rect 4214 37776 4216 37785
rect 8540 37808 8592 37814
rect 4268 37776 4270 37785
rect 8540 37750 8592 37756
rect 4214 37711 4270 37720
rect 6618 37564 6926 37573
rect 6618 37562 6624 37564
rect 6680 37562 6704 37564
rect 6760 37562 6784 37564
rect 6840 37562 6864 37564
rect 6920 37562 6926 37564
rect 6680 37510 6682 37562
rect 6862 37510 6864 37562
rect 6618 37508 6624 37510
rect 6680 37508 6704 37510
rect 6760 37508 6784 37510
rect 6840 37508 6864 37510
rect 6920 37508 6926 37510
rect 6618 37499 6926 37508
rect 8540 37332 8592 37338
rect 8540 37274 8592 37280
rect 4124 37128 4176 37134
rect 4122 37096 4124 37105
rect 8552 37105 8580 37274
rect 4176 37096 4178 37105
rect 4122 37031 4178 37040
rect 8538 37096 8594 37105
rect 8538 37031 8594 37040
rect 5882 37020 6190 37029
rect 5882 37018 5888 37020
rect 5944 37018 5968 37020
rect 6024 37018 6048 37020
rect 6104 37018 6128 37020
rect 6184 37018 6190 37020
rect 5944 36966 5946 37018
rect 6126 36966 6128 37018
rect 5882 36964 5888 36966
rect 5944 36964 5968 36966
rect 6024 36964 6048 36966
rect 6104 36964 6128 36966
rect 6184 36964 6190 36966
rect 5882 36955 6190 36964
rect 6618 36476 6926 36485
rect 6618 36474 6624 36476
rect 6680 36474 6704 36476
rect 6760 36474 6784 36476
rect 6840 36474 6864 36476
rect 6920 36474 6926 36476
rect 6680 36422 6682 36474
rect 6862 36422 6864 36474
rect 6618 36420 6624 36422
rect 6680 36420 6704 36422
rect 6760 36420 6784 36422
rect 6840 36420 6864 36422
rect 6920 36420 6926 36422
rect 6618 36411 6926 36420
rect 5412 36244 5464 36250
rect 5412 36186 5464 36192
rect 4124 36176 4176 36182
rect 5424 36153 5452 36186
rect 4124 36118 4176 36124
rect 5410 36144 5466 36153
rect 4136 35745 4164 36118
rect 5410 36079 5466 36088
rect 5882 35932 6190 35941
rect 5882 35930 5888 35932
rect 5944 35930 5968 35932
rect 6024 35930 6048 35932
rect 6104 35930 6128 35932
rect 6184 35930 6190 35932
rect 5944 35878 5946 35930
rect 6126 35878 6128 35930
rect 5882 35876 5888 35878
rect 5944 35876 5968 35878
rect 6024 35876 6048 35878
rect 6104 35876 6128 35878
rect 6184 35876 6190 35878
rect 5882 35867 6190 35876
rect 4122 35736 4178 35745
rect 4122 35671 4178 35680
rect 6618 35388 6926 35397
rect 6618 35386 6624 35388
rect 6680 35386 6704 35388
rect 6760 35386 6784 35388
rect 6840 35386 6864 35388
rect 6920 35386 6926 35388
rect 6680 35334 6682 35386
rect 6862 35334 6864 35386
rect 6618 35332 6624 35334
rect 6680 35332 6704 35334
rect 6760 35332 6784 35334
rect 6840 35332 6864 35334
rect 6920 35332 6926 35334
rect 6618 35323 6926 35332
rect 8540 35156 8592 35162
rect 8540 35098 8592 35104
rect 4216 35088 4268 35094
rect 4214 35056 4216 35065
rect 4268 35056 4270 35065
rect 4214 34991 4270 35000
rect 8552 34929 8580 35098
rect 8538 34920 8594 34929
rect 8538 34855 8594 34864
rect 5882 34844 6190 34853
rect 5882 34842 5888 34844
rect 5944 34842 5968 34844
rect 6024 34842 6048 34844
rect 6104 34842 6128 34844
rect 6184 34842 6190 34844
rect 5944 34790 5946 34842
rect 6126 34790 6128 34842
rect 5882 34788 5888 34790
rect 5944 34788 5968 34790
rect 6024 34788 6048 34790
rect 6104 34788 6128 34790
rect 6184 34788 6190 34790
rect 5882 34779 6190 34788
rect 6618 34300 6926 34309
rect 6618 34298 6624 34300
rect 6680 34298 6704 34300
rect 6760 34298 6784 34300
rect 6840 34298 6864 34300
rect 6920 34298 6926 34300
rect 6680 34246 6682 34298
rect 6862 34246 6864 34298
rect 6618 34244 6624 34246
rect 6680 34244 6704 34246
rect 6760 34244 6784 34246
rect 6840 34244 6864 34246
rect 6920 34244 6926 34246
rect 6618 34235 6926 34244
rect 8540 34068 8592 34074
rect 8540 34010 8592 34016
rect 4216 33864 4268 33870
rect 8552 33841 8580 34010
rect 4216 33806 4268 33812
rect 8538 33832 8594 33841
rect 4228 33705 4256 33806
rect 8538 33767 8594 33776
rect 5882 33756 6190 33765
rect 5882 33754 5888 33756
rect 5944 33754 5968 33756
rect 6024 33754 6048 33756
rect 6104 33754 6128 33756
rect 6184 33754 6190 33756
rect 4214 33696 4270 33705
rect 5944 33702 5946 33754
rect 6126 33702 6128 33754
rect 5882 33700 5888 33702
rect 5944 33700 5968 33702
rect 6024 33700 6048 33702
rect 6104 33700 6128 33702
rect 6184 33700 6190 33702
rect 5882 33691 6190 33700
rect 4214 33631 4270 33640
rect 6618 33212 6926 33221
rect 6618 33210 6624 33212
rect 6680 33210 6704 33212
rect 6760 33210 6784 33212
rect 6840 33210 6864 33212
rect 6920 33210 6926 33212
rect 6680 33158 6682 33210
rect 6862 33158 6864 33210
rect 6618 33156 6624 33158
rect 6680 33156 6704 33158
rect 6760 33156 6784 33158
rect 6840 33156 6864 33158
rect 6920 33156 6926 33158
rect 6618 33147 6926 33156
rect 5882 32668 6190 32677
rect 5882 32666 5888 32668
rect 5944 32666 5968 32668
rect 6024 32666 6048 32668
rect 6104 32666 6128 32668
rect 6184 32666 6190 32668
rect 5944 32614 5946 32666
rect 6126 32614 6128 32666
rect 5882 32612 5888 32614
rect 5944 32612 5968 32614
rect 6024 32612 6048 32614
rect 6104 32612 6128 32614
rect 6184 32612 6190 32614
rect 5882 32603 6190 32612
rect 8538 32608 8594 32617
rect 8538 32543 8594 32552
rect 8552 32374 8580 32543
rect 4216 32368 4268 32374
rect 4214 32336 4216 32345
rect 8540 32368 8592 32374
rect 4268 32336 4270 32345
rect 8540 32310 8592 32316
rect 4214 32271 4270 32280
rect 6618 32124 6926 32133
rect 6618 32122 6624 32124
rect 6680 32122 6704 32124
rect 6760 32122 6784 32124
rect 6840 32122 6864 32124
rect 6920 32122 6926 32124
rect 6680 32070 6682 32122
rect 6862 32070 6864 32122
rect 6618 32068 6624 32070
rect 6680 32068 6704 32070
rect 6760 32068 6784 32070
rect 6840 32068 6864 32070
rect 6920 32068 6926 32070
rect 6618 32059 6926 32068
rect 8540 31892 8592 31898
rect 8540 31834 8592 31840
rect 4124 31688 4176 31694
rect 4122 31656 4124 31665
rect 8552 31665 8580 31834
rect 4176 31656 4178 31665
rect 4122 31591 4178 31600
rect 8538 31656 8594 31665
rect 8538 31591 8594 31600
rect 5882 31580 6190 31589
rect 5882 31578 5888 31580
rect 5944 31578 5968 31580
rect 6024 31578 6048 31580
rect 6104 31578 6128 31580
rect 6184 31578 6190 31580
rect 5944 31526 5946 31578
rect 6126 31526 6128 31578
rect 5882 31524 5888 31526
rect 5944 31524 5968 31526
rect 6024 31524 6048 31526
rect 6104 31524 6128 31526
rect 6184 31524 6190 31526
rect 5882 31515 6190 31524
rect 6618 31036 6926 31045
rect 6618 31034 6624 31036
rect 6680 31034 6704 31036
rect 6760 31034 6784 31036
rect 6840 31034 6864 31036
rect 6920 31034 6926 31036
rect 6680 30982 6682 31034
rect 6862 30982 6864 31034
rect 6618 30980 6624 30982
rect 6680 30980 6704 30982
rect 6760 30980 6784 30982
rect 6840 30980 6864 30982
rect 6920 30980 6926 30982
rect 6618 30971 6926 30980
rect 5412 30804 5464 30810
rect 5412 30746 5464 30752
rect 4124 30668 4176 30674
rect 4124 30610 4176 30616
rect 4136 30305 4164 30610
rect 5424 30305 5452 30746
rect 5882 30492 6190 30501
rect 5882 30490 5888 30492
rect 5944 30490 5968 30492
rect 6024 30490 6048 30492
rect 6104 30490 6128 30492
rect 6184 30490 6190 30492
rect 5944 30438 5946 30490
rect 6126 30438 6128 30490
rect 5882 30436 5888 30438
rect 5944 30436 5968 30438
rect 6024 30436 6048 30438
rect 6104 30436 6128 30438
rect 6184 30436 6190 30438
rect 5882 30427 6190 30436
rect 4122 30296 4178 30305
rect 4122 30231 4178 30240
rect 5410 30296 5466 30305
rect 5410 30231 5466 30240
rect 6618 29948 6926 29957
rect 6618 29946 6624 29948
rect 6680 29946 6704 29948
rect 6760 29946 6784 29948
rect 6840 29946 6864 29948
rect 6920 29946 6926 29948
rect 6680 29894 6682 29946
rect 6862 29894 6864 29946
rect 6618 29892 6624 29894
rect 6680 29892 6704 29894
rect 6760 29892 6784 29894
rect 6840 29892 6864 29894
rect 6920 29892 6926 29894
rect 6618 29883 6926 29892
rect 4308 29716 4360 29722
rect 4308 29658 4360 29664
rect 4320 29625 4348 29658
rect 4306 29616 4362 29625
rect 4306 29551 4362 29560
rect 8540 29580 8592 29586
rect 8540 29522 8592 29528
rect 8552 29489 8580 29522
rect 8538 29480 8594 29489
rect 8538 29415 8594 29424
rect 5882 29404 6190 29413
rect 5882 29402 5888 29404
rect 5944 29402 5968 29404
rect 6024 29402 6048 29404
rect 6104 29402 6128 29404
rect 6184 29402 6190 29404
rect 5944 29350 5946 29402
rect 6126 29350 6128 29402
rect 5882 29348 5888 29350
rect 5944 29348 5968 29350
rect 6024 29348 6048 29350
rect 6104 29348 6128 29350
rect 6184 29348 6190 29350
rect 5882 29339 6190 29348
rect 6618 28860 6926 28869
rect 6618 28858 6624 28860
rect 6680 28858 6704 28860
rect 6760 28858 6784 28860
rect 6840 28858 6864 28860
rect 6920 28858 6926 28860
rect 6680 28806 6682 28858
rect 6862 28806 6864 28858
rect 6618 28804 6624 28806
rect 6680 28804 6704 28806
rect 6760 28804 6784 28806
rect 6840 28804 6864 28806
rect 6920 28804 6926 28806
rect 6618 28795 6926 28804
rect 4308 28628 4360 28634
rect 4308 28570 4360 28576
rect 4320 28265 4348 28570
rect 8540 28492 8592 28498
rect 8540 28434 8592 28440
rect 8552 28401 8580 28434
rect 8538 28392 8594 28401
rect 8538 28327 8594 28336
rect 5882 28316 6190 28325
rect 5882 28314 5888 28316
rect 5944 28314 5968 28316
rect 6024 28314 6048 28316
rect 6104 28314 6128 28316
rect 6184 28314 6190 28316
rect 4306 28256 4362 28265
rect 5944 28262 5946 28314
rect 6126 28262 6128 28314
rect 5882 28260 5888 28262
rect 5944 28260 5968 28262
rect 6024 28260 6048 28262
rect 6104 28260 6128 28262
rect 6184 28260 6190 28262
rect 5882 28251 6190 28260
rect 4306 28191 4362 28200
rect 6618 27772 6926 27781
rect 6618 27770 6624 27772
rect 6680 27770 6704 27772
rect 6760 27770 6784 27772
rect 6840 27770 6864 27772
rect 6920 27770 6926 27772
rect 6680 27718 6682 27770
rect 6862 27718 6864 27770
rect 6618 27716 6624 27718
rect 6680 27716 6704 27718
rect 6760 27716 6784 27718
rect 6840 27716 6864 27718
rect 6920 27716 6926 27718
rect 6618 27707 6926 27716
rect 5882 27228 6190 27237
rect 5882 27226 5888 27228
rect 5944 27226 5968 27228
rect 6024 27226 6048 27228
rect 6104 27226 6128 27228
rect 6184 27226 6190 27228
rect 5944 27174 5946 27226
rect 6126 27174 6128 27226
rect 5882 27172 5888 27174
rect 5944 27172 5968 27174
rect 6024 27172 6048 27174
rect 6104 27172 6128 27174
rect 6184 27172 6190 27174
rect 5882 27163 6190 27172
rect 8538 27168 8594 27177
rect 8538 27103 8594 27112
rect 8552 27070 8580 27103
rect 8540 27064 8592 27070
rect 8540 27006 8592 27012
rect 4308 26928 4360 26934
rect 4306 26896 4308 26905
rect 4360 26896 4362 26905
rect 4306 26831 4362 26840
rect 6618 26684 6926 26693
rect 6618 26682 6624 26684
rect 6680 26682 6704 26684
rect 6760 26682 6784 26684
rect 6840 26682 6864 26684
rect 6920 26682 6926 26684
rect 6680 26630 6682 26682
rect 6862 26630 6864 26682
rect 6618 26628 6624 26630
rect 6680 26628 6704 26630
rect 6760 26628 6784 26630
rect 6840 26628 6864 26630
rect 6920 26628 6926 26630
rect 6618 26619 6926 26628
rect 4308 26452 4360 26458
rect 4308 26394 4360 26400
rect 4320 26225 4348 26394
rect 8540 26316 8592 26322
rect 8540 26258 8592 26264
rect 8552 26225 8580 26258
rect 4306 26216 4362 26225
rect 4306 26151 4362 26160
rect 8538 26216 8594 26225
rect 8538 26151 8594 26160
rect 5882 26140 6190 26149
rect 5882 26138 5888 26140
rect 5944 26138 5968 26140
rect 6024 26138 6048 26140
rect 6104 26138 6128 26140
rect 6184 26138 6190 26140
rect 5944 26086 5946 26138
rect 6126 26086 6128 26138
rect 5882 26084 5888 26086
rect 5944 26084 5968 26086
rect 6024 26084 6048 26086
rect 6104 26084 6128 26086
rect 6184 26084 6190 26086
rect 5882 26075 6190 26084
rect 6618 25596 6926 25605
rect 6618 25594 6624 25596
rect 6680 25594 6704 25596
rect 6760 25594 6784 25596
rect 6840 25594 6864 25596
rect 6920 25594 6926 25596
rect 6680 25542 6682 25594
rect 6862 25542 6864 25594
rect 6618 25540 6624 25542
rect 6680 25540 6704 25542
rect 6760 25540 6784 25542
rect 6840 25540 6864 25542
rect 6920 25540 6926 25542
rect 6618 25531 6926 25540
rect 4308 25364 4360 25370
rect 4308 25306 4360 25312
rect 4320 24865 4348 25306
rect 5412 25160 5464 25166
rect 5412 25102 5464 25108
rect 5424 24865 5452 25102
rect 5882 25052 6190 25061
rect 5882 25050 5888 25052
rect 5944 25050 5968 25052
rect 6024 25050 6048 25052
rect 6104 25050 6128 25052
rect 6184 25050 6190 25052
rect 5944 24998 5946 25050
rect 6126 24998 6128 25050
rect 5882 24996 5888 24998
rect 5944 24996 5968 24998
rect 6024 24996 6048 24998
rect 6104 24996 6128 24998
rect 6184 24996 6190 24998
rect 5882 24987 6190 24996
rect 4306 24856 4362 24865
rect 4306 24791 4362 24800
rect 5410 24856 5466 24865
rect 5410 24791 5466 24800
rect 6618 24508 6926 24517
rect 6618 24506 6624 24508
rect 6680 24506 6704 24508
rect 6760 24506 6784 24508
rect 6840 24506 6864 24508
rect 6920 24506 6926 24508
rect 6680 24454 6682 24506
rect 6862 24454 6864 24506
rect 6618 24452 6624 24454
rect 6680 24452 6704 24454
rect 6760 24452 6784 24454
rect 6840 24452 6864 24454
rect 6920 24452 6926 24454
rect 6618 24443 6926 24452
rect 4308 24276 4360 24282
rect 4308 24218 4360 24224
rect 4320 24185 4348 24218
rect 4306 24176 4362 24185
rect 4306 24111 4362 24120
rect 8540 24140 8592 24146
rect 8540 24082 8592 24088
rect 8552 24049 8580 24082
rect 8538 24040 8594 24049
rect 8538 23975 8594 23984
rect 5882 23964 6190 23973
rect 5882 23962 5888 23964
rect 5944 23962 5968 23964
rect 6024 23962 6048 23964
rect 6104 23962 6128 23964
rect 6184 23962 6190 23964
rect 5944 23910 5946 23962
rect 6126 23910 6128 23962
rect 5882 23908 5888 23910
rect 5944 23908 5968 23910
rect 6024 23908 6048 23910
rect 6104 23908 6128 23910
rect 6184 23908 6190 23910
rect 5882 23899 6190 23908
rect 6618 23420 6926 23429
rect 6618 23418 6624 23420
rect 6680 23418 6704 23420
rect 6760 23418 6784 23420
rect 6840 23418 6864 23420
rect 6920 23418 6926 23420
rect 6680 23366 6682 23418
rect 6862 23366 6864 23418
rect 6618 23364 6624 23366
rect 6680 23364 6704 23366
rect 6760 23364 6784 23366
rect 6840 23364 6864 23366
rect 6920 23364 6926 23366
rect 6618 23355 6926 23364
rect 4308 23188 4360 23194
rect 4308 23130 4360 23136
rect 4320 22825 4348 23130
rect 8540 23052 8592 23058
rect 8540 22994 8592 23000
rect 8552 22961 8580 22994
rect 8538 22952 8594 22961
rect 8538 22887 8594 22896
rect 5882 22876 6190 22885
rect 5882 22874 5888 22876
rect 5944 22874 5968 22876
rect 6024 22874 6048 22876
rect 6104 22874 6128 22876
rect 6184 22874 6190 22876
rect 4306 22816 4362 22825
rect 5944 22822 5946 22874
rect 6126 22822 6128 22874
rect 5882 22820 5888 22822
rect 5944 22820 5968 22822
rect 6024 22820 6048 22822
rect 6104 22820 6128 22822
rect 6184 22820 6190 22822
rect 5882 22811 6190 22820
rect 4306 22751 4362 22760
rect 6618 22332 6926 22341
rect 6618 22330 6624 22332
rect 6680 22330 6704 22332
rect 6760 22330 6784 22332
rect 6840 22330 6864 22332
rect 6920 22330 6926 22332
rect 6680 22278 6682 22330
rect 6862 22278 6864 22330
rect 6618 22276 6624 22278
rect 6680 22276 6704 22278
rect 6760 22276 6784 22278
rect 6840 22276 6864 22278
rect 6920 22276 6926 22278
rect 6618 22267 6926 22276
rect 5882 21788 6190 21797
rect 5882 21786 5888 21788
rect 5944 21786 5968 21788
rect 6024 21786 6048 21788
rect 6104 21786 6128 21788
rect 6184 21786 6190 21788
rect 5944 21734 5946 21786
rect 6126 21734 6128 21786
rect 5882 21732 5888 21734
rect 5944 21732 5968 21734
rect 6024 21732 6048 21734
rect 6104 21732 6128 21734
rect 6184 21732 6190 21734
rect 5882 21723 6190 21732
rect 8538 21728 8594 21737
rect 8538 21663 8594 21672
rect 8552 21630 8580 21663
rect 8540 21624 8592 21630
rect 8540 21566 8592 21572
rect 4308 21488 4360 21494
rect 4306 21456 4308 21465
rect 4360 21456 4362 21465
rect 4306 21391 4362 21400
rect 6618 21244 6926 21253
rect 6618 21242 6624 21244
rect 6680 21242 6704 21244
rect 6760 21242 6784 21244
rect 6840 21242 6864 21244
rect 6920 21242 6926 21244
rect 6680 21190 6682 21242
rect 6862 21190 6864 21242
rect 6618 21188 6624 21190
rect 6680 21188 6704 21190
rect 6760 21188 6784 21190
rect 6840 21188 6864 21190
rect 6920 21188 6926 21190
rect 6618 21179 6926 21188
rect 5688 21080 5740 21086
rect 5688 21022 5740 21028
rect 4308 21012 4360 21018
rect 4308 20954 4360 20960
rect 4320 20785 4348 20954
rect 5700 20921 5728 21022
rect 5686 20912 5742 20921
rect 5686 20847 5742 20856
rect 4306 20776 4362 20785
rect 4306 20711 4362 20720
rect 5882 20700 6190 20709
rect 5882 20698 5888 20700
rect 5944 20698 5968 20700
rect 6024 20698 6048 20700
rect 6104 20698 6128 20700
rect 6184 20698 6190 20700
rect 5944 20646 5946 20698
rect 6126 20646 6128 20698
rect 5882 20644 5888 20646
rect 5944 20644 5968 20646
rect 6024 20644 6048 20646
rect 6104 20644 6128 20646
rect 6184 20644 6190 20646
rect 5882 20635 6190 20644
rect 6618 20156 6926 20165
rect 6618 20154 6624 20156
rect 6680 20154 6704 20156
rect 6760 20154 6784 20156
rect 6840 20154 6864 20156
rect 6920 20154 6926 20156
rect 6680 20102 6682 20154
rect 6862 20102 6864 20154
rect 6618 20100 6624 20102
rect 6680 20100 6704 20102
rect 6760 20100 6784 20102
rect 6840 20100 6864 20102
rect 6920 20100 6926 20102
rect 6618 20091 6926 20100
rect 4308 19924 4360 19930
rect 4308 19866 4360 19872
rect 4320 19425 4348 19866
rect 8540 19788 8592 19794
rect 8540 19730 8592 19736
rect 8552 19697 8580 19730
rect 8538 19688 8594 19697
rect 8538 19623 8594 19632
rect 5882 19612 6190 19621
rect 5882 19610 5888 19612
rect 5944 19610 5968 19612
rect 6024 19610 6048 19612
rect 6104 19610 6128 19612
rect 6184 19610 6190 19612
rect 5944 19558 5946 19610
rect 6126 19558 6128 19610
rect 5882 19556 5888 19558
rect 5944 19556 5968 19558
rect 6024 19556 6048 19558
rect 6104 19556 6128 19558
rect 6184 19556 6190 19558
rect 5882 19547 6190 19556
rect 4306 19416 4362 19425
rect 4306 19351 4362 19360
rect 6618 19068 6926 19077
rect 6618 19066 6624 19068
rect 6680 19066 6704 19068
rect 6760 19066 6784 19068
rect 6840 19066 6864 19068
rect 6920 19066 6926 19068
rect 6680 19014 6682 19066
rect 6862 19014 6864 19066
rect 6618 19012 6624 19014
rect 6680 19012 6704 19014
rect 6760 19012 6784 19014
rect 6840 19012 6864 19014
rect 6920 19012 6926 19014
rect 6618 19003 6926 19012
rect 4308 18836 4360 18842
rect 4308 18778 4360 18784
rect 4320 18745 4348 18778
rect 4306 18736 4362 18745
rect 4306 18671 4362 18680
rect 8540 18700 8592 18706
rect 8540 18642 8592 18648
rect 8552 18609 8580 18642
rect 8538 18600 8594 18609
rect 8538 18535 8594 18544
rect 5882 18524 6190 18533
rect 5882 18522 5888 18524
rect 5944 18522 5968 18524
rect 6024 18522 6048 18524
rect 6104 18522 6128 18524
rect 6184 18522 6190 18524
rect 5944 18470 5946 18522
rect 6126 18470 6128 18522
rect 5882 18468 5888 18470
rect 5944 18468 5968 18470
rect 6024 18468 6048 18470
rect 6104 18468 6128 18470
rect 6184 18468 6190 18470
rect 5882 18459 6190 18468
rect 6618 17980 6926 17989
rect 6618 17978 6624 17980
rect 6680 17978 6704 17980
rect 6760 17978 6784 17980
rect 6840 17978 6864 17980
rect 6920 17978 6926 17980
rect 6680 17926 6682 17978
rect 6862 17926 6864 17978
rect 6618 17924 6624 17926
rect 6680 17924 6704 17926
rect 6760 17924 6784 17926
rect 6840 17924 6864 17926
rect 6920 17924 6926 17926
rect 6618 17915 6926 17924
rect 4308 17748 4360 17754
rect 4308 17690 4360 17696
rect 4320 17385 4348 17690
rect 8540 17612 8592 17618
rect 8540 17554 8592 17560
rect 8552 17521 8580 17554
rect 8538 17512 8594 17521
rect 8538 17447 8594 17456
rect 5882 17436 6190 17445
rect 5882 17434 5888 17436
rect 5944 17434 5968 17436
rect 6024 17434 6048 17436
rect 6104 17434 6128 17436
rect 6184 17434 6190 17436
rect 4306 17376 4362 17385
rect 5944 17382 5946 17434
rect 6126 17382 6128 17434
rect 5882 17380 5888 17382
rect 5944 17380 5968 17382
rect 6024 17380 6048 17382
rect 6104 17380 6128 17382
rect 6184 17380 6190 17382
rect 5882 17371 6190 17380
rect 4306 17311 4362 17320
rect 6618 16892 6926 16901
rect 6618 16890 6624 16892
rect 6680 16890 6704 16892
rect 6760 16890 6784 16892
rect 6840 16890 6864 16892
rect 6920 16890 6926 16892
rect 6680 16838 6682 16890
rect 6862 16838 6864 16890
rect 6618 16836 6624 16838
rect 6680 16836 6704 16838
rect 6760 16836 6784 16838
rect 6840 16836 6864 16838
rect 6920 16836 6926 16838
rect 6618 16827 6926 16836
rect 5882 16348 6190 16357
rect 5882 16346 5888 16348
rect 5944 16346 5968 16348
rect 6024 16346 6048 16348
rect 6104 16346 6128 16348
rect 6184 16346 6190 16348
rect 5944 16294 5946 16346
rect 6126 16294 6128 16346
rect 5882 16292 5888 16294
rect 5944 16292 5968 16294
rect 6024 16292 6048 16294
rect 6104 16292 6128 16294
rect 6184 16292 6190 16294
rect 5882 16283 6190 16292
rect 8538 16288 8594 16297
rect 8538 16223 8594 16232
rect 8552 16190 8580 16223
rect 8540 16184 8592 16190
rect 8540 16126 8592 16132
rect 4308 16048 4360 16054
rect 4306 16016 4308 16025
rect 4360 16016 4362 16025
rect 4306 15951 4362 15960
rect 6618 15804 6926 15813
rect 6618 15802 6624 15804
rect 6680 15802 6704 15804
rect 6760 15802 6784 15804
rect 6840 15802 6864 15804
rect 6920 15802 6926 15804
rect 6680 15750 6682 15802
rect 6862 15750 6864 15802
rect 6618 15748 6624 15750
rect 6680 15748 6704 15750
rect 6760 15748 6784 15750
rect 6840 15748 6864 15750
rect 6920 15748 6926 15750
rect 6618 15739 6926 15748
rect 5688 15640 5740 15646
rect 5688 15582 5740 15588
rect 4308 15572 4360 15578
rect 4308 15514 4360 15520
rect 4320 15345 4348 15514
rect 4306 15336 4362 15345
rect 4306 15271 4362 15280
rect 5700 15073 5728 15582
rect 5882 15260 6190 15269
rect 5882 15258 5888 15260
rect 5944 15258 5968 15260
rect 6024 15258 6048 15260
rect 6104 15258 6128 15260
rect 6184 15258 6190 15260
rect 5944 15206 5946 15258
rect 6126 15206 6128 15258
rect 5882 15204 5888 15206
rect 5944 15204 5968 15206
rect 6024 15204 6048 15206
rect 6104 15204 6128 15206
rect 6184 15204 6190 15206
rect 5882 15195 6190 15204
rect 5686 15064 5742 15073
rect 5686 14999 5742 15008
rect 6618 14716 6926 14725
rect 6618 14714 6624 14716
rect 6680 14714 6704 14716
rect 6760 14714 6784 14716
rect 6840 14714 6864 14716
rect 6920 14714 6926 14716
rect 6680 14662 6682 14714
rect 6862 14662 6864 14714
rect 6618 14660 6624 14662
rect 6680 14660 6704 14662
rect 6760 14660 6784 14662
rect 6840 14660 6864 14662
rect 6920 14660 6926 14662
rect 6618 14651 6926 14660
rect 5882 14172 6190 14181
rect 5882 14170 5888 14172
rect 5944 14170 5968 14172
rect 6024 14170 6048 14172
rect 6104 14170 6128 14172
rect 6184 14170 6190 14172
rect 5944 14118 5946 14170
rect 6126 14118 6128 14170
rect 5882 14116 5888 14118
rect 5944 14116 5968 14118
rect 6024 14116 6048 14118
rect 6104 14116 6128 14118
rect 6184 14116 6190 14118
rect 5882 14107 6190 14116
rect 6618 13628 6926 13637
rect 6618 13626 6624 13628
rect 6680 13626 6704 13628
rect 6760 13626 6784 13628
rect 6840 13626 6864 13628
rect 6920 13626 6926 13628
rect 6680 13574 6682 13626
rect 6862 13574 6864 13626
rect 6618 13572 6624 13574
rect 6680 13572 6704 13574
rect 6760 13572 6784 13574
rect 6840 13572 6864 13574
rect 6920 13572 6926 13574
rect 6618 13563 6926 13572
rect 45904 13101 45932 49407
rect 45996 14189 46024 50495
rect 46088 48393 46116 84534
rect 46074 48384 46130 48393
rect 46074 48319 46130 48328
rect 45982 14180 46038 14189
rect 45982 14115 46038 14124
rect 5882 13084 6190 13093
rect 5882 13082 5888 13084
rect 5944 13082 5968 13084
rect 6024 13082 6048 13084
rect 6104 13082 6128 13084
rect 6184 13082 6190 13084
rect 5944 13030 5946 13082
rect 6126 13030 6128 13082
rect 5882 13028 5888 13030
rect 5944 13028 5968 13030
rect 6024 13028 6048 13030
rect 6104 13028 6128 13030
rect 6184 13028 6190 13030
rect 5882 13019 6190 13028
rect 45890 13092 45946 13101
rect 45890 13027 45946 13036
rect 6618 12540 6926 12549
rect 6618 12538 6624 12540
rect 6680 12538 6704 12540
rect 6760 12538 6784 12540
rect 6840 12538 6864 12540
rect 6920 12538 6926 12540
rect 6680 12486 6682 12538
rect 6862 12486 6864 12538
rect 6618 12484 6624 12486
rect 6680 12484 6704 12486
rect 6760 12484 6784 12486
rect 6840 12484 6864 12486
rect 6920 12484 6926 12486
rect 6618 12475 6926 12484
rect 5882 11996 6190 12005
rect 5882 11994 5888 11996
rect 5944 11994 5968 11996
rect 6024 11994 6048 11996
rect 6104 11994 6128 11996
rect 6184 11994 6190 11996
rect 5944 11942 5946 11994
rect 6126 11942 6128 11994
rect 5882 11940 5888 11942
rect 5944 11940 5968 11942
rect 6024 11940 6048 11942
rect 6104 11940 6128 11942
rect 6184 11940 6190 11942
rect 5882 11931 6190 11940
rect 6618 11452 6926 11461
rect 6618 11450 6624 11452
rect 6680 11450 6704 11452
rect 6760 11450 6784 11452
rect 6840 11450 6864 11452
rect 6920 11450 6926 11452
rect 6680 11398 6682 11450
rect 6862 11398 6864 11450
rect 6618 11396 6624 11398
rect 6680 11396 6704 11398
rect 6760 11396 6784 11398
rect 6840 11396 6864 11398
rect 6920 11396 6926 11398
rect 6618 11387 6926 11396
rect 5882 10908 6190 10917
rect 5882 10906 5888 10908
rect 5944 10906 5968 10908
rect 6024 10906 6048 10908
rect 6104 10906 6128 10908
rect 6184 10906 6190 10908
rect 5944 10854 5946 10906
rect 6126 10854 6128 10906
rect 5882 10852 5888 10854
rect 5944 10852 5968 10854
rect 6024 10852 6048 10854
rect 6104 10852 6128 10854
rect 6184 10852 6190 10854
rect 5882 10843 6190 10852
rect 6618 10364 6926 10373
rect 6618 10362 6624 10364
rect 6680 10362 6704 10364
rect 6760 10362 6784 10364
rect 6840 10362 6864 10364
rect 6920 10362 6926 10364
rect 6680 10310 6682 10362
rect 6862 10310 6864 10362
rect 6618 10308 6624 10310
rect 6680 10308 6704 10310
rect 6760 10308 6784 10310
rect 6840 10308 6864 10310
rect 6920 10308 6926 10310
rect 6618 10299 6926 10308
rect 45708 10200 45760 10206
rect 45430 10168 45486 10177
rect 5882 9820 6190 9829
rect 5882 9818 5888 9820
rect 5944 9818 5968 9820
rect 6024 9818 6048 9820
rect 6104 9818 6128 9820
rect 6184 9818 6190 9820
rect 5944 9766 5946 9818
rect 6126 9766 6128 9818
rect 5882 9764 5888 9766
rect 5944 9764 5968 9766
rect 6024 9764 6048 9766
rect 6104 9764 6128 9766
rect 6184 9764 6190 9766
rect 5882 9755 6190 9764
rect 6618 9276 6926 9285
rect 6618 9274 6624 9276
rect 6680 9274 6704 9276
rect 6760 9274 6784 9276
rect 6840 9274 6864 9276
rect 6920 9274 6926 9276
rect 6680 9222 6682 9274
rect 6862 9222 6864 9274
rect 6618 9220 6624 9222
rect 6680 9220 6704 9222
rect 6760 9220 6784 9222
rect 6840 9220 6864 9222
rect 6920 9220 6926 9222
rect 6618 9211 6926 9220
rect 5882 8732 6190 8741
rect 5882 8730 5888 8732
rect 5944 8730 5968 8732
rect 6024 8730 6048 8732
rect 6104 8730 6128 8732
rect 6184 8730 6190 8732
rect 5944 8678 5946 8730
rect 6126 8678 6128 8730
rect 5882 8676 5888 8678
rect 5944 8676 5968 8678
rect 6024 8676 6048 8678
rect 6104 8676 6128 8678
rect 6184 8676 6190 8678
rect 5882 8667 6190 8676
rect 6618 8188 6926 8197
rect 6618 8186 6624 8188
rect 6680 8186 6704 8188
rect 6760 8186 6784 8188
rect 6840 8186 6864 8188
rect 6920 8186 6926 8188
rect 6680 8134 6682 8186
rect 6862 8134 6864 8186
rect 6618 8132 6624 8134
rect 6680 8132 6704 8134
rect 6760 8132 6784 8134
rect 6840 8132 6864 8134
rect 6920 8132 6926 8134
rect 6618 8123 6926 8132
rect 5882 7644 6190 7653
rect 5882 7642 5888 7644
rect 5944 7642 5968 7644
rect 6024 7642 6048 7644
rect 6104 7642 6128 7644
rect 6184 7642 6190 7644
rect 5944 7590 5946 7642
rect 6126 7590 6128 7642
rect 5882 7588 5888 7590
rect 5944 7588 5968 7590
rect 6024 7588 6048 7590
rect 6104 7588 6128 7590
rect 6184 7588 6190 7590
rect 5882 7579 6190 7588
rect 6618 7100 6926 7109
rect 6618 7098 6624 7100
rect 6680 7098 6704 7100
rect 6760 7098 6784 7100
rect 6840 7098 6864 7100
rect 6920 7098 6926 7100
rect 6680 7046 6682 7098
rect 6862 7046 6864 7098
rect 6618 7044 6624 7046
rect 6680 7044 6704 7046
rect 6760 7044 6784 7046
rect 6840 7044 6864 7046
rect 6920 7044 6926 7046
rect 6618 7035 6926 7044
rect 14992 5174 15020 10140
rect 16110 10126 16216 10154
rect 16188 5174 16216 10126
rect 17200 5174 17228 10140
rect 17722 7644 18030 7653
rect 17722 7642 17728 7644
rect 17784 7642 17808 7644
rect 17864 7642 17888 7644
rect 17944 7642 17968 7644
rect 18024 7642 18030 7644
rect 17784 7590 17786 7642
rect 17966 7590 17968 7642
rect 17722 7588 17728 7590
rect 17784 7588 17808 7590
rect 17864 7588 17888 7590
rect 17944 7588 17968 7590
rect 18024 7588 18030 7590
rect 17722 7579 18030 7588
rect 17722 6556 18030 6565
rect 17722 6554 17728 6556
rect 17784 6554 17808 6556
rect 17864 6554 17888 6556
rect 17944 6554 17968 6556
rect 18024 6554 18030 6556
rect 17784 6502 17786 6554
rect 17966 6502 17968 6554
rect 17722 6500 17728 6502
rect 17784 6500 17808 6502
rect 17864 6500 17888 6502
rect 17944 6500 17968 6502
rect 18024 6500 18030 6502
rect 17722 6491 18030 6500
rect 17722 5468 18030 5477
rect 17722 5466 17728 5468
rect 17784 5466 17808 5468
rect 17864 5466 17888 5468
rect 17944 5466 17968 5468
rect 18024 5466 18030 5468
rect 17784 5414 17786 5466
rect 17966 5414 17968 5466
rect 17722 5412 17728 5414
rect 17784 5412 17808 5414
rect 17864 5412 17888 5414
rect 17944 5412 17968 5414
rect 18024 5412 18030 5414
rect 17722 5403 18030 5412
rect 18304 5174 18332 10140
rect 18382 7100 18690 7109
rect 18382 7098 18388 7100
rect 18444 7098 18468 7100
rect 18524 7098 18548 7100
rect 18604 7098 18628 7100
rect 18684 7098 18690 7100
rect 18444 7046 18446 7098
rect 18626 7046 18628 7098
rect 18382 7044 18388 7046
rect 18444 7044 18468 7046
rect 18524 7044 18548 7046
rect 18604 7044 18628 7046
rect 18684 7044 18690 7046
rect 18382 7035 18690 7044
rect 18382 6012 18690 6021
rect 18382 6010 18388 6012
rect 18444 6010 18468 6012
rect 18524 6010 18548 6012
rect 18604 6010 18628 6012
rect 18684 6010 18690 6012
rect 18444 5958 18446 6010
rect 18626 5958 18628 6010
rect 18382 5956 18388 5958
rect 18444 5956 18468 5958
rect 18524 5956 18548 5958
rect 18604 5956 18628 5958
rect 18684 5956 18690 5958
rect 18382 5947 18690 5956
rect 19408 5174 19436 10140
rect 20512 5174 20540 10140
rect 21616 5174 21644 10140
rect 22720 5174 22748 10140
rect 23838 10126 23944 10154
rect 23916 5174 23944 10126
rect 24928 5174 24956 10140
rect 26032 5174 26060 10140
rect 27136 5174 27164 10140
rect 28240 5174 28268 10140
rect 29344 5174 29372 10140
rect 30448 5310 30476 10140
rect 31552 5310 31580 10140
rect 32656 5310 32684 10140
rect 33760 5310 33788 10140
rect 34864 5310 34892 10140
rect 35968 5310 35996 10140
rect 37086 10126 37192 10154
rect 36122 7644 36430 7653
rect 36122 7642 36128 7644
rect 36184 7642 36208 7644
rect 36264 7642 36288 7644
rect 36344 7642 36368 7644
rect 36424 7642 36430 7644
rect 36184 7590 36186 7642
rect 36366 7590 36368 7642
rect 36122 7588 36128 7590
rect 36184 7588 36208 7590
rect 36264 7588 36288 7590
rect 36344 7588 36368 7590
rect 36424 7588 36430 7590
rect 36122 7579 36430 7588
rect 36782 7100 37090 7109
rect 36782 7098 36788 7100
rect 36844 7098 36868 7100
rect 36924 7098 36948 7100
rect 37004 7098 37028 7100
rect 37084 7098 37090 7100
rect 36844 7046 36846 7098
rect 37026 7046 37028 7098
rect 36782 7044 36788 7046
rect 36844 7044 36868 7046
rect 36924 7044 36948 7046
rect 37004 7044 37028 7046
rect 37084 7044 37090 7046
rect 36782 7035 37090 7044
rect 36122 6556 36430 6565
rect 36122 6554 36128 6556
rect 36184 6554 36208 6556
rect 36264 6554 36288 6556
rect 36344 6554 36368 6556
rect 36424 6554 36430 6556
rect 36184 6502 36186 6554
rect 36366 6502 36368 6554
rect 36122 6500 36128 6502
rect 36184 6500 36208 6502
rect 36264 6500 36288 6502
rect 36344 6500 36368 6502
rect 36424 6500 36430 6502
rect 36122 6491 36430 6500
rect 36782 6012 37090 6021
rect 36782 6010 36788 6012
rect 36844 6010 36868 6012
rect 36924 6010 36948 6012
rect 37004 6010 37028 6012
rect 37084 6010 37090 6012
rect 36844 5958 36846 6010
rect 37026 5958 37028 6010
rect 36782 5956 36788 5958
rect 36844 5956 36868 5958
rect 36924 5956 36948 5958
rect 37004 5956 37028 5958
rect 37084 5956 37090 5958
rect 36782 5947 37090 5956
rect 36122 5468 36430 5477
rect 36122 5466 36128 5468
rect 36184 5466 36208 5468
rect 36264 5466 36288 5468
rect 36344 5466 36368 5468
rect 36424 5466 36430 5468
rect 36184 5414 36186 5466
rect 36366 5414 36368 5466
rect 36122 5412 36128 5414
rect 36184 5412 36208 5414
rect 36264 5412 36288 5414
rect 36344 5412 36368 5414
rect 36424 5412 36430 5414
rect 36122 5403 36430 5412
rect 37164 5310 37192 10126
rect 38176 5310 38204 10140
rect 39280 5310 39308 10140
rect 40384 5310 40412 10140
rect 41488 5310 41516 10140
rect 42592 5310 42620 10140
rect 43696 5310 43724 10140
rect 44800 5310 44828 10140
rect 45708 10142 45760 10148
rect 45430 10103 45486 10112
rect 45444 7486 45472 10103
rect 45720 7486 45748 10142
rect 45904 7486 45932 13027
rect 45996 7486 46024 14115
rect 46088 12013 46116 48319
rect 46180 47305 46208 84670
rect 46166 47296 46222 47305
rect 46166 47231 46222 47240
rect 47008 46042 47036 86574
rect 50320 84734 50348 86574
rect 50308 84728 50360 84734
rect 50308 84670 50360 84676
rect 49112 84660 49164 84666
rect 49112 84602 49164 84608
rect 49124 84462 49152 84602
rect 48008 84456 48060 84462
rect 48008 84398 48060 84404
rect 49112 84456 49164 84462
rect 49112 84398 49164 84404
rect 48020 82370 48048 84398
rect 49124 82370 49152 84398
rect 50320 82370 50348 84670
rect 51320 84660 51372 84666
rect 51320 84602 51372 84608
rect 51332 84462 51360 84602
rect 51320 84456 51372 84462
rect 51320 84398 51372 84404
rect 51332 82370 51360 84398
rect 47974 82342 48048 82370
rect 49078 82342 49152 82370
rect 50182 82342 50348 82370
rect 51286 82342 51360 82370
rect 52896 82354 52924 87186
rect 53540 82370 53568 87186
rect 52378 82348 52430 82354
rect 47974 81713 48002 82342
rect 49078 82084 49106 82342
rect 50182 82084 50210 82342
rect 51286 82084 51314 82342
rect 52378 82290 52430 82296
rect 52884 82348 52936 82354
rect 52884 82290 52936 82296
rect 53494 82342 53568 82370
rect 54460 82370 54488 87186
rect 54522 87068 54830 87077
rect 54522 87066 54528 87068
rect 54584 87066 54608 87068
rect 54664 87066 54688 87068
rect 54744 87066 54768 87068
rect 54824 87066 54830 87068
rect 54584 87014 54586 87066
rect 54766 87014 54768 87066
rect 54522 87012 54528 87014
rect 54584 87012 54608 87014
rect 54664 87012 54688 87014
rect 54744 87012 54768 87014
rect 54824 87012 54830 87014
rect 54522 87003 54830 87012
rect 55182 86524 55490 86533
rect 55182 86522 55188 86524
rect 55244 86522 55268 86524
rect 55324 86522 55348 86524
rect 55404 86522 55428 86524
rect 55484 86522 55490 86524
rect 55244 86470 55246 86522
rect 55426 86470 55428 86522
rect 55182 86468 55188 86470
rect 55244 86468 55268 86470
rect 55324 86468 55348 86470
rect 55404 86468 55428 86470
rect 55484 86468 55490 86470
rect 55182 86459 55490 86468
rect 54522 85980 54830 85989
rect 54522 85978 54528 85980
rect 54584 85978 54608 85980
rect 54664 85978 54688 85980
rect 54744 85978 54768 85980
rect 54824 85978 54830 85980
rect 54584 85926 54586 85978
rect 54766 85926 54768 85978
rect 54522 85924 54528 85926
rect 54584 85924 54608 85926
rect 54664 85924 54688 85926
rect 54744 85924 54768 85926
rect 54824 85924 54830 85926
rect 54522 85915 54830 85924
rect 55182 85436 55490 85445
rect 55182 85434 55188 85436
rect 55244 85434 55268 85436
rect 55324 85434 55348 85436
rect 55404 85434 55428 85436
rect 55484 85434 55490 85436
rect 55244 85382 55246 85434
rect 55426 85382 55428 85434
rect 55182 85380 55188 85382
rect 55244 85380 55268 85382
rect 55324 85380 55348 85382
rect 55404 85380 55428 85382
rect 55484 85380 55490 85382
rect 55182 85371 55490 85380
rect 54522 84892 54830 84901
rect 54522 84890 54528 84892
rect 54584 84890 54608 84892
rect 54664 84890 54688 84892
rect 54744 84890 54768 84892
rect 54824 84890 54830 84892
rect 54584 84838 54586 84890
rect 54766 84838 54768 84890
rect 54522 84836 54528 84838
rect 54584 84836 54608 84838
rect 54664 84836 54688 84838
rect 54744 84836 54768 84838
rect 54824 84836 54830 84838
rect 54522 84827 54830 84836
rect 55182 84348 55490 84357
rect 55182 84346 55188 84348
rect 55244 84346 55268 84348
rect 55324 84346 55348 84348
rect 55404 84346 55428 84348
rect 55484 84346 55490 84348
rect 55244 84294 55246 84346
rect 55426 84294 55428 84346
rect 55182 84292 55188 84294
rect 55244 84292 55268 84294
rect 55324 84292 55348 84294
rect 55404 84292 55428 84294
rect 55484 84292 55490 84294
rect 55182 84283 55490 84292
rect 55748 82370 55776 87186
rect 56852 82370 56880 87186
rect 57956 82370 57984 87186
rect 59060 82370 59088 87186
rect 60164 82370 60192 87186
rect 54460 82342 54626 82370
rect 52390 82084 52418 82290
rect 53494 82084 53522 82342
rect 54598 82084 54626 82342
rect 55702 82342 55776 82370
rect 56806 82342 56880 82370
rect 57910 82342 57984 82370
rect 59014 82342 59088 82370
rect 60118 82342 60192 82370
rect 61176 82370 61204 87186
rect 62372 87166 62492 87186
rect 62372 82370 62400 87166
rect 63476 82370 63504 87186
rect 64580 82370 64608 87186
rect 65684 82370 65712 87186
rect 66788 82370 66816 87186
rect 67892 82370 67920 87322
rect 68076 87250 68104 88000
rect 68720 87454 68748 88000
rect 70008 87538 70036 88000
rect 70008 87510 70128 87538
rect 68708 87448 68760 87454
rect 68708 87390 68760 87396
rect 68984 87380 69036 87386
rect 68984 87322 69036 87328
rect 69996 87380 70048 87386
rect 69996 87322 70048 87328
rect 68064 87244 68116 87250
rect 68064 87186 68116 87192
rect 68996 82370 69024 87322
rect 61176 82342 61250 82370
rect 55702 82084 55730 82342
rect 56806 82084 56834 82342
rect 57910 82084 57938 82342
rect 59014 82084 59042 82342
rect 60118 82084 60146 82342
rect 61222 82084 61250 82342
rect 62326 82342 62400 82370
rect 63430 82342 63504 82370
rect 64534 82342 64608 82370
rect 65638 82342 65712 82370
rect 66742 82342 66816 82370
rect 67846 82342 67920 82370
rect 68950 82342 69024 82370
rect 70008 82370 70036 87322
rect 70100 87250 70128 87510
rect 71192 87380 71244 87386
rect 71192 87322 71244 87328
rect 70088 87244 70140 87250
rect 70088 87186 70140 87192
rect 71204 82370 71232 87322
rect 71296 87250 71324 88000
rect 72296 87380 72348 87386
rect 72296 87322 72348 87328
rect 71284 87244 71336 87250
rect 71284 87186 71336 87192
rect 72308 82370 72336 87322
rect 72584 87250 72612 88000
rect 73228 87250 73256 88000
rect 73582 87612 73890 87621
rect 73582 87610 73588 87612
rect 73644 87610 73668 87612
rect 73724 87610 73748 87612
rect 73804 87610 73828 87612
rect 73884 87610 73890 87612
rect 73644 87558 73646 87610
rect 73826 87558 73828 87610
rect 73582 87556 73588 87558
rect 73644 87556 73668 87558
rect 73724 87556 73748 87558
rect 73804 87556 73828 87558
rect 73884 87556 73890 87558
rect 73582 87547 73890 87556
rect 74516 87538 74544 88000
rect 74516 87510 74636 87538
rect 73400 87380 73452 87386
rect 73400 87322 73452 87328
rect 74504 87380 74556 87386
rect 74504 87322 74556 87328
rect 72572 87244 72624 87250
rect 72572 87186 72624 87192
rect 73216 87244 73268 87250
rect 73216 87186 73268 87192
rect 72922 87068 73230 87077
rect 72922 87066 72928 87068
rect 72984 87066 73008 87068
rect 73064 87066 73088 87068
rect 73144 87066 73168 87068
rect 73224 87066 73230 87068
rect 72984 87014 72986 87066
rect 73166 87014 73168 87066
rect 72922 87012 72928 87014
rect 72984 87012 73008 87014
rect 73064 87012 73088 87014
rect 73144 87012 73168 87014
rect 73224 87012 73230 87014
rect 72922 87003 73230 87012
rect 72922 85980 73230 85989
rect 72922 85978 72928 85980
rect 72984 85978 73008 85980
rect 73064 85978 73088 85980
rect 73144 85978 73168 85980
rect 73224 85978 73230 85980
rect 72984 85926 72986 85978
rect 73166 85926 73168 85978
rect 72922 85924 72928 85926
rect 72984 85924 73008 85926
rect 73064 85924 73088 85926
rect 73144 85924 73168 85926
rect 73224 85924 73230 85926
rect 72922 85915 73230 85924
rect 72922 84892 73230 84901
rect 72922 84890 72928 84892
rect 72984 84890 73008 84892
rect 73064 84890 73088 84892
rect 73144 84890 73168 84892
rect 73224 84890 73230 84892
rect 72984 84838 72986 84890
rect 73166 84838 73168 84890
rect 72922 84836 72928 84838
rect 72984 84836 73008 84838
rect 73064 84836 73088 84838
rect 73144 84836 73168 84838
rect 73224 84836 73230 84838
rect 72922 84827 73230 84836
rect 73412 82370 73440 87322
rect 73582 86524 73890 86533
rect 73582 86522 73588 86524
rect 73644 86522 73668 86524
rect 73724 86522 73748 86524
rect 73804 86522 73828 86524
rect 73884 86522 73890 86524
rect 73644 86470 73646 86522
rect 73826 86470 73828 86522
rect 73582 86468 73588 86470
rect 73644 86468 73668 86470
rect 73724 86468 73748 86470
rect 73804 86468 73828 86470
rect 73884 86468 73890 86470
rect 73582 86459 73890 86468
rect 73582 85436 73890 85445
rect 73582 85434 73588 85436
rect 73644 85434 73668 85436
rect 73724 85434 73748 85436
rect 73804 85434 73828 85436
rect 73884 85434 73890 85436
rect 73644 85382 73646 85434
rect 73826 85382 73828 85434
rect 73582 85380 73588 85382
rect 73644 85380 73668 85382
rect 73724 85380 73748 85382
rect 73804 85380 73828 85382
rect 73884 85380 73890 85382
rect 73582 85371 73890 85380
rect 73582 84348 73890 84357
rect 73582 84346 73588 84348
rect 73644 84346 73668 84348
rect 73724 84346 73748 84348
rect 73804 84346 73828 84348
rect 73884 84346 73890 84348
rect 73644 84294 73646 84346
rect 73826 84294 73828 84346
rect 73582 84292 73588 84294
rect 73644 84292 73668 84294
rect 73724 84292 73748 84294
rect 73804 84292 73828 84294
rect 73884 84292 73890 84294
rect 73582 84283 73890 84292
rect 74516 82370 74544 87322
rect 74608 87250 74636 87510
rect 75608 87380 75660 87386
rect 75608 87322 75660 87328
rect 74596 87244 74648 87250
rect 74596 87186 74648 87192
rect 75620 82370 75648 87322
rect 75804 87250 75832 88000
rect 76448 87454 76476 88000
rect 77736 87538 77764 88000
rect 77736 87510 77856 87538
rect 76436 87448 76488 87454
rect 76436 87390 76488 87396
rect 76712 87380 76764 87386
rect 76712 87322 76764 87328
rect 77724 87380 77776 87386
rect 77724 87322 77776 87328
rect 75792 87244 75844 87250
rect 75792 87186 75844 87192
rect 76724 82370 76752 87322
rect 70008 82342 70082 82370
rect 62326 82084 62354 82342
rect 63430 82084 63458 82342
rect 64534 82084 64562 82342
rect 65638 82084 65666 82342
rect 66742 82084 66770 82342
rect 67846 82084 67874 82342
rect 68950 82084 68978 82342
rect 70054 82084 70082 82342
rect 71158 82342 71232 82370
rect 72262 82342 72336 82370
rect 73366 82342 73440 82370
rect 74470 82342 74544 82370
rect 75574 82342 75648 82370
rect 76678 82342 76752 82370
rect 77736 82370 77764 87322
rect 77828 87250 77856 87510
rect 78920 87380 78972 87386
rect 78920 87322 78972 87328
rect 77816 87244 77868 87250
rect 77816 87186 77868 87192
rect 78932 82370 78960 87322
rect 79024 87250 79052 88000
rect 80312 87250 80340 88000
rect 80392 87380 80444 87386
rect 80392 87322 80444 87328
rect 79012 87244 79064 87250
rect 79012 87186 79064 87192
rect 80300 87244 80352 87250
rect 80300 87186 80352 87192
rect 77736 82342 77810 82370
rect 71158 82084 71186 82342
rect 72262 82084 72290 82342
rect 73366 82084 73394 82342
rect 74470 82084 74498 82342
rect 75574 82084 75602 82342
rect 76678 82084 76706 82342
rect 77782 82084 77810 82342
rect 78886 82342 78960 82370
rect 80404 82354 80432 87322
rect 80956 87250 80984 88000
rect 82244 87538 82272 88000
rect 82244 87510 82364 87538
rect 81128 87380 81180 87386
rect 81128 87322 81180 87328
rect 82232 87380 82284 87386
rect 82232 87322 82284 87328
rect 80944 87244 80996 87250
rect 80944 87186 80996 87192
rect 81140 82370 81168 87322
rect 82244 82370 82272 87322
rect 82336 87250 82364 87510
rect 82324 87244 82376 87250
rect 82324 87186 82376 87192
rect 86474 84892 86782 84901
rect 86474 84890 86480 84892
rect 86536 84890 86560 84892
rect 86616 84890 86640 84892
rect 86696 84890 86720 84892
rect 86776 84890 86782 84892
rect 86536 84838 86538 84890
rect 86718 84838 86720 84890
rect 86474 84836 86480 84838
rect 86536 84836 86560 84838
rect 86616 84836 86640 84838
rect 86696 84836 86720 84838
rect 86776 84836 86782 84838
rect 86474 84827 86782 84836
rect 87210 84348 87518 84357
rect 87210 84346 87216 84348
rect 87272 84346 87296 84348
rect 87352 84346 87376 84348
rect 87432 84346 87456 84348
rect 87512 84346 87518 84348
rect 87272 84294 87274 84346
rect 87454 84294 87456 84346
rect 87210 84292 87216 84294
rect 87272 84292 87296 84294
rect 87352 84292 87376 84294
rect 87432 84292 87456 84294
rect 87512 84292 87518 84294
rect 87210 84283 87518 84292
rect 86474 83804 86782 83813
rect 86474 83802 86480 83804
rect 86536 83802 86560 83804
rect 86616 83802 86640 83804
rect 86696 83802 86720 83804
rect 86776 83802 86782 83804
rect 86536 83750 86538 83802
rect 86718 83750 86720 83802
rect 86474 83748 86480 83750
rect 86536 83748 86560 83750
rect 86616 83748 86640 83750
rect 86696 83748 86720 83750
rect 86776 83748 86782 83750
rect 86474 83739 86782 83748
rect 87210 83260 87518 83269
rect 87210 83258 87216 83260
rect 87272 83258 87296 83260
rect 87352 83258 87376 83260
rect 87432 83258 87456 83260
rect 87512 83258 87518 83260
rect 87272 83206 87274 83258
rect 87454 83206 87456 83258
rect 87210 83204 87216 83206
rect 87272 83204 87296 83206
rect 87352 83204 87376 83206
rect 87432 83204 87456 83206
rect 87512 83204 87518 83206
rect 87210 83195 87518 83204
rect 83244 83164 83296 83170
rect 83244 83106 83296 83112
rect 79978 82348 80030 82354
rect 78886 82084 78914 82342
rect 79978 82290 80030 82296
rect 80392 82348 80444 82354
rect 80392 82290 80444 82296
rect 81094 82342 81168 82370
rect 82198 82342 82272 82370
rect 79990 82084 80018 82290
rect 81094 82084 81122 82342
rect 82198 82084 82226 82342
rect 47086 81704 47142 81713
rect 47086 81639 47142 81648
rect 47960 81704 48016 81713
rect 47960 81639 48016 81648
rect 46996 46036 47048 46042
rect 46996 45978 47048 45984
rect 46444 45900 46496 45906
rect 46444 45842 46496 45848
rect 46074 12004 46130 12013
rect 46074 11939 46130 11948
rect 46088 10206 46116 11939
rect 46456 10993 46484 45842
rect 47100 45673 47128 81639
rect 50170 45968 50222 45974
rect 49064 45936 49120 45945
rect 51136 45968 51188 45974
rect 50170 45910 50222 45916
rect 51134 45936 51136 45945
rect 51188 45936 51190 45945
rect 49064 45871 49120 45880
rect 49078 45772 49106 45871
rect 50182 45772 50210 45910
rect 51134 45871 51190 45880
rect 51274 45900 51326 45906
rect 51274 45842 51326 45848
rect 51286 45772 51314 45842
rect 52390 45772 52418 46452
rect 53494 45772 53522 46452
rect 54598 45772 54626 46452
rect 55702 45772 55730 46452
rect 56806 45772 56834 46452
rect 57910 45772 57938 46452
rect 59014 45772 59042 46452
rect 60118 45772 60146 46452
rect 61222 45772 61250 46452
rect 62326 45772 62354 46452
rect 63430 45772 63458 46452
rect 64534 45772 64562 46452
rect 65638 45772 65666 46452
rect 66742 45772 66770 46452
rect 67846 45772 67874 46452
rect 68950 45772 68978 46452
rect 70054 45772 70082 46452
rect 71158 45772 71186 46452
rect 72262 45772 72290 46452
rect 73366 45772 73394 46452
rect 74470 45772 74498 46452
rect 75574 45772 75602 46452
rect 76678 45772 76706 46452
rect 77782 45772 77810 46452
rect 78886 45772 78914 46452
rect 79990 45772 80018 46452
rect 81094 45772 81122 46452
rect 82198 45772 82226 46452
rect 47086 45664 47142 45673
rect 47086 45599 47142 45608
rect 47960 45664 48016 45673
rect 47960 45599 48016 45608
rect 83256 11294 83284 83106
rect 86474 82716 86782 82725
rect 86474 82714 86480 82716
rect 86536 82714 86560 82716
rect 86616 82714 86640 82716
rect 86696 82714 86720 82716
rect 86776 82714 86782 82716
rect 86536 82662 86538 82714
rect 86718 82662 86720 82714
rect 86474 82660 86480 82662
rect 86536 82660 86560 82662
rect 86616 82660 86640 82662
rect 86696 82660 86720 82662
rect 86776 82660 86782 82662
rect 86474 82651 86782 82660
rect 87210 82172 87518 82181
rect 87210 82170 87216 82172
rect 87272 82170 87296 82172
rect 87352 82170 87376 82172
rect 87432 82170 87456 82172
rect 87512 82170 87518 82172
rect 87272 82118 87274 82170
rect 87454 82118 87456 82170
rect 87210 82116 87216 82118
rect 87272 82116 87296 82118
rect 87352 82116 87376 82118
rect 87432 82116 87456 82118
rect 87512 82116 87518 82118
rect 87210 82107 87518 82116
rect 86474 81628 86782 81637
rect 86474 81626 86480 81628
rect 86536 81626 86560 81628
rect 86616 81626 86640 81628
rect 86696 81626 86720 81628
rect 86776 81626 86782 81628
rect 86536 81574 86538 81626
rect 86718 81574 86720 81626
rect 86474 81572 86480 81574
rect 86536 81572 86560 81574
rect 86616 81572 86640 81574
rect 86696 81572 86720 81574
rect 86776 81572 86782 81574
rect 86474 81563 86782 81572
rect 88212 81328 88264 81334
rect 88210 81296 88212 81305
rect 88264 81296 88266 81305
rect 84348 81260 84400 81266
rect 88210 81231 88266 81240
rect 84348 81202 84400 81208
rect 84360 81033 84388 81202
rect 87210 81084 87518 81093
rect 87210 81082 87216 81084
rect 87272 81082 87296 81084
rect 87352 81082 87376 81084
rect 87432 81082 87456 81084
rect 87512 81082 87518 81084
rect 84346 81024 84402 81033
rect 87272 81030 87274 81082
rect 87454 81030 87456 81082
rect 87210 81028 87216 81030
rect 87272 81028 87296 81030
rect 87352 81028 87376 81030
rect 87432 81028 87456 81030
rect 87512 81028 87518 81030
rect 87210 81019 87518 81028
rect 84346 80959 84402 80968
rect 86474 80540 86782 80549
rect 86474 80538 86480 80540
rect 86536 80538 86560 80540
rect 86616 80538 86640 80540
rect 86696 80538 86720 80540
rect 86776 80538 86782 80540
rect 86536 80486 86538 80538
rect 86718 80486 86720 80538
rect 86474 80484 86480 80486
rect 86536 80484 86560 80486
rect 86616 80484 86640 80486
rect 86696 80484 86720 80486
rect 86776 80484 86782 80486
rect 86474 80475 86782 80484
rect 88212 80240 88264 80246
rect 88212 80182 88264 80188
rect 85820 80172 85872 80178
rect 85820 80114 85872 80120
rect 85832 79945 85860 80114
rect 87210 79996 87518 80005
rect 87210 79994 87216 79996
rect 87272 79994 87296 79996
rect 87352 79994 87376 79996
rect 87432 79994 87456 79996
rect 87512 79994 87518 79996
rect 85818 79936 85874 79945
rect 87272 79942 87274 79994
rect 87454 79942 87456 79994
rect 88224 79945 88252 80182
rect 87210 79940 87216 79942
rect 87272 79940 87296 79942
rect 87352 79940 87376 79942
rect 87432 79940 87456 79942
rect 87512 79940 87518 79942
rect 87210 79931 87518 79940
rect 88210 79936 88266 79945
rect 85818 79871 85874 79880
rect 88210 79871 88266 79880
rect 86474 79452 86782 79461
rect 86474 79450 86480 79452
rect 86536 79450 86560 79452
rect 86616 79450 86640 79452
rect 86696 79450 86720 79452
rect 86776 79450 86782 79452
rect 86536 79398 86538 79450
rect 86718 79398 86720 79450
rect 86474 79396 86480 79398
rect 86536 79396 86560 79398
rect 86616 79396 86640 79398
rect 86696 79396 86720 79398
rect 86776 79396 86782 79398
rect 86474 79387 86782 79396
rect 87210 78908 87518 78917
rect 87210 78906 87216 78908
rect 87272 78906 87296 78908
rect 87352 78906 87376 78908
rect 87432 78906 87456 78908
rect 87512 78906 87518 78908
rect 85818 78848 85874 78857
rect 87272 78854 87274 78906
rect 87454 78854 87456 78906
rect 87210 78852 87216 78854
rect 87272 78852 87296 78854
rect 87352 78852 87376 78854
rect 87432 78852 87456 78854
rect 87512 78852 87518 78854
rect 87210 78843 87518 78852
rect 85818 78783 85874 78792
rect 85832 78750 85860 78783
rect 85820 78744 85872 78750
rect 85820 78686 85872 78692
rect 88212 78676 88264 78682
rect 88212 78618 88264 78624
rect 88224 78585 88252 78618
rect 88210 78576 88266 78585
rect 88210 78511 88266 78520
rect 86474 78364 86782 78373
rect 86474 78362 86480 78364
rect 86536 78362 86560 78364
rect 86616 78362 86640 78364
rect 86696 78362 86720 78364
rect 86776 78362 86782 78364
rect 86536 78310 86538 78362
rect 86718 78310 86720 78362
rect 86474 78308 86480 78310
rect 86536 78308 86560 78310
rect 86616 78308 86640 78310
rect 86696 78308 86720 78310
rect 86776 78308 86782 78310
rect 86474 78299 86782 78308
rect 88212 78064 88264 78070
rect 88212 78006 88264 78012
rect 85820 77996 85872 78002
rect 85820 77938 85872 77944
rect 85832 77769 85860 77938
rect 88224 77905 88252 78006
rect 88210 77896 88266 77905
rect 88210 77831 88266 77840
rect 87210 77820 87518 77829
rect 87210 77818 87216 77820
rect 87272 77818 87296 77820
rect 87352 77818 87376 77820
rect 87432 77818 87456 77820
rect 87512 77818 87518 77820
rect 85818 77760 85874 77769
rect 87272 77766 87274 77818
rect 87454 77766 87456 77818
rect 87210 77764 87216 77766
rect 87272 77764 87296 77766
rect 87352 77764 87376 77766
rect 87432 77764 87456 77766
rect 87512 77764 87518 77766
rect 87210 77755 87518 77764
rect 85818 77695 85874 77704
rect 86474 77276 86782 77285
rect 86474 77274 86480 77276
rect 86536 77274 86560 77276
rect 86616 77274 86640 77276
rect 86696 77274 86720 77276
rect 86776 77274 86782 77276
rect 86536 77222 86538 77274
rect 86718 77222 86720 77274
rect 86474 77220 86480 77222
rect 86536 77220 86560 77222
rect 86616 77220 86640 77222
rect 86696 77220 86720 77222
rect 86776 77220 86782 77222
rect 86474 77211 86782 77220
rect 85820 76840 85872 76846
rect 85820 76782 85872 76788
rect 88028 76840 88080 76846
rect 88028 76782 88080 76788
rect 85832 76681 85860 76782
rect 87210 76732 87518 76741
rect 87210 76730 87216 76732
rect 87272 76730 87296 76732
rect 87352 76730 87376 76732
rect 87432 76730 87456 76732
rect 87512 76730 87518 76732
rect 85818 76672 85874 76681
rect 87272 76678 87274 76730
rect 87454 76678 87456 76730
rect 87210 76676 87216 76678
rect 87272 76676 87296 76678
rect 87352 76676 87376 76678
rect 87432 76676 87456 76678
rect 87512 76676 87518 76678
rect 87210 76667 87518 76676
rect 85818 76607 85874 76616
rect 88040 76545 88068 76782
rect 88026 76536 88082 76545
rect 88026 76471 88082 76480
rect 86474 76188 86782 76197
rect 86474 76186 86480 76188
rect 86536 76186 86560 76188
rect 86616 76186 86640 76188
rect 86696 76186 86720 76188
rect 86776 76186 86782 76188
rect 86536 76134 86538 76186
rect 86718 76134 86720 76186
rect 86474 76132 86480 76134
rect 86536 76132 86560 76134
rect 86616 76132 86640 76134
rect 86696 76132 86720 76134
rect 86776 76132 86782 76134
rect 86474 76123 86782 76132
rect 88212 75888 88264 75894
rect 88210 75856 88212 75865
rect 88264 75856 88266 75865
rect 85820 75820 85872 75826
rect 88210 75791 88266 75800
rect 85820 75762 85872 75768
rect 85832 75593 85860 75762
rect 87210 75644 87518 75653
rect 87210 75642 87216 75644
rect 87272 75642 87296 75644
rect 87352 75642 87376 75644
rect 87432 75642 87456 75644
rect 87512 75642 87518 75644
rect 85818 75584 85874 75593
rect 87272 75590 87274 75642
rect 87454 75590 87456 75642
rect 87210 75588 87216 75590
rect 87272 75588 87296 75590
rect 87352 75588 87376 75590
rect 87432 75588 87456 75590
rect 87512 75588 87518 75590
rect 87210 75579 87518 75588
rect 85818 75519 85874 75528
rect 86474 75100 86782 75109
rect 86474 75098 86480 75100
rect 86536 75098 86560 75100
rect 86616 75098 86640 75100
rect 86696 75098 86720 75100
rect 86776 75098 86782 75100
rect 86536 75046 86538 75098
rect 86718 75046 86720 75098
rect 86474 75044 86480 75046
rect 86536 75044 86560 75046
rect 86616 75044 86640 75046
rect 86696 75044 86720 75046
rect 86776 75044 86782 75046
rect 86474 75035 86782 75044
rect 84532 74800 84584 74806
rect 84532 74742 84584 74748
rect 88580 74800 88632 74806
rect 88580 74742 88632 74748
rect 84544 74505 84572 74742
rect 87210 74556 87518 74565
rect 87210 74554 87216 74556
rect 87272 74554 87296 74556
rect 87352 74554 87376 74556
rect 87432 74554 87456 74556
rect 87512 74554 87518 74556
rect 84530 74496 84586 74505
rect 87272 74502 87274 74554
rect 87454 74502 87456 74554
rect 88592 74505 88620 74742
rect 87210 74500 87216 74502
rect 87272 74500 87296 74502
rect 87352 74500 87376 74502
rect 87432 74500 87456 74502
rect 87512 74500 87518 74502
rect 87210 74491 87518 74500
rect 88578 74496 88634 74505
rect 84530 74431 84586 74440
rect 88578 74431 88634 74440
rect 86474 74012 86782 74021
rect 86474 74010 86480 74012
rect 86536 74010 86560 74012
rect 86616 74010 86640 74012
rect 86696 74010 86720 74012
rect 86776 74010 86782 74012
rect 86536 73958 86538 74010
rect 86718 73958 86720 74010
rect 86474 73956 86480 73958
rect 86536 73956 86560 73958
rect 86616 73956 86640 73958
rect 86696 73956 86720 73958
rect 86776 73956 86782 73958
rect 86474 73947 86782 73956
rect 87210 73468 87518 73477
rect 87210 73466 87216 73468
rect 87272 73466 87296 73468
rect 87352 73466 87376 73468
rect 87432 73466 87456 73468
rect 87512 73466 87518 73468
rect 84806 73408 84862 73417
rect 87272 73414 87274 73466
rect 87454 73414 87456 73466
rect 87210 73412 87216 73414
rect 87272 73412 87296 73414
rect 87352 73412 87376 73414
rect 87432 73412 87456 73414
rect 87512 73412 87518 73414
rect 87210 73403 87518 73412
rect 84806 73343 84862 73352
rect 84820 73310 84848 73343
rect 84808 73304 84860 73310
rect 84808 73246 84860 73252
rect 88212 73236 88264 73242
rect 88212 73178 88264 73184
rect 88224 73145 88252 73178
rect 88210 73136 88266 73145
rect 88210 73071 88266 73080
rect 86474 72924 86782 72933
rect 86474 72922 86480 72924
rect 86536 72922 86560 72924
rect 86616 72922 86640 72924
rect 86696 72922 86720 72924
rect 86776 72922 86782 72924
rect 86536 72870 86538 72922
rect 86718 72870 86720 72922
rect 86474 72868 86480 72870
rect 86536 72868 86560 72870
rect 86616 72868 86640 72870
rect 86696 72868 86720 72870
rect 86776 72868 86782 72870
rect 86474 72859 86782 72868
rect 88212 72624 88264 72630
rect 88212 72566 88264 72572
rect 87844 72488 87896 72494
rect 88224 72465 88252 72566
rect 87844 72430 87896 72436
rect 88210 72456 88266 72465
rect 87210 72380 87518 72389
rect 87210 72378 87216 72380
rect 87272 72378 87296 72380
rect 87352 72378 87376 72380
rect 87432 72378 87456 72380
rect 87512 72378 87518 72380
rect 87272 72326 87274 72378
rect 87454 72326 87456 72378
rect 87210 72324 87216 72326
rect 87272 72324 87296 72326
rect 87352 72324 87376 72326
rect 87432 72324 87456 72326
rect 87512 72324 87518 72326
rect 87210 72315 87518 72324
rect 87856 72193 87884 72430
rect 88210 72391 88266 72400
rect 87842 72184 87898 72193
rect 87842 72119 87898 72128
rect 86474 71836 86782 71845
rect 86474 71834 86480 71836
rect 86536 71834 86560 71836
rect 86616 71834 86640 71836
rect 86696 71834 86720 71836
rect 86776 71834 86782 71836
rect 86536 71782 86538 71834
rect 86718 71782 86720 71834
rect 86474 71780 86480 71782
rect 86536 71780 86560 71782
rect 86616 71780 86640 71782
rect 86696 71780 86720 71782
rect 86776 71780 86782 71782
rect 86474 71771 86782 71780
rect 88212 71536 88264 71542
rect 88212 71478 88264 71484
rect 85820 71468 85872 71474
rect 85820 71410 85872 71416
rect 85832 71241 85860 71410
rect 87210 71292 87518 71301
rect 87210 71290 87216 71292
rect 87272 71290 87296 71292
rect 87352 71290 87376 71292
rect 87432 71290 87456 71292
rect 87512 71290 87518 71292
rect 85818 71232 85874 71241
rect 87272 71238 87274 71290
rect 87454 71238 87456 71290
rect 87210 71236 87216 71238
rect 87272 71236 87296 71238
rect 87352 71236 87376 71238
rect 87432 71236 87456 71238
rect 87512 71236 87518 71238
rect 87210 71227 87518 71236
rect 85818 71167 85874 71176
rect 88224 71105 88252 71478
rect 88210 71096 88266 71105
rect 88210 71031 88266 71040
rect 86474 70748 86782 70757
rect 86474 70746 86480 70748
rect 86536 70746 86560 70748
rect 86616 70746 86640 70748
rect 86696 70746 86720 70748
rect 86776 70746 86782 70748
rect 86536 70694 86538 70746
rect 86718 70694 86720 70746
rect 86474 70692 86480 70694
rect 86536 70692 86560 70694
rect 86616 70692 86640 70694
rect 86696 70692 86720 70694
rect 86776 70692 86782 70694
rect 86474 70683 86782 70692
rect 88212 70448 88264 70454
rect 88210 70416 88212 70425
rect 88264 70416 88266 70425
rect 85820 70380 85872 70386
rect 88210 70351 88266 70360
rect 85820 70322 85872 70328
rect 85832 70153 85860 70322
rect 87210 70204 87518 70213
rect 87210 70202 87216 70204
rect 87272 70202 87296 70204
rect 87352 70202 87376 70204
rect 87432 70202 87456 70204
rect 87512 70202 87518 70204
rect 85818 70144 85874 70153
rect 87272 70150 87274 70202
rect 87454 70150 87456 70202
rect 87210 70148 87216 70150
rect 87272 70148 87296 70150
rect 87352 70148 87376 70150
rect 87432 70148 87456 70150
rect 87512 70148 87518 70150
rect 87210 70139 87518 70148
rect 85818 70079 85874 70088
rect 86474 69660 86782 69669
rect 86474 69658 86480 69660
rect 86536 69658 86560 69660
rect 86616 69658 86640 69660
rect 86696 69658 86720 69660
rect 86776 69658 86782 69660
rect 86536 69606 86538 69658
rect 86718 69606 86720 69658
rect 86474 69604 86480 69606
rect 86536 69604 86560 69606
rect 86616 69604 86640 69606
rect 86696 69604 86720 69606
rect 86776 69604 86782 69606
rect 86474 69595 86782 69604
rect 88580 69360 88632 69366
rect 88580 69302 88632 69308
rect 84808 69292 84860 69298
rect 84808 69234 84860 69240
rect 84820 69065 84848 69234
rect 87210 69116 87518 69125
rect 87210 69114 87216 69116
rect 87272 69114 87296 69116
rect 87352 69114 87376 69116
rect 87432 69114 87456 69116
rect 87512 69114 87518 69116
rect 84806 69056 84862 69065
rect 87272 69062 87274 69114
rect 87454 69062 87456 69114
rect 88592 69065 88620 69302
rect 87210 69060 87216 69062
rect 87272 69060 87296 69062
rect 87352 69060 87376 69062
rect 87432 69060 87456 69062
rect 87512 69060 87518 69062
rect 87210 69051 87518 69060
rect 88578 69056 88634 69065
rect 84806 68991 84862 69000
rect 88578 68991 88634 69000
rect 86474 68572 86782 68581
rect 86474 68570 86480 68572
rect 86536 68570 86560 68572
rect 86616 68570 86640 68572
rect 86696 68570 86720 68572
rect 86776 68570 86782 68572
rect 86536 68518 86538 68570
rect 86718 68518 86720 68570
rect 86474 68516 86480 68518
rect 86536 68516 86560 68518
rect 86616 68516 86640 68518
rect 86696 68516 86720 68518
rect 86776 68516 86782 68518
rect 86474 68507 86782 68516
rect 87210 68028 87518 68037
rect 87210 68026 87216 68028
rect 87272 68026 87296 68028
rect 87352 68026 87376 68028
rect 87432 68026 87456 68028
rect 87512 68026 87518 68028
rect 85266 67968 85322 67977
rect 87272 67974 87274 68026
rect 87454 67974 87456 68026
rect 87210 67972 87216 67974
rect 87272 67972 87296 67974
rect 87352 67972 87376 67974
rect 87432 67972 87456 67974
rect 87512 67972 87518 67974
rect 87210 67963 87518 67972
rect 85266 67903 85322 67912
rect 85280 67870 85308 67903
rect 85268 67864 85320 67870
rect 85268 67806 85320 67812
rect 88212 67796 88264 67802
rect 88212 67738 88264 67744
rect 88224 67705 88252 67738
rect 88210 67696 88266 67705
rect 88210 67631 88266 67640
rect 86474 67484 86782 67493
rect 86474 67482 86480 67484
rect 86536 67482 86560 67484
rect 86616 67482 86640 67484
rect 86696 67482 86720 67484
rect 86776 67482 86782 67484
rect 86536 67430 86538 67482
rect 86718 67430 86720 67482
rect 86474 67428 86480 67430
rect 86536 67428 86560 67430
rect 86616 67428 86640 67430
rect 86696 67428 86720 67430
rect 86776 67428 86782 67430
rect 86474 67419 86782 67428
rect 88212 67184 88264 67190
rect 88212 67126 88264 67132
rect 85820 67116 85872 67122
rect 85820 67058 85872 67064
rect 85832 66889 85860 67058
rect 88224 67025 88252 67126
rect 88210 67016 88266 67025
rect 88210 66951 88266 66960
rect 87210 66940 87518 66949
rect 87210 66938 87216 66940
rect 87272 66938 87296 66940
rect 87352 66938 87376 66940
rect 87432 66938 87456 66940
rect 87512 66938 87518 66940
rect 85818 66880 85874 66889
rect 87272 66886 87274 66938
rect 87454 66886 87456 66938
rect 87210 66884 87216 66886
rect 87272 66884 87296 66886
rect 87352 66884 87376 66886
rect 87432 66884 87456 66886
rect 87512 66884 87518 66886
rect 87210 66875 87518 66884
rect 85818 66815 85874 66824
rect 86474 66396 86782 66405
rect 86474 66394 86480 66396
rect 86536 66394 86560 66396
rect 86616 66394 86640 66396
rect 86696 66394 86720 66396
rect 86776 66394 86782 66396
rect 86536 66342 86538 66394
rect 86718 66342 86720 66394
rect 86474 66340 86480 66342
rect 86536 66340 86560 66342
rect 86616 66340 86640 66342
rect 86696 66340 86720 66342
rect 86776 66340 86782 66342
rect 86474 66331 86782 66340
rect 85820 66096 85872 66102
rect 85820 66038 85872 66044
rect 85832 65801 85860 66038
rect 88212 65960 88264 65966
rect 88212 65902 88264 65908
rect 87210 65852 87518 65861
rect 87210 65850 87216 65852
rect 87272 65850 87296 65852
rect 87352 65850 87376 65852
rect 87432 65850 87456 65852
rect 87512 65850 87518 65852
rect 85818 65792 85874 65801
rect 87272 65798 87274 65850
rect 87454 65798 87456 65850
rect 87210 65796 87216 65798
rect 87272 65796 87296 65798
rect 87352 65796 87376 65798
rect 87432 65796 87456 65798
rect 87512 65796 87518 65798
rect 87210 65787 87518 65796
rect 85818 65727 85874 65736
rect 88224 65665 88252 65902
rect 88210 65656 88266 65665
rect 88210 65591 88266 65600
rect 86474 65308 86782 65317
rect 86474 65306 86480 65308
rect 86536 65306 86560 65308
rect 86616 65306 86640 65308
rect 86696 65306 86720 65308
rect 86776 65306 86782 65308
rect 86536 65254 86538 65306
rect 86718 65254 86720 65306
rect 86474 65252 86480 65254
rect 86536 65252 86560 65254
rect 86616 65252 86640 65254
rect 86696 65252 86720 65254
rect 86776 65252 86782 65254
rect 86474 65243 86782 65252
rect 85820 65008 85872 65014
rect 85820 64950 85872 64956
rect 88394 64976 88450 64985
rect 85832 64713 85860 64950
rect 88394 64911 88450 64920
rect 88408 64878 88436 64911
rect 88396 64872 88448 64878
rect 88396 64814 88448 64820
rect 87210 64764 87518 64773
rect 87210 64762 87216 64764
rect 87272 64762 87296 64764
rect 87352 64762 87376 64764
rect 87432 64762 87456 64764
rect 87512 64762 87518 64764
rect 85818 64704 85874 64713
rect 87272 64710 87274 64762
rect 87454 64710 87456 64762
rect 87210 64708 87216 64710
rect 87272 64708 87296 64710
rect 87352 64708 87376 64710
rect 87432 64708 87456 64710
rect 87512 64708 87518 64710
rect 87210 64699 87518 64708
rect 85818 64639 85874 64648
rect 86474 64220 86782 64229
rect 86474 64218 86480 64220
rect 86536 64218 86560 64220
rect 86616 64218 86640 64220
rect 86696 64218 86720 64220
rect 86776 64218 86782 64220
rect 86536 64166 86538 64218
rect 86718 64166 86720 64218
rect 86474 64164 86480 64166
rect 86536 64164 86560 64166
rect 86616 64164 86640 64166
rect 86696 64164 86720 64166
rect 86776 64164 86782 64166
rect 86474 64155 86782 64164
rect 84532 63920 84584 63926
rect 84532 63862 84584 63868
rect 84544 63625 84572 63862
rect 88580 63784 88632 63790
rect 88580 63726 88632 63732
rect 87210 63676 87518 63685
rect 87210 63674 87216 63676
rect 87272 63674 87296 63676
rect 87352 63674 87376 63676
rect 87432 63674 87456 63676
rect 87512 63674 87518 63676
rect 84530 63616 84586 63625
rect 87272 63622 87274 63674
rect 87454 63622 87456 63674
rect 88592 63625 88620 63726
rect 87210 63620 87216 63622
rect 87272 63620 87296 63622
rect 87352 63620 87376 63622
rect 87432 63620 87456 63622
rect 87512 63620 87518 63622
rect 87210 63611 87518 63620
rect 88578 63616 88634 63625
rect 84530 63551 84586 63560
rect 88578 63551 88634 63560
rect 86474 63132 86782 63141
rect 86474 63130 86480 63132
rect 86536 63130 86560 63132
rect 86616 63130 86640 63132
rect 86696 63130 86720 63132
rect 86776 63130 86782 63132
rect 86536 63078 86538 63130
rect 86718 63078 86720 63130
rect 86474 63076 86480 63078
rect 86536 63076 86560 63078
rect 86616 63076 86640 63078
rect 86696 63076 86720 63078
rect 86776 63076 86782 63078
rect 86474 63067 86782 63076
rect 87210 62588 87518 62597
rect 87210 62586 87216 62588
rect 87272 62586 87296 62588
rect 87352 62586 87376 62588
rect 87432 62586 87456 62588
rect 87512 62586 87518 62588
rect 84806 62528 84862 62537
rect 87272 62534 87274 62586
rect 87454 62534 87456 62586
rect 87210 62532 87216 62534
rect 87272 62532 87296 62534
rect 87352 62532 87376 62534
rect 87432 62532 87456 62534
rect 87512 62532 87518 62534
rect 87210 62523 87518 62532
rect 84806 62463 84862 62472
rect 84820 62362 84848 62463
rect 84808 62356 84860 62362
rect 84808 62298 84860 62304
rect 88394 62256 88450 62265
rect 88394 62191 88450 62200
rect 88408 62158 88436 62191
rect 88396 62152 88448 62158
rect 88396 62094 88448 62100
rect 86474 62044 86782 62053
rect 86474 62042 86480 62044
rect 86536 62042 86560 62044
rect 86616 62042 86640 62044
rect 86696 62042 86720 62044
rect 86776 62042 86782 62044
rect 86536 61990 86538 62042
rect 86718 61990 86720 62042
rect 86474 61988 86480 61990
rect 86536 61988 86560 61990
rect 86616 61988 86640 61990
rect 86696 61988 86720 61990
rect 86776 61988 86782 61990
rect 86474 61979 86782 61988
rect 85820 61744 85872 61750
rect 85820 61686 85872 61692
rect 85832 61449 85860 61686
rect 88212 61608 88264 61614
rect 88210 61576 88212 61585
rect 88264 61576 88266 61585
rect 88210 61511 88266 61520
rect 87210 61500 87518 61509
rect 87210 61498 87216 61500
rect 87272 61498 87296 61500
rect 87352 61498 87376 61500
rect 87432 61498 87456 61500
rect 87512 61498 87518 61500
rect 85818 61440 85874 61449
rect 87272 61446 87274 61498
rect 87454 61446 87456 61498
rect 87210 61444 87216 61446
rect 87272 61444 87296 61446
rect 87352 61444 87376 61446
rect 87432 61444 87456 61446
rect 87512 61444 87518 61446
rect 87210 61435 87518 61444
rect 85818 61375 85874 61384
rect 86474 60956 86782 60965
rect 86474 60954 86480 60956
rect 86536 60954 86560 60956
rect 86616 60954 86640 60956
rect 86696 60954 86720 60956
rect 86776 60954 86782 60956
rect 86536 60902 86538 60954
rect 86718 60902 86720 60954
rect 86474 60900 86480 60902
rect 86536 60900 86560 60902
rect 86616 60900 86640 60902
rect 86696 60900 86720 60902
rect 86776 60900 86782 60902
rect 86474 60891 86782 60900
rect 85820 60656 85872 60662
rect 85820 60598 85872 60604
rect 85832 60361 85860 60598
rect 88212 60520 88264 60526
rect 88212 60462 88264 60468
rect 87210 60412 87518 60421
rect 87210 60410 87216 60412
rect 87272 60410 87296 60412
rect 87352 60410 87376 60412
rect 87432 60410 87456 60412
rect 87512 60410 87518 60412
rect 85818 60352 85874 60361
rect 87272 60358 87274 60410
rect 87454 60358 87456 60410
rect 87210 60356 87216 60358
rect 87272 60356 87296 60358
rect 87352 60356 87376 60358
rect 87432 60356 87456 60358
rect 87512 60356 87518 60358
rect 87210 60347 87518 60356
rect 85818 60287 85874 60296
rect 88224 60225 88252 60462
rect 88210 60216 88266 60225
rect 88210 60151 88266 60160
rect 86474 59868 86782 59877
rect 86474 59866 86480 59868
rect 86536 59866 86560 59868
rect 86616 59866 86640 59868
rect 86696 59866 86720 59868
rect 86776 59866 86782 59868
rect 86536 59814 86538 59866
rect 86718 59814 86720 59866
rect 86474 59812 86480 59814
rect 86536 59812 86560 59814
rect 86616 59812 86640 59814
rect 86696 59812 86720 59814
rect 86776 59812 86782 59814
rect 86474 59803 86782 59812
rect 87476 59568 87528 59574
rect 87474 59536 87476 59545
rect 87528 59536 87530 59545
rect 87474 59471 87530 59480
rect 88210 59536 88266 59545
rect 88210 59471 88266 59480
rect 88224 59438 88252 59471
rect 88212 59432 88264 59438
rect 88212 59374 88264 59380
rect 87210 59324 87518 59333
rect 87210 59322 87216 59324
rect 87272 59322 87296 59324
rect 87352 59322 87376 59324
rect 87432 59322 87456 59324
rect 87512 59322 87518 59324
rect 87272 59270 87274 59322
rect 87454 59270 87456 59322
rect 87210 59268 87216 59270
rect 87272 59268 87296 59270
rect 87352 59268 87376 59270
rect 87432 59268 87456 59270
rect 87512 59268 87518 59270
rect 87210 59259 87518 59268
rect 86474 58780 86782 58789
rect 86474 58778 86480 58780
rect 86536 58778 86560 58780
rect 86616 58778 86640 58780
rect 86696 58778 86720 58780
rect 86776 58778 86782 58780
rect 86536 58726 86538 58778
rect 86718 58726 86720 58778
rect 86474 58724 86480 58726
rect 86536 58724 86560 58726
rect 86616 58724 86640 58726
rect 86696 58724 86720 58726
rect 86776 58724 86782 58726
rect 86474 58715 86782 58724
rect 85084 58480 85136 58486
rect 85084 58422 85136 58428
rect 85096 58185 85124 58422
rect 88580 58344 88632 58350
rect 88580 58286 88632 58292
rect 87210 58236 87518 58245
rect 87210 58234 87216 58236
rect 87272 58234 87296 58236
rect 87352 58234 87376 58236
rect 87432 58234 87456 58236
rect 87512 58234 87518 58236
rect 85082 58176 85138 58185
rect 87272 58182 87274 58234
rect 87454 58182 87456 58234
rect 88592 58185 88620 58286
rect 87210 58180 87216 58182
rect 87272 58180 87296 58182
rect 87352 58180 87376 58182
rect 87432 58180 87456 58182
rect 87512 58180 87518 58182
rect 87210 58171 87518 58180
rect 88578 58176 88634 58185
rect 85082 58111 85138 58120
rect 88578 58111 88634 58120
rect 86474 57692 86782 57701
rect 86474 57690 86480 57692
rect 86536 57690 86560 57692
rect 86616 57690 86640 57692
rect 86696 57690 86720 57692
rect 86776 57690 86782 57692
rect 86536 57638 86538 57690
rect 86718 57638 86720 57690
rect 86474 57636 86480 57638
rect 86536 57636 86560 57638
rect 86616 57636 86640 57638
rect 86696 57636 86720 57638
rect 86776 57636 86782 57638
rect 86474 57627 86782 57636
rect 87210 57148 87518 57157
rect 87210 57146 87216 57148
rect 87272 57146 87296 57148
rect 87352 57146 87376 57148
rect 87432 57146 87456 57148
rect 87512 57146 87518 57148
rect 87272 57094 87274 57146
rect 87454 57094 87456 57146
rect 87210 57092 87216 57094
rect 87272 57092 87296 57094
rect 87352 57092 87376 57094
rect 87432 57092 87456 57094
rect 87512 57092 87518 57094
rect 87210 57083 87518 57092
rect 88580 56984 88632 56990
rect 87566 56952 87622 56961
rect 88580 56926 88632 56932
rect 87566 56887 87568 56896
rect 87620 56887 87622 56896
rect 87568 56858 87620 56864
rect 88592 56825 88620 56926
rect 88578 56816 88634 56825
rect 88578 56751 88634 56760
rect 86474 56604 86782 56613
rect 86474 56602 86480 56604
rect 86536 56602 86560 56604
rect 86616 56602 86640 56604
rect 86696 56602 86720 56604
rect 86776 56602 86782 56604
rect 86536 56550 86538 56602
rect 86718 56550 86720 56602
rect 86474 56548 86480 56550
rect 86536 56548 86560 56550
rect 86616 56548 86640 56550
rect 86696 56548 86720 56550
rect 86776 56548 86782 56550
rect 86474 56539 86782 56548
rect 85820 56304 85872 56310
rect 85820 56246 85872 56252
rect 85832 56009 85860 56246
rect 88212 56168 88264 56174
rect 88210 56136 88212 56145
rect 88264 56136 88266 56145
rect 88210 56071 88266 56080
rect 87210 56060 87518 56069
rect 87210 56058 87216 56060
rect 87272 56058 87296 56060
rect 87352 56058 87376 56060
rect 87432 56058 87456 56060
rect 87512 56058 87518 56060
rect 85818 56000 85874 56009
rect 87272 56006 87274 56058
rect 87454 56006 87456 56058
rect 87210 56004 87216 56006
rect 87272 56004 87296 56006
rect 87352 56004 87376 56006
rect 87432 56004 87456 56006
rect 87512 56004 87518 56006
rect 87210 55995 87518 56004
rect 85818 55935 85874 55944
rect 86474 55516 86782 55525
rect 86474 55514 86480 55516
rect 86536 55514 86560 55516
rect 86616 55514 86640 55516
rect 86696 55514 86720 55516
rect 86776 55514 86782 55516
rect 86536 55462 86538 55514
rect 86718 55462 86720 55514
rect 86474 55460 86480 55462
rect 86536 55460 86560 55462
rect 86616 55460 86640 55462
rect 86696 55460 86720 55462
rect 86776 55460 86782 55462
rect 86474 55451 86782 55460
rect 85820 55216 85872 55222
rect 85820 55158 85872 55164
rect 85832 54921 85860 55158
rect 88212 55080 88264 55086
rect 88212 55022 88264 55028
rect 87210 54972 87518 54981
rect 87210 54970 87216 54972
rect 87272 54970 87296 54972
rect 87352 54970 87376 54972
rect 87432 54970 87456 54972
rect 87512 54970 87518 54972
rect 85818 54912 85874 54921
rect 87272 54918 87274 54970
rect 87454 54918 87456 54970
rect 87210 54916 87216 54918
rect 87272 54916 87296 54918
rect 87352 54916 87376 54918
rect 87432 54916 87456 54918
rect 87512 54916 87518 54918
rect 87210 54907 87518 54916
rect 85818 54847 85874 54856
rect 88224 54785 88252 55022
rect 88210 54776 88266 54785
rect 88210 54711 88266 54720
rect 86474 54428 86782 54437
rect 86474 54426 86480 54428
rect 86536 54426 86560 54428
rect 86616 54426 86640 54428
rect 86696 54426 86720 54428
rect 86776 54426 86782 54428
rect 86536 54374 86538 54426
rect 86718 54374 86720 54426
rect 86474 54372 86480 54374
rect 86536 54372 86560 54374
rect 86616 54372 86640 54374
rect 86696 54372 86720 54374
rect 86776 54372 86782 54374
rect 86474 54363 86782 54372
rect 84532 54128 84584 54134
rect 88212 54128 88264 54134
rect 84532 54070 84584 54076
rect 88210 54096 88212 54105
rect 88264 54096 88266 54105
rect 84544 53833 84572 54070
rect 88210 54031 88266 54040
rect 87210 53884 87518 53893
rect 87210 53882 87216 53884
rect 87272 53882 87296 53884
rect 87352 53882 87376 53884
rect 87432 53882 87456 53884
rect 87512 53882 87518 53884
rect 84530 53824 84586 53833
rect 87272 53830 87274 53882
rect 87454 53830 87456 53882
rect 87210 53828 87216 53830
rect 87272 53828 87296 53830
rect 87352 53828 87376 53830
rect 87432 53828 87456 53830
rect 87512 53828 87518 53830
rect 87210 53819 87518 53828
rect 84530 53759 84586 53768
rect 86474 53340 86782 53349
rect 86474 53338 86480 53340
rect 86536 53338 86560 53340
rect 86616 53338 86640 53340
rect 86696 53338 86720 53340
rect 86776 53338 86782 53340
rect 86536 53286 86538 53338
rect 86718 53286 86720 53338
rect 86474 53284 86480 53286
rect 86536 53284 86560 53286
rect 86616 53284 86640 53286
rect 86696 53284 86720 53286
rect 86776 53284 86782 53286
rect 86474 53275 86782 53284
rect 87568 53040 87620 53046
rect 87566 53008 87568 53017
rect 87620 53008 87622 53017
rect 87566 52943 87622 52952
rect 88212 52904 88264 52910
rect 88212 52846 88264 52852
rect 87210 52796 87518 52805
rect 87210 52794 87216 52796
rect 87272 52794 87296 52796
rect 87352 52794 87376 52796
rect 87432 52794 87456 52796
rect 87512 52794 87518 52796
rect 87272 52742 87274 52794
rect 87454 52742 87456 52794
rect 88224 52745 88252 52846
rect 87210 52740 87216 52742
rect 87272 52740 87296 52742
rect 87352 52740 87376 52742
rect 87432 52740 87456 52742
rect 87512 52740 87518 52742
rect 87210 52731 87518 52740
rect 88210 52736 88266 52745
rect 88210 52671 88266 52680
rect 86474 52252 86782 52261
rect 86474 52250 86480 52252
rect 86536 52250 86560 52252
rect 86616 52250 86640 52252
rect 86696 52250 86720 52252
rect 86776 52250 86782 52252
rect 86536 52198 86538 52250
rect 86718 52198 86720 52250
rect 86474 52196 86480 52198
rect 86536 52196 86560 52198
rect 86616 52196 86640 52198
rect 86696 52196 86720 52198
rect 86776 52196 86782 52198
rect 86474 52187 86782 52196
rect 87210 51708 87518 51717
rect 87210 51706 87216 51708
rect 87272 51706 87296 51708
rect 87352 51706 87376 51708
rect 87432 51706 87456 51708
rect 87512 51706 87518 51708
rect 87272 51654 87274 51706
rect 87454 51654 87456 51706
rect 87210 51652 87216 51654
rect 87272 51652 87296 51654
rect 87352 51652 87376 51654
rect 87432 51652 87456 51654
rect 87512 51652 87518 51654
rect 87210 51643 87518 51652
rect 87566 51512 87622 51521
rect 87566 51447 87568 51456
rect 87620 51447 87622 51456
rect 87568 51418 87620 51424
rect 88210 51376 88266 51385
rect 88210 51311 88212 51320
rect 88264 51311 88266 51320
rect 88212 51282 88264 51288
rect 86474 51164 86782 51173
rect 86474 51162 86480 51164
rect 86536 51162 86560 51164
rect 86616 51162 86640 51164
rect 86696 51162 86720 51164
rect 86776 51162 86782 51164
rect 86536 51110 86538 51162
rect 86718 51110 86720 51162
rect 86474 51108 86480 51110
rect 86536 51108 86560 51110
rect 86616 51108 86640 51110
rect 86696 51108 86720 51110
rect 86776 51108 86782 51110
rect 86474 51099 86782 51108
rect 85636 50728 85688 50734
rect 85636 50670 85688 50676
rect 85648 50569 85676 50670
rect 87210 50620 87518 50629
rect 87210 50618 87216 50620
rect 87272 50618 87296 50620
rect 87352 50618 87376 50620
rect 87432 50618 87456 50620
rect 87512 50618 87518 50620
rect 85450 50560 85506 50569
rect 85450 50495 85506 50504
rect 85634 50560 85690 50569
rect 87272 50566 87274 50618
rect 87454 50566 87456 50618
rect 87210 50564 87216 50566
rect 87272 50564 87296 50566
rect 87352 50564 87376 50566
rect 87432 50564 87456 50566
rect 87512 50564 87518 50566
rect 87210 50555 87518 50564
rect 85634 50495 85690 50504
rect 85360 48620 85412 48626
rect 85360 48562 85412 48568
rect 85372 48393 85400 48562
rect 85358 48384 85414 48393
rect 85358 48319 85414 48328
rect 83610 44644 83666 44653
rect 83610 44579 83666 44588
rect 83624 44410 83652 44579
rect 83612 44404 83664 44410
rect 83612 44346 83664 44352
rect 84808 36176 84860 36182
rect 84808 36118 84860 36124
rect 84820 36017 84848 36118
rect 84806 36008 84862 36017
rect 84806 35943 84862 35952
rect 84808 30668 84860 30674
rect 84808 30610 84860 30616
rect 84820 30577 84848 30610
rect 84806 30568 84862 30577
rect 84806 30503 84862 30512
rect 84808 25364 84860 25370
rect 84808 25306 84860 25312
rect 84820 25001 84848 25306
rect 84806 24992 84862 25001
rect 84806 24927 84862 24936
rect 84808 21012 84860 21018
rect 84808 20954 84860 20960
rect 84820 20785 84848 20954
rect 84806 20776 84862 20785
rect 84806 20711 84862 20720
rect 84808 15572 84860 15578
rect 84808 15514 84860 15520
rect 84820 15345 84848 15514
rect 84806 15336 84862 15345
rect 84806 15271 84862 15280
rect 83428 14280 83480 14286
rect 83428 14222 83480 14228
rect 83440 14189 83468 14222
rect 83426 14180 83482 14189
rect 83426 14115 83482 14124
rect 83244 11288 83296 11294
rect 83244 11230 83296 11236
rect 46442 10984 46498 10993
rect 46442 10919 46498 10928
rect 46076 10200 46128 10206
rect 46456 10177 46484 10919
rect 83256 10902 83284 11230
rect 83334 10916 83390 10925
rect 83256 10874 83334 10902
rect 83334 10851 83390 10860
rect 82508 10200 82560 10206
rect 46076 10142 46128 10148
rect 46442 10168 46498 10177
rect 52404 10126 52648 10154
rect 53508 10126 53568 10154
rect 46442 10103 46498 10112
rect 45432 7480 45484 7486
rect 45432 7422 45484 7428
rect 45708 7480 45760 7486
rect 45708 7422 45760 7428
rect 45892 7480 45944 7486
rect 45892 7422 45944 7428
rect 45984 7480 46036 7486
rect 45984 7422 46036 7428
rect 45720 7214 45748 7422
rect 45996 7282 46024 7422
rect 45984 7276 46036 7282
rect 45984 7218 46036 7224
rect 45708 7208 45760 7214
rect 45708 7150 45760 7156
rect 30436 5304 30488 5310
rect 30436 5246 30488 5252
rect 31540 5304 31592 5310
rect 31540 5246 31592 5252
rect 32644 5304 32696 5310
rect 32644 5246 32696 5252
rect 33748 5304 33800 5310
rect 33748 5246 33800 5252
rect 34852 5304 34904 5310
rect 34852 5246 34904 5252
rect 35956 5304 36008 5310
rect 35956 5246 36008 5252
rect 37152 5304 37204 5310
rect 37152 5246 37204 5252
rect 38164 5304 38216 5310
rect 38164 5246 38216 5252
rect 39268 5304 39320 5310
rect 39268 5246 39320 5252
rect 40372 5304 40424 5310
rect 40372 5246 40424 5252
rect 41476 5304 41528 5310
rect 41476 5246 41528 5252
rect 42580 5304 42632 5310
rect 42580 5246 42632 5252
rect 43684 5304 43736 5310
rect 43684 5246 43736 5252
rect 44788 5304 44840 5310
rect 44788 5246 44840 5252
rect 52620 5174 52648 10126
rect 53540 5174 53568 10126
rect 54460 10126 54612 10154
rect 55716 10126 55868 10154
rect 56820 10126 57064 10154
rect 57924 10126 58076 10154
rect 59028 10126 59088 10154
rect 60132 10126 60376 10154
rect 61236 10126 61296 10154
rect 62340 10126 62400 10154
rect 63444 10126 63596 10154
rect 64548 10126 64792 10154
rect 65652 10126 65804 10154
rect 66756 10126 66816 10154
rect 67860 10126 68104 10154
rect 68964 10126 69024 10154
rect 54460 5174 54488 10126
rect 54522 7644 54830 7653
rect 54522 7642 54528 7644
rect 54584 7642 54608 7644
rect 54664 7642 54688 7644
rect 54744 7642 54768 7644
rect 54824 7642 54830 7644
rect 54584 7590 54586 7642
rect 54766 7590 54768 7642
rect 54522 7588 54528 7590
rect 54584 7588 54608 7590
rect 54664 7588 54688 7590
rect 54744 7588 54768 7590
rect 54824 7588 54830 7590
rect 54522 7579 54830 7588
rect 55182 7100 55490 7109
rect 55182 7098 55188 7100
rect 55244 7098 55268 7100
rect 55324 7098 55348 7100
rect 55404 7098 55428 7100
rect 55484 7098 55490 7100
rect 55244 7046 55246 7098
rect 55426 7046 55428 7098
rect 55182 7044 55188 7046
rect 55244 7044 55268 7046
rect 55324 7044 55348 7046
rect 55404 7044 55428 7046
rect 55484 7044 55490 7046
rect 55182 7035 55490 7044
rect 54522 6556 54830 6565
rect 54522 6554 54528 6556
rect 54584 6554 54608 6556
rect 54664 6554 54688 6556
rect 54744 6554 54768 6556
rect 54824 6554 54830 6556
rect 54584 6502 54586 6554
rect 54766 6502 54768 6554
rect 54522 6500 54528 6502
rect 54584 6500 54608 6502
rect 54664 6500 54688 6502
rect 54744 6500 54768 6502
rect 54824 6500 54830 6502
rect 54522 6491 54830 6500
rect 55182 6012 55490 6021
rect 55182 6010 55188 6012
rect 55244 6010 55268 6012
rect 55324 6010 55348 6012
rect 55404 6010 55428 6012
rect 55484 6010 55490 6012
rect 55244 5958 55246 6010
rect 55426 5958 55428 6010
rect 55182 5956 55188 5958
rect 55244 5956 55268 5958
rect 55324 5956 55348 5958
rect 55404 5956 55428 5958
rect 55484 5956 55490 5958
rect 55182 5947 55490 5956
rect 54522 5468 54830 5477
rect 54522 5466 54528 5468
rect 54584 5466 54608 5468
rect 54664 5466 54688 5468
rect 54744 5466 54768 5468
rect 54824 5466 54830 5468
rect 54584 5414 54586 5466
rect 54766 5414 54768 5466
rect 54522 5412 54528 5414
rect 54584 5412 54608 5414
rect 54664 5412 54688 5414
rect 54744 5412 54768 5414
rect 54824 5412 54830 5414
rect 54522 5403 54830 5412
rect 55840 5174 55868 10126
rect 57036 5174 57064 10126
rect 58048 5174 58076 10126
rect 59060 5174 59088 10126
rect 60348 5174 60376 10126
rect 61268 5174 61296 10126
rect 62372 5174 62400 10126
rect 63568 5174 63596 10126
rect 64764 5174 64792 10126
rect 65776 5174 65804 10126
rect 66788 5174 66816 10126
rect 68076 5310 68104 10126
rect 68996 5310 69024 10126
rect 70054 9914 70082 10140
rect 71172 10126 71324 10154
rect 72276 10126 72612 10154
rect 73380 10126 73440 10154
rect 74484 10126 74544 10154
rect 75588 10126 75832 10154
rect 76692 10126 76752 10154
rect 70008 9886 70082 9914
rect 70008 5310 70036 9886
rect 71296 5310 71324 10126
rect 72584 5310 72612 10126
rect 72922 7644 73230 7653
rect 72922 7642 72928 7644
rect 72984 7642 73008 7644
rect 73064 7642 73088 7644
rect 73144 7642 73168 7644
rect 73224 7642 73230 7644
rect 72984 7590 72986 7642
rect 73166 7590 73168 7642
rect 72922 7588 72928 7590
rect 72984 7588 73008 7590
rect 73064 7588 73088 7590
rect 73144 7588 73168 7590
rect 73224 7588 73230 7590
rect 72922 7579 73230 7588
rect 72922 6556 73230 6565
rect 72922 6554 72928 6556
rect 72984 6554 73008 6556
rect 73064 6554 73088 6556
rect 73144 6554 73168 6556
rect 73224 6554 73230 6556
rect 72984 6502 72986 6554
rect 73166 6502 73168 6554
rect 72922 6500 72928 6502
rect 72984 6500 73008 6502
rect 73064 6500 73088 6502
rect 73144 6500 73168 6502
rect 73224 6500 73230 6502
rect 72922 6491 73230 6500
rect 72922 5468 73230 5477
rect 72922 5466 72928 5468
rect 72984 5466 73008 5468
rect 73064 5466 73088 5468
rect 73144 5466 73168 5468
rect 73224 5466 73230 5468
rect 72984 5414 72986 5466
rect 73166 5414 73168 5466
rect 72922 5412 72928 5414
rect 72984 5412 73008 5414
rect 73064 5412 73088 5414
rect 73144 5412 73168 5414
rect 73224 5412 73230 5414
rect 72922 5403 73230 5412
rect 73412 5310 73440 10126
rect 73582 7100 73890 7109
rect 73582 7098 73588 7100
rect 73644 7098 73668 7100
rect 73724 7098 73748 7100
rect 73804 7098 73828 7100
rect 73884 7098 73890 7100
rect 73644 7046 73646 7098
rect 73826 7046 73828 7098
rect 73582 7044 73588 7046
rect 73644 7044 73668 7046
rect 73724 7044 73748 7046
rect 73804 7044 73828 7046
rect 73884 7044 73890 7046
rect 73582 7035 73890 7044
rect 73582 6012 73890 6021
rect 73582 6010 73588 6012
rect 73644 6010 73668 6012
rect 73724 6010 73748 6012
rect 73804 6010 73828 6012
rect 73884 6010 73890 6012
rect 73644 5958 73646 6010
rect 73826 5958 73828 6010
rect 73582 5956 73588 5958
rect 73644 5956 73668 5958
rect 73724 5956 73748 5958
rect 73804 5956 73828 5958
rect 73884 5956 73890 5958
rect 73582 5947 73890 5956
rect 74516 5310 74544 10126
rect 75804 5310 75832 10126
rect 76724 5310 76752 10126
rect 77782 9914 77810 10140
rect 78900 10126 79052 10154
rect 80004 10126 80156 10154
rect 81108 10126 81168 10154
rect 82212 10148 82508 10154
rect 82212 10142 82560 10148
rect 82212 10126 82548 10142
rect 77736 9886 77810 9914
rect 77736 5310 77764 9886
rect 79024 5310 79052 10126
rect 80128 5310 80156 10126
rect 81140 5310 81168 10126
rect 83440 9914 83468 14115
rect 83612 13464 83664 13470
rect 83612 13406 83664 13412
rect 83624 13101 83652 13406
rect 83610 13092 83666 13101
rect 83348 9886 83468 9914
rect 83532 13050 83610 13078
rect 83348 7282 83376 9886
rect 83532 7350 83560 13050
rect 83610 13027 83666 13036
rect 85372 12654 85400 48319
rect 85464 15034 85492 50495
rect 86474 50076 86782 50085
rect 86474 50074 86480 50076
rect 86536 50074 86560 50076
rect 86616 50074 86640 50076
rect 86696 50074 86720 50076
rect 86776 50074 86782 50076
rect 86536 50022 86538 50074
rect 86718 50022 86720 50074
rect 86474 50020 86480 50022
rect 86536 50020 86560 50022
rect 86616 50020 86640 50022
rect 86696 50020 86720 50022
rect 86776 50020 86782 50022
rect 86474 50011 86782 50020
rect 85636 49640 85688 49646
rect 85636 49582 85688 49588
rect 85648 49481 85676 49582
rect 87210 49532 87518 49541
rect 87210 49530 87216 49532
rect 87272 49530 87296 49532
rect 87352 49530 87376 49532
rect 87432 49530 87456 49532
rect 87512 49530 87518 49532
rect 85634 49472 85690 49481
rect 87272 49478 87274 49530
rect 87454 49478 87456 49530
rect 87210 49476 87216 49478
rect 87272 49476 87296 49478
rect 87352 49476 87376 49478
rect 87432 49476 87456 49478
rect 87512 49476 87518 49478
rect 87210 49467 87518 49476
rect 85634 49407 85690 49416
rect 85648 48554 85676 49407
rect 86474 48988 86782 48997
rect 86474 48986 86480 48988
rect 86536 48986 86560 48988
rect 86616 48986 86640 48988
rect 86696 48986 86720 48988
rect 86776 48986 86782 48988
rect 86536 48934 86538 48986
rect 86718 48934 86720 48986
rect 86474 48932 86480 48934
rect 86536 48932 86560 48934
rect 86616 48932 86640 48934
rect 86696 48932 86720 48934
rect 86776 48932 86782 48934
rect 86474 48923 86782 48932
rect 88212 48688 88264 48694
rect 88210 48656 88212 48665
rect 88264 48656 88266 48665
rect 88210 48591 88266 48600
rect 85556 48526 85676 48554
rect 85452 15028 85504 15034
rect 85452 14970 85504 14976
rect 85556 13470 85584 48526
rect 87210 48444 87518 48453
rect 87210 48442 87216 48444
rect 87272 48442 87296 48444
rect 87352 48442 87376 48444
rect 87432 48442 87456 48444
rect 87512 48442 87518 48444
rect 87272 48390 87274 48442
rect 87454 48390 87456 48442
rect 87210 48388 87216 48390
rect 87272 48388 87296 48390
rect 87352 48388 87376 48390
rect 87432 48388 87456 48390
rect 87512 48388 87518 48390
rect 87210 48379 87518 48388
rect 88212 48008 88264 48014
rect 88210 47976 88212 47985
rect 88264 47976 88266 47985
rect 88210 47911 88266 47920
rect 86474 47900 86782 47909
rect 86474 47898 86480 47900
rect 86536 47898 86560 47900
rect 86616 47898 86640 47900
rect 86696 47898 86720 47900
rect 86776 47898 86782 47900
rect 86536 47846 86538 47898
rect 86718 47846 86720 47898
rect 86474 47844 86480 47846
rect 86536 47844 86560 47846
rect 86616 47844 86640 47846
rect 86696 47844 86720 47846
rect 86776 47844 86782 47846
rect 86474 47835 86782 47844
rect 85820 47600 85872 47606
rect 85820 47542 85872 47548
rect 85832 47305 85860 47542
rect 88212 47464 88264 47470
rect 88212 47406 88264 47412
rect 87210 47356 87518 47365
rect 87210 47354 87216 47356
rect 87272 47354 87296 47356
rect 87352 47354 87376 47356
rect 87432 47354 87456 47356
rect 87512 47354 87518 47356
rect 85818 47296 85874 47305
rect 87272 47302 87274 47354
rect 87454 47302 87456 47354
rect 88224 47305 88252 47406
rect 87210 47300 87216 47302
rect 87272 47300 87296 47302
rect 87352 47300 87376 47302
rect 87432 47300 87456 47302
rect 87512 47300 87518 47302
rect 87210 47291 87518 47300
rect 88210 47296 88266 47305
rect 85818 47231 85874 47240
rect 88210 47231 88266 47240
rect 88212 46920 88264 46926
rect 88212 46862 88264 46868
rect 86474 46812 86782 46821
rect 86474 46810 86480 46812
rect 86536 46810 86560 46812
rect 86616 46810 86640 46812
rect 86696 46810 86720 46812
rect 86776 46810 86782 46812
rect 86536 46758 86538 46810
rect 86718 46758 86720 46810
rect 86474 46756 86480 46758
rect 86536 46756 86560 46758
rect 86616 46756 86640 46758
rect 86696 46756 86720 46758
rect 86776 46756 86782 46758
rect 86474 46747 86782 46756
rect 88224 46625 88252 46862
rect 88210 46616 88266 46625
rect 88210 46551 88266 46560
rect 87210 46268 87518 46277
rect 87210 46266 87216 46268
rect 87272 46266 87296 46268
rect 87352 46266 87376 46268
rect 87432 46266 87456 46268
rect 87512 46266 87518 46268
rect 87272 46214 87274 46266
rect 87454 46214 87456 46266
rect 87210 46212 87216 46214
rect 87272 46212 87296 46214
rect 87352 46212 87376 46214
rect 87432 46212 87456 46214
rect 87512 46212 87518 46214
rect 87210 46203 87518 46212
rect 85820 45900 85872 45906
rect 85820 45842 85872 45848
rect 85832 45566 85860 45842
rect 86474 45724 86782 45733
rect 86474 45722 86480 45724
rect 86536 45722 86560 45724
rect 86616 45722 86640 45724
rect 86696 45722 86720 45724
rect 86776 45722 86782 45724
rect 86536 45670 86538 45722
rect 86718 45670 86720 45722
rect 86474 45668 86480 45670
rect 86536 45668 86560 45670
rect 86616 45668 86640 45670
rect 86696 45668 86720 45670
rect 86776 45668 86782 45670
rect 86474 45659 86782 45668
rect 85820 45560 85872 45566
rect 85820 45502 85872 45508
rect 86004 45424 86056 45430
rect 86002 45392 86004 45401
rect 88212 45424 88264 45430
rect 86056 45392 86058 45401
rect 88212 45366 88264 45372
rect 86002 45327 86058 45336
rect 85636 45288 85688 45294
rect 86188 45288 86240 45294
rect 85636 45230 85688 45236
rect 86186 45256 86188 45265
rect 88224 45265 88252 45366
rect 86240 45256 86242 45265
rect 85648 45129 85676 45230
rect 86186 45191 86242 45200
rect 88210 45256 88266 45265
rect 88210 45191 88266 45200
rect 87210 45180 87518 45189
rect 87210 45178 87216 45180
rect 87272 45178 87296 45180
rect 87352 45178 87376 45180
rect 87432 45178 87456 45180
rect 87512 45178 87518 45180
rect 85634 45120 85690 45129
rect 87272 45126 87274 45178
rect 87454 45126 87456 45178
rect 87210 45124 87216 45126
rect 87272 45124 87296 45126
rect 87352 45124 87376 45126
rect 87432 45124 87456 45126
rect 87512 45124 87518 45126
rect 87210 45115 87518 45124
rect 85634 45055 85690 45064
rect 88212 44744 88264 44750
rect 88212 44686 88264 44692
rect 86474 44636 86782 44645
rect 86474 44634 86480 44636
rect 86536 44634 86560 44636
rect 86616 44634 86640 44636
rect 86696 44634 86720 44636
rect 86776 44634 86782 44636
rect 86536 44582 86538 44634
rect 86718 44582 86720 44634
rect 88224 44585 88252 44686
rect 86474 44580 86480 44582
rect 86536 44580 86560 44582
rect 86616 44580 86640 44582
rect 86696 44580 86720 44582
rect 86776 44580 86782 44582
rect 86474 44571 86782 44580
rect 88210 44576 88266 44585
rect 88210 44511 88266 44520
rect 88212 44336 88264 44342
rect 88212 44278 88264 44284
rect 87210 44092 87518 44101
rect 87210 44090 87216 44092
rect 87272 44090 87296 44092
rect 87352 44090 87376 44092
rect 87432 44090 87456 44092
rect 87512 44090 87518 44092
rect 87272 44038 87274 44090
rect 87454 44038 87456 44090
rect 87210 44036 87216 44038
rect 87272 44036 87296 44038
rect 87352 44036 87376 44038
rect 87432 44036 87456 44038
rect 87512 44036 87518 44038
rect 87210 44027 87518 44036
rect 88224 43905 88252 44278
rect 88210 43896 88266 43905
rect 88210 43831 88266 43840
rect 86474 43548 86782 43557
rect 86474 43546 86480 43548
rect 86536 43546 86560 43548
rect 86616 43546 86640 43548
rect 86696 43546 86720 43548
rect 86776 43546 86782 43548
rect 85818 43488 85874 43497
rect 86536 43494 86538 43546
rect 86718 43494 86720 43546
rect 86474 43492 86480 43494
rect 86536 43492 86560 43494
rect 86616 43492 86640 43494
rect 86696 43492 86720 43494
rect 86776 43492 86782 43494
rect 86474 43483 86782 43492
rect 85818 43423 85874 43432
rect 85832 43390 85860 43423
rect 85820 43384 85872 43390
rect 85820 43326 85872 43332
rect 88212 43248 88264 43254
rect 88210 43216 88212 43225
rect 88264 43216 88266 43225
rect 88210 43151 88266 43160
rect 87210 43004 87518 43013
rect 87210 43002 87216 43004
rect 87272 43002 87296 43004
rect 87352 43002 87376 43004
rect 87432 43002 87456 43004
rect 87512 43002 87518 43004
rect 87272 42950 87274 43002
rect 87454 42950 87456 43002
rect 87210 42948 87216 42950
rect 87272 42948 87296 42950
rect 87352 42948 87376 42950
rect 87432 42948 87456 42950
rect 87512 42948 87518 42950
rect 87210 42939 87518 42948
rect 88212 42772 88264 42778
rect 88212 42714 88264 42720
rect 85820 42636 85872 42642
rect 85820 42578 85872 42584
rect 85832 42545 85860 42578
rect 88224 42545 88252 42714
rect 85818 42536 85874 42545
rect 85818 42471 85874 42480
rect 88210 42536 88266 42545
rect 88210 42471 88266 42480
rect 86474 42460 86782 42469
rect 86474 42458 86480 42460
rect 86536 42458 86560 42460
rect 86616 42458 86640 42460
rect 86696 42458 86720 42460
rect 86776 42458 86782 42460
rect 86536 42406 86538 42458
rect 86718 42406 86720 42458
rect 86474 42404 86480 42406
rect 86536 42404 86560 42406
rect 86616 42404 86640 42406
rect 86696 42404 86720 42406
rect 86776 42404 86782 42406
rect 86474 42395 86782 42404
rect 87210 41916 87518 41925
rect 87210 41914 87216 41916
rect 87272 41914 87296 41916
rect 87352 41914 87376 41916
rect 87432 41914 87456 41916
rect 87512 41914 87518 41916
rect 87272 41862 87274 41914
rect 87454 41862 87456 41914
rect 87210 41860 87216 41862
rect 87272 41860 87296 41862
rect 87352 41860 87376 41862
rect 87432 41860 87456 41862
rect 87512 41860 87518 41862
rect 87210 41851 87518 41860
rect 87568 41684 87620 41690
rect 87568 41626 87620 41632
rect 88212 41684 88264 41690
rect 88212 41626 88264 41632
rect 87580 41593 87608 41626
rect 87566 41584 87622 41593
rect 87566 41519 87622 41528
rect 86474 41372 86782 41381
rect 86474 41370 86480 41372
rect 86536 41370 86560 41372
rect 86616 41370 86640 41372
rect 86696 41370 86720 41372
rect 86776 41370 86782 41372
rect 86536 41318 86538 41370
rect 86718 41318 86720 41370
rect 86474 41316 86480 41318
rect 86536 41316 86560 41318
rect 86616 41316 86640 41318
rect 86696 41316 86720 41318
rect 86776 41316 86782 41318
rect 86474 41307 86782 41316
rect 88224 41185 88252 41626
rect 88210 41176 88266 41185
rect 88210 41111 88266 41120
rect 87210 40828 87518 40837
rect 87210 40826 87216 40828
rect 87272 40826 87296 40828
rect 87352 40826 87376 40828
rect 87432 40826 87456 40828
rect 87512 40826 87518 40828
rect 87272 40774 87274 40826
rect 87454 40774 87456 40826
rect 87210 40772 87216 40774
rect 87272 40772 87296 40774
rect 87352 40772 87376 40774
rect 87432 40772 87456 40774
rect 87512 40772 87518 40774
rect 87210 40763 87518 40772
rect 87936 40528 87988 40534
rect 87934 40496 87936 40505
rect 88212 40528 88264 40534
rect 87988 40496 87990 40505
rect 87934 40431 87990 40440
rect 88210 40496 88212 40505
rect 88264 40496 88266 40505
rect 88210 40431 88266 40440
rect 86474 40284 86782 40293
rect 86474 40282 86480 40284
rect 86536 40282 86560 40284
rect 86616 40282 86640 40284
rect 86696 40282 86720 40284
rect 86776 40282 86782 40284
rect 86536 40230 86538 40282
rect 86718 40230 86720 40282
rect 86474 40228 86480 40230
rect 86536 40228 86560 40230
rect 86616 40228 86640 40230
rect 86696 40228 86720 40230
rect 86776 40228 86782 40230
rect 86474 40219 86782 40228
rect 88224 40126 88252 40431
rect 88212 40120 88264 40126
rect 88212 40062 88264 40068
rect 87210 39740 87518 39749
rect 87210 39738 87216 39740
rect 87272 39738 87296 39740
rect 87352 39738 87376 39740
rect 87432 39738 87456 39740
rect 87512 39738 87518 39740
rect 87272 39686 87274 39738
rect 87454 39686 87456 39738
rect 87210 39684 87216 39686
rect 87272 39684 87296 39686
rect 87352 39684 87376 39686
rect 87432 39684 87456 39686
rect 87512 39684 87518 39686
rect 87210 39675 87518 39684
rect 88212 39508 88264 39514
rect 88212 39450 88264 39456
rect 87566 39408 87622 39417
rect 87566 39343 87568 39352
rect 87620 39343 87622 39352
rect 87568 39314 87620 39320
rect 86474 39196 86782 39205
rect 86474 39194 86480 39196
rect 86536 39194 86560 39196
rect 86616 39194 86640 39196
rect 86696 39194 86720 39196
rect 86776 39194 86782 39196
rect 86536 39142 86538 39194
rect 86718 39142 86720 39194
rect 88224 39145 88252 39450
rect 86474 39140 86480 39142
rect 86536 39140 86560 39142
rect 86616 39140 86640 39142
rect 86696 39140 86720 39142
rect 86776 39140 86782 39142
rect 86474 39131 86782 39140
rect 88210 39136 88266 39145
rect 88210 39071 88266 39080
rect 87210 38652 87518 38661
rect 87210 38650 87216 38652
rect 87272 38650 87296 38652
rect 87352 38650 87376 38652
rect 87432 38650 87456 38652
rect 87512 38650 87518 38652
rect 87272 38598 87274 38650
rect 87454 38598 87456 38650
rect 87210 38596 87216 38598
rect 87272 38596 87296 38598
rect 87352 38596 87376 38598
rect 87432 38596 87456 38598
rect 87512 38596 87518 38598
rect 87210 38587 87518 38596
rect 86474 38108 86782 38117
rect 86474 38106 86480 38108
rect 86536 38106 86560 38108
rect 86616 38106 86640 38108
rect 86696 38106 86720 38108
rect 86776 38106 86782 38108
rect 85818 38048 85874 38057
rect 86536 38054 86538 38106
rect 86718 38054 86720 38106
rect 86474 38052 86480 38054
rect 86536 38052 86560 38054
rect 86616 38052 86640 38054
rect 86696 38052 86720 38054
rect 86776 38052 86782 38054
rect 86474 38043 86782 38052
rect 85818 37983 85874 37992
rect 85832 37950 85860 37983
rect 85820 37944 85872 37950
rect 85820 37886 85872 37892
rect 88212 37808 88264 37814
rect 88210 37776 88212 37785
rect 88264 37776 88266 37785
rect 88210 37711 88266 37720
rect 87210 37564 87518 37573
rect 87210 37562 87216 37564
rect 87272 37562 87296 37564
rect 87352 37562 87376 37564
rect 87432 37562 87456 37564
rect 87512 37562 87518 37564
rect 87272 37510 87274 37562
rect 87454 37510 87456 37562
rect 87210 37508 87216 37510
rect 87272 37508 87296 37510
rect 87352 37508 87376 37510
rect 87432 37508 87456 37510
rect 87512 37508 87518 37510
rect 87210 37499 87518 37508
rect 88212 37332 88264 37338
rect 88212 37274 88264 37280
rect 85820 37196 85872 37202
rect 85820 37138 85872 37144
rect 85832 37105 85860 37138
rect 88224 37105 88252 37274
rect 85818 37096 85874 37105
rect 85818 37031 85874 37040
rect 88210 37096 88266 37105
rect 88210 37031 88266 37040
rect 86474 37020 86782 37029
rect 86474 37018 86480 37020
rect 86536 37018 86560 37020
rect 86616 37018 86640 37020
rect 86696 37018 86720 37020
rect 86776 37018 86782 37020
rect 86536 36966 86538 37018
rect 86718 36966 86720 37018
rect 86474 36964 86480 36966
rect 86536 36964 86560 36966
rect 86616 36964 86640 36966
rect 86696 36964 86720 36966
rect 86776 36964 86782 36966
rect 86474 36955 86782 36964
rect 87210 36476 87518 36485
rect 87210 36474 87216 36476
rect 87272 36474 87296 36476
rect 87352 36474 87376 36476
rect 87432 36474 87456 36476
rect 87512 36474 87518 36476
rect 87272 36422 87274 36474
rect 87454 36422 87456 36474
rect 87210 36420 87216 36422
rect 87272 36420 87296 36422
rect 87352 36420 87376 36422
rect 87432 36420 87456 36422
rect 87512 36420 87518 36422
rect 87210 36411 87518 36420
rect 88580 36244 88632 36250
rect 88580 36186 88632 36192
rect 86474 35932 86782 35941
rect 86474 35930 86480 35932
rect 86536 35930 86560 35932
rect 86616 35930 86640 35932
rect 86696 35930 86720 35932
rect 86776 35930 86782 35932
rect 86536 35878 86538 35930
rect 86718 35878 86720 35930
rect 86474 35876 86480 35878
rect 86536 35876 86560 35878
rect 86616 35876 86640 35878
rect 86696 35876 86720 35878
rect 86776 35876 86782 35878
rect 86474 35867 86782 35876
rect 88592 35745 88620 36186
rect 88578 35736 88634 35745
rect 88578 35671 88634 35680
rect 87210 35388 87518 35397
rect 87210 35386 87216 35388
rect 87272 35386 87296 35388
rect 87352 35386 87376 35388
rect 87432 35386 87456 35388
rect 87512 35386 87518 35388
rect 87272 35334 87274 35386
rect 87454 35334 87456 35386
rect 87210 35332 87216 35334
rect 87272 35332 87296 35334
rect 87352 35332 87376 35334
rect 87432 35332 87456 35334
rect 87512 35332 87518 35334
rect 87210 35323 87518 35332
rect 88212 35156 88264 35162
rect 88212 35098 88264 35104
rect 88224 35065 88252 35098
rect 88210 35056 88266 35065
rect 85820 35020 85872 35026
rect 88210 34991 88266 35000
rect 85820 34962 85872 34968
rect 85832 34929 85860 34962
rect 85818 34920 85874 34929
rect 85818 34855 85874 34864
rect 86474 34844 86782 34853
rect 86474 34842 86480 34844
rect 86536 34842 86560 34844
rect 86616 34842 86640 34844
rect 86696 34842 86720 34844
rect 86776 34842 86782 34844
rect 86536 34790 86538 34842
rect 86718 34790 86720 34842
rect 86474 34788 86480 34790
rect 86536 34788 86560 34790
rect 86616 34788 86640 34790
rect 86696 34788 86720 34790
rect 86776 34788 86782 34790
rect 86474 34779 86782 34788
rect 87210 34300 87518 34309
rect 87210 34298 87216 34300
rect 87272 34298 87296 34300
rect 87352 34298 87376 34300
rect 87432 34298 87456 34300
rect 87512 34298 87518 34300
rect 87272 34246 87274 34298
rect 87454 34246 87456 34298
rect 87210 34244 87216 34246
rect 87272 34244 87296 34246
rect 87352 34244 87376 34246
rect 87432 34244 87456 34246
rect 87512 34244 87518 34246
rect 87210 34235 87518 34244
rect 88212 34068 88264 34074
rect 88212 34010 88264 34016
rect 85820 33932 85872 33938
rect 85820 33874 85872 33880
rect 85832 33841 85860 33874
rect 85818 33832 85874 33841
rect 85818 33767 85874 33776
rect 86474 33756 86782 33765
rect 86474 33754 86480 33756
rect 86536 33754 86560 33756
rect 86616 33754 86640 33756
rect 86696 33754 86720 33756
rect 86776 33754 86782 33756
rect 86536 33702 86538 33754
rect 86718 33702 86720 33754
rect 88224 33705 88252 34010
rect 86474 33700 86480 33702
rect 86536 33700 86560 33702
rect 86616 33700 86640 33702
rect 86696 33700 86720 33702
rect 86776 33700 86782 33702
rect 86474 33691 86782 33700
rect 88210 33696 88266 33705
rect 88210 33631 88266 33640
rect 87210 33212 87518 33221
rect 87210 33210 87216 33212
rect 87272 33210 87296 33212
rect 87352 33210 87376 33212
rect 87432 33210 87456 33212
rect 87512 33210 87518 33212
rect 87272 33158 87274 33210
rect 87454 33158 87456 33210
rect 87210 33156 87216 33158
rect 87272 33156 87296 33158
rect 87352 33156 87376 33158
rect 87432 33156 87456 33158
rect 87512 33156 87518 33158
rect 87210 33147 87518 33156
rect 86474 32668 86782 32677
rect 86474 32666 86480 32668
rect 86536 32666 86560 32668
rect 86616 32666 86640 32668
rect 86696 32666 86720 32668
rect 86776 32666 86782 32668
rect 85818 32608 85874 32617
rect 86536 32614 86538 32666
rect 86718 32614 86720 32666
rect 86474 32612 86480 32614
rect 86536 32612 86560 32614
rect 86616 32612 86640 32614
rect 86696 32612 86720 32614
rect 86776 32612 86782 32614
rect 86474 32603 86782 32612
rect 85818 32543 85874 32552
rect 85832 32510 85860 32543
rect 85820 32504 85872 32510
rect 85820 32446 85872 32452
rect 88212 32368 88264 32374
rect 88210 32336 88212 32345
rect 88264 32336 88266 32345
rect 88210 32271 88266 32280
rect 87210 32124 87518 32133
rect 87210 32122 87216 32124
rect 87272 32122 87296 32124
rect 87352 32122 87376 32124
rect 87432 32122 87456 32124
rect 87512 32122 87518 32124
rect 87272 32070 87274 32122
rect 87454 32070 87456 32122
rect 87210 32068 87216 32070
rect 87272 32068 87296 32070
rect 87352 32068 87376 32070
rect 87432 32068 87456 32070
rect 87512 32068 87518 32070
rect 87210 32059 87518 32068
rect 88212 31892 88264 31898
rect 88212 31834 88264 31840
rect 85820 31756 85872 31762
rect 85820 31698 85872 31704
rect 85832 31665 85860 31698
rect 88224 31665 88252 31834
rect 85818 31656 85874 31665
rect 85818 31591 85874 31600
rect 88210 31656 88266 31665
rect 88210 31591 88266 31600
rect 86474 31580 86782 31589
rect 86474 31578 86480 31580
rect 86536 31578 86560 31580
rect 86616 31578 86640 31580
rect 86696 31578 86720 31580
rect 86776 31578 86782 31580
rect 86536 31526 86538 31578
rect 86718 31526 86720 31578
rect 86474 31524 86480 31526
rect 86536 31524 86560 31526
rect 86616 31524 86640 31526
rect 86696 31524 86720 31526
rect 86776 31524 86782 31526
rect 86474 31515 86782 31524
rect 87210 31036 87518 31045
rect 87210 31034 87216 31036
rect 87272 31034 87296 31036
rect 87352 31034 87376 31036
rect 87432 31034 87456 31036
rect 87512 31034 87518 31036
rect 87272 30982 87274 31034
rect 87454 30982 87456 31034
rect 87210 30980 87216 30982
rect 87272 30980 87296 30982
rect 87352 30980 87376 30982
rect 87432 30980 87456 30982
rect 87512 30980 87518 30982
rect 87210 30971 87518 30980
rect 88580 30804 88632 30810
rect 88580 30746 88632 30752
rect 86474 30492 86782 30501
rect 86474 30490 86480 30492
rect 86536 30490 86560 30492
rect 86616 30490 86640 30492
rect 86696 30490 86720 30492
rect 86776 30490 86782 30492
rect 86536 30438 86538 30490
rect 86718 30438 86720 30490
rect 86474 30436 86480 30438
rect 86536 30436 86560 30438
rect 86616 30436 86640 30438
rect 86696 30436 86720 30438
rect 86776 30436 86782 30438
rect 86474 30427 86782 30436
rect 88592 30305 88620 30746
rect 88578 30296 88634 30305
rect 88578 30231 88634 30240
rect 87210 29948 87518 29957
rect 87210 29946 87216 29948
rect 87272 29946 87296 29948
rect 87352 29946 87376 29948
rect 87432 29946 87456 29948
rect 87512 29946 87518 29948
rect 87272 29894 87274 29946
rect 87454 29894 87456 29946
rect 87210 29892 87216 29894
rect 87272 29892 87296 29894
rect 87352 29892 87376 29894
rect 87432 29892 87456 29894
rect 87512 29892 87518 29894
rect 87210 29883 87518 29892
rect 85820 29716 85872 29722
rect 85820 29658 85872 29664
rect 85832 29489 85860 29658
rect 88394 29616 88450 29625
rect 88394 29551 88450 29560
rect 88408 29518 88436 29551
rect 88396 29512 88448 29518
rect 85818 29480 85874 29489
rect 88396 29454 88448 29460
rect 85818 29415 85874 29424
rect 86474 29404 86782 29413
rect 86474 29402 86480 29404
rect 86536 29402 86560 29404
rect 86616 29402 86640 29404
rect 86696 29402 86720 29404
rect 86776 29402 86782 29404
rect 86536 29350 86538 29402
rect 86718 29350 86720 29402
rect 86474 29348 86480 29350
rect 86536 29348 86560 29350
rect 86616 29348 86640 29350
rect 86696 29348 86720 29350
rect 86776 29348 86782 29350
rect 86474 29339 86782 29348
rect 87210 28860 87518 28869
rect 87210 28858 87216 28860
rect 87272 28858 87296 28860
rect 87352 28858 87376 28860
rect 87432 28858 87456 28860
rect 87512 28858 87518 28860
rect 87272 28806 87274 28858
rect 87454 28806 87456 28858
rect 87210 28804 87216 28806
rect 87272 28804 87296 28806
rect 87352 28804 87376 28806
rect 87432 28804 87456 28806
rect 87512 28804 87518 28806
rect 87210 28795 87518 28804
rect 85820 28628 85872 28634
rect 85820 28570 85872 28576
rect 85832 28401 85860 28570
rect 88212 28424 88264 28430
rect 85818 28392 85874 28401
rect 88212 28366 88264 28372
rect 85818 28327 85874 28336
rect 86474 28316 86782 28325
rect 86474 28314 86480 28316
rect 86536 28314 86560 28316
rect 86616 28314 86640 28316
rect 86696 28314 86720 28316
rect 86776 28314 86782 28316
rect 86536 28262 86538 28314
rect 86718 28262 86720 28314
rect 88224 28265 88252 28366
rect 86474 28260 86480 28262
rect 86536 28260 86560 28262
rect 86616 28260 86640 28262
rect 86696 28260 86720 28262
rect 86776 28260 86782 28262
rect 86474 28251 86782 28260
rect 88210 28256 88266 28265
rect 88210 28191 88266 28200
rect 87210 27772 87518 27781
rect 87210 27770 87216 27772
rect 87272 27770 87296 27772
rect 87352 27770 87376 27772
rect 87432 27770 87456 27772
rect 87512 27770 87518 27772
rect 87272 27718 87274 27770
rect 87454 27718 87456 27770
rect 87210 27716 87216 27718
rect 87272 27716 87296 27718
rect 87352 27716 87376 27718
rect 87432 27716 87456 27718
rect 87512 27716 87518 27718
rect 87210 27707 87518 27716
rect 86474 27228 86782 27237
rect 86474 27226 86480 27228
rect 86536 27226 86560 27228
rect 86616 27226 86640 27228
rect 86696 27226 86720 27228
rect 86776 27226 86782 27228
rect 85818 27168 85874 27177
rect 86536 27174 86538 27226
rect 86718 27174 86720 27226
rect 86474 27172 86480 27174
rect 86536 27172 86560 27174
rect 86616 27172 86640 27174
rect 86696 27172 86720 27174
rect 86776 27172 86782 27174
rect 86474 27163 86782 27172
rect 85818 27103 85874 27112
rect 85832 26934 85860 27103
rect 85820 26928 85872 26934
rect 85820 26870 85872 26876
rect 88394 26896 88450 26905
rect 88394 26831 88450 26840
rect 88408 26798 88436 26831
rect 88396 26792 88448 26798
rect 88396 26734 88448 26740
rect 87210 26684 87518 26693
rect 87210 26682 87216 26684
rect 87272 26682 87296 26684
rect 87352 26682 87376 26684
rect 87432 26682 87456 26684
rect 87512 26682 87518 26684
rect 87272 26630 87274 26682
rect 87454 26630 87456 26682
rect 87210 26628 87216 26630
rect 87272 26628 87296 26630
rect 87352 26628 87376 26630
rect 87432 26628 87456 26630
rect 87512 26628 87518 26630
rect 87210 26619 87518 26628
rect 87568 26452 87620 26458
rect 87568 26394 87620 26400
rect 87580 26361 87608 26394
rect 87566 26352 87622 26361
rect 87566 26287 87622 26296
rect 88212 26248 88264 26254
rect 88210 26216 88212 26225
rect 88264 26216 88266 26225
rect 88210 26151 88266 26160
rect 86474 26140 86782 26149
rect 86474 26138 86480 26140
rect 86536 26138 86560 26140
rect 86616 26138 86640 26140
rect 86696 26138 86720 26140
rect 86776 26138 86782 26140
rect 86536 26086 86538 26138
rect 86718 26086 86720 26138
rect 86474 26084 86480 26086
rect 86536 26084 86560 26086
rect 86616 26084 86640 26086
rect 86696 26084 86720 26086
rect 86776 26084 86782 26086
rect 86474 26075 86782 26084
rect 87210 25596 87518 25605
rect 87210 25594 87216 25596
rect 87272 25594 87296 25596
rect 87352 25594 87376 25596
rect 87432 25594 87456 25596
rect 87512 25594 87518 25596
rect 87272 25542 87274 25594
rect 87454 25542 87456 25594
rect 87210 25540 87216 25542
rect 87272 25540 87296 25542
rect 87352 25540 87376 25542
rect 87432 25540 87456 25542
rect 87512 25540 87518 25542
rect 87210 25531 87518 25540
rect 88580 25160 88632 25166
rect 88580 25102 88632 25108
rect 86474 25052 86782 25061
rect 86474 25050 86480 25052
rect 86536 25050 86560 25052
rect 86616 25050 86640 25052
rect 86696 25050 86720 25052
rect 86776 25050 86782 25052
rect 86536 24998 86538 25050
rect 86718 24998 86720 25050
rect 86474 24996 86480 24998
rect 86536 24996 86560 24998
rect 86616 24996 86640 24998
rect 86696 24996 86720 24998
rect 86776 24996 86782 24998
rect 86474 24987 86782 24996
rect 88592 24865 88620 25102
rect 88578 24856 88634 24865
rect 88578 24791 88634 24800
rect 87210 24508 87518 24517
rect 87210 24506 87216 24508
rect 87272 24506 87296 24508
rect 87352 24506 87376 24508
rect 87432 24506 87456 24508
rect 87512 24506 87518 24508
rect 87272 24454 87274 24506
rect 87454 24454 87456 24506
rect 87210 24452 87216 24454
rect 87272 24452 87296 24454
rect 87352 24452 87376 24454
rect 87432 24452 87456 24454
rect 87512 24452 87518 24454
rect 87210 24443 87518 24452
rect 87568 24276 87620 24282
rect 87568 24218 87620 24224
rect 87580 24185 87608 24218
rect 87566 24176 87622 24185
rect 87566 24111 87622 24120
rect 88486 24176 88542 24185
rect 88486 24111 88488 24120
rect 88540 24111 88542 24120
rect 88488 24082 88540 24088
rect 86474 23964 86782 23973
rect 86474 23962 86480 23964
rect 86536 23962 86560 23964
rect 86616 23962 86640 23964
rect 86696 23962 86720 23964
rect 86776 23962 86782 23964
rect 86536 23910 86538 23962
rect 86718 23910 86720 23962
rect 86474 23908 86480 23910
rect 86536 23908 86560 23910
rect 86616 23908 86640 23910
rect 86696 23908 86720 23910
rect 86776 23908 86782 23910
rect 86474 23899 86782 23908
rect 87210 23420 87518 23429
rect 87210 23418 87216 23420
rect 87272 23418 87296 23420
rect 87352 23418 87376 23420
rect 87432 23418 87456 23420
rect 87512 23418 87518 23420
rect 87272 23366 87274 23418
rect 87454 23366 87456 23418
rect 87210 23364 87216 23366
rect 87272 23364 87296 23366
rect 87352 23364 87376 23366
rect 87432 23364 87456 23366
rect 87512 23364 87518 23366
rect 87210 23355 87518 23364
rect 85820 23188 85872 23194
rect 85820 23130 85872 23136
rect 85832 22961 85860 23130
rect 88212 22984 88264 22990
rect 85818 22952 85874 22961
rect 88212 22926 88264 22932
rect 85818 22887 85874 22896
rect 86474 22876 86782 22885
rect 86474 22874 86480 22876
rect 86536 22874 86560 22876
rect 86616 22874 86640 22876
rect 86696 22874 86720 22876
rect 86776 22874 86782 22876
rect 86536 22822 86538 22874
rect 86718 22822 86720 22874
rect 88224 22825 88252 22926
rect 86474 22820 86480 22822
rect 86536 22820 86560 22822
rect 86616 22820 86640 22822
rect 86696 22820 86720 22822
rect 86776 22820 86782 22822
rect 86474 22811 86782 22820
rect 88210 22816 88266 22825
rect 88210 22751 88266 22760
rect 87210 22332 87518 22341
rect 87210 22330 87216 22332
rect 87272 22330 87296 22332
rect 87352 22330 87376 22332
rect 87432 22330 87456 22332
rect 87512 22330 87518 22332
rect 87272 22278 87274 22330
rect 87454 22278 87456 22330
rect 87210 22276 87216 22278
rect 87272 22276 87296 22278
rect 87352 22276 87376 22278
rect 87432 22276 87456 22278
rect 87512 22276 87518 22278
rect 87210 22267 87518 22276
rect 86474 21788 86782 21797
rect 86474 21786 86480 21788
rect 86536 21786 86560 21788
rect 86616 21786 86640 21788
rect 86696 21786 86720 21788
rect 86776 21786 86782 21788
rect 85818 21728 85874 21737
rect 86536 21734 86538 21786
rect 86718 21734 86720 21786
rect 86474 21732 86480 21734
rect 86536 21732 86560 21734
rect 86616 21732 86640 21734
rect 86696 21732 86720 21734
rect 86776 21732 86782 21734
rect 86474 21723 86782 21732
rect 85818 21663 85874 21672
rect 85832 21494 85860 21663
rect 85820 21488 85872 21494
rect 85820 21430 85872 21436
rect 88394 21456 88450 21465
rect 88394 21391 88450 21400
rect 88408 21358 88436 21391
rect 88396 21352 88448 21358
rect 88396 21294 88448 21300
rect 87210 21244 87518 21253
rect 87210 21242 87216 21244
rect 87272 21242 87296 21244
rect 87352 21242 87376 21244
rect 87432 21242 87456 21244
rect 87512 21242 87518 21244
rect 87272 21190 87274 21242
rect 87454 21190 87456 21242
rect 87210 21188 87216 21190
rect 87272 21188 87296 21190
rect 87352 21188 87376 21190
rect 87432 21188 87456 21190
rect 87512 21188 87518 21190
rect 87210 21179 87518 21188
rect 88580 21080 88632 21086
rect 88580 21022 88632 21028
rect 88592 20785 88620 21022
rect 88578 20776 88634 20785
rect 88578 20711 88634 20720
rect 86474 20700 86782 20709
rect 86474 20698 86480 20700
rect 86536 20698 86560 20700
rect 86616 20698 86640 20700
rect 86696 20698 86720 20700
rect 86776 20698 86782 20700
rect 86536 20646 86538 20698
rect 86718 20646 86720 20698
rect 86474 20644 86480 20646
rect 86536 20644 86560 20646
rect 86616 20644 86640 20646
rect 86696 20644 86720 20646
rect 86776 20644 86782 20646
rect 86474 20635 86782 20644
rect 87210 20156 87518 20165
rect 87210 20154 87216 20156
rect 87272 20154 87296 20156
rect 87352 20154 87376 20156
rect 87432 20154 87456 20156
rect 87512 20154 87518 20156
rect 87272 20102 87274 20154
rect 87454 20102 87456 20154
rect 87210 20100 87216 20102
rect 87272 20100 87296 20102
rect 87352 20100 87376 20102
rect 87432 20100 87456 20102
rect 87512 20100 87518 20102
rect 87210 20091 87518 20100
rect 87568 19924 87620 19930
rect 87568 19866 87620 19872
rect 87580 19833 87608 19866
rect 87566 19824 87622 19833
rect 87566 19759 87622 19768
rect 88672 19720 88724 19726
rect 88672 19662 88724 19668
rect 86474 19612 86782 19621
rect 86474 19610 86480 19612
rect 86536 19610 86560 19612
rect 86616 19610 86640 19612
rect 86696 19610 86720 19612
rect 86776 19610 86782 19612
rect 86536 19558 86538 19610
rect 86718 19558 86720 19610
rect 86474 19556 86480 19558
rect 86536 19556 86560 19558
rect 86616 19556 86640 19558
rect 86696 19556 86720 19558
rect 86776 19556 86782 19558
rect 86474 19547 86782 19556
rect 88684 19425 88712 19662
rect 88670 19416 88726 19425
rect 88670 19351 88726 19360
rect 87210 19068 87518 19077
rect 87210 19066 87216 19068
rect 87272 19066 87296 19068
rect 87352 19066 87376 19068
rect 87432 19066 87456 19068
rect 87512 19066 87518 19068
rect 87272 19014 87274 19066
rect 87454 19014 87456 19066
rect 87210 19012 87216 19014
rect 87272 19012 87296 19014
rect 87352 19012 87376 19014
rect 87432 19012 87456 19014
rect 87512 19012 87518 19014
rect 87210 19003 87518 19012
rect 87292 18836 87344 18842
rect 87292 18778 87344 18784
rect 87304 18745 87332 18778
rect 87290 18736 87346 18745
rect 87290 18671 87346 18680
rect 88210 18736 88266 18745
rect 88210 18671 88212 18680
rect 88264 18671 88266 18680
rect 88212 18642 88264 18648
rect 86474 18524 86782 18533
rect 86474 18522 86480 18524
rect 86536 18522 86560 18524
rect 86616 18522 86640 18524
rect 86696 18522 86720 18524
rect 86776 18522 86782 18524
rect 86536 18470 86538 18522
rect 86718 18470 86720 18522
rect 86474 18468 86480 18470
rect 86536 18468 86560 18470
rect 86616 18468 86640 18470
rect 86696 18468 86720 18470
rect 86776 18468 86782 18470
rect 86474 18459 86782 18468
rect 87210 17980 87518 17989
rect 87210 17978 87216 17980
rect 87272 17978 87296 17980
rect 87352 17978 87376 17980
rect 87432 17978 87456 17980
rect 87512 17978 87518 17980
rect 87272 17926 87274 17978
rect 87454 17926 87456 17978
rect 87210 17924 87216 17926
rect 87272 17924 87296 17926
rect 87352 17924 87376 17926
rect 87432 17924 87456 17926
rect 87512 17924 87518 17926
rect 87210 17915 87518 17924
rect 85820 17748 85872 17754
rect 85820 17690 85872 17696
rect 85832 17521 85860 17690
rect 88212 17544 88264 17550
rect 85818 17512 85874 17521
rect 88212 17486 88264 17492
rect 85818 17447 85874 17456
rect 86474 17436 86782 17445
rect 86474 17434 86480 17436
rect 86536 17434 86560 17436
rect 86616 17434 86640 17436
rect 86696 17434 86720 17436
rect 86776 17434 86782 17436
rect 86536 17382 86538 17434
rect 86718 17382 86720 17434
rect 88224 17385 88252 17486
rect 86474 17380 86480 17382
rect 86536 17380 86560 17382
rect 86616 17380 86640 17382
rect 86696 17380 86720 17382
rect 86776 17380 86782 17382
rect 86474 17371 86782 17380
rect 88210 17376 88266 17385
rect 88210 17311 88266 17320
rect 87210 16892 87518 16901
rect 87210 16890 87216 16892
rect 87272 16890 87296 16892
rect 87352 16890 87376 16892
rect 87432 16890 87456 16892
rect 87512 16890 87518 16892
rect 87272 16838 87274 16890
rect 87454 16838 87456 16890
rect 87210 16836 87216 16838
rect 87272 16836 87296 16838
rect 87352 16836 87376 16838
rect 87432 16836 87456 16838
rect 87512 16836 87518 16838
rect 87210 16827 87518 16836
rect 86474 16348 86782 16357
rect 86474 16346 86480 16348
rect 86536 16346 86560 16348
rect 86616 16346 86640 16348
rect 86696 16346 86720 16348
rect 86776 16346 86782 16348
rect 85818 16288 85874 16297
rect 86536 16294 86538 16346
rect 86718 16294 86720 16346
rect 86474 16292 86480 16294
rect 86536 16292 86560 16294
rect 86616 16292 86640 16294
rect 86696 16292 86720 16294
rect 86776 16292 86782 16294
rect 86474 16283 86782 16292
rect 85818 16223 85874 16232
rect 85832 16054 85860 16223
rect 85820 16048 85872 16054
rect 85820 15990 85872 15996
rect 88210 16016 88266 16025
rect 88210 15951 88266 15960
rect 88224 15918 88252 15951
rect 88212 15912 88264 15918
rect 88212 15854 88264 15860
rect 87210 15804 87518 15813
rect 87210 15802 87216 15804
rect 87272 15802 87296 15804
rect 87352 15802 87376 15804
rect 87432 15802 87456 15804
rect 87512 15802 87518 15804
rect 87272 15750 87274 15802
rect 87454 15750 87456 15802
rect 87210 15748 87216 15750
rect 87272 15748 87296 15750
rect 87352 15748 87376 15750
rect 87432 15748 87456 15750
rect 87512 15748 87518 15750
rect 87210 15739 87518 15748
rect 88580 15640 88632 15646
rect 88580 15582 88632 15588
rect 88592 15345 88620 15582
rect 88578 15336 88634 15345
rect 88578 15271 88634 15280
rect 86474 15260 86782 15269
rect 86474 15258 86480 15260
rect 86536 15258 86560 15260
rect 86616 15258 86640 15260
rect 86696 15258 86720 15260
rect 86776 15258 86782 15260
rect 86536 15206 86538 15258
rect 86718 15206 86720 15258
rect 86474 15204 86480 15206
rect 86536 15204 86560 15206
rect 86616 15204 86640 15206
rect 86696 15204 86720 15206
rect 86776 15204 86782 15206
rect 86474 15195 86782 15204
rect 85636 15028 85688 15034
rect 85636 14970 85688 14976
rect 85648 14286 85676 14970
rect 88028 14824 88080 14830
rect 88028 14766 88080 14772
rect 87210 14716 87518 14725
rect 87210 14714 87216 14716
rect 87272 14714 87296 14716
rect 87352 14714 87376 14716
rect 87432 14714 87456 14716
rect 87512 14714 87518 14716
rect 87272 14662 87274 14714
rect 87454 14662 87456 14714
rect 88040 14665 88068 14766
rect 87210 14660 87216 14662
rect 87272 14660 87296 14662
rect 87352 14660 87376 14662
rect 87432 14660 87456 14662
rect 87512 14660 87518 14662
rect 87210 14651 87518 14660
rect 88026 14656 88082 14665
rect 88026 14591 88082 14600
rect 85636 14280 85688 14286
rect 85636 14222 85688 14228
rect 86474 14172 86782 14181
rect 86474 14170 86480 14172
rect 86536 14170 86560 14172
rect 86616 14170 86640 14172
rect 86696 14170 86720 14172
rect 86776 14170 86782 14172
rect 86536 14118 86538 14170
rect 86718 14118 86720 14170
rect 86474 14116 86480 14118
rect 86536 14116 86560 14118
rect 86616 14116 86640 14118
rect 86696 14116 86720 14118
rect 86776 14116 86782 14118
rect 86474 14107 86782 14116
rect 87210 13628 87518 13637
rect 87210 13626 87216 13628
rect 87272 13626 87296 13628
rect 87352 13626 87376 13628
rect 87432 13626 87456 13628
rect 87512 13626 87518 13628
rect 87272 13574 87274 13626
rect 87454 13574 87456 13626
rect 87210 13572 87216 13574
rect 87272 13572 87296 13574
rect 87352 13572 87376 13574
rect 87432 13572 87456 13574
rect 87512 13572 87518 13574
rect 87210 13563 87518 13572
rect 85544 13464 85596 13470
rect 85544 13406 85596 13412
rect 88212 13396 88264 13402
rect 88212 13338 88264 13344
rect 87936 13328 87988 13334
rect 88224 13305 88252 13338
rect 87936 13270 87988 13276
rect 88210 13296 88266 13305
rect 86474 13084 86782 13093
rect 86474 13082 86480 13084
rect 86536 13082 86560 13084
rect 86616 13082 86640 13084
rect 86696 13082 86720 13084
rect 86776 13082 86782 13084
rect 86536 13030 86538 13082
rect 86718 13030 86720 13082
rect 86474 13028 86480 13030
rect 86536 13028 86560 13030
rect 86616 13028 86640 13030
rect 86696 13028 86720 13030
rect 86776 13028 86782 13030
rect 86474 13019 86782 13028
rect 87948 12926 87976 13270
rect 88210 13231 88266 13240
rect 87936 12920 87988 12926
rect 87936 12862 87988 12868
rect 87568 12716 87620 12722
rect 87568 12658 87620 12664
rect 88580 12716 88632 12722
rect 88580 12658 88632 12664
rect 85360 12648 85412 12654
rect 85360 12590 85412 12596
rect 85372 12382 85400 12590
rect 87210 12540 87518 12549
rect 87210 12538 87216 12540
rect 87272 12538 87296 12540
rect 87352 12538 87376 12540
rect 87432 12538 87456 12540
rect 87512 12538 87518 12540
rect 87272 12486 87274 12538
rect 87454 12486 87456 12538
rect 87210 12484 87216 12486
rect 87272 12484 87296 12486
rect 87352 12484 87376 12486
rect 87432 12484 87456 12486
rect 87512 12484 87518 12486
rect 87210 12475 87518 12484
rect 87580 12382 87608 12658
rect 88592 12625 88620 12658
rect 88578 12616 88634 12625
rect 88578 12551 88634 12560
rect 83612 12376 83664 12382
rect 83612 12318 83664 12324
rect 85360 12376 85412 12382
rect 85360 12318 85412 12324
rect 87568 12376 87620 12382
rect 87568 12318 87620 12324
rect 83624 12013 83652 12318
rect 83610 12004 83666 12013
rect 83610 11939 83666 11948
rect 86474 11996 86782 12005
rect 86474 11994 86480 11996
rect 86536 11994 86560 11996
rect 86616 11994 86640 11996
rect 86696 11994 86720 11996
rect 86776 11994 86782 11996
rect 86536 11942 86538 11994
rect 86718 11942 86720 11994
rect 86474 11940 86480 11942
rect 86536 11940 86560 11942
rect 86616 11940 86640 11942
rect 86696 11940 86720 11942
rect 86776 11940 86782 11942
rect 83520 7344 83572 7350
rect 83520 7286 83572 7292
rect 83336 7276 83388 7282
rect 83336 7218 83388 7224
rect 83624 7214 83652 11939
rect 86474 11931 86782 11940
rect 87210 11452 87518 11461
rect 87210 11450 87216 11452
rect 87272 11450 87296 11452
rect 87352 11450 87376 11452
rect 87432 11450 87456 11452
rect 87512 11450 87518 11452
rect 87272 11398 87274 11450
rect 87454 11398 87456 11450
rect 87210 11396 87216 11398
rect 87272 11396 87296 11398
rect 87352 11396 87376 11398
rect 87432 11396 87456 11398
rect 87512 11396 87518 11398
rect 87210 11387 87518 11396
rect 86474 10908 86782 10917
rect 86474 10906 86480 10908
rect 86536 10906 86560 10908
rect 86616 10906 86640 10908
rect 86696 10906 86720 10908
rect 86776 10906 86782 10908
rect 86536 10854 86538 10906
rect 86718 10854 86720 10906
rect 86474 10852 86480 10854
rect 86536 10852 86560 10854
rect 86616 10852 86640 10854
rect 86696 10852 86720 10854
rect 86776 10852 86782 10854
rect 86474 10843 86782 10852
rect 88212 10608 88264 10614
rect 88210 10576 88212 10585
rect 88264 10576 88266 10585
rect 88210 10511 88266 10520
rect 87210 10364 87518 10373
rect 87210 10362 87216 10364
rect 87272 10362 87296 10364
rect 87352 10362 87376 10364
rect 87432 10362 87456 10364
rect 87512 10362 87518 10364
rect 87272 10310 87274 10362
rect 87454 10310 87456 10362
rect 87210 10308 87216 10310
rect 87272 10308 87296 10310
rect 87352 10308 87376 10310
rect 87432 10308 87456 10310
rect 87512 10308 87518 10310
rect 87210 10299 87518 10308
rect 86474 9820 86782 9829
rect 86474 9818 86480 9820
rect 86536 9818 86560 9820
rect 86616 9818 86640 9820
rect 86696 9818 86720 9820
rect 86776 9818 86782 9820
rect 86536 9766 86538 9818
rect 86718 9766 86720 9818
rect 86474 9764 86480 9766
rect 86536 9764 86560 9766
rect 86616 9764 86640 9766
rect 86696 9764 86720 9766
rect 86776 9764 86782 9766
rect 86474 9755 86782 9764
rect 87210 9276 87518 9285
rect 87210 9274 87216 9276
rect 87272 9274 87296 9276
rect 87352 9274 87376 9276
rect 87432 9274 87456 9276
rect 87512 9274 87518 9276
rect 87272 9222 87274 9274
rect 87454 9222 87456 9274
rect 87210 9220 87216 9222
rect 87272 9220 87296 9222
rect 87352 9220 87376 9222
rect 87432 9220 87456 9222
rect 87512 9220 87518 9222
rect 87210 9211 87518 9220
rect 86474 8732 86782 8741
rect 86474 8730 86480 8732
rect 86536 8730 86560 8732
rect 86616 8730 86640 8732
rect 86696 8730 86720 8732
rect 86776 8730 86782 8732
rect 86536 8678 86538 8730
rect 86718 8678 86720 8730
rect 86474 8676 86480 8678
rect 86536 8676 86560 8678
rect 86616 8676 86640 8678
rect 86696 8676 86720 8678
rect 86776 8676 86782 8678
rect 86474 8667 86782 8676
rect 87210 8188 87518 8197
rect 87210 8186 87216 8188
rect 87272 8186 87296 8188
rect 87352 8186 87376 8188
rect 87432 8186 87456 8188
rect 87512 8186 87518 8188
rect 87272 8134 87274 8186
rect 87454 8134 87456 8186
rect 87210 8132 87216 8134
rect 87272 8132 87296 8134
rect 87352 8132 87376 8134
rect 87432 8132 87456 8134
rect 87512 8132 87518 8134
rect 87210 8123 87518 8132
rect 86474 7644 86782 7653
rect 86474 7642 86480 7644
rect 86536 7642 86560 7644
rect 86616 7642 86640 7644
rect 86696 7642 86720 7644
rect 86776 7642 86782 7644
rect 86536 7590 86538 7642
rect 86718 7590 86720 7642
rect 86474 7588 86480 7590
rect 86536 7588 86560 7590
rect 86616 7588 86640 7590
rect 86696 7588 86720 7590
rect 86776 7588 86782 7590
rect 86474 7579 86782 7588
rect 83612 7208 83664 7214
rect 83612 7150 83664 7156
rect 87210 7100 87518 7109
rect 87210 7098 87216 7100
rect 87272 7098 87296 7100
rect 87352 7098 87376 7100
rect 87432 7098 87456 7100
rect 87512 7098 87518 7100
rect 87272 7046 87274 7098
rect 87454 7046 87456 7098
rect 87210 7044 87216 7046
rect 87272 7044 87296 7046
rect 87352 7044 87376 7046
rect 87432 7044 87456 7046
rect 87512 7044 87518 7046
rect 87210 7035 87518 7044
rect 68064 5304 68116 5310
rect 68064 5246 68116 5252
rect 68984 5304 69036 5310
rect 68984 5246 69036 5252
rect 69996 5304 70048 5310
rect 69996 5246 70048 5252
rect 71284 5304 71336 5310
rect 71284 5246 71336 5252
rect 72572 5304 72624 5310
rect 72572 5246 72624 5252
rect 73400 5304 73452 5310
rect 73400 5246 73452 5252
rect 74504 5304 74556 5310
rect 74504 5246 74556 5252
rect 75792 5304 75844 5310
rect 75792 5246 75844 5252
rect 76712 5304 76764 5310
rect 76712 5246 76764 5252
rect 77724 5304 77776 5310
rect 77724 5246 77776 5252
rect 79012 5304 79064 5310
rect 79012 5246 79064 5252
rect 80116 5304 80168 5310
rect 80116 5246 80168 5252
rect 81128 5304 81180 5310
rect 81128 5246 81180 5252
rect 14980 5168 15032 5174
rect 14980 5110 15032 5116
rect 16176 5168 16228 5174
rect 16176 5110 16228 5116
rect 17188 5168 17240 5174
rect 17188 5110 17240 5116
rect 18292 5168 18344 5174
rect 18292 5110 18344 5116
rect 19396 5168 19448 5174
rect 19396 5110 19448 5116
rect 20500 5168 20552 5174
rect 20500 5110 20552 5116
rect 21604 5168 21656 5174
rect 21604 5110 21656 5116
rect 22708 5168 22760 5174
rect 22708 5110 22760 5116
rect 23904 5168 23956 5174
rect 23904 5110 23956 5116
rect 24916 5168 24968 5174
rect 24916 5110 24968 5116
rect 26020 5168 26072 5174
rect 26020 5110 26072 5116
rect 27124 5168 27176 5174
rect 27124 5110 27176 5116
rect 28228 5168 28280 5174
rect 28228 5110 28280 5116
rect 29332 5168 29384 5174
rect 29332 5110 29384 5116
rect 30712 5168 30764 5174
rect 30712 5110 30764 5116
rect 31356 5168 31408 5174
rect 31356 5110 31408 5116
rect 32644 5168 32696 5174
rect 32644 5110 32696 5116
rect 33932 5168 33984 5174
rect 33932 5110 33984 5116
rect 34576 5168 34628 5174
rect 34576 5110 34628 5116
rect 35864 5168 35916 5174
rect 35864 5110 35916 5116
rect 37152 5168 37204 5174
rect 37152 5110 37204 5116
rect 38440 5168 38492 5174
rect 38440 5110 38492 5116
rect 39084 5168 39136 5174
rect 39084 5110 39136 5116
rect 40372 5168 40424 5174
rect 40372 5110 40424 5116
rect 41660 5168 41712 5174
rect 41660 5110 41712 5116
rect 42304 5168 42356 5174
rect 42304 5110 42356 5116
rect 43592 5168 43644 5174
rect 43592 5110 43644 5116
rect 44880 5168 44932 5174
rect 44880 5110 44932 5116
rect 52608 5168 52660 5174
rect 52608 5110 52660 5116
rect 53528 5168 53580 5174
rect 53528 5110 53580 5116
rect 54448 5168 54500 5174
rect 54448 5110 54500 5116
rect 55828 5168 55880 5174
rect 55828 5110 55880 5116
rect 57024 5168 57076 5174
rect 57024 5110 57076 5116
rect 58036 5168 58088 5174
rect 58036 5110 58088 5116
rect 59048 5168 59100 5174
rect 59048 5110 59100 5116
rect 60336 5168 60388 5174
rect 60336 5110 60388 5116
rect 61256 5168 61308 5174
rect 61256 5110 61308 5116
rect 62360 5168 62412 5174
rect 62360 5110 62412 5116
rect 63556 5168 63608 5174
rect 63556 5110 63608 5116
rect 64752 5168 64804 5174
rect 64752 5110 64804 5116
rect 65764 5168 65816 5174
rect 65764 5110 65816 5116
rect 66776 5168 66828 5174
rect 66776 5110 66828 5116
rect 68064 5168 68116 5174
rect 68064 5110 68116 5116
rect 68708 5168 68760 5174
rect 68708 5110 68760 5116
rect 69996 5168 70048 5174
rect 69996 5110 70048 5116
rect 71284 5168 71336 5174
rect 71284 5110 71336 5116
rect 72572 5168 72624 5174
rect 72572 5110 72624 5116
rect 73216 5168 73268 5174
rect 73216 5110 73268 5116
rect 74504 5168 74556 5174
rect 74504 5110 74556 5116
rect 75792 5168 75844 5174
rect 75792 5110 75844 5116
rect 76436 5168 76488 5174
rect 76436 5110 76488 5116
rect 77724 5168 77776 5174
rect 77724 5110 77776 5116
rect 79012 5168 79064 5174
rect 79012 5110 79064 5116
rect 80300 5168 80352 5174
rect 80300 5110 80352 5116
rect 80944 5168 80996 5174
rect 80944 5110 80996 5116
rect 15256 5032 15308 5038
rect 15256 4974 15308 4980
rect 15900 5032 15952 5038
rect 15900 4974 15952 4980
rect 17188 5032 17240 5038
rect 17188 4974 17240 4980
rect 18752 5032 18804 5038
rect 18752 4974 18804 4980
rect 19120 5032 19172 5038
rect 19120 4974 19172 4980
rect 20408 5032 20460 5038
rect 20408 4974 20460 4980
rect 21696 5032 21748 5038
rect 21696 4974 21748 4980
rect 22984 5032 23036 5038
rect 22984 4974 23036 4980
rect 23628 5032 23680 5038
rect 23628 4974 23680 4980
rect 24916 5032 24968 5038
rect 24916 4974 24968 4980
rect 26204 5032 26256 5038
rect 26204 4974 26256 4980
rect 26848 5032 26900 5038
rect 26848 4974 26900 4980
rect 28136 5032 28188 5038
rect 28136 4974 28188 4980
rect 29424 5032 29476 5038
rect 29424 4974 29476 4980
rect 15268 3800 15296 4974
rect 15912 3800 15940 4974
rect 17200 3800 17228 4974
rect 18382 4924 18690 4933
rect 18382 4922 18388 4924
rect 18444 4922 18468 4924
rect 18524 4922 18548 4924
rect 18604 4922 18628 4924
rect 18684 4922 18690 4924
rect 18444 4870 18446 4922
rect 18626 4870 18628 4922
rect 18382 4868 18388 4870
rect 18444 4868 18468 4870
rect 18524 4868 18548 4870
rect 18604 4868 18628 4870
rect 18684 4868 18690 4870
rect 18382 4859 18690 4868
rect 18488 3870 18608 3898
rect 18488 3800 18516 3870
rect 3018 3000 3074 3800
rect 3662 3000 3718 3800
rect 4306 3000 4362 3800
rect 4950 3000 5006 3800
rect 5594 3000 5650 3800
rect 6238 3000 6294 3800
rect 6882 3000 6938 3800
rect 7526 3000 7582 3800
rect 8170 3000 8226 3800
rect 8814 3000 8870 3800
rect 9458 3000 9514 3800
rect 10102 3000 10158 3800
rect 10746 3000 10802 3800
rect 11390 3000 11446 3800
rect 12034 3000 12090 3800
rect 12678 3000 12734 3800
rect 15254 3000 15310 3800
rect 15898 3000 15954 3800
rect 17186 3000 17242 3800
rect 18474 3000 18530 3800
rect 18580 3762 18608 3870
rect 18764 3762 18792 4974
rect 19132 3800 19160 4974
rect 20420 3800 20448 4974
rect 21708 3800 21736 4974
rect 22996 3800 23024 4974
rect 23640 3800 23668 4974
rect 24928 3800 24956 4974
rect 26216 3800 26244 4974
rect 26860 3800 26888 4974
rect 28148 3800 28176 4974
rect 29436 3800 29464 4974
rect 30724 3800 30752 5110
rect 31368 3800 31396 5110
rect 32656 3800 32684 5110
rect 33944 3800 33972 5110
rect 34588 3800 34616 5110
rect 35876 3800 35904 5110
rect 36782 4924 37090 4933
rect 36782 4922 36788 4924
rect 36844 4922 36868 4924
rect 36924 4922 36948 4924
rect 37004 4922 37028 4924
rect 37084 4922 37090 4924
rect 36844 4870 36846 4922
rect 37026 4870 37028 4922
rect 36782 4868 36788 4870
rect 36844 4868 36868 4870
rect 36924 4868 36948 4870
rect 37004 4868 37028 4870
rect 37084 4868 37090 4870
rect 36782 4859 37090 4868
rect 37164 3800 37192 5110
rect 38452 3800 38480 5110
rect 39096 3800 39124 5110
rect 40384 3800 40412 5110
rect 41672 3800 41700 5110
rect 42316 3800 42344 5110
rect 43604 3800 43632 5110
rect 44892 3800 44920 5110
rect 52608 5032 52660 5038
rect 52608 4974 52660 4980
rect 53252 5032 53304 5038
rect 53252 4974 53304 4980
rect 54540 5032 54592 5038
rect 54540 4974 54592 4980
rect 55828 5032 55880 5038
rect 55828 4974 55880 4980
rect 57116 5032 57168 5038
rect 57116 4974 57168 4980
rect 57760 5032 57812 5038
rect 57760 4974 57812 4980
rect 59048 5032 59100 5038
rect 59048 4974 59100 4980
rect 60336 5032 60388 5038
rect 60336 4974 60388 4980
rect 60980 5032 61032 5038
rect 60980 4974 61032 4980
rect 62268 5032 62320 5038
rect 62268 4974 62320 4980
rect 63556 5032 63608 5038
rect 63556 4974 63608 4980
rect 64844 5032 64896 5038
rect 64844 4974 64896 4980
rect 65488 5032 65540 5038
rect 65488 4974 65540 4980
rect 66776 5032 66828 5038
rect 66776 4974 66828 4980
rect 52620 3800 52648 4974
rect 53264 3800 53292 4974
rect 54552 3800 54580 4974
rect 55182 4924 55490 4933
rect 55182 4922 55188 4924
rect 55244 4922 55268 4924
rect 55324 4922 55348 4924
rect 55404 4922 55428 4924
rect 55484 4922 55490 4924
rect 55244 4870 55246 4922
rect 55426 4870 55428 4922
rect 55182 4868 55188 4870
rect 55244 4868 55268 4870
rect 55324 4868 55348 4870
rect 55404 4868 55428 4870
rect 55484 4868 55490 4870
rect 55182 4859 55490 4868
rect 55840 3800 55868 4974
rect 57128 3800 57156 4974
rect 57772 3800 57800 4974
rect 59060 3800 59088 4974
rect 60348 3800 60376 4974
rect 60992 3800 61020 4974
rect 62280 3800 62308 4974
rect 63568 3800 63596 4974
rect 64856 3800 64884 4974
rect 65500 3800 65528 4974
rect 66788 3800 66816 4974
rect 68076 3800 68104 5110
rect 68720 3800 68748 5110
rect 70008 3800 70036 5110
rect 71296 3800 71324 5110
rect 72584 3800 72612 5110
rect 73228 3800 73256 5110
rect 73582 4924 73890 4933
rect 73582 4922 73588 4924
rect 73644 4922 73668 4924
rect 73724 4922 73748 4924
rect 73804 4922 73828 4924
rect 73884 4922 73890 4924
rect 73644 4870 73646 4922
rect 73826 4870 73828 4922
rect 73582 4868 73588 4870
rect 73644 4868 73668 4870
rect 73724 4868 73748 4870
rect 73804 4868 73828 4870
rect 73884 4868 73890 4870
rect 73582 4859 73890 4868
rect 74516 3800 74544 5110
rect 75804 3800 75832 5110
rect 76448 3800 76476 5110
rect 77736 3800 77764 5110
rect 79024 3800 79052 5110
rect 80312 3800 80340 5110
rect 80956 3800 80984 5110
rect 18580 3734 18792 3762
rect 19118 3000 19174 3800
rect 20406 3000 20462 3800
rect 21694 3000 21750 3800
rect 22982 3000 23038 3800
rect 23626 3000 23682 3800
rect 24914 3000 24970 3800
rect 26202 3000 26258 3800
rect 26846 3000 26902 3800
rect 28134 3000 28190 3800
rect 29422 3000 29478 3800
rect 30710 3000 30766 3800
rect 31354 3000 31410 3800
rect 32642 3000 32698 3800
rect 33930 3000 33986 3800
rect 34574 3000 34630 3800
rect 35862 3000 35918 3800
rect 37150 3000 37206 3800
rect 38438 3000 38494 3800
rect 39082 3000 39138 3800
rect 40370 3000 40426 3800
rect 41658 3000 41714 3800
rect 42302 3000 42358 3800
rect 43590 3000 43646 3800
rect 44878 3000 44934 3800
rect 52606 3000 52662 3800
rect 53250 3000 53306 3800
rect 54538 3000 54594 3800
rect 55826 3000 55882 3800
rect 57114 3000 57170 3800
rect 57758 3000 57814 3800
rect 59046 3000 59102 3800
rect 60334 3000 60390 3800
rect 60978 3000 61034 3800
rect 62266 3000 62322 3800
rect 63554 3000 63610 3800
rect 64842 3000 64898 3800
rect 65486 3000 65542 3800
rect 66774 3000 66830 3800
rect 68062 3000 68118 3800
rect 68706 3000 68762 3800
rect 69994 3000 70050 3800
rect 71282 3000 71338 3800
rect 72570 3000 72626 3800
rect 73214 3000 73270 3800
rect 74502 3000 74558 3800
rect 75790 3000 75846 3800
rect 76434 3000 76490 3800
rect 77722 3000 77778 3800
rect 79010 3000 79066 3800
rect 80298 3000 80354 3800
rect 80942 3000 80998 3800
<< via2 >>
rect 18388 87610 18444 87612
rect 18468 87610 18524 87612
rect 18548 87610 18604 87612
rect 18628 87610 18684 87612
rect 18388 87558 18434 87610
rect 18434 87558 18444 87610
rect 18468 87558 18498 87610
rect 18498 87558 18510 87610
rect 18510 87558 18524 87610
rect 18548 87558 18562 87610
rect 18562 87558 18574 87610
rect 18574 87558 18604 87610
rect 18628 87558 18638 87610
rect 18638 87558 18684 87610
rect 18388 87556 18444 87558
rect 18468 87556 18524 87558
rect 18548 87556 18604 87558
rect 18628 87556 18684 87558
rect 5888 84890 5944 84892
rect 5968 84890 6024 84892
rect 6048 84890 6104 84892
rect 6128 84890 6184 84892
rect 5888 84838 5934 84890
rect 5934 84838 5944 84890
rect 5968 84838 5998 84890
rect 5998 84838 6010 84890
rect 6010 84838 6024 84890
rect 6048 84838 6062 84890
rect 6062 84838 6074 84890
rect 6074 84838 6104 84890
rect 6128 84838 6138 84890
rect 6138 84838 6184 84890
rect 5888 84836 5944 84838
rect 5968 84836 6024 84838
rect 6048 84836 6104 84838
rect 6128 84836 6184 84838
rect 6624 84346 6680 84348
rect 6704 84346 6760 84348
rect 6784 84346 6840 84348
rect 6864 84346 6920 84348
rect 6624 84294 6670 84346
rect 6670 84294 6680 84346
rect 6704 84294 6734 84346
rect 6734 84294 6746 84346
rect 6746 84294 6760 84346
rect 6784 84294 6798 84346
rect 6798 84294 6810 84346
rect 6810 84294 6840 84346
rect 6864 84294 6874 84346
rect 6874 84294 6920 84346
rect 6624 84292 6680 84294
rect 6704 84292 6760 84294
rect 6784 84292 6840 84294
rect 6864 84292 6920 84294
rect 5888 83802 5944 83804
rect 5968 83802 6024 83804
rect 6048 83802 6104 83804
rect 6128 83802 6184 83804
rect 5888 83750 5934 83802
rect 5934 83750 5944 83802
rect 5968 83750 5998 83802
rect 5998 83750 6010 83802
rect 6010 83750 6024 83802
rect 6048 83750 6062 83802
rect 6062 83750 6074 83802
rect 6074 83750 6104 83802
rect 6128 83750 6138 83802
rect 6138 83750 6184 83802
rect 5888 83748 5944 83750
rect 5968 83748 6024 83750
rect 6048 83748 6104 83750
rect 6128 83748 6184 83750
rect 6624 83258 6680 83260
rect 6704 83258 6760 83260
rect 6784 83258 6840 83260
rect 6864 83258 6920 83260
rect 6624 83206 6670 83258
rect 6670 83206 6680 83258
rect 6704 83206 6734 83258
rect 6734 83206 6746 83258
rect 6746 83206 6760 83258
rect 6784 83206 6798 83258
rect 6798 83206 6810 83258
rect 6810 83206 6840 83258
rect 6864 83206 6874 83258
rect 6874 83206 6920 83258
rect 6624 83204 6680 83206
rect 6704 83204 6760 83206
rect 6784 83204 6840 83206
rect 6864 83204 6920 83206
rect 5888 82714 5944 82716
rect 5968 82714 6024 82716
rect 6048 82714 6104 82716
rect 6128 82714 6184 82716
rect 5888 82662 5934 82714
rect 5934 82662 5944 82714
rect 5968 82662 5998 82714
rect 5998 82662 6010 82714
rect 6010 82662 6024 82714
rect 6048 82662 6062 82714
rect 6062 82662 6074 82714
rect 6074 82662 6104 82714
rect 6128 82662 6138 82714
rect 6138 82662 6184 82714
rect 5888 82660 5944 82662
rect 5968 82660 6024 82662
rect 6048 82660 6104 82662
rect 6128 82660 6184 82662
rect 6624 82170 6680 82172
rect 6704 82170 6760 82172
rect 6784 82170 6840 82172
rect 6864 82170 6920 82172
rect 6624 82118 6670 82170
rect 6670 82118 6680 82170
rect 6704 82118 6734 82170
rect 6734 82118 6746 82170
rect 6746 82118 6760 82170
rect 6784 82118 6798 82170
rect 6798 82118 6810 82170
rect 6810 82118 6840 82170
rect 6864 82118 6874 82170
rect 6874 82118 6920 82170
rect 6624 82116 6680 82118
rect 6704 82116 6760 82118
rect 6784 82116 6840 82118
rect 6864 82116 6920 82118
rect 5888 81626 5944 81628
rect 5968 81626 6024 81628
rect 6048 81626 6104 81628
rect 6128 81626 6184 81628
rect 5888 81574 5934 81626
rect 5934 81574 5944 81626
rect 5968 81574 5998 81626
rect 5998 81574 6010 81626
rect 6010 81574 6024 81626
rect 6048 81574 6062 81626
rect 6062 81574 6074 81626
rect 6074 81574 6104 81626
rect 6128 81574 6138 81626
rect 6138 81574 6184 81626
rect 5888 81572 5944 81574
rect 5968 81572 6024 81574
rect 6048 81572 6104 81574
rect 6128 81572 6184 81574
rect 4122 81276 4124 81296
rect 4124 81276 4176 81296
rect 4176 81276 4178 81296
rect 4122 81240 4178 81276
rect 6624 81082 6680 81084
rect 6704 81082 6760 81084
rect 6784 81082 6840 81084
rect 6864 81082 6920 81084
rect 6624 81030 6670 81082
rect 6670 81030 6680 81082
rect 6704 81030 6734 81082
rect 6734 81030 6746 81082
rect 6746 81030 6760 81082
rect 6784 81030 6798 81082
rect 6798 81030 6810 81082
rect 6810 81030 6840 81082
rect 6864 81030 6874 81082
rect 6874 81030 6920 81082
rect 6624 81028 6680 81030
rect 6704 81028 6760 81030
rect 6784 81028 6840 81030
rect 6864 81028 6920 81030
rect 5888 80538 5944 80540
rect 5968 80538 6024 80540
rect 6048 80538 6104 80540
rect 6128 80538 6184 80540
rect 5888 80486 5934 80538
rect 5934 80486 5944 80538
rect 5968 80486 5998 80538
rect 5998 80486 6010 80538
rect 6010 80486 6024 80538
rect 6048 80486 6062 80538
rect 6062 80486 6074 80538
rect 6074 80486 6104 80538
rect 6128 80486 6138 80538
rect 6138 80486 6184 80538
rect 5888 80484 5944 80486
rect 5968 80484 6024 80486
rect 6048 80484 6104 80486
rect 6128 80484 6184 80486
rect 6624 79994 6680 79996
rect 6704 79994 6760 79996
rect 6784 79994 6840 79996
rect 6864 79994 6920 79996
rect 4122 79880 4178 79936
rect 6624 79942 6670 79994
rect 6670 79942 6680 79994
rect 6704 79942 6734 79994
rect 6734 79942 6746 79994
rect 6746 79942 6760 79994
rect 6784 79942 6798 79994
rect 6798 79942 6810 79994
rect 6810 79942 6840 79994
rect 6864 79942 6874 79994
rect 6874 79942 6920 79994
rect 6624 79940 6680 79942
rect 6704 79940 6760 79942
rect 6784 79940 6840 79942
rect 6864 79940 6920 79942
rect 5888 79450 5944 79452
rect 5968 79450 6024 79452
rect 6048 79450 6104 79452
rect 6128 79450 6184 79452
rect 5888 79398 5934 79450
rect 5934 79398 5944 79450
rect 5968 79398 5998 79450
rect 5998 79398 6010 79450
rect 6010 79398 6024 79450
rect 6048 79398 6062 79450
rect 6062 79398 6074 79450
rect 6074 79398 6104 79450
rect 6128 79398 6138 79450
rect 6138 79398 6184 79450
rect 5888 79396 5944 79398
rect 5968 79396 6024 79398
rect 6048 79396 6104 79398
rect 6128 79396 6184 79398
rect 6624 78906 6680 78908
rect 6704 78906 6760 78908
rect 6784 78906 6840 78908
rect 6864 78906 6920 78908
rect 6624 78854 6670 78906
rect 6670 78854 6680 78906
rect 6704 78854 6734 78906
rect 6734 78854 6746 78906
rect 6746 78854 6760 78906
rect 6784 78854 6798 78906
rect 6798 78854 6810 78906
rect 6810 78854 6840 78906
rect 6864 78854 6874 78906
rect 6874 78854 6920 78906
rect 6624 78852 6680 78854
rect 6704 78852 6760 78854
rect 6784 78852 6840 78854
rect 6864 78852 6920 78854
rect 4122 78540 4178 78576
rect 4122 78520 4124 78540
rect 4124 78520 4176 78540
rect 4176 78520 4178 78540
rect 5888 78362 5944 78364
rect 5968 78362 6024 78364
rect 6048 78362 6104 78364
rect 6128 78362 6184 78364
rect 5888 78310 5934 78362
rect 5934 78310 5944 78362
rect 5968 78310 5998 78362
rect 5998 78310 6010 78362
rect 6010 78310 6024 78362
rect 6048 78310 6062 78362
rect 6062 78310 6074 78362
rect 6074 78310 6104 78362
rect 6128 78310 6138 78362
rect 6138 78310 6184 78362
rect 5888 78308 5944 78310
rect 5968 78308 6024 78310
rect 6048 78308 6104 78310
rect 6128 78308 6184 78310
rect 4122 77876 4124 77896
rect 4124 77876 4176 77896
rect 4176 77876 4178 77896
rect 4122 77840 4178 77876
rect 6624 77818 6680 77820
rect 6704 77818 6760 77820
rect 6784 77818 6840 77820
rect 6864 77818 6920 77820
rect 6624 77766 6670 77818
rect 6670 77766 6680 77818
rect 6704 77766 6734 77818
rect 6734 77766 6746 77818
rect 6746 77766 6760 77818
rect 6784 77766 6798 77818
rect 6798 77766 6810 77818
rect 6810 77766 6840 77818
rect 6864 77766 6874 77818
rect 6874 77766 6920 77818
rect 6624 77764 6680 77766
rect 6704 77764 6760 77766
rect 6784 77764 6840 77766
rect 6864 77764 6920 77766
rect 5888 77274 5944 77276
rect 5968 77274 6024 77276
rect 6048 77274 6104 77276
rect 6128 77274 6184 77276
rect 5888 77222 5934 77274
rect 5934 77222 5944 77274
rect 5968 77222 5998 77274
rect 5998 77222 6010 77274
rect 6010 77222 6024 77274
rect 6048 77222 6062 77274
rect 6062 77222 6074 77274
rect 6074 77222 6104 77274
rect 6128 77222 6138 77274
rect 6138 77222 6184 77274
rect 5888 77220 5944 77222
rect 5968 77220 6024 77222
rect 6048 77220 6104 77222
rect 6128 77220 6184 77222
rect 6624 76730 6680 76732
rect 6704 76730 6760 76732
rect 6784 76730 6840 76732
rect 6864 76730 6920 76732
rect 6624 76678 6670 76730
rect 6670 76678 6680 76730
rect 6704 76678 6734 76730
rect 6734 76678 6746 76730
rect 6746 76678 6760 76730
rect 6784 76678 6798 76730
rect 6798 76678 6810 76730
rect 6810 76678 6840 76730
rect 6864 76678 6874 76730
rect 6874 76678 6920 76730
rect 6624 76676 6680 76678
rect 6704 76676 6760 76678
rect 6784 76676 6840 76678
rect 6864 76676 6920 76678
rect 4214 76480 4270 76536
rect 5888 76186 5944 76188
rect 5968 76186 6024 76188
rect 6048 76186 6104 76188
rect 6128 76186 6184 76188
rect 5888 76134 5934 76186
rect 5934 76134 5944 76186
rect 5968 76134 5998 76186
rect 5998 76134 6010 76186
rect 6010 76134 6024 76186
rect 6048 76134 6062 76186
rect 6062 76134 6074 76186
rect 6074 76134 6104 76186
rect 6128 76134 6138 76186
rect 6138 76134 6184 76186
rect 5888 76132 5944 76134
rect 5968 76132 6024 76134
rect 6048 76132 6104 76134
rect 6128 76132 6184 76134
rect 4122 75820 4178 75856
rect 4122 75800 4124 75820
rect 4124 75800 4176 75820
rect 4176 75800 4178 75820
rect 6624 75642 6680 75644
rect 6704 75642 6760 75644
rect 6784 75642 6840 75644
rect 6864 75642 6920 75644
rect 6624 75590 6670 75642
rect 6670 75590 6680 75642
rect 6704 75590 6734 75642
rect 6734 75590 6746 75642
rect 6746 75590 6760 75642
rect 6784 75590 6798 75642
rect 6798 75590 6810 75642
rect 6810 75590 6840 75642
rect 6864 75590 6874 75642
rect 6874 75590 6920 75642
rect 6624 75588 6680 75590
rect 6704 75588 6760 75590
rect 6784 75588 6840 75590
rect 6864 75588 6920 75590
rect 5888 75098 5944 75100
rect 5968 75098 6024 75100
rect 6048 75098 6104 75100
rect 6128 75098 6184 75100
rect 5888 75046 5934 75098
rect 5934 75046 5944 75098
rect 5968 75046 5998 75098
rect 5998 75046 6010 75098
rect 6010 75046 6024 75098
rect 6048 75046 6062 75098
rect 6062 75046 6074 75098
rect 6074 75046 6104 75098
rect 6128 75046 6138 75098
rect 6138 75046 6184 75098
rect 5888 75044 5944 75046
rect 5968 75044 6024 75046
rect 6048 75044 6104 75046
rect 6128 75044 6184 75046
rect 5410 74748 5412 74768
rect 5412 74748 5464 74768
rect 5464 74748 5466 74768
rect 5410 74712 5466 74748
rect 6624 74554 6680 74556
rect 6704 74554 6760 74556
rect 6784 74554 6840 74556
rect 6864 74554 6920 74556
rect 4122 74440 4178 74496
rect 6624 74502 6670 74554
rect 6670 74502 6680 74554
rect 6704 74502 6734 74554
rect 6734 74502 6746 74554
rect 6746 74502 6760 74554
rect 6784 74502 6798 74554
rect 6798 74502 6810 74554
rect 6810 74502 6840 74554
rect 6864 74502 6874 74554
rect 6874 74502 6920 74554
rect 6624 74500 6680 74502
rect 6704 74500 6760 74502
rect 6784 74500 6840 74502
rect 6864 74500 6920 74502
rect 5888 74010 5944 74012
rect 5968 74010 6024 74012
rect 6048 74010 6104 74012
rect 6128 74010 6184 74012
rect 5888 73958 5934 74010
rect 5934 73958 5944 74010
rect 5968 73958 5998 74010
rect 5998 73958 6010 74010
rect 6010 73958 6024 74010
rect 6048 73958 6062 74010
rect 6062 73958 6074 74010
rect 6074 73958 6104 74010
rect 6128 73958 6138 74010
rect 6138 73958 6184 74010
rect 5888 73956 5944 73958
rect 5968 73956 6024 73958
rect 6048 73956 6104 73958
rect 6128 73956 6184 73958
rect 5410 73624 5466 73680
rect 6624 73466 6680 73468
rect 6704 73466 6760 73468
rect 6784 73466 6840 73468
rect 6864 73466 6920 73468
rect 6624 73414 6670 73466
rect 6670 73414 6680 73466
rect 6704 73414 6734 73466
rect 6734 73414 6746 73466
rect 6746 73414 6760 73466
rect 6784 73414 6798 73466
rect 6798 73414 6810 73466
rect 6810 73414 6840 73466
rect 6864 73414 6874 73466
rect 6874 73414 6920 73466
rect 6624 73412 6680 73414
rect 6704 73412 6760 73414
rect 6784 73412 6840 73414
rect 6864 73412 6920 73414
rect 4122 73100 4178 73136
rect 4122 73080 4124 73100
rect 4124 73080 4176 73100
rect 4176 73080 4178 73100
rect 5888 72922 5944 72924
rect 5968 72922 6024 72924
rect 6048 72922 6104 72924
rect 6128 72922 6184 72924
rect 5888 72870 5934 72922
rect 5934 72870 5944 72922
rect 5968 72870 5998 72922
rect 5998 72870 6010 72922
rect 6010 72870 6024 72922
rect 6048 72870 6062 72922
rect 6062 72870 6074 72922
rect 6074 72870 6104 72922
rect 6128 72870 6138 72922
rect 6138 72870 6184 72922
rect 5888 72868 5944 72870
rect 5968 72868 6024 72870
rect 6048 72868 6104 72870
rect 6128 72868 6184 72870
rect 4122 72436 4124 72456
rect 4124 72436 4176 72456
rect 4176 72436 4178 72456
rect 4122 72400 4178 72436
rect 6624 72378 6680 72380
rect 6704 72378 6760 72380
rect 6784 72378 6840 72380
rect 6864 72378 6920 72380
rect 6624 72326 6670 72378
rect 6670 72326 6680 72378
rect 6704 72326 6734 72378
rect 6734 72326 6746 72378
rect 6746 72326 6760 72378
rect 6784 72326 6798 72378
rect 6798 72326 6810 72378
rect 6810 72326 6840 72378
rect 6864 72326 6874 72378
rect 6874 72326 6920 72378
rect 6624 72324 6680 72326
rect 6704 72324 6760 72326
rect 6784 72324 6840 72326
rect 6864 72324 6920 72326
rect 5888 71834 5944 71836
rect 5968 71834 6024 71836
rect 6048 71834 6104 71836
rect 6128 71834 6184 71836
rect 5888 71782 5934 71834
rect 5934 71782 5944 71834
rect 5968 71782 5998 71834
rect 5998 71782 6010 71834
rect 6010 71782 6024 71834
rect 6048 71782 6062 71834
rect 6062 71782 6074 71834
rect 6074 71782 6104 71834
rect 6128 71782 6138 71834
rect 6138 71782 6184 71834
rect 5888 71780 5944 71782
rect 5968 71780 6024 71782
rect 6048 71780 6104 71782
rect 6128 71780 6184 71782
rect 6624 71290 6680 71292
rect 6704 71290 6760 71292
rect 6784 71290 6840 71292
rect 6864 71290 6920 71292
rect 6624 71238 6670 71290
rect 6670 71238 6680 71290
rect 6704 71238 6734 71290
rect 6734 71238 6746 71290
rect 6746 71238 6760 71290
rect 6784 71238 6798 71290
rect 6798 71238 6810 71290
rect 6810 71238 6840 71290
rect 6864 71238 6874 71290
rect 6874 71238 6920 71290
rect 6624 71236 6680 71238
rect 6704 71236 6760 71238
rect 6784 71236 6840 71238
rect 6864 71236 6920 71238
rect 4214 71040 4270 71096
rect 5888 70746 5944 70748
rect 5968 70746 6024 70748
rect 6048 70746 6104 70748
rect 6128 70746 6184 70748
rect 5888 70694 5934 70746
rect 5934 70694 5944 70746
rect 5968 70694 5998 70746
rect 5998 70694 6010 70746
rect 6010 70694 6024 70746
rect 6048 70694 6062 70746
rect 6062 70694 6074 70746
rect 6074 70694 6104 70746
rect 6128 70694 6138 70746
rect 6138 70694 6184 70746
rect 5888 70692 5944 70694
rect 5968 70692 6024 70694
rect 6048 70692 6104 70694
rect 6128 70692 6184 70694
rect 4122 70380 4178 70416
rect 4122 70360 4124 70380
rect 4124 70360 4176 70380
rect 4176 70360 4178 70380
rect 6624 70202 6680 70204
rect 6704 70202 6760 70204
rect 6784 70202 6840 70204
rect 6864 70202 6920 70204
rect 6624 70150 6670 70202
rect 6670 70150 6680 70202
rect 6704 70150 6734 70202
rect 6734 70150 6746 70202
rect 6746 70150 6760 70202
rect 6784 70150 6798 70202
rect 6798 70150 6810 70202
rect 6810 70150 6840 70202
rect 6864 70150 6874 70202
rect 6874 70150 6920 70202
rect 6624 70148 6680 70150
rect 6704 70148 6760 70150
rect 6784 70148 6840 70150
rect 6864 70148 6920 70150
rect 5888 69658 5944 69660
rect 5968 69658 6024 69660
rect 6048 69658 6104 69660
rect 6128 69658 6184 69660
rect 5888 69606 5934 69658
rect 5934 69606 5944 69658
rect 5968 69606 5998 69658
rect 5998 69606 6010 69658
rect 6010 69606 6024 69658
rect 6048 69606 6062 69658
rect 6062 69606 6074 69658
rect 6074 69606 6104 69658
rect 6128 69606 6138 69658
rect 6138 69606 6184 69658
rect 5888 69604 5944 69606
rect 5968 69604 6024 69606
rect 6048 69604 6104 69606
rect 6128 69604 6184 69606
rect 4122 69000 4178 69056
rect 6624 69114 6680 69116
rect 6704 69114 6760 69116
rect 6784 69114 6840 69116
rect 6864 69114 6920 69116
rect 6624 69062 6670 69114
rect 6670 69062 6680 69114
rect 6704 69062 6734 69114
rect 6734 69062 6746 69114
rect 6746 69062 6760 69114
rect 6784 69062 6798 69114
rect 6798 69062 6810 69114
rect 6810 69062 6840 69114
rect 6864 69062 6874 69114
rect 6874 69062 6920 69114
rect 6624 69060 6680 69062
rect 6704 69060 6760 69062
rect 6784 69060 6840 69062
rect 6864 69060 6920 69062
rect 5410 68864 5466 68920
rect 5888 68570 5944 68572
rect 5968 68570 6024 68572
rect 6048 68570 6104 68572
rect 6128 68570 6184 68572
rect 5888 68518 5934 68570
rect 5934 68518 5944 68570
rect 5968 68518 5998 68570
rect 5998 68518 6010 68570
rect 6010 68518 6024 68570
rect 6048 68518 6062 68570
rect 6062 68518 6074 68570
rect 6074 68518 6104 68570
rect 6128 68518 6138 68570
rect 6138 68518 6184 68570
rect 5888 68516 5944 68518
rect 5968 68516 6024 68518
rect 6048 68516 6104 68518
rect 6128 68516 6184 68518
rect 5410 68184 5466 68240
rect 6624 68026 6680 68028
rect 6704 68026 6760 68028
rect 6784 68026 6840 68028
rect 6864 68026 6920 68028
rect 6624 67974 6670 68026
rect 6670 67974 6680 68026
rect 6704 67974 6734 68026
rect 6734 67974 6746 68026
rect 6746 67974 6760 68026
rect 6784 67974 6798 68026
rect 6798 67974 6810 68026
rect 6810 67974 6840 68026
rect 6864 67974 6874 68026
rect 6874 67974 6920 68026
rect 6624 67972 6680 67974
rect 6704 67972 6760 67974
rect 6784 67972 6840 67974
rect 6864 67972 6920 67974
rect 4030 67660 4086 67696
rect 4030 67640 4032 67660
rect 4032 67640 4084 67660
rect 4084 67640 4086 67660
rect 5888 67482 5944 67484
rect 5968 67482 6024 67484
rect 6048 67482 6104 67484
rect 6128 67482 6184 67484
rect 5888 67430 5934 67482
rect 5934 67430 5944 67482
rect 5968 67430 5998 67482
rect 5998 67430 6010 67482
rect 6010 67430 6024 67482
rect 6048 67430 6062 67482
rect 6062 67430 6074 67482
rect 6074 67430 6104 67482
rect 6128 67430 6138 67482
rect 6138 67430 6184 67482
rect 5888 67428 5944 67430
rect 5968 67428 6024 67430
rect 6048 67428 6104 67430
rect 6128 67428 6184 67430
rect 4122 66996 4124 67016
rect 4124 66996 4176 67016
rect 4176 66996 4178 67016
rect 4122 66960 4178 66996
rect 6624 66938 6680 66940
rect 6704 66938 6760 66940
rect 6784 66938 6840 66940
rect 6864 66938 6920 66940
rect 6624 66886 6670 66938
rect 6670 66886 6680 66938
rect 6704 66886 6734 66938
rect 6734 66886 6746 66938
rect 6746 66886 6760 66938
rect 6784 66886 6798 66938
rect 6798 66886 6810 66938
rect 6810 66886 6840 66938
rect 6864 66886 6874 66938
rect 6874 66886 6920 66938
rect 6624 66884 6680 66886
rect 6704 66884 6760 66886
rect 6784 66884 6840 66886
rect 6864 66884 6920 66886
rect 5888 66394 5944 66396
rect 5968 66394 6024 66396
rect 6048 66394 6104 66396
rect 6128 66394 6184 66396
rect 5888 66342 5934 66394
rect 5934 66342 5944 66394
rect 5968 66342 5998 66394
rect 5998 66342 6010 66394
rect 6010 66342 6024 66394
rect 6048 66342 6062 66394
rect 6062 66342 6074 66394
rect 6074 66342 6104 66394
rect 6128 66342 6138 66394
rect 6138 66342 6184 66394
rect 5888 66340 5944 66342
rect 5968 66340 6024 66342
rect 6048 66340 6104 66342
rect 6128 66340 6184 66342
rect 6624 65850 6680 65852
rect 6704 65850 6760 65852
rect 6784 65850 6840 65852
rect 6864 65850 6920 65852
rect 6624 65798 6670 65850
rect 6670 65798 6680 65850
rect 6704 65798 6734 65850
rect 6734 65798 6746 65850
rect 6746 65798 6760 65850
rect 6784 65798 6798 65850
rect 6798 65798 6810 65850
rect 6810 65798 6840 65850
rect 6864 65798 6874 65850
rect 6874 65798 6920 65850
rect 6624 65796 6680 65798
rect 6704 65796 6760 65798
rect 6784 65796 6840 65798
rect 6864 65796 6920 65798
rect 4306 65600 4362 65656
rect 5888 65306 5944 65308
rect 5968 65306 6024 65308
rect 6048 65306 6104 65308
rect 6128 65306 6184 65308
rect 5888 65254 5934 65306
rect 5934 65254 5944 65306
rect 5968 65254 5998 65306
rect 5998 65254 6010 65306
rect 6010 65254 6024 65306
rect 6048 65254 6062 65306
rect 6062 65254 6074 65306
rect 6074 65254 6104 65306
rect 6128 65254 6138 65306
rect 6138 65254 6184 65306
rect 5888 65252 5944 65254
rect 5968 65252 6024 65254
rect 6048 65252 6104 65254
rect 6128 65252 6184 65254
rect 4306 64956 4308 64976
rect 4308 64956 4360 64976
rect 4360 64956 4362 64976
rect 4306 64920 4362 64956
rect 6624 64762 6680 64764
rect 6704 64762 6760 64764
rect 6784 64762 6840 64764
rect 6864 64762 6920 64764
rect 6624 64710 6670 64762
rect 6670 64710 6680 64762
rect 6704 64710 6734 64762
rect 6734 64710 6746 64762
rect 6746 64710 6760 64762
rect 6784 64710 6798 64762
rect 6798 64710 6810 64762
rect 6810 64710 6840 64762
rect 6864 64710 6874 64762
rect 6874 64710 6920 64762
rect 6624 64708 6680 64710
rect 6704 64708 6760 64710
rect 6784 64708 6840 64710
rect 6864 64708 6920 64710
rect 5888 64218 5944 64220
rect 5968 64218 6024 64220
rect 6048 64218 6104 64220
rect 6128 64218 6184 64220
rect 5888 64166 5934 64218
rect 5934 64166 5944 64218
rect 5968 64166 5998 64218
rect 5998 64166 6010 64218
rect 6010 64166 6024 64218
rect 6048 64166 6062 64218
rect 6062 64166 6074 64218
rect 6074 64166 6104 64218
rect 6128 64166 6138 64218
rect 6138 64166 6184 64218
rect 5888 64164 5944 64166
rect 5968 64164 6024 64166
rect 6048 64164 6104 64166
rect 6128 64164 6184 64166
rect 4306 63560 4362 63616
rect 6624 63674 6680 63676
rect 6704 63674 6760 63676
rect 6784 63674 6840 63676
rect 6864 63674 6920 63676
rect 6624 63622 6670 63674
rect 6670 63622 6680 63674
rect 6704 63622 6734 63674
rect 6734 63622 6746 63674
rect 6746 63622 6760 63674
rect 6784 63622 6798 63674
rect 6798 63622 6810 63674
rect 6810 63622 6840 63674
rect 6864 63622 6874 63674
rect 6874 63622 6920 63674
rect 6624 63620 6680 63622
rect 6704 63620 6760 63622
rect 6784 63620 6840 63622
rect 6864 63620 6920 63622
rect 5686 63424 5742 63480
rect 5888 63130 5944 63132
rect 5968 63130 6024 63132
rect 6048 63130 6104 63132
rect 6128 63130 6184 63132
rect 5888 63078 5934 63130
rect 5934 63078 5944 63130
rect 5968 63078 5998 63130
rect 5998 63078 6010 63130
rect 6010 63078 6024 63130
rect 6048 63078 6062 63130
rect 6062 63078 6074 63130
rect 6074 63078 6104 63130
rect 6128 63078 6138 63130
rect 6138 63078 6184 63130
rect 5888 63076 5944 63078
rect 5968 63076 6024 63078
rect 6048 63076 6104 63078
rect 6128 63076 6184 63078
rect 6624 62586 6680 62588
rect 6704 62586 6760 62588
rect 6784 62586 6840 62588
rect 6864 62586 6920 62588
rect 6624 62534 6670 62586
rect 6670 62534 6680 62586
rect 6704 62534 6734 62586
rect 6734 62534 6746 62586
rect 6746 62534 6760 62586
rect 6784 62534 6798 62586
rect 6798 62534 6810 62586
rect 6810 62534 6840 62586
rect 6864 62534 6874 62586
rect 6874 62534 6920 62586
rect 6624 62532 6680 62534
rect 6704 62532 6760 62534
rect 6784 62532 6840 62534
rect 6864 62532 6920 62534
rect 5686 62336 5742 62392
rect 4306 62200 4362 62256
rect 5888 62042 5944 62044
rect 5968 62042 6024 62044
rect 6048 62042 6104 62044
rect 6128 62042 6184 62044
rect 5888 61990 5934 62042
rect 5934 61990 5944 62042
rect 5968 61990 5998 62042
rect 5998 61990 6010 62042
rect 6010 61990 6024 62042
rect 6048 61990 6062 62042
rect 6062 61990 6074 62042
rect 6074 61990 6104 62042
rect 6128 61990 6138 62042
rect 6138 61990 6184 62042
rect 5888 61988 5944 61990
rect 5968 61988 6024 61990
rect 6048 61988 6104 61990
rect 6128 61988 6184 61990
rect 4306 61520 4362 61576
rect 6624 61498 6680 61500
rect 6704 61498 6760 61500
rect 6784 61498 6840 61500
rect 6864 61498 6920 61500
rect 6624 61446 6670 61498
rect 6670 61446 6680 61498
rect 6704 61446 6734 61498
rect 6734 61446 6746 61498
rect 6746 61446 6760 61498
rect 6784 61446 6798 61498
rect 6798 61446 6810 61498
rect 6810 61446 6840 61498
rect 6864 61446 6874 61498
rect 6874 61446 6920 61498
rect 6624 61444 6680 61446
rect 6704 61444 6760 61446
rect 6784 61444 6840 61446
rect 6864 61444 6920 61446
rect 5888 60954 5944 60956
rect 5968 60954 6024 60956
rect 6048 60954 6104 60956
rect 6128 60954 6184 60956
rect 5888 60902 5934 60954
rect 5934 60902 5944 60954
rect 5968 60902 5998 60954
rect 5998 60902 6010 60954
rect 6010 60902 6024 60954
rect 6048 60902 6062 60954
rect 6062 60902 6074 60954
rect 6074 60902 6104 60954
rect 6128 60902 6138 60954
rect 6138 60902 6184 60954
rect 5888 60900 5944 60902
rect 5968 60900 6024 60902
rect 6048 60900 6104 60902
rect 6128 60900 6184 60902
rect 6624 60410 6680 60412
rect 6704 60410 6760 60412
rect 6784 60410 6840 60412
rect 6864 60410 6920 60412
rect 6624 60358 6670 60410
rect 6670 60358 6680 60410
rect 6704 60358 6734 60410
rect 6734 60358 6746 60410
rect 6746 60358 6760 60410
rect 6784 60358 6798 60410
rect 6798 60358 6810 60410
rect 6810 60358 6840 60410
rect 6864 60358 6874 60410
rect 6874 60358 6920 60410
rect 6624 60356 6680 60358
rect 6704 60356 6760 60358
rect 6784 60356 6840 60358
rect 6864 60356 6920 60358
rect 4306 60160 4362 60216
rect 5888 59866 5944 59868
rect 5968 59866 6024 59868
rect 6048 59866 6104 59868
rect 6128 59866 6184 59868
rect 5888 59814 5934 59866
rect 5934 59814 5944 59866
rect 5968 59814 5998 59866
rect 5998 59814 6010 59866
rect 6010 59814 6024 59866
rect 6048 59814 6062 59866
rect 6062 59814 6074 59866
rect 6074 59814 6104 59866
rect 6128 59814 6138 59866
rect 6138 59814 6184 59866
rect 5888 59812 5944 59814
rect 5968 59812 6024 59814
rect 6048 59812 6104 59814
rect 6128 59812 6184 59814
rect 4306 59516 4308 59536
rect 4308 59516 4360 59536
rect 4360 59516 4362 59536
rect 4306 59480 4362 59516
rect 6624 59322 6680 59324
rect 6704 59322 6760 59324
rect 6784 59322 6840 59324
rect 6864 59322 6920 59324
rect 6624 59270 6670 59322
rect 6670 59270 6680 59322
rect 6704 59270 6734 59322
rect 6734 59270 6746 59322
rect 6746 59270 6760 59322
rect 6784 59270 6798 59322
rect 6798 59270 6810 59322
rect 6810 59270 6840 59322
rect 6864 59270 6874 59322
rect 6874 59270 6920 59322
rect 6624 59268 6680 59270
rect 6704 59268 6760 59270
rect 6784 59268 6840 59270
rect 6864 59268 6920 59270
rect 5888 58778 5944 58780
rect 5968 58778 6024 58780
rect 6048 58778 6104 58780
rect 6128 58778 6184 58780
rect 5888 58726 5934 58778
rect 5934 58726 5944 58778
rect 5968 58726 5998 58778
rect 5998 58726 6010 58778
rect 6010 58726 6024 58778
rect 6048 58726 6062 58778
rect 6062 58726 6074 58778
rect 6074 58726 6104 58778
rect 6128 58726 6138 58778
rect 6138 58726 6184 58778
rect 5888 58724 5944 58726
rect 5968 58724 6024 58726
rect 6048 58724 6104 58726
rect 6128 58724 6184 58726
rect 4306 58120 4362 58176
rect 6624 58234 6680 58236
rect 6704 58234 6760 58236
rect 6784 58234 6840 58236
rect 6864 58234 6920 58236
rect 6624 58182 6670 58234
rect 6670 58182 6680 58234
rect 6704 58182 6734 58234
rect 6734 58182 6746 58234
rect 6746 58182 6760 58234
rect 6784 58182 6798 58234
rect 6798 58182 6810 58234
rect 6810 58182 6840 58234
rect 6864 58182 6874 58234
rect 6874 58182 6920 58234
rect 6624 58180 6680 58182
rect 6704 58180 6760 58182
rect 6784 58180 6840 58182
rect 6864 58180 6920 58182
rect 5410 57984 5466 58040
rect 5888 57690 5944 57692
rect 5968 57690 6024 57692
rect 6048 57690 6104 57692
rect 6128 57690 6184 57692
rect 5888 57638 5934 57690
rect 5934 57638 5944 57690
rect 5968 57638 5998 57690
rect 5998 57638 6010 57690
rect 6010 57638 6024 57690
rect 6048 57638 6062 57690
rect 6062 57638 6074 57690
rect 6074 57638 6104 57690
rect 6128 57638 6138 57690
rect 6138 57638 6184 57690
rect 5888 57636 5944 57638
rect 5968 57636 6024 57638
rect 6048 57636 6104 57638
rect 6128 57636 6184 57638
rect 6624 57146 6680 57148
rect 6704 57146 6760 57148
rect 6784 57146 6840 57148
rect 6864 57146 6920 57148
rect 6624 57094 6670 57146
rect 6670 57094 6680 57146
rect 6704 57094 6734 57146
rect 6734 57094 6746 57146
rect 6746 57094 6760 57146
rect 6784 57094 6798 57146
rect 6798 57094 6810 57146
rect 6810 57094 6840 57146
rect 6864 57094 6874 57146
rect 6874 57094 6920 57146
rect 6624 57092 6680 57094
rect 6704 57092 6760 57094
rect 6784 57092 6840 57094
rect 6864 57092 6920 57094
rect 4306 56760 4362 56816
rect 5888 56602 5944 56604
rect 5968 56602 6024 56604
rect 6048 56602 6104 56604
rect 6128 56602 6184 56604
rect 5888 56550 5934 56602
rect 5934 56550 5944 56602
rect 5968 56550 5998 56602
rect 5998 56550 6010 56602
rect 6010 56550 6024 56602
rect 6048 56550 6062 56602
rect 6062 56550 6074 56602
rect 6074 56550 6104 56602
rect 6128 56550 6138 56602
rect 6138 56550 6184 56602
rect 5888 56548 5944 56550
rect 5968 56548 6024 56550
rect 6048 56548 6104 56550
rect 6128 56548 6184 56550
rect 4306 56080 4362 56136
rect 6624 56058 6680 56060
rect 6704 56058 6760 56060
rect 6784 56058 6840 56060
rect 6864 56058 6920 56060
rect 6624 56006 6670 56058
rect 6670 56006 6680 56058
rect 6704 56006 6734 56058
rect 6734 56006 6746 56058
rect 6746 56006 6760 56058
rect 6784 56006 6798 56058
rect 6798 56006 6810 56058
rect 6810 56006 6840 56058
rect 6864 56006 6874 56058
rect 6874 56006 6920 56058
rect 6624 56004 6680 56006
rect 6704 56004 6760 56006
rect 6784 56004 6840 56006
rect 6864 56004 6920 56006
rect 5888 55514 5944 55516
rect 5968 55514 6024 55516
rect 6048 55514 6104 55516
rect 6128 55514 6184 55516
rect 5888 55462 5934 55514
rect 5934 55462 5944 55514
rect 5968 55462 5998 55514
rect 5998 55462 6010 55514
rect 6010 55462 6024 55514
rect 6048 55462 6062 55514
rect 6062 55462 6074 55514
rect 6074 55462 6104 55514
rect 6128 55462 6138 55514
rect 6138 55462 6184 55514
rect 5888 55460 5944 55462
rect 5968 55460 6024 55462
rect 6048 55460 6104 55462
rect 6128 55460 6184 55462
rect 6624 54970 6680 54972
rect 6704 54970 6760 54972
rect 6784 54970 6840 54972
rect 6864 54970 6920 54972
rect 6624 54918 6670 54970
rect 6670 54918 6680 54970
rect 6704 54918 6734 54970
rect 6734 54918 6746 54970
rect 6746 54918 6760 54970
rect 6784 54918 6798 54970
rect 6798 54918 6810 54970
rect 6810 54918 6840 54970
rect 6864 54918 6874 54970
rect 6874 54918 6920 54970
rect 6624 54916 6680 54918
rect 6704 54916 6760 54918
rect 6784 54916 6840 54918
rect 6864 54916 6920 54918
rect 4306 54720 4362 54776
rect 5888 54426 5944 54428
rect 5968 54426 6024 54428
rect 6048 54426 6104 54428
rect 6128 54426 6184 54428
rect 5888 54374 5934 54426
rect 5934 54374 5944 54426
rect 5968 54374 5998 54426
rect 5998 54374 6010 54426
rect 6010 54374 6024 54426
rect 6048 54374 6062 54426
rect 6062 54374 6074 54426
rect 6074 54374 6104 54426
rect 6128 54374 6138 54426
rect 6138 54374 6184 54426
rect 5888 54372 5944 54374
rect 5968 54372 6024 54374
rect 6048 54372 6104 54374
rect 6128 54372 6184 54374
rect 4306 54076 4308 54096
rect 4308 54076 4360 54096
rect 4360 54076 4362 54096
rect 4306 54040 4362 54076
rect 6624 53882 6680 53884
rect 6704 53882 6760 53884
rect 6784 53882 6840 53884
rect 6864 53882 6920 53884
rect 6624 53830 6670 53882
rect 6670 53830 6680 53882
rect 6704 53830 6734 53882
rect 6734 53830 6746 53882
rect 6746 53830 6760 53882
rect 6784 53830 6798 53882
rect 6798 53830 6810 53882
rect 6810 53830 6840 53882
rect 6864 53830 6874 53882
rect 6874 53830 6920 53882
rect 6624 53828 6680 53830
rect 6704 53828 6760 53830
rect 6784 53828 6840 53830
rect 6864 53828 6920 53830
rect 5686 53632 5742 53688
rect 5888 53338 5944 53340
rect 5968 53338 6024 53340
rect 6048 53338 6104 53340
rect 6128 53338 6184 53340
rect 5888 53286 5934 53338
rect 5934 53286 5944 53338
rect 5968 53286 5998 53338
rect 5998 53286 6010 53338
rect 6010 53286 6024 53338
rect 6048 53286 6062 53338
rect 6062 53286 6074 53338
rect 6074 53286 6104 53338
rect 6128 53286 6138 53338
rect 6138 53286 6184 53338
rect 5888 53284 5944 53286
rect 5968 53284 6024 53286
rect 6048 53284 6104 53286
rect 6128 53284 6184 53286
rect 6624 52794 6680 52796
rect 6704 52794 6760 52796
rect 6784 52794 6840 52796
rect 6864 52794 6920 52796
rect 4306 52680 4362 52736
rect 6624 52742 6670 52794
rect 6670 52742 6680 52794
rect 6704 52742 6734 52794
rect 6734 52742 6746 52794
rect 6746 52742 6760 52794
rect 6784 52742 6798 52794
rect 6798 52742 6810 52794
rect 6810 52742 6840 52794
rect 6864 52742 6874 52794
rect 6874 52742 6920 52794
rect 6624 52740 6680 52742
rect 6704 52740 6760 52742
rect 6784 52740 6840 52742
rect 6864 52740 6920 52742
rect 5888 52250 5944 52252
rect 5968 52250 6024 52252
rect 6048 52250 6104 52252
rect 6128 52250 6184 52252
rect 5888 52198 5934 52250
rect 5934 52198 5944 52250
rect 5968 52198 5998 52250
rect 5998 52198 6010 52250
rect 6010 52198 6024 52250
rect 6048 52198 6062 52250
rect 6062 52198 6074 52250
rect 6074 52198 6104 52250
rect 6128 52198 6138 52250
rect 6138 52198 6184 52250
rect 5888 52196 5944 52198
rect 5968 52196 6024 52198
rect 6048 52196 6104 52198
rect 6128 52196 6184 52198
rect 6624 51706 6680 51708
rect 6704 51706 6760 51708
rect 6784 51706 6840 51708
rect 6864 51706 6920 51708
rect 6624 51654 6670 51706
rect 6670 51654 6680 51706
rect 6704 51654 6734 51706
rect 6734 51654 6746 51706
rect 6746 51654 6760 51706
rect 6784 51654 6798 51706
rect 6798 51654 6810 51706
rect 6810 51654 6840 51706
rect 6864 51654 6874 51706
rect 6874 51654 6920 51706
rect 6624 51652 6680 51654
rect 6704 51652 6760 51654
rect 6784 51652 6840 51654
rect 6864 51652 6920 51654
rect 4306 51320 4362 51376
rect 5888 51162 5944 51164
rect 5968 51162 6024 51164
rect 6048 51162 6104 51164
rect 6128 51162 6184 51164
rect 5888 51110 5934 51162
rect 5934 51110 5944 51162
rect 5968 51110 5998 51162
rect 5998 51110 6010 51162
rect 6010 51110 6024 51162
rect 6048 51110 6062 51162
rect 6062 51110 6074 51162
rect 6074 51110 6104 51162
rect 6128 51110 6138 51162
rect 6138 51110 6184 51162
rect 5888 51108 5944 51110
rect 5968 51108 6024 51110
rect 6048 51108 6104 51110
rect 6128 51108 6184 51110
rect 6624 50618 6680 50620
rect 6704 50618 6760 50620
rect 6784 50618 6840 50620
rect 6864 50618 6920 50620
rect 6624 50566 6670 50618
rect 6670 50566 6680 50618
rect 6704 50566 6734 50618
rect 6734 50566 6746 50618
rect 6746 50566 6760 50618
rect 6784 50566 6798 50618
rect 6798 50566 6810 50618
rect 6810 50566 6840 50618
rect 6864 50566 6874 50618
rect 6874 50566 6920 50618
rect 6624 50564 6680 50566
rect 6704 50564 6760 50566
rect 6784 50564 6840 50566
rect 6864 50564 6920 50566
rect 5888 50074 5944 50076
rect 5968 50074 6024 50076
rect 6048 50074 6104 50076
rect 6128 50074 6184 50076
rect 5888 50022 5934 50074
rect 5934 50022 5944 50074
rect 5968 50022 5998 50074
rect 5998 50022 6010 50074
rect 6010 50022 6024 50074
rect 6048 50022 6062 50074
rect 6062 50022 6074 50074
rect 6074 50022 6104 50074
rect 6128 50022 6138 50074
rect 6138 50022 6184 50074
rect 5888 50020 5944 50022
rect 5968 50020 6024 50022
rect 6048 50020 6104 50022
rect 6128 50020 6184 50022
rect 6624 49530 6680 49532
rect 6704 49530 6760 49532
rect 6784 49530 6840 49532
rect 6864 49530 6920 49532
rect 6624 49478 6670 49530
rect 6670 49478 6680 49530
rect 6704 49478 6734 49530
rect 6734 49478 6746 49530
rect 6746 49478 6760 49530
rect 6784 49478 6798 49530
rect 6798 49478 6810 49530
rect 6810 49478 6840 49530
rect 6864 49478 6874 49530
rect 6874 49478 6920 49530
rect 6624 49476 6680 49478
rect 6704 49476 6760 49478
rect 6784 49476 6840 49478
rect 6864 49476 6920 49478
rect 5888 48986 5944 48988
rect 5968 48986 6024 48988
rect 6048 48986 6104 48988
rect 6128 48986 6184 48988
rect 5888 48934 5934 48986
rect 5934 48934 5944 48986
rect 5968 48934 5998 48986
rect 5998 48934 6010 48986
rect 6010 48934 6024 48986
rect 6048 48934 6062 48986
rect 6062 48934 6074 48986
rect 6074 48934 6104 48986
rect 6128 48934 6138 48986
rect 6138 48934 6184 48986
rect 5888 48932 5944 48934
rect 5968 48932 6024 48934
rect 6048 48932 6104 48934
rect 6128 48932 6184 48934
rect 6624 48442 6680 48444
rect 6704 48442 6760 48444
rect 6784 48442 6840 48444
rect 6864 48442 6920 48444
rect 6624 48390 6670 48442
rect 6670 48390 6680 48442
rect 6704 48390 6734 48442
rect 6734 48390 6746 48442
rect 6746 48390 6760 48442
rect 6784 48390 6798 48442
rect 6798 48390 6810 48442
rect 6810 48390 6840 48442
rect 6864 48390 6874 48442
rect 6874 48390 6920 48442
rect 6624 48388 6680 48390
rect 6704 48388 6760 48390
rect 6784 48388 6840 48390
rect 6864 48388 6920 48390
rect 5888 47898 5944 47900
rect 5968 47898 6024 47900
rect 6048 47898 6104 47900
rect 6128 47898 6184 47900
rect 5888 47846 5934 47898
rect 5934 47846 5944 47898
rect 5968 47846 5998 47898
rect 5998 47846 6010 47898
rect 6010 47846 6024 47898
rect 6048 47846 6062 47898
rect 6062 47846 6074 47898
rect 6074 47846 6104 47898
rect 6128 47846 6138 47898
rect 6138 47846 6184 47898
rect 5888 47844 5944 47846
rect 5968 47844 6024 47846
rect 6048 47844 6104 47846
rect 6128 47844 6184 47846
rect 6624 47354 6680 47356
rect 6704 47354 6760 47356
rect 6784 47354 6840 47356
rect 6864 47354 6920 47356
rect 6624 47302 6670 47354
rect 6670 47302 6680 47354
rect 6704 47302 6734 47354
rect 6734 47302 6746 47354
rect 6746 47302 6760 47354
rect 6784 47302 6798 47354
rect 6798 47302 6810 47354
rect 6810 47302 6840 47354
rect 6864 47302 6874 47354
rect 6874 47302 6920 47354
rect 6624 47300 6680 47302
rect 6704 47300 6760 47302
rect 6784 47300 6840 47302
rect 6864 47300 6920 47302
rect 5888 46810 5944 46812
rect 5968 46810 6024 46812
rect 6048 46810 6104 46812
rect 6128 46810 6184 46812
rect 5888 46758 5934 46810
rect 5934 46758 5944 46810
rect 5968 46758 5998 46810
rect 5998 46758 6010 46810
rect 6010 46758 6024 46810
rect 6048 46758 6062 46810
rect 6062 46758 6074 46810
rect 6074 46758 6104 46810
rect 6128 46758 6138 46810
rect 6138 46758 6184 46810
rect 5888 46756 5944 46758
rect 5968 46756 6024 46758
rect 6048 46756 6104 46758
rect 6128 46756 6184 46758
rect 6624 46266 6680 46268
rect 6704 46266 6760 46268
rect 6784 46266 6840 46268
rect 6864 46266 6920 46268
rect 6624 46214 6670 46266
rect 6670 46214 6680 46266
rect 6704 46214 6734 46266
rect 6734 46214 6746 46266
rect 6746 46214 6760 46266
rect 6784 46214 6798 46266
rect 6798 46214 6810 46266
rect 6810 46214 6840 46266
rect 6864 46214 6874 46266
rect 6874 46214 6920 46266
rect 6624 46212 6680 46214
rect 6704 46212 6760 46214
rect 6784 46212 6840 46214
rect 6864 46212 6920 46214
rect 5888 45722 5944 45724
rect 5968 45722 6024 45724
rect 6048 45722 6104 45724
rect 6128 45722 6184 45724
rect 5888 45670 5934 45722
rect 5934 45670 5944 45722
rect 5968 45670 5998 45722
rect 5998 45670 6010 45722
rect 6010 45670 6024 45722
rect 6048 45670 6062 45722
rect 6062 45670 6074 45722
rect 6074 45670 6104 45722
rect 6128 45670 6138 45722
rect 6138 45670 6184 45722
rect 5888 45668 5944 45670
rect 5968 45668 6024 45670
rect 6048 45668 6104 45670
rect 6128 45668 6184 45670
rect 8538 80968 8594 81024
rect 8538 79880 8594 79936
rect 8538 78792 8594 78848
rect 8538 77704 8594 77760
rect 8538 76616 8594 76672
rect 8538 75528 8594 75584
rect 8538 72264 8594 72320
rect 8538 71176 8594 71232
rect 8538 70088 8594 70144
rect 8538 66824 8594 66880
rect 8538 65736 8594 65792
rect 8538 64648 8594 64704
rect 8538 61384 8594 61440
rect 8538 60296 8594 60352
rect 8538 59208 8594 59264
rect 8538 54856 8594 54912
rect 8538 52680 8594 52736
rect 8538 51592 8594 51648
rect 7618 45744 7674 45800
rect 5686 45356 5742 45392
rect 5686 45336 5688 45356
rect 5688 45336 5740 45356
rect 5740 45336 5742 45356
rect 4306 45200 4362 45256
rect 6624 45178 6680 45180
rect 6704 45178 6760 45180
rect 6784 45178 6840 45180
rect 6864 45178 6920 45180
rect 6624 45126 6670 45178
rect 6670 45126 6680 45178
rect 6704 45126 6734 45178
rect 6734 45126 6746 45178
rect 6746 45126 6760 45178
rect 6784 45126 6798 45178
rect 6798 45126 6810 45178
rect 6810 45126 6840 45178
rect 6864 45126 6874 45178
rect 6874 45126 6920 45178
rect 6624 45124 6680 45126
rect 6704 45124 6760 45126
rect 6784 45124 6840 45126
rect 6864 45124 6920 45126
rect 17728 87066 17784 87068
rect 17808 87066 17864 87068
rect 17888 87066 17944 87068
rect 17968 87066 18024 87068
rect 17728 87014 17774 87066
rect 17774 87014 17784 87066
rect 17808 87014 17838 87066
rect 17838 87014 17850 87066
rect 17850 87014 17864 87066
rect 17888 87014 17902 87066
rect 17902 87014 17914 87066
rect 17914 87014 17944 87066
rect 17968 87014 17978 87066
rect 17978 87014 18024 87066
rect 17728 87012 17784 87014
rect 17808 87012 17864 87014
rect 17888 87012 17944 87014
rect 17968 87012 18024 87014
rect 17728 85978 17784 85980
rect 17808 85978 17864 85980
rect 17888 85978 17944 85980
rect 17968 85978 18024 85980
rect 17728 85926 17774 85978
rect 17774 85926 17784 85978
rect 17808 85926 17838 85978
rect 17838 85926 17850 85978
rect 17850 85926 17864 85978
rect 17888 85926 17902 85978
rect 17902 85926 17914 85978
rect 17914 85926 17944 85978
rect 17968 85926 17978 85978
rect 17978 85926 18024 85978
rect 17728 85924 17784 85926
rect 17808 85924 17864 85926
rect 17888 85924 17944 85926
rect 17968 85924 18024 85926
rect 17728 84890 17784 84892
rect 17808 84890 17864 84892
rect 17888 84890 17944 84892
rect 17968 84890 18024 84892
rect 17728 84838 17774 84890
rect 17774 84838 17784 84890
rect 17808 84838 17838 84890
rect 17838 84838 17850 84890
rect 17850 84838 17864 84890
rect 17888 84838 17902 84890
rect 17902 84838 17914 84890
rect 17914 84838 17944 84890
rect 17968 84838 17978 84890
rect 17978 84838 18024 84890
rect 17728 84836 17784 84838
rect 17808 84836 17864 84838
rect 17888 84836 17944 84838
rect 17968 84836 18024 84838
rect 18388 86522 18444 86524
rect 18468 86522 18524 86524
rect 18548 86522 18604 86524
rect 18628 86522 18684 86524
rect 18388 86470 18434 86522
rect 18434 86470 18444 86522
rect 18468 86470 18498 86522
rect 18498 86470 18510 86522
rect 18510 86470 18524 86522
rect 18548 86470 18562 86522
rect 18562 86470 18574 86522
rect 18574 86470 18604 86522
rect 18628 86470 18638 86522
rect 18638 86470 18684 86522
rect 18388 86468 18444 86470
rect 18468 86468 18524 86470
rect 18548 86468 18604 86470
rect 18628 86468 18684 86470
rect 18388 85434 18444 85436
rect 18468 85434 18524 85436
rect 18548 85434 18604 85436
rect 18628 85434 18684 85436
rect 18388 85382 18434 85434
rect 18434 85382 18444 85434
rect 18468 85382 18498 85434
rect 18498 85382 18510 85434
rect 18510 85382 18524 85434
rect 18548 85382 18562 85434
rect 18562 85382 18574 85434
rect 18574 85382 18604 85434
rect 18628 85382 18638 85434
rect 18638 85382 18684 85434
rect 18388 85380 18444 85382
rect 18468 85380 18524 85382
rect 18548 85380 18604 85382
rect 18628 85380 18684 85382
rect 18388 84346 18444 84348
rect 18468 84346 18524 84348
rect 18548 84346 18604 84348
rect 18628 84346 18684 84348
rect 18388 84294 18434 84346
rect 18434 84294 18444 84346
rect 18468 84294 18498 84346
rect 18498 84294 18510 84346
rect 18510 84294 18524 84346
rect 18548 84294 18562 84346
rect 18562 84294 18574 84346
rect 18574 84294 18604 84346
rect 18628 84294 18638 84346
rect 18638 84294 18684 84346
rect 18388 84292 18444 84294
rect 18468 84292 18524 84294
rect 18548 84292 18604 84294
rect 18628 84292 18684 84294
rect 36788 87610 36844 87612
rect 36868 87610 36924 87612
rect 36948 87610 37004 87612
rect 37028 87610 37084 87612
rect 36788 87558 36834 87610
rect 36834 87558 36844 87610
rect 36868 87558 36898 87610
rect 36898 87558 36910 87610
rect 36910 87558 36924 87610
rect 36948 87558 36962 87610
rect 36962 87558 36974 87610
rect 36974 87558 37004 87610
rect 37028 87558 37038 87610
rect 37038 87558 37084 87610
rect 36788 87556 36844 87558
rect 36868 87556 36924 87558
rect 36948 87556 37004 87558
rect 37028 87556 37084 87558
rect 36128 87066 36184 87068
rect 36208 87066 36264 87068
rect 36288 87066 36344 87068
rect 36368 87066 36424 87068
rect 36128 87014 36174 87066
rect 36174 87014 36184 87066
rect 36208 87014 36238 87066
rect 36238 87014 36250 87066
rect 36250 87014 36264 87066
rect 36288 87014 36302 87066
rect 36302 87014 36314 87066
rect 36314 87014 36344 87066
rect 36368 87014 36378 87066
rect 36378 87014 36424 87066
rect 36128 87012 36184 87014
rect 36208 87012 36264 87014
rect 36288 87012 36344 87014
rect 36368 87012 36424 87014
rect 36128 85978 36184 85980
rect 36208 85978 36264 85980
rect 36288 85978 36344 85980
rect 36368 85978 36424 85980
rect 36128 85926 36174 85978
rect 36174 85926 36184 85978
rect 36208 85926 36238 85978
rect 36238 85926 36250 85978
rect 36250 85926 36264 85978
rect 36288 85926 36302 85978
rect 36302 85926 36314 85978
rect 36314 85926 36344 85978
rect 36368 85926 36378 85978
rect 36378 85926 36424 85978
rect 36128 85924 36184 85926
rect 36208 85924 36264 85926
rect 36288 85924 36344 85926
rect 36368 85924 36424 85926
rect 36128 84890 36184 84892
rect 36208 84890 36264 84892
rect 36288 84890 36344 84892
rect 36368 84890 36424 84892
rect 36128 84838 36174 84890
rect 36174 84838 36184 84890
rect 36208 84838 36238 84890
rect 36238 84838 36250 84890
rect 36250 84838 36264 84890
rect 36288 84838 36302 84890
rect 36302 84838 36314 84890
rect 36314 84838 36344 84890
rect 36368 84838 36378 84890
rect 36378 84838 36424 84890
rect 36128 84836 36184 84838
rect 36208 84836 36264 84838
rect 36288 84836 36344 84838
rect 36368 84836 36424 84838
rect 36788 86522 36844 86524
rect 36868 86522 36924 86524
rect 36948 86522 37004 86524
rect 37028 86522 37084 86524
rect 36788 86470 36834 86522
rect 36834 86470 36844 86522
rect 36868 86470 36898 86522
rect 36898 86470 36910 86522
rect 36910 86470 36924 86522
rect 36948 86470 36962 86522
rect 36962 86470 36974 86522
rect 36974 86470 37004 86522
rect 37028 86470 37038 86522
rect 37038 86470 37084 86522
rect 36788 86468 36844 86470
rect 36868 86468 36924 86470
rect 36948 86468 37004 86470
rect 37028 86468 37084 86470
rect 36788 85434 36844 85436
rect 36868 85434 36924 85436
rect 36948 85434 37004 85436
rect 37028 85434 37084 85436
rect 36788 85382 36834 85434
rect 36834 85382 36844 85434
rect 36868 85382 36898 85434
rect 36898 85382 36910 85434
rect 36910 85382 36924 85434
rect 36948 85382 36962 85434
rect 36962 85382 36974 85434
rect 36974 85382 37004 85434
rect 37028 85382 37038 85434
rect 37038 85382 37084 85434
rect 36788 85380 36844 85382
rect 36868 85380 36924 85382
rect 36948 85380 37004 85382
rect 37028 85380 37084 85382
rect 36788 84346 36844 84348
rect 36868 84346 36924 84348
rect 36948 84346 37004 84348
rect 37028 84346 37084 84348
rect 36788 84294 36834 84346
rect 36834 84294 36844 84346
rect 36868 84294 36898 84346
rect 36898 84294 36910 84346
rect 36910 84294 36924 84346
rect 36948 84294 36962 84346
rect 36962 84294 36974 84346
rect 36974 84294 37004 84346
rect 37028 84294 37038 84346
rect 37038 84294 37084 84346
rect 36788 84292 36844 84294
rect 36868 84292 36924 84294
rect 36948 84292 37004 84294
rect 37028 84292 37084 84294
rect 55188 87610 55244 87612
rect 55268 87610 55324 87612
rect 55348 87610 55404 87612
rect 55428 87610 55484 87612
rect 55188 87558 55234 87610
rect 55234 87558 55244 87610
rect 55268 87558 55298 87610
rect 55298 87558 55310 87610
rect 55310 87558 55324 87610
rect 55348 87558 55362 87610
rect 55362 87558 55374 87610
rect 55374 87558 55404 87610
rect 55428 87558 55438 87610
rect 55438 87558 55484 87610
rect 55188 87556 55244 87558
rect 55268 87556 55324 87558
rect 55348 87556 55404 87558
rect 55428 87556 55484 87558
rect 9918 56932 9920 56952
rect 9920 56932 9972 56952
rect 9972 56932 9974 56952
rect 9918 56896 9974 56932
rect 9918 56216 9974 56272
rect 45982 50504 46038 50560
rect 45890 49416 45946 49472
rect 11666 45880 11722 45936
rect 12770 45880 12826 45936
rect 13874 45880 13930 45936
rect 8998 45492 9054 45528
rect 8998 45472 9000 45492
rect 9000 45472 9052 45492
rect 9052 45472 9054 45492
rect 9826 45472 9882 45528
rect 8538 44656 8594 44712
rect 5888 44634 5944 44636
rect 5968 44634 6024 44636
rect 6048 44634 6104 44636
rect 6128 44634 6184 44636
rect 4214 44520 4270 44576
rect 5888 44582 5934 44634
rect 5934 44582 5944 44634
rect 5968 44582 5998 44634
rect 5998 44582 6010 44634
rect 6010 44582 6024 44634
rect 6048 44582 6062 44634
rect 6062 44582 6074 44634
rect 6074 44582 6104 44634
rect 6128 44582 6138 44634
rect 6138 44582 6184 44634
rect 5888 44580 5944 44582
rect 5968 44580 6024 44582
rect 6048 44580 6104 44582
rect 6128 44580 6184 44582
rect 6624 44090 6680 44092
rect 6704 44090 6760 44092
rect 6784 44090 6840 44092
rect 6864 44090 6920 44092
rect 6624 44038 6670 44090
rect 6670 44038 6680 44090
rect 6704 44038 6734 44090
rect 6734 44038 6746 44090
rect 6746 44038 6760 44090
rect 6784 44038 6798 44090
rect 6798 44038 6810 44090
rect 6810 44038 6840 44090
rect 6864 44038 6874 44090
rect 6874 44038 6920 44090
rect 6624 44036 6680 44038
rect 6704 44036 6760 44038
rect 6784 44036 6840 44038
rect 6864 44036 6920 44038
rect 5888 43546 5944 43548
rect 5968 43546 6024 43548
rect 6048 43546 6104 43548
rect 6128 43546 6184 43548
rect 5888 43494 5934 43546
rect 5934 43494 5944 43546
rect 5968 43494 5998 43546
rect 5998 43494 6010 43546
rect 6010 43494 6024 43546
rect 6048 43494 6062 43546
rect 6062 43494 6074 43546
rect 6074 43494 6104 43546
rect 6128 43494 6138 43546
rect 6138 43494 6184 43546
rect 5888 43492 5944 43494
rect 5968 43492 6024 43494
rect 6048 43492 6104 43494
rect 6128 43492 6184 43494
rect 8538 43432 8594 43488
rect 4122 43196 4124 43216
rect 4124 43196 4176 43216
rect 4176 43196 4178 43216
rect 4122 43160 4178 43196
rect 6624 43002 6680 43004
rect 6704 43002 6760 43004
rect 6784 43002 6840 43004
rect 6864 43002 6920 43004
rect 6624 42950 6670 43002
rect 6670 42950 6680 43002
rect 6704 42950 6734 43002
rect 6734 42950 6746 43002
rect 6746 42950 6760 43002
rect 6784 42950 6798 43002
rect 6798 42950 6810 43002
rect 6810 42950 6840 43002
rect 6864 42950 6874 43002
rect 6874 42950 6920 43002
rect 6624 42948 6680 42950
rect 6704 42948 6760 42950
rect 6784 42948 6840 42950
rect 6864 42948 6920 42950
rect 4122 42516 4124 42536
rect 4124 42516 4176 42536
rect 4176 42516 4178 42536
rect 4122 42480 4178 42516
rect 8538 42480 8594 42536
rect 5888 42458 5944 42460
rect 5968 42458 6024 42460
rect 6048 42458 6104 42460
rect 6128 42458 6184 42460
rect 5888 42406 5934 42458
rect 5934 42406 5944 42458
rect 5968 42406 5998 42458
rect 5998 42406 6010 42458
rect 6010 42406 6024 42458
rect 6048 42406 6062 42458
rect 6062 42406 6074 42458
rect 6074 42406 6104 42458
rect 6128 42406 6138 42458
rect 6138 42406 6184 42458
rect 5888 42404 5944 42406
rect 5968 42404 6024 42406
rect 6048 42404 6104 42406
rect 6128 42404 6184 42406
rect 6624 41914 6680 41916
rect 6704 41914 6760 41916
rect 6784 41914 6840 41916
rect 6864 41914 6920 41916
rect 6624 41862 6670 41914
rect 6670 41862 6680 41914
rect 6704 41862 6734 41914
rect 6734 41862 6746 41914
rect 6746 41862 6760 41914
rect 6784 41862 6798 41914
rect 6798 41862 6810 41914
rect 6810 41862 6840 41914
rect 6864 41862 6874 41914
rect 6874 41862 6920 41914
rect 6624 41860 6680 41862
rect 6704 41860 6760 41862
rect 6784 41860 6840 41862
rect 6864 41860 6920 41862
rect 5410 41528 5466 41584
rect 5888 41370 5944 41372
rect 5968 41370 6024 41372
rect 6048 41370 6104 41372
rect 6128 41370 6184 41372
rect 5888 41318 5934 41370
rect 5934 41318 5944 41370
rect 5968 41318 5998 41370
rect 5998 41318 6010 41370
rect 6010 41318 6024 41370
rect 6048 41318 6062 41370
rect 6062 41318 6074 41370
rect 6074 41318 6104 41370
rect 6128 41318 6138 41370
rect 6138 41318 6184 41370
rect 5888 41316 5944 41318
rect 5968 41316 6024 41318
rect 6048 41316 6104 41318
rect 6128 41316 6184 41318
rect 4122 41120 4178 41176
rect 6624 40826 6680 40828
rect 6704 40826 6760 40828
rect 6784 40826 6840 40828
rect 6864 40826 6920 40828
rect 6624 40774 6670 40826
rect 6670 40774 6680 40826
rect 6704 40774 6734 40826
rect 6734 40774 6746 40826
rect 6746 40774 6760 40826
rect 6784 40774 6798 40826
rect 6798 40774 6810 40826
rect 6810 40774 6840 40826
rect 6864 40774 6874 40826
rect 6874 40774 6920 40826
rect 6624 40772 6680 40774
rect 6704 40772 6760 40774
rect 6784 40772 6840 40774
rect 6864 40772 6920 40774
rect 3938 40460 3994 40496
rect 3938 40440 3940 40460
rect 3940 40440 3992 40460
rect 3992 40440 3994 40460
rect 8538 40304 8594 40360
rect 5888 40282 5944 40284
rect 5968 40282 6024 40284
rect 6048 40282 6104 40284
rect 6128 40282 6184 40284
rect 5888 40230 5934 40282
rect 5934 40230 5944 40282
rect 5968 40230 5998 40282
rect 5998 40230 6010 40282
rect 6010 40230 6024 40282
rect 6048 40230 6062 40282
rect 6062 40230 6074 40282
rect 6074 40230 6104 40282
rect 6128 40230 6138 40282
rect 6138 40230 6184 40282
rect 5888 40228 5944 40230
rect 5968 40228 6024 40230
rect 6048 40228 6104 40230
rect 6128 40228 6184 40230
rect 6624 39738 6680 39740
rect 6704 39738 6760 39740
rect 6784 39738 6840 39740
rect 6864 39738 6920 39740
rect 6624 39686 6670 39738
rect 6670 39686 6680 39738
rect 6704 39686 6734 39738
rect 6734 39686 6746 39738
rect 6746 39686 6760 39738
rect 6784 39686 6798 39738
rect 6798 39686 6810 39738
rect 6810 39686 6840 39738
rect 6864 39686 6874 39738
rect 6874 39686 6920 39738
rect 6624 39684 6680 39686
rect 6704 39684 6760 39686
rect 6784 39684 6840 39686
rect 6864 39684 6920 39686
rect 8538 39216 8594 39272
rect 5888 39194 5944 39196
rect 5968 39194 6024 39196
rect 6048 39194 6104 39196
rect 6128 39194 6184 39196
rect 4214 39080 4270 39136
rect 5888 39142 5934 39194
rect 5934 39142 5944 39194
rect 5968 39142 5998 39194
rect 5998 39142 6010 39194
rect 6010 39142 6024 39194
rect 6048 39142 6062 39194
rect 6062 39142 6074 39194
rect 6074 39142 6104 39194
rect 6128 39142 6138 39194
rect 6138 39142 6184 39194
rect 5888 39140 5944 39142
rect 5968 39140 6024 39142
rect 6048 39140 6104 39142
rect 6128 39140 6184 39142
rect 6624 38650 6680 38652
rect 6704 38650 6760 38652
rect 6784 38650 6840 38652
rect 6864 38650 6920 38652
rect 6624 38598 6670 38650
rect 6670 38598 6680 38650
rect 6704 38598 6734 38650
rect 6734 38598 6746 38650
rect 6746 38598 6760 38650
rect 6784 38598 6798 38650
rect 6798 38598 6810 38650
rect 6810 38598 6840 38650
rect 6864 38598 6874 38650
rect 6874 38598 6920 38650
rect 6624 38596 6680 38598
rect 6704 38596 6760 38598
rect 6784 38596 6840 38598
rect 6864 38596 6920 38598
rect 5888 38106 5944 38108
rect 5968 38106 6024 38108
rect 6048 38106 6104 38108
rect 6128 38106 6184 38108
rect 5888 38054 5934 38106
rect 5934 38054 5944 38106
rect 5968 38054 5998 38106
rect 5998 38054 6010 38106
rect 6010 38054 6024 38106
rect 6048 38054 6062 38106
rect 6062 38054 6074 38106
rect 6074 38054 6104 38106
rect 6128 38054 6138 38106
rect 6138 38054 6184 38106
rect 5888 38052 5944 38054
rect 5968 38052 6024 38054
rect 6048 38052 6104 38054
rect 6128 38052 6184 38054
rect 8538 37992 8594 38048
rect 4214 37756 4216 37776
rect 4216 37756 4268 37776
rect 4268 37756 4270 37776
rect 4214 37720 4270 37756
rect 6624 37562 6680 37564
rect 6704 37562 6760 37564
rect 6784 37562 6840 37564
rect 6864 37562 6920 37564
rect 6624 37510 6670 37562
rect 6670 37510 6680 37562
rect 6704 37510 6734 37562
rect 6734 37510 6746 37562
rect 6746 37510 6760 37562
rect 6784 37510 6798 37562
rect 6798 37510 6810 37562
rect 6810 37510 6840 37562
rect 6864 37510 6874 37562
rect 6874 37510 6920 37562
rect 6624 37508 6680 37510
rect 6704 37508 6760 37510
rect 6784 37508 6840 37510
rect 6864 37508 6920 37510
rect 4122 37076 4124 37096
rect 4124 37076 4176 37096
rect 4176 37076 4178 37096
rect 4122 37040 4178 37076
rect 8538 37040 8594 37096
rect 5888 37018 5944 37020
rect 5968 37018 6024 37020
rect 6048 37018 6104 37020
rect 6128 37018 6184 37020
rect 5888 36966 5934 37018
rect 5934 36966 5944 37018
rect 5968 36966 5998 37018
rect 5998 36966 6010 37018
rect 6010 36966 6024 37018
rect 6048 36966 6062 37018
rect 6062 36966 6074 37018
rect 6074 36966 6104 37018
rect 6128 36966 6138 37018
rect 6138 36966 6184 37018
rect 5888 36964 5944 36966
rect 5968 36964 6024 36966
rect 6048 36964 6104 36966
rect 6128 36964 6184 36966
rect 6624 36474 6680 36476
rect 6704 36474 6760 36476
rect 6784 36474 6840 36476
rect 6864 36474 6920 36476
rect 6624 36422 6670 36474
rect 6670 36422 6680 36474
rect 6704 36422 6734 36474
rect 6734 36422 6746 36474
rect 6746 36422 6760 36474
rect 6784 36422 6798 36474
rect 6798 36422 6810 36474
rect 6810 36422 6840 36474
rect 6864 36422 6874 36474
rect 6874 36422 6920 36474
rect 6624 36420 6680 36422
rect 6704 36420 6760 36422
rect 6784 36420 6840 36422
rect 6864 36420 6920 36422
rect 5410 36088 5466 36144
rect 5888 35930 5944 35932
rect 5968 35930 6024 35932
rect 6048 35930 6104 35932
rect 6128 35930 6184 35932
rect 5888 35878 5934 35930
rect 5934 35878 5944 35930
rect 5968 35878 5998 35930
rect 5998 35878 6010 35930
rect 6010 35878 6024 35930
rect 6048 35878 6062 35930
rect 6062 35878 6074 35930
rect 6074 35878 6104 35930
rect 6128 35878 6138 35930
rect 6138 35878 6184 35930
rect 5888 35876 5944 35878
rect 5968 35876 6024 35878
rect 6048 35876 6104 35878
rect 6128 35876 6184 35878
rect 4122 35680 4178 35736
rect 6624 35386 6680 35388
rect 6704 35386 6760 35388
rect 6784 35386 6840 35388
rect 6864 35386 6920 35388
rect 6624 35334 6670 35386
rect 6670 35334 6680 35386
rect 6704 35334 6734 35386
rect 6734 35334 6746 35386
rect 6746 35334 6760 35386
rect 6784 35334 6798 35386
rect 6798 35334 6810 35386
rect 6810 35334 6840 35386
rect 6864 35334 6874 35386
rect 6874 35334 6920 35386
rect 6624 35332 6680 35334
rect 6704 35332 6760 35334
rect 6784 35332 6840 35334
rect 6864 35332 6920 35334
rect 4214 35036 4216 35056
rect 4216 35036 4268 35056
rect 4268 35036 4270 35056
rect 4214 35000 4270 35036
rect 8538 34864 8594 34920
rect 5888 34842 5944 34844
rect 5968 34842 6024 34844
rect 6048 34842 6104 34844
rect 6128 34842 6184 34844
rect 5888 34790 5934 34842
rect 5934 34790 5944 34842
rect 5968 34790 5998 34842
rect 5998 34790 6010 34842
rect 6010 34790 6024 34842
rect 6048 34790 6062 34842
rect 6062 34790 6074 34842
rect 6074 34790 6104 34842
rect 6128 34790 6138 34842
rect 6138 34790 6184 34842
rect 5888 34788 5944 34790
rect 5968 34788 6024 34790
rect 6048 34788 6104 34790
rect 6128 34788 6184 34790
rect 6624 34298 6680 34300
rect 6704 34298 6760 34300
rect 6784 34298 6840 34300
rect 6864 34298 6920 34300
rect 6624 34246 6670 34298
rect 6670 34246 6680 34298
rect 6704 34246 6734 34298
rect 6734 34246 6746 34298
rect 6746 34246 6760 34298
rect 6784 34246 6798 34298
rect 6798 34246 6810 34298
rect 6810 34246 6840 34298
rect 6864 34246 6874 34298
rect 6874 34246 6920 34298
rect 6624 34244 6680 34246
rect 6704 34244 6760 34246
rect 6784 34244 6840 34246
rect 6864 34244 6920 34246
rect 8538 33776 8594 33832
rect 5888 33754 5944 33756
rect 5968 33754 6024 33756
rect 6048 33754 6104 33756
rect 6128 33754 6184 33756
rect 4214 33640 4270 33696
rect 5888 33702 5934 33754
rect 5934 33702 5944 33754
rect 5968 33702 5998 33754
rect 5998 33702 6010 33754
rect 6010 33702 6024 33754
rect 6048 33702 6062 33754
rect 6062 33702 6074 33754
rect 6074 33702 6104 33754
rect 6128 33702 6138 33754
rect 6138 33702 6184 33754
rect 5888 33700 5944 33702
rect 5968 33700 6024 33702
rect 6048 33700 6104 33702
rect 6128 33700 6184 33702
rect 6624 33210 6680 33212
rect 6704 33210 6760 33212
rect 6784 33210 6840 33212
rect 6864 33210 6920 33212
rect 6624 33158 6670 33210
rect 6670 33158 6680 33210
rect 6704 33158 6734 33210
rect 6734 33158 6746 33210
rect 6746 33158 6760 33210
rect 6784 33158 6798 33210
rect 6798 33158 6810 33210
rect 6810 33158 6840 33210
rect 6864 33158 6874 33210
rect 6874 33158 6920 33210
rect 6624 33156 6680 33158
rect 6704 33156 6760 33158
rect 6784 33156 6840 33158
rect 6864 33156 6920 33158
rect 5888 32666 5944 32668
rect 5968 32666 6024 32668
rect 6048 32666 6104 32668
rect 6128 32666 6184 32668
rect 5888 32614 5934 32666
rect 5934 32614 5944 32666
rect 5968 32614 5998 32666
rect 5998 32614 6010 32666
rect 6010 32614 6024 32666
rect 6048 32614 6062 32666
rect 6062 32614 6074 32666
rect 6074 32614 6104 32666
rect 6128 32614 6138 32666
rect 6138 32614 6184 32666
rect 5888 32612 5944 32614
rect 5968 32612 6024 32614
rect 6048 32612 6104 32614
rect 6128 32612 6184 32614
rect 8538 32552 8594 32608
rect 4214 32316 4216 32336
rect 4216 32316 4268 32336
rect 4268 32316 4270 32336
rect 4214 32280 4270 32316
rect 6624 32122 6680 32124
rect 6704 32122 6760 32124
rect 6784 32122 6840 32124
rect 6864 32122 6920 32124
rect 6624 32070 6670 32122
rect 6670 32070 6680 32122
rect 6704 32070 6734 32122
rect 6734 32070 6746 32122
rect 6746 32070 6760 32122
rect 6784 32070 6798 32122
rect 6798 32070 6810 32122
rect 6810 32070 6840 32122
rect 6864 32070 6874 32122
rect 6874 32070 6920 32122
rect 6624 32068 6680 32070
rect 6704 32068 6760 32070
rect 6784 32068 6840 32070
rect 6864 32068 6920 32070
rect 4122 31636 4124 31656
rect 4124 31636 4176 31656
rect 4176 31636 4178 31656
rect 4122 31600 4178 31636
rect 8538 31600 8594 31656
rect 5888 31578 5944 31580
rect 5968 31578 6024 31580
rect 6048 31578 6104 31580
rect 6128 31578 6184 31580
rect 5888 31526 5934 31578
rect 5934 31526 5944 31578
rect 5968 31526 5998 31578
rect 5998 31526 6010 31578
rect 6010 31526 6024 31578
rect 6048 31526 6062 31578
rect 6062 31526 6074 31578
rect 6074 31526 6104 31578
rect 6128 31526 6138 31578
rect 6138 31526 6184 31578
rect 5888 31524 5944 31526
rect 5968 31524 6024 31526
rect 6048 31524 6104 31526
rect 6128 31524 6184 31526
rect 6624 31034 6680 31036
rect 6704 31034 6760 31036
rect 6784 31034 6840 31036
rect 6864 31034 6920 31036
rect 6624 30982 6670 31034
rect 6670 30982 6680 31034
rect 6704 30982 6734 31034
rect 6734 30982 6746 31034
rect 6746 30982 6760 31034
rect 6784 30982 6798 31034
rect 6798 30982 6810 31034
rect 6810 30982 6840 31034
rect 6864 30982 6874 31034
rect 6874 30982 6920 31034
rect 6624 30980 6680 30982
rect 6704 30980 6760 30982
rect 6784 30980 6840 30982
rect 6864 30980 6920 30982
rect 5888 30490 5944 30492
rect 5968 30490 6024 30492
rect 6048 30490 6104 30492
rect 6128 30490 6184 30492
rect 5888 30438 5934 30490
rect 5934 30438 5944 30490
rect 5968 30438 5998 30490
rect 5998 30438 6010 30490
rect 6010 30438 6024 30490
rect 6048 30438 6062 30490
rect 6062 30438 6074 30490
rect 6074 30438 6104 30490
rect 6128 30438 6138 30490
rect 6138 30438 6184 30490
rect 5888 30436 5944 30438
rect 5968 30436 6024 30438
rect 6048 30436 6104 30438
rect 6128 30436 6184 30438
rect 4122 30240 4178 30296
rect 5410 30240 5466 30296
rect 6624 29946 6680 29948
rect 6704 29946 6760 29948
rect 6784 29946 6840 29948
rect 6864 29946 6920 29948
rect 6624 29894 6670 29946
rect 6670 29894 6680 29946
rect 6704 29894 6734 29946
rect 6734 29894 6746 29946
rect 6746 29894 6760 29946
rect 6784 29894 6798 29946
rect 6798 29894 6810 29946
rect 6810 29894 6840 29946
rect 6864 29894 6874 29946
rect 6874 29894 6920 29946
rect 6624 29892 6680 29894
rect 6704 29892 6760 29894
rect 6784 29892 6840 29894
rect 6864 29892 6920 29894
rect 4306 29560 4362 29616
rect 8538 29424 8594 29480
rect 5888 29402 5944 29404
rect 5968 29402 6024 29404
rect 6048 29402 6104 29404
rect 6128 29402 6184 29404
rect 5888 29350 5934 29402
rect 5934 29350 5944 29402
rect 5968 29350 5998 29402
rect 5998 29350 6010 29402
rect 6010 29350 6024 29402
rect 6048 29350 6062 29402
rect 6062 29350 6074 29402
rect 6074 29350 6104 29402
rect 6128 29350 6138 29402
rect 6138 29350 6184 29402
rect 5888 29348 5944 29350
rect 5968 29348 6024 29350
rect 6048 29348 6104 29350
rect 6128 29348 6184 29350
rect 6624 28858 6680 28860
rect 6704 28858 6760 28860
rect 6784 28858 6840 28860
rect 6864 28858 6920 28860
rect 6624 28806 6670 28858
rect 6670 28806 6680 28858
rect 6704 28806 6734 28858
rect 6734 28806 6746 28858
rect 6746 28806 6760 28858
rect 6784 28806 6798 28858
rect 6798 28806 6810 28858
rect 6810 28806 6840 28858
rect 6864 28806 6874 28858
rect 6874 28806 6920 28858
rect 6624 28804 6680 28806
rect 6704 28804 6760 28806
rect 6784 28804 6840 28806
rect 6864 28804 6920 28806
rect 8538 28336 8594 28392
rect 5888 28314 5944 28316
rect 5968 28314 6024 28316
rect 6048 28314 6104 28316
rect 6128 28314 6184 28316
rect 4306 28200 4362 28256
rect 5888 28262 5934 28314
rect 5934 28262 5944 28314
rect 5968 28262 5998 28314
rect 5998 28262 6010 28314
rect 6010 28262 6024 28314
rect 6048 28262 6062 28314
rect 6062 28262 6074 28314
rect 6074 28262 6104 28314
rect 6128 28262 6138 28314
rect 6138 28262 6184 28314
rect 5888 28260 5944 28262
rect 5968 28260 6024 28262
rect 6048 28260 6104 28262
rect 6128 28260 6184 28262
rect 6624 27770 6680 27772
rect 6704 27770 6760 27772
rect 6784 27770 6840 27772
rect 6864 27770 6920 27772
rect 6624 27718 6670 27770
rect 6670 27718 6680 27770
rect 6704 27718 6734 27770
rect 6734 27718 6746 27770
rect 6746 27718 6760 27770
rect 6784 27718 6798 27770
rect 6798 27718 6810 27770
rect 6810 27718 6840 27770
rect 6864 27718 6874 27770
rect 6874 27718 6920 27770
rect 6624 27716 6680 27718
rect 6704 27716 6760 27718
rect 6784 27716 6840 27718
rect 6864 27716 6920 27718
rect 5888 27226 5944 27228
rect 5968 27226 6024 27228
rect 6048 27226 6104 27228
rect 6128 27226 6184 27228
rect 5888 27174 5934 27226
rect 5934 27174 5944 27226
rect 5968 27174 5998 27226
rect 5998 27174 6010 27226
rect 6010 27174 6024 27226
rect 6048 27174 6062 27226
rect 6062 27174 6074 27226
rect 6074 27174 6104 27226
rect 6128 27174 6138 27226
rect 6138 27174 6184 27226
rect 5888 27172 5944 27174
rect 5968 27172 6024 27174
rect 6048 27172 6104 27174
rect 6128 27172 6184 27174
rect 8538 27112 8594 27168
rect 4306 26876 4308 26896
rect 4308 26876 4360 26896
rect 4360 26876 4362 26896
rect 4306 26840 4362 26876
rect 6624 26682 6680 26684
rect 6704 26682 6760 26684
rect 6784 26682 6840 26684
rect 6864 26682 6920 26684
rect 6624 26630 6670 26682
rect 6670 26630 6680 26682
rect 6704 26630 6734 26682
rect 6734 26630 6746 26682
rect 6746 26630 6760 26682
rect 6784 26630 6798 26682
rect 6798 26630 6810 26682
rect 6810 26630 6840 26682
rect 6864 26630 6874 26682
rect 6874 26630 6920 26682
rect 6624 26628 6680 26630
rect 6704 26628 6760 26630
rect 6784 26628 6840 26630
rect 6864 26628 6920 26630
rect 4306 26160 4362 26216
rect 8538 26160 8594 26216
rect 5888 26138 5944 26140
rect 5968 26138 6024 26140
rect 6048 26138 6104 26140
rect 6128 26138 6184 26140
rect 5888 26086 5934 26138
rect 5934 26086 5944 26138
rect 5968 26086 5998 26138
rect 5998 26086 6010 26138
rect 6010 26086 6024 26138
rect 6048 26086 6062 26138
rect 6062 26086 6074 26138
rect 6074 26086 6104 26138
rect 6128 26086 6138 26138
rect 6138 26086 6184 26138
rect 5888 26084 5944 26086
rect 5968 26084 6024 26086
rect 6048 26084 6104 26086
rect 6128 26084 6184 26086
rect 6624 25594 6680 25596
rect 6704 25594 6760 25596
rect 6784 25594 6840 25596
rect 6864 25594 6920 25596
rect 6624 25542 6670 25594
rect 6670 25542 6680 25594
rect 6704 25542 6734 25594
rect 6734 25542 6746 25594
rect 6746 25542 6760 25594
rect 6784 25542 6798 25594
rect 6798 25542 6810 25594
rect 6810 25542 6840 25594
rect 6864 25542 6874 25594
rect 6874 25542 6920 25594
rect 6624 25540 6680 25542
rect 6704 25540 6760 25542
rect 6784 25540 6840 25542
rect 6864 25540 6920 25542
rect 5888 25050 5944 25052
rect 5968 25050 6024 25052
rect 6048 25050 6104 25052
rect 6128 25050 6184 25052
rect 5888 24998 5934 25050
rect 5934 24998 5944 25050
rect 5968 24998 5998 25050
rect 5998 24998 6010 25050
rect 6010 24998 6024 25050
rect 6048 24998 6062 25050
rect 6062 24998 6074 25050
rect 6074 24998 6104 25050
rect 6128 24998 6138 25050
rect 6138 24998 6184 25050
rect 5888 24996 5944 24998
rect 5968 24996 6024 24998
rect 6048 24996 6104 24998
rect 6128 24996 6184 24998
rect 4306 24800 4362 24856
rect 5410 24800 5466 24856
rect 6624 24506 6680 24508
rect 6704 24506 6760 24508
rect 6784 24506 6840 24508
rect 6864 24506 6920 24508
rect 6624 24454 6670 24506
rect 6670 24454 6680 24506
rect 6704 24454 6734 24506
rect 6734 24454 6746 24506
rect 6746 24454 6760 24506
rect 6784 24454 6798 24506
rect 6798 24454 6810 24506
rect 6810 24454 6840 24506
rect 6864 24454 6874 24506
rect 6874 24454 6920 24506
rect 6624 24452 6680 24454
rect 6704 24452 6760 24454
rect 6784 24452 6840 24454
rect 6864 24452 6920 24454
rect 4306 24120 4362 24176
rect 8538 23984 8594 24040
rect 5888 23962 5944 23964
rect 5968 23962 6024 23964
rect 6048 23962 6104 23964
rect 6128 23962 6184 23964
rect 5888 23910 5934 23962
rect 5934 23910 5944 23962
rect 5968 23910 5998 23962
rect 5998 23910 6010 23962
rect 6010 23910 6024 23962
rect 6048 23910 6062 23962
rect 6062 23910 6074 23962
rect 6074 23910 6104 23962
rect 6128 23910 6138 23962
rect 6138 23910 6184 23962
rect 5888 23908 5944 23910
rect 5968 23908 6024 23910
rect 6048 23908 6104 23910
rect 6128 23908 6184 23910
rect 6624 23418 6680 23420
rect 6704 23418 6760 23420
rect 6784 23418 6840 23420
rect 6864 23418 6920 23420
rect 6624 23366 6670 23418
rect 6670 23366 6680 23418
rect 6704 23366 6734 23418
rect 6734 23366 6746 23418
rect 6746 23366 6760 23418
rect 6784 23366 6798 23418
rect 6798 23366 6810 23418
rect 6810 23366 6840 23418
rect 6864 23366 6874 23418
rect 6874 23366 6920 23418
rect 6624 23364 6680 23366
rect 6704 23364 6760 23366
rect 6784 23364 6840 23366
rect 6864 23364 6920 23366
rect 8538 22896 8594 22952
rect 5888 22874 5944 22876
rect 5968 22874 6024 22876
rect 6048 22874 6104 22876
rect 6128 22874 6184 22876
rect 4306 22760 4362 22816
rect 5888 22822 5934 22874
rect 5934 22822 5944 22874
rect 5968 22822 5998 22874
rect 5998 22822 6010 22874
rect 6010 22822 6024 22874
rect 6048 22822 6062 22874
rect 6062 22822 6074 22874
rect 6074 22822 6104 22874
rect 6128 22822 6138 22874
rect 6138 22822 6184 22874
rect 5888 22820 5944 22822
rect 5968 22820 6024 22822
rect 6048 22820 6104 22822
rect 6128 22820 6184 22822
rect 6624 22330 6680 22332
rect 6704 22330 6760 22332
rect 6784 22330 6840 22332
rect 6864 22330 6920 22332
rect 6624 22278 6670 22330
rect 6670 22278 6680 22330
rect 6704 22278 6734 22330
rect 6734 22278 6746 22330
rect 6746 22278 6760 22330
rect 6784 22278 6798 22330
rect 6798 22278 6810 22330
rect 6810 22278 6840 22330
rect 6864 22278 6874 22330
rect 6874 22278 6920 22330
rect 6624 22276 6680 22278
rect 6704 22276 6760 22278
rect 6784 22276 6840 22278
rect 6864 22276 6920 22278
rect 5888 21786 5944 21788
rect 5968 21786 6024 21788
rect 6048 21786 6104 21788
rect 6128 21786 6184 21788
rect 5888 21734 5934 21786
rect 5934 21734 5944 21786
rect 5968 21734 5998 21786
rect 5998 21734 6010 21786
rect 6010 21734 6024 21786
rect 6048 21734 6062 21786
rect 6062 21734 6074 21786
rect 6074 21734 6104 21786
rect 6128 21734 6138 21786
rect 6138 21734 6184 21786
rect 5888 21732 5944 21734
rect 5968 21732 6024 21734
rect 6048 21732 6104 21734
rect 6128 21732 6184 21734
rect 8538 21672 8594 21728
rect 4306 21436 4308 21456
rect 4308 21436 4360 21456
rect 4360 21436 4362 21456
rect 4306 21400 4362 21436
rect 6624 21242 6680 21244
rect 6704 21242 6760 21244
rect 6784 21242 6840 21244
rect 6864 21242 6920 21244
rect 6624 21190 6670 21242
rect 6670 21190 6680 21242
rect 6704 21190 6734 21242
rect 6734 21190 6746 21242
rect 6746 21190 6760 21242
rect 6784 21190 6798 21242
rect 6798 21190 6810 21242
rect 6810 21190 6840 21242
rect 6864 21190 6874 21242
rect 6874 21190 6920 21242
rect 6624 21188 6680 21190
rect 6704 21188 6760 21190
rect 6784 21188 6840 21190
rect 6864 21188 6920 21190
rect 5686 20856 5742 20912
rect 4306 20720 4362 20776
rect 5888 20698 5944 20700
rect 5968 20698 6024 20700
rect 6048 20698 6104 20700
rect 6128 20698 6184 20700
rect 5888 20646 5934 20698
rect 5934 20646 5944 20698
rect 5968 20646 5998 20698
rect 5998 20646 6010 20698
rect 6010 20646 6024 20698
rect 6048 20646 6062 20698
rect 6062 20646 6074 20698
rect 6074 20646 6104 20698
rect 6128 20646 6138 20698
rect 6138 20646 6184 20698
rect 5888 20644 5944 20646
rect 5968 20644 6024 20646
rect 6048 20644 6104 20646
rect 6128 20644 6184 20646
rect 6624 20154 6680 20156
rect 6704 20154 6760 20156
rect 6784 20154 6840 20156
rect 6864 20154 6920 20156
rect 6624 20102 6670 20154
rect 6670 20102 6680 20154
rect 6704 20102 6734 20154
rect 6734 20102 6746 20154
rect 6746 20102 6760 20154
rect 6784 20102 6798 20154
rect 6798 20102 6810 20154
rect 6810 20102 6840 20154
rect 6864 20102 6874 20154
rect 6874 20102 6920 20154
rect 6624 20100 6680 20102
rect 6704 20100 6760 20102
rect 6784 20100 6840 20102
rect 6864 20100 6920 20102
rect 8538 19632 8594 19688
rect 5888 19610 5944 19612
rect 5968 19610 6024 19612
rect 6048 19610 6104 19612
rect 6128 19610 6184 19612
rect 5888 19558 5934 19610
rect 5934 19558 5944 19610
rect 5968 19558 5998 19610
rect 5998 19558 6010 19610
rect 6010 19558 6024 19610
rect 6048 19558 6062 19610
rect 6062 19558 6074 19610
rect 6074 19558 6104 19610
rect 6128 19558 6138 19610
rect 6138 19558 6184 19610
rect 5888 19556 5944 19558
rect 5968 19556 6024 19558
rect 6048 19556 6104 19558
rect 6128 19556 6184 19558
rect 4306 19360 4362 19416
rect 6624 19066 6680 19068
rect 6704 19066 6760 19068
rect 6784 19066 6840 19068
rect 6864 19066 6920 19068
rect 6624 19014 6670 19066
rect 6670 19014 6680 19066
rect 6704 19014 6734 19066
rect 6734 19014 6746 19066
rect 6746 19014 6760 19066
rect 6784 19014 6798 19066
rect 6798 19014 6810 19066
rect 6810 19014 6840 19066
rect 6864 19014 6874 19066
rect 6874 19014 6920 19066
rect 6624 19012 6680 19014
rect 6704 19012 6760 19014
rect 6784 19012 6840 19014
rect 6864 19012 6920 19014
rect 4306 18680 4362 18736
rect 8538 18544 8594 18600
rect 5888 18522 5944 18524
rect 5968 18522 6024 18524
rect 6048 18522 6104 18524
rect 6128 18522 6184 18524
rect 5888 18470 5934 18522
rect 5934 18470 5944 18522
rect 5968 18470 5998 18522
rect 5998 18470 6010 18522
rect 6010 18470 6024 18522
rect 6048 18470 6062 18522
rect 6062 18470 6074 18522
rect 6074 18470 6104 18522
rect 6128 18470 6138 18522
rect 6138 18470 6184 18522
rect 5888 18468 5944 18470
rect 5968 18468 6024 18470
rect 6048 18468 6104 18470
rect 6128 18468 6184 18470
rect 6624 17978 6680 17980
rect 6704 17978 6760 17980
rect 6784 17978 6840 17980
rect 6864 17978 6920 17980
rect 6624 17926 6670 17978
rect 6670 17926 6680 17978
rect 6704 17926 6734 17978
rect 6734 17926 6746 17978
rect 6746 17926 6760 17978
rect 6784 17926 6798 17978
rect 6798 17926 6810 17978
rect 6810 17926 6840 17978
rect 6864 17926 6874 17978
rect 6874 17926 6920 17978
rect 6624 17924 6680 17926
rect 6704 17924 6760 17926
rect 6784 17924 6840 17926
rect 6864 17924 6920 17926
rect 8538 17456 8594 17512
rect 5888 17434 5944 17436
rect 5968 17434 6024 17436
rect 6048 17434 6104 17436
rect 6128 17434 6184 17436
rect 4306 17320 4362 17376
rect 5888 17382 5934 17434
rect 5934 17382 5944 17434
rect 5968 17382 5998 17434
rect 5998 17382 6010 17434
rect 6010 17382 6024 17434
rect 6048 17382 6062 17434
rect 6062 17382 6074 17434
rect 6074 17382 6104 17434
rect 6128 17382 6138 17434
rect 6138 17382 6184 17434
rect 5888 17380 5944 17382
rect 5968 17380 6024 17382
rect 6048 17380 6104 17382
rect 6128 17380 6184 17382
rect 6624 16890 6680 16892
rect 6704 16890 6760 16892
rect 6784 16890 6840 16892
rect 6864 16890 6920 16892
rect 6624 16838 6670 16890
rect 6670 16838 6680 16890
rect 6704 16838 6734 16890
rect 6734 16838 6746 16890
rect 6746 16838 6760 16890
rect 6784 16838 6798 16890
rect 6798 16838 6810 16890
rect 6810 16838 6840 16890
rect 6864 16838 6874 16890
rect 6874 16838 6920 16890
rect 6624 16836 6680 16838
rect 6704 16836 6760 16838
rect 6784 16836 6840 16838
rect 6864 16836 6920 16838
rect 5888 16346 5944 16348
rect 5968 16346 6024 16348
rect 6048 16346 6104 16348
rect 6128 16346 6184 16348
rect 5888 16294 5934 16346
rect 5934 16294 5944 16346
rect 5968 16294 5998 16346
rect 5998 16294 6010 16346
rect 6010 16294 6024 16346
rect 6048 16294 6062 16346
rect 6062 16294 6074 16346
rect 6074 16294 6104 16346
rect 6128 16294 6138 16346
rect 6138 16294 6184 16346
rect 5888 16292 5944 16294
rect 5968 16292 6024 16294
rect 6048 16292 6104 16294
rect 6128 16292 6184 16294
rect 8538 16232 8594 16288
rect 4306 15996 4308 16016
rect 4308 15996 4360 16016
rect 4360 15996 4362 16016
rect 4306 15960 4362 15996
rect 6624 15802 6680 15804
rect 6704 15802 6760 15804
rect 6784 15802 6840 15804
rect 6864 15802 6920 15804
rect 6624 15750 6670 15802
rect 6670 15750 6680 15802
rect 6704 15750 6734 15802
rect 6734 15750 6746 15802
rect 6746 15750 6760 15802
rect 6784 15750 6798 15802
rect 6798 15750 6810 15802
rect 6810 15750 6840 15802
rect 6864 15750 6874 15802
rect 6874 15750 6920 15802
rect 6624 15748 6680 15750
rect 6704 15748 6760 15750
rect 6784 15748 6840 15750
rect 6864 15748 6920 15750
rect 4306 15280 4362 15336
rect 5888 15258 5944 15260
rect 5968 15258 6024 15260
rect 6048 15258 6104 15260
rect 6128 15258 6184 15260
rect 5888 15206 5934 15258
rect 5934 15206 5944 15258
rect 5968 15206 5998 15258
rect 5998 15206 6010 15258
rect 6010 15206 6024 15258
rect 6048 15206 6062 15258
rect 6062 15206 6074 15258
rect 6074 15206 6104 15258
rect 6128 15206 6138 15258
rect 6138 15206 6184 15258
rect 5888 15204 5944 15206
rect 5968 15204 6024 15206
rect 6048 15204 6104 15206
rect 6128 15204 6184 15206
rect 5686 15008 5742 15064
rect 6624 14714 6680 14716
rect 6704 14714 6760 14716
rect 6784 14714 6840 14716
rect 6864 14714 6920 14716
rect 6624 14662 6670 14714
rect 6670 14662 6680 14714
rect 6704 14662 6734 14714
rect 6734 14662 6746 14714
rect 6746 14662 6760 14714
rect 6784 14662 6798 14714
rect 6798 14662 6810 14714
rect 6810 14662 6840 14714
rect 6864 14662 6874 14714
rect 6874 14662 6920 14714
rect 6624 14660 6680 14662
rect 6704 14660 6760 14662
rect 6784 14660 6840 14662
rect 6864 14660 6920 14662
rect 5888 14170 5944 14172
rect 5968 14170 6024 14172
rect 6048 14170 6104 14172
rect 6128 14170 6184 14172
rect 5888 14118 5934 14170
rect 5934 14118 5944 14170
rect 5968 14118 5998 14170
rect 5998 14118 6010 14170
rect 6010 14118 6024 14170
rect 6048 14118 6062 14170
rect 6062 14118 6074 14170
rect 6074 14118 6104 14170
rect 6128 14118 6138 14170
rect 6138 14118 6184 14170
rect 5888 14116 5944 14118
rect 5968 14116 6024 14118
rect 6048 14116 6104 14118
rect 6128 14116 6184 14118
rect 6624 13626 6680 13628
rect 6704 13626 6760 13628
rect 6784 13626 6840 13628
rect 6864 13626 6920 13628
rect 6624 13574 6670 13626
rect 6670 13574 6680 13626
rect 6704 13574 6734 13626
rect 6734 13574 6746 13626
rect 6746 13574 6760 13626
rect 6784 13574 6798 13626
rect 6798 13574 6810 13626
rect 6810 13574 6840 13626
rect 6864 13574 6874 13626
rect 6874 13574 6920 13626
rect 6624 13572 6680 13574
rect 6704 13572 6760 13574
rect 6784 13572 6840 13574
rect 6864 13572 6920 13574
rect 46074 48328 46130 48384
rect 45982 14124 46038 14180
rect 5888 13082 5944 13084
rect 5968 13082 6024 13084
rect 6048 13082 6104 13084
rect 6128 13082 6184 13084
rect 5888 13030 5934 13082
rect 5934 13030 5944 13082
rect 5968 13030 5998 13082
rect 5998 13030 6010 13082
rect 6010 13030 6024 13082
rect 6048 13030 6062 13082
rect 6062 13030 6074 13082
rect 6074 13030 6104 13082
rect 6128 13030 6138 13082
rect 6138 13030 6184 13082
rect 5888 13028 5944 13030
rect 5968 13028 6024 13030
rect 6048 13028 6104 13030
rect 6128 13028 6184 13030
rect 45890 13036 45946 13092
rect 6624 12538 6680 12540
rect 6704 12538 6760 12540
rect 6784 12538 6840 12540
rect 6864 12538 6920 12540
rect 6624 12486 6670 12538
rect 6670 12486 6680 12538
rect 6704 12486 6734 12538
rect 6734 12486 6746 12538
rect 6746 12486 6760 12538
rect 6784 12486 6798 12538
rect 6798 12486 6810 12538
rect 6810 12486 6840 12538
rect 6864 12486 6874 12538
rect 6874 12486 6920 12538
rect 6624 12484 6680 12486
rect 6704 12484 6760 12486
rect 6784 12484 6840 12486
rect 6864 12484 6920 12486
rect 5888 11994 5944 11996
rect 5968 11994 6024 11996
rect 6048 11994 6104 11996
rect 6128 11994 6184 11996
rect 5888 11942 5934 11994
rect 5934 11942 5944 11994
rect 5968 11942 5998 11994
rect 5998 11942 6010 11994
rect 6010 11942 6024 11994
rect 6048 11942 6062 11994
rect 6062 11942 6074 11994
rect 6074 11942 6104 11994
rect 6128 11942 6138 11994
rect 6138 11942 6184 11994
rect 5888 11940 5944 11942
rect 5968 11940 6024 11942
rect 6048 11940 6104 11942
rect 6128 11940 6184 11942
rect 6624 11450 6680 11452
rect 6704 11450 6760 11452
rect 6784 11450 6840 11452
rect 6864 11450 6920 11452
rect 6624 11398 6670 11450
rect 6670 11398 6680 11450
rect 6704 11398 6734 11450
rect 6734 11398 6746 11450
rect 6746 11398 6760 11450
rect 6784 11398 6798 11450
rect 6798 11398 6810 11450
rect 6810 11398 6840 11450
rect 6864 11398 6874 11450
rect 6874 11398 6920 11450
rect 6624 11396 6680 11398
rect 6704 11396 6760 11398
rect 6784 11396 6840 11398
rect 6864 11396 6920 11398
rect 5888 10906 5944 10908
rect 5968 10906 6024 10908
rect 6048 10906 6104 10908
rect 6128 10906 6184 10908
rect 5888 10854 5934 10906
rect 5934 10854 5944 10906
rect 5968 10854 5998 10906
rect 5998 10854 6010 10906
rect 6010 10854 6024 10906
rect 6048 10854 6062 10906
rect 6062 10854 6074 10906
rect 6074 10854 6104 10906
rect 6128 10854 6138 10906
rect 6138 10854 6184 10906
rect 5888 10852 5944 10854
rect 5968 10852 6024 10854
rect 6048 10852 6104 10854
rect 6128 10852 6184 10854
rect 6624 10362 6680 10364
rect 6704 10362 6760 10364
rect 6784 10362 6840 10364
rect 6864 10362 6920 10364
rect 6624 10310 6670 10362
rect 6670 10310 6680 10362
rect 6704 10310 6734 10362
rect 6734 10310 6746 10362
rect 6746 10310 6760 10362
rect 6784 10310 6798 10362
rect 6798 10310 6810 10362
rect 6810 10310 6840 10362
rect 6864 10310 6874 10362
rect 6874 10310 6920 10362
rect 6624 10308 6680 10310
rect 6704 10308 6760 10310
rect 6784 10308 6840 10310
rect 6864 10308 6920 10310
rect 5888 9818 5944 9820
rect 5968 9818 6024 9820
rect 6048 9818 6104 9820
rect 6128 9818 6184 9820
rect 5888 9766 5934 9818
rect 5934 9766 5944 9818
rect 5968 9766 5998 9818
rect 5998 9766 6010 9818
rect 6010 9766 6024 9818
rect 6048 9766 6062 9818
rect 6062 9766 6074 9818
rect 6074 9766 6104 9818
rect 6128 9766 6138 9818
rect 6138 9766 6184 9818
rect 5888 9764 5944 9766
rect 5968 9764 6024 9766
rect 6048 9764 6104 9766
rect 6128 9764 6184 9766
rect 6624 9274 6680 9276
rect 6704 9274 6760 9276
rect 6784 9274 6840 9276
rect 6864 9274 6920 9276
rect 6624 9222 6670 9274
rect 6670 9222 6680 9274
rect 6704 9222 6734 9274
rect 6734 9222 6746 9274
rect 6746 9222 6760 9274
rect 6784 9222 6798 9274
rect 6798 9222 6810 9274
rect 6810 9222 6840 9274
rect 6864 9222 6874 9274
rect 6874 9222 6920 9274
rect 6624 9220 6680 9222
rect 6704 9220 6760 9222
rect 6784 9220 6840 9222
rect 6864 9220 6920 9222
rect 5888 8730 5944 8732
rect 5968 8730 6024 8732
rect 6048 8730 6104 8732
rect 6128 8730 6184 8732
rect 5888 8678 5934 8730
rect 5934 8678 5944 8730
rect 5968 8678 5998 8730
rect 5998 8678 6010 8730
rect 6010 8678 6024 8730
rect 6048 8678 6062 8730
rect 6062 8678 6074 8730
rect 6074 8678 6104 8730
rect 6128 8678 6138 8730
rect 6138 8678 6184 8730
rect 5888 8676 5944 8678
rect 5968 8676 6024 8678
rect 6048 8676 6104 8678
rect 6128 8676 6184 8678
rect 6624 8186 6680 8188
rect 6704 8186 6760 8188
rect 6784 8186 6840 8188
rect 6864 8186 6920 8188
rect 6624 8134 6670 8186
rect 6670 8134 6680 8186
rect 6704 8134 6734 8186
rect 6734 8134 6746 8186
rect 6746 8134 6760 8186
rect 6784 8134 6798 8186
rect 6798 8134 6810 8186
rect 6810 8134 6840 8186
rect 6864 8134 6874 8186
rect 6874 8134 6920 8186
rect 6624 8132 6680 8134
rect 6704 8132 6760 8134
rect 6784 8132 6840 8134
rect 6864 8132 6920 8134
rect 5888 7642 5944 7644
rect 5968 7642 6024 7644
rect 6048 7642 6104 7644
rect 6128 7642 6184 7644
rect 5888 7590 5934 7642
rect 5934 7590 5944 7642
rect 5968 7590 5998 7642
rect 5998 7590 6010 7642
rect 6010 7590 6024 7642
rect 6048 7590 6062 7642
rect 6062 7590 6074 7642
rect 6074 7590 6104 7642
rect 6128 7590 6138 7642
rect 6138 7590 6184 7642
rect 5888 7588 5944 7590
rect 5968 7588 6024 7590
rect 6048 7588 6104 7590
rect 6128 7588 6184 7590
rect 6624 7098 6680 7100
rect 6704 7098 6760 7100
rect 6784 7098 6840 7100
rect 6864 7098 6920 7100
rect 6624 7046 6670 7098
rect 6670 7046 6680 7098
rect 6704 7046 6734 7098
rect 6734 7046 6746 7098
rect 6746 7046 6760 7098
rect 6784 7046 6798 7098
rect 6798 7046 6810 7098
rect 6810 7046 6840 7098
rect 6864 7046 6874 7098
rect 6874 7046 6920 7098
rect 6624 7044 6680 7046
rect 6704 7044 6760 7046
rect 6784 7044 6840 7046
rect 6864 7044 6920 7046
rect 17728 7642 17784 7644
rect 17808 7642 17864 7644
rect 17888 7642 17944 7644
rect 17968 7642 18024 7644
rect 17728 7590 17774 7642
rect 17774 7590 17784 7642
rect 17808 7590 17838 7642
rect 17838 7590 17850 7642
rect 17850 7590 17864 7642
rect 17888 7590 17902 7642
rect 17902 7590 17914 7642
rect 17914 7590 17944 7642
rect 17968 7590 17978 7642
rect 17978 7590 18024 7642
rect 17728 7588 17784 7590
rect 17808 7588 17864 7590
rect 17888 7588 17944 7590
rect 17968 7588 18024 7590
rect 17728 6554 17784 6556
rect 17808 6554 17864 6556
rect 17888 6554 17944 6556
rect 17968 6554 18024 6556
rect 17728 6502 17774 6554
rect 17774 6502 17784 6554
rect 17808 6502 17838 6554
rect 17838 6502 17850 6554
rect 17850 6502 17864 6554
rect 17888 6502 17902 6554
rect 17902 6502 17914 6554
rect 17914 6502 17944 6554
rect 17968 6502 17978 6554
rect 17978 6502 18024 6554
rect 17728 6500 17784 6502
rect 17808 6500 17864 6502
rect 17888 6500 17944 6502
rect 17968 6500 18024 6502
rect 17728 5466 17784 5468
rect 17808 5466 17864 5468
rect 17888 5466 17944 5468
rect 17968 5466 18024 5468
rect 17728 5414 17774 5466
rect 17774 5414 17784 5466
rect 17808 5414 17838 5466
rect 17838 5414 17850 5466
rect 17850 5414 17864 5466
rect 17888 5414 17902 5466
rect 17902 5414 17914 5466
rect 17914 5414 17944 5466
rect 17968 5414 17978 5466
rect 17978 5414 18024 5466
rect 17728 5412 17784 5414
rect 17808 5412 17864 5414
rect 17888 5412 17944 5414
rect 17968 5412 18024 5414
rect 18388 7098 18444 7100
rect 18468 7098 18524 7100
rect 18548 7098 18604 7100
rect 18628 7098 18684 7100
rect 18388 7046 18434 7098
rect 18434 7046 18444 7098
rect 18468 7046 18498 7098
rect 18498 7046 18510 7098
rect 18510 7046 18524 7098
rect 18548 7046 18562 7098
rect 18562 7046 18574 7098
rect 18574 7046 18604 7098
rect 18628 7046 18638 7098
rect 18638 7046 18684 7098
rect 18388 7044 18444 7046
rect 18468 7044 18524 7046
rect 18548 7044 18604 7046
rect 18628 7044 18684 7046
rect 18388 6010 18444 6012
rect 18468 6010 18524 6012
rect 18548 6010 18604 6012
rect 18628 6010 18684 6012
rect 18388 5958 18434 6010
rect 18434 5958 18444 6010
rect 18468 5958 18498 6010
rect 18498 5958 18510 6010
rect 18510 5958 18524 6010
rect 18548 5958 18562 6010
rect 18562 5958 18574 6010
rect 18574 5958 18604 6010
rect 18628 5958 18638 6010
rect 18638 5958 18684 6010
rect 18388 5956 18444 5958
rect 18468 5956 18524 5958
rect 18548 5956 18604 5958
rect 18628 5956 18684 5958
rect 36128 7642 36184 7644
rect 36208 7642 36264 7644
rect 36288 7642 36344 7644
rect 36368 7642 36424 7644
rect 36128 7590 36174 7642
rect 36174 7590 36184 7642
rect 36208 7590 36238 7642
rect 36238 7590 36250 7642
rect 36250 7590 36264 7642
rect 36288 7590 36302 7642
rect 36302 7590 36314 7642
rect 36314 7590 36344 7642
rect 36368 7590 36378 7642
rect 36378 7590 36424 7642
rect 36128 7588 36184 7590
rect 36208 7588 36264 7590
rect 36288 7588 36344 7590
rect 36368 7588 36424 7590
rect 36788 7098 36844 7100
rect 36868 7098 36924 7100
rect 36948 7098 37004 7100
rect 37028 7098 37084 7100
rect 36788 7046 36834 7098
rect 36834 7046 36844 7098
rect 36868 7046 36898 7098
rect 36898 7046 36910 7098
rect 36910 7046 36924 7098
rect 36948 7046 36962 7098
rect 36962 7046 36974 7098
rect 36974 7046 37004 7098
rect 37028 7046 37038 7098
rect 37038 7046 37084 7098
rect 36788 7044 36844 7046
rect 36868 7044 36924 7046
rect 36948 7044 37004 7046
rect 37028 7044 37084 7046
rect 36128 6554 36184 6556
rect 36208 6554 36264 6556
rect 36288 6554 36344 6556
rect 36368 6554 36424 6556
rect 36128 6502 36174 6554
rect 36174 6502 36184 6554
rect 36208 6502 36238 6554
rect 36238 6502 36250 6554
rect 36250 6502 36264 6554
rect 36288 6502 36302 6554
rect 36302 6502 36314 6554
rect 36314 6502 36344 6554
rect 36368 6502 36378 6554
rect 36378 6502 36424 6554
rect 36128 6500 36184 6502
rect 36208 6500 36264 6502
rect 36288 6500 36344 6502
rect 36368 6500 36424 6502
rect 36788 6010 36844 6012
rect 36868 6010 36924 6012
rect 36948 6010 37004 6012
rect 37028 6010 37084 6012
rect 36788 5958 36834 6010
rect 36834 5958 36844 6010
rect 36868 5958 36898 6010
rect 36898 5958 36910 6010
rect 36910 5958 36924 6010
rect 36948 5958 36962 6010
rect 36962 5958 36974 6010
rect 36974 5958 37004 6010
rect 37028 5958 37038 6010
rect 37038 5958 37084 6010
rect 36788 5956 36844 5958
rect 36868 5956 36924 5958
rect 36948 5956 37004 5958
rect 37028 5956 37084 5958
rect 36128 5466 36184 5468
rect 36208 5466 36264 5468
rect 36288 5466 36344 5468
rect 36368 5466 36424 5468
rect 36128 5414 36174 5466
rect 36174 5414 36184 5466
rect 36208 5414 36238 5466
rect 36238 5414 36250 5466
rect 36250 5414 36264 5466
rect 36288 5414 36302 5466
rect 36302 5414 36314 5466
rect 36314 5414 36344 5466
rect 36368 5414 36378 5466
rect 36378 5414 36424 5466
rect 36128 5412 36184 5414
rect 36208 5412 36264 5414
rect 36288 5412 36344 5414
rect 36368 5412 36424 5414
rect 45430 10112 45486 10168
rect 46166 47240 46222 47296
rect 54528 87066 54584 87068
rect 54608 87066 54664 87068
rect 54688 87066 54744 87068
rect 54768 87066 54824 87068
rect 54528 87014 54574 87066
rect 54574 87014 54584 87066
rect 54608 87014 54638 87066
rect 54638 87014 54650 87066
rect 54650 87014 54664 87066
rect 54688 87014 54702 87066
rect 54702 87014 54714 87066
rect 54714 87014 54744 87066
rect 54768 87014 54778 87066
rect 54778 87014 54824 87066
rect 54528 87012 54584 87014
rect 54608 87012 54664 87014
rect 54688 87012 54744 87014
rect 54768 87012 54824 87014
rect 55188 86522 55244 86524
rect 55268 86522 55324 86524
rect 55348 86522 55404 86524
rect 55428 86522 55484 86524
rect 55188 86470 55234 86522
rect 55234 86470 55244 86522
rect 55268 86470 55298 86522
rect 55298 86470 55310 86522
rect 55310 86470 55324 86522
rect 55348 86470 55362 86522
rect 55362 86470 55374 86522
rect 55374 86470 55404 86522
rect 55428 86470 55438 86522
rect 55438 86470 55484 86522
rect 55188 86468 55244 86470
rect 55268 86468 55324 86470
rect 55348 86468 55404 86470
rect 55428 86468 55484 86470
rect 54528 85978 54584 85980
rect 54608 85978 54664 85980
rect 54688 85978 54744 85980
rect 54768 85978 54824 85980
rect 54528 85926 54574 85978
rect 54574 85926 54584 85978
rect 54608 85926 54638 85978
rect 54638 85926 54650 85978
rect 54650 85926 54664 85978
rect 54688 85926 54702 85978
rect 54702 85926 54714 85978
rect 54714 85926 54744 85978
rect 54768 85926 54778 85978
rect 54778 85926 54824 85978
rect 54528 85924 54584 85926
rect 54608 85924 54664 85926
rect 54688 85924 54744 85926
rect 54768 85924 54824 85926
rect 55188 85434 55244 85436
rect 55268 85434 55324 85436
rect 55348 85434 55404 85436
rect 55428 85434 55484 85436
rect 55188 85382 55234 85434
rect 55234 85382 55244 85434
rect 55268 85382 55298 85434
rect 55298 85382 55310 85434
rect 55310 85382 55324 85434
rect 55348 85382 55362 85434
rect 55362 85382 55374 85434
rect 55374 85382 55404 85434
rect 55428 85382 55438 85434
rect 55438 85382 55484 85434
rect 55188 85380 55244 85382
rect 55268 85380 55324 85382
rect 55348 85380 55404 85382
rect 55428 85380 55484 85382
rect 54528 84890 54584 84892
rect 54608 84890 54664 84892
rect 54688 84890 54744 84892
rect 54768 84890 54824 84892
rect 54528 84838 54574 84890
rect 54574 84838 54584 84890
rect 54608 84838 54638 84890
rect 54638 84838 54650 84890
rect 54650 84838 54664 84890
rect 54688 84838 54702 84890
rect 54702 84838 54714 84890
rect 54714 84838 54744 84890
rect 54768 84838 54778 84890
rect 54778 84838 54824 84890
rect 54528 84836 54584 84838
rect 54608 84836 54664 84838
rect 54688 84836 54744 84838
rect 54768 84836 54824 84838
rect 55188 84346 55244 84348
rect 55268 84346 55324 84348
rect 55348 84346 55404 84348
rect 55428 84346 55484 84348
rect 55188 84294 55234 84346
rect 55234 84294 55244 84346
rect 55268 84294 55298 84346
rect 55298 84294 55310 84346
rect 55310 84294 55324 84346
rect 55348 84294 55362 84346
rect 55362 84294 55374 84346
rect 55374 84294 55404 84346
rect 55428 84294 55438 84346
rect 55438 84294 55484 84346
rect 55188 84292 55244 84294
rect 55268 84292 55324 84294
rect 55348 84292 55404 84294
rect 55428 84292 55484 84294
rect 73588 87610 73644 87612
rect 73668 87610 73724 87612
rect 73748 87610 73804 87612
rect 73828 87610 73884 87612
rect 73588 87558 73634 87610
rect 73634 87558 73644 87610
rect 73668 87558 73698 87610
rect 73698 87558 73710 87610
rect 73710 87558 73724 87610
rect 73748 87558 73762 87610
rect 73762 87558 73774 87610
rect 73774 87558 73804 87610
rect 73828 87558 73838 87610
rect 73838 87558 73884 87610
rect 73588 87556 73644 87558
rect 73668 87556 73724 87558
rect 73748 87556 73804 87558
rect 73828 87556 73884 87558
rect 72928 87066 72984 87068
rect 73008 87066 73064 87068
rect 73088 87066 73144 87068
rect 73168 87066 73224 87068
rect 72928 87014 72974 87066
rect 72974 87014 72984 87066
rect 73008 87014 73038 87066
rect 73038 87014 73050 87066
rect 73050 87014 73064 87066
rect 73088 87014 73102 87066
rect 73102 87014 73114 87066
rect 73114 87014 73144 87066
rect 73168 87014 73178 87066
rect 73178 87014 73224 87066
rect 72928 87012 72984 87014
rect 73008 87012 73064 87014
rect 73088 87012 73144 87014
rect 73168 87012 73224 87014
rect 72928 85978 72984 85980
rect 73008 85978 73064 85980
rect 73088 85978 73144 85980
rect 73168 85978 73224 85980
rect 72928 85926 72974 85978
rect 72974 85926 72984 85978
rect 73008 85926 73038 85978
rect 73038 85926 73050 85978
rect 73050 85926 73064 85978
rect 73088 85926 73102 85978
rect 73102 85926 73114 85978
rect 73114 85926 73144 85978
rect 73168 85926 73178 85978
rect 73178 85926 73224 85978
rect 72928 85924 72984 85926
rect 73008 85924 73064 85926
rect 73088 85924 73144 85926
rect 73168 85924 73224 85926
rect 72928 84890 72984 84892
rect 73008 84890 73064 84892
rect 73088 84890 73144 84892
rect 73168 84890 73224 84892
rect 72928 84838 72974 84890
rect 72974 84838 72984 84890
rect 73008 84838 73038 84890
rect 73038 84838 73050 84890
rect 73050 84838 73064 84890
rect 73088 84838 73102 84890
rect 73102 84838 73114 84890
rect 73114 84838 73144 84890
rect 73168 84838 73178 84890
rect 73178 84838 73224 84890
rect 72928 84836 72984 84838
rect 73008 84836 73064 84838
rect 73088 84836 73144 84838
rect 73168 84836 73224 84838
rect 73588 86522 73644 86524
rect 73668 86522 73724 86524
rect 73748 86522 73804 86524
rect 73828 86522 73884 86524
rect 73588 86470 73634 86522
rect 73634 86470 73644 86522
rect 73668 86470 73698 86522
rect 73698 86470 73710 86522
rect 73710 86470 73724 86522
rect 73748 86470 73762 86522
rect 73762 86470 73774 86522
rect 73774 86470 73804 86522
rect 73828 86470 73838 86522
rect 73838 86470 73884 86522
rect 73588 86468 73644 86470
rect 73668 86468 73724 86470
rect 73748 86468 73804 86470
rect 73828 86468 73884 86470
rect 73588 85434 73644 85436
rect 73668 85434 73724 85436
rect 73748 85434 73804 85436
rect 73828 85434 73884 85436
rect 73588 85382 73634 85434
rect 73634 85382 73644 85434
rect 73668 85382 73698 85434
rect 73698 85382 73710 85434
rect 73710 85382 73724 85434
rect 73748 85382 73762 85434
rect 73762 85382 73774 85434
rect 73774 85382 73804 85434
rect 73828 85382 73838 85434
rect 73838 85382 73884 85434
rect 73588 85380 73644 85382
rect 73668 85380 73724 85382
rect 73748 85380 73804 85382
rect 73828 85380 73884 85382
rect 73588 84346 73644 84348
rect 73668 84346 73724 84348
rect 73748 84346 73804 84348
rect 73828 84346 73884 84348
rect 73588 84294 73634 84346
rect 73634 84294 73644 84346
rect 73668 84294 73698 84346
rect 73698 84294 73710 84346
rect 73710 84294 73724 84346
rect 73748 84294 73762 84346
rect 73762 84294 73774 84346
rect 73774 84294 73804 84346
rect 73828 84294 73838 84346
rect 73838 84294 73884 84346
rect 73588 84292 73644 84294
rect 73668 84292 73724 84294
rect 73748 84292 73804 84294
rect 73828 84292 73884 84294
rect 86480 84890 86536 84892
rect 86560 84890 86616 84892
rect 86640 84890 86696 84892
rect 86720 84890 86776 84892
rect 86480 84838 86526 84890
rect 86526 84838 86536 84890
rect 86560 84838 86590 84890
rect 86590 84838 86602 84890
rect 86602 84838 86616 84890
rect 86640 84838 86654 84890
rect 86654 84838 86666 84890
rect 86666 84838 86696 84890
rect 86720 84838 86730 84890
rect 86730 84838 86776 84890
rect 86480 84836 86536 84838
rect 86560 84836 86616 84838
rect 86640 84836 86696 84838
rect 86720 84836 86776 84838
rect 87216 84346 87272 84348
rect 87296 84346 87352 84348
rect 87376 84346 87432 84348
rect 87456 84346 87512 84348
rect 87216 84294 87262 84346
rect 87262 84294 87272 84346
rect 87296 84294 87326 84346
rect 87326 84294 87338 84346
rect 87338 84294 87352 84346
rect 87376 84294 87390 84346
rect 87390 84294 87402 84346
rect 87402 84294 87432 84346
rect 87456 84294 87466 84346
rect 87466 84294 87512 84346
rect 87216 84292 87272 84294
rect 87296 84292 87352 84294
rect 87376 84292 87432 84294
rect 87456 84292 87512 84294
rect 86480 83802 86536 83804
rect 86560 83802 86616 83804
rect 86640 83802 86696 83804
rect 86720 83802 86776 83804
rect 86480 83750 86526 83802
rect 86526 83750 86536 83802
rect 86560 83750 86590 83802
rect 86590 83750 86602 83802
rect 86602 83750 86616 83802
rect 86640 83750 86654 83802
rect 86654 83750 86666 83802
rect 86666 83750 86696 83802
rect 86720 83750 86730 83802
rect 86730 83750 86776 83802
rect 86480 83748 86536 83750
rect 86560 83748 86616 83750
rect 86640 83748 86696 83750
rect 86720 83748 86776 83750
rect 87216 83258 87272 83260
rect 87296 83258 87352 83260
rect 87376 83258 87432 83260
rect 87456 83258 87512 83260
rect 87216 83206 87262 83258
rect 87262 83206 87272 83258
rect 87296 83206 87326 83258
rect 87326 83206 87338 83258
rect 87338 83206 87352 83258
rect 87376 83206 87390 83258
rect 87390 83206 87402 83258
rect 87402 83206 87432 83258
rect 87456 83206 87466 83258
rect 87466 83206 87512 83258
rect 87216 83204 87272 83206
rect 87296 83204 87352 83206
rect 87376 83204 87432 83206
rect 87456 83204 87512 83206
rect 47086 81648 47142 81704
rect 47960 81648 48016 81704
rect 46074 11948 46130 12004
rect 49064 45880 49120 45936
rect 51134 45916 51136 45936
rect 51136 45916 51188 45936
rect 51188 45916 51190 45936
rect 51134 45880 51190 45916
rect 47086 45608 47142 45664
rect 47960 45608 48016 45664
rect 86480 82714 86536 82716
rect 86560 82714 86616 82716
rect 86640 82714 86696 82716
rect 86720 82714 86776 82716
rect 86480 82662 86526 82714
rect 86526 82662 86536 82714
rect 86560 82662 86590 82714
rect 86590 82662 86602 82714
rect 86602 82662 86616 82714
rect 86640 82662 86654 82714
rect 86654 82662 86666 82714
rect 86666 82662 86696 82714
rect 86720 82662 86730 82714
rect 86730 82662 86776 82714
rect 86480 82660 86536 82662
rect 86560 82660 86616 82662
rect 86640 82660 86696 82662
rect 86720 82660 86776 82662
rect 87216 82170 87272 82172
rect 87296 82170 87352 82172
rect 87376 82170 87432 82172
rect 87456 82170 87512 82172
rect 87216 82118 87262 82170
rect 87262 82118 87272 82170
rect 87296 82118 87326 82170
rect 87326 82118 87338 82170
rect 87338 82118 87352 82170
rect 87376 82118 87390 82170
rect 87390 82118 87402 82170
rect 87402 82118 87432 82170
rect 87456 82118 87466 82170
rect 87466 82118 87512 82170
rect 87216 82116 87272 82118
rect 87296 82116 87352 82118
rect 87376 82116 87432 82118
rect 87456 82116 87512 82118
rect 86480 81626 86536 81628
rect 86560 81626 86616 81628
rect 86640 81626 86696 81628
rect 86720 81626 86776 81628
rect 86480 81574 86526 81626
rect 86526 81574 86536 81626
rect 86560 81574 86590 81626
rect 86590 81574 86602 81626
rect 86602 81574 86616 81626
rect 86640 81574 86654 81626
rect 86654 81574 86666 81626
rect 86666 81574 86696 81626
rect 86720 81574 86730 81626
rect 86730 81574 86776 81626
rect 86480 81572 86536 81574
rect 86560 81572 86616 81574
rect 86640 81572 86696 81574
rect 86720 81572 86776 81574
rect 88210 81276 88212 81296
rect 88212 81276 88264 81296
rect 88264 81276 88266 81296
rect 88210 81240 88266 81276
rect 87216 81082 87272 81084
rect 87296 81082 87352 81084
rect 87376 81082 87432 81084
rect 87456 81082 87512 81084
rect 84346 80968 84402 81024
rect 87216 81030 87262 81082
rect 87262 81030 87272 81082
rect 87296 81030 87326 81082
rect 87326 81030 87338 81082
rect 87338 81030 87352 81082
rect 87376 81030 87390 81082
rect 87390 81030 87402 81082
rect 87402 81030 87432 81082
rect 87456 81030 87466 81082
rect 87466 81030 87512 81082
rect 87216 81028 87272 81030
rect 87296 81028 87352 81030
rect 87376 81028 87432 81030
rect 87456 81028 87512 81030
rect 86480 80538 86536 80540
rect 86560 80538 86616 80540
rect 86640 80538 86696 80540
rect 86720 80538 86776 80540
rect 86480 80486 86526 80538
rect 86526 80486 86536 80538
rect 86560 80486 86590 80538
rect 86590 80486 86602 80538
rect 86602 80486 86616 80538
rect 86640 80486 86654 80538
rect 86654 80486 86666 80538
rect 86666 80486 86696 80538
rect 86720 80486 86730 80538
rect 86730 80486 86776 80538
rect 86480 80484 86536 80486
rect 86560 80484 86616 80486
rect 86640 80484 86696 80486
rect 86720 80484 86776 80486
rect 87216 79994 87272 79996
rect 87296 79994 87352 79996
rect 87376 79994 87432 79996
rect 87456 79994 87512 79996
rect 85818 79880 85874 79936
rect 87216 79942 87262 79994
rect 87262 79942 87272 79994
rect 87296 79942 87326 79994
rect 87326 79942 87338 79994
rect 87338 79942 87352 79994
rect 87376 79942 87390 79994
rect 87390 79942 87402 79994
rect 87402 79942 87432 79994
rect 87456 79942 87466 79994
rect 87466 79942 87512 79994
rect 87216 79940 87272 79942
rect 87296 79940 87352 79942
rect 87376 79940 87432 79942
rect 87456 79940 87512 79942
rect 88210 79880 88266 79936
rect 86480 79450 86536 79452
rect 86560 79450 86616 79452
rect 86640 79450 86696 79452
rect 86720 79450 86776 79452
rect 86480 79398 86526 79450
rect 86526 79398 86536 79450
rect 86560 79398 86590 79450
rect 86590 79398 86602 79450
rect 86602 79398 86616 79450
rect 86640 79398 86654 79450
rect 86654 79398 86666 79450
rect 86666 79398 86696 79450
rect 86720 79398 86730 79450
rect 86730 79398 86776 79450
rect 86480 79396 86536 79398
rect 86560 79396 86616 79398
rect 86640 79396 86696 79398
rect 86720 79396 86776 79398
rect 87216 78906 87272 78908
rect 87296 78906 87352 78908
rect 87376 78906 87432 78908
rect 87456 78906 87512 78908
rect 85818 78792 85874 78848
rect 87216 78854 87262 78906
rect 87262 78854 87272 78906
rect 87296 78854 87326 78906
rect 87326 78854 87338 78906
rect 87338 78854 87352 78906
rect 87376 78854 87390 78906
rect 87390 78854 87402 78906
rect 87402 78854 87432 78906
rect 87456 78854 87466 78906
rect 87466 78854 87512 78906
rect 87216 78852 87272 78854
rect 87296 78852 87352 78854
rect 87376 78852 87432 78854
rect 87456 78852 87512 78854
rect 88210 78520 88266 78576
rect 86480 78362 86536 78364
rect 86560 78362 86616 78364
rect 86640 78362 86696 78364
rect 86720 78362 86776 78364
rect 86480 78310 86526 78362
rect 86526 78310 86536 78362
rect 86560 78310 86590 78362
rect 86590 78310 86602 78362
rect 86602 78310 86616 78362
rect 86640 78310 86654 78362
rect 86654 78310 86666 78362
rect 86666 78310 86696 78362
rect 86720 78310 86730 78362
rect 86730 78310 86776 78362
rect 86480 78308 86536 78310
rect 86560 78308 86616 78310
rect 86640 78308 86696 78310
rect 86720 78308 86776 78310
rect 88210 77840 88266 77896
rect 87216 77818 87272 77820
rect 87296 77818 87352 77820
rect 87376 77818 87432 77820
rect 87456 77818 87512 77820
rect 85818 77704 85874 77760
rect 87216 77766 87262 77818
rect 87262 77766 87272 77818
rect 87296 77766 87326 77818
rect 87326 77766 87338 77818
rect 87338 77766 87352 77818
rect 87376 77766 87390 77818
rect 87390 77766 87402 77818
rect 87402 77766 87432 77818
rect 87456 77766 87466 77818
rect 87466 77766 87512 77818
rect 87216 77764 87272 77766
rect 87296 77764 87352 77766
rect 87376 77764 87432 77766
rect 87456 77764 87512 77766
rect 86480 77274 86536 77276
rect 86560 77274 86616 77276
rect 86640 77274 86696 77276
rect 86720 77274 86776 77276
rect 86480 77222 86526 77274
rect 86526 77222 86536 77274
rect 86560 77222 86590 77274
rect 86590 77222 86602 77274
rect 86602 77222 86616 77274
rect 86640 77222 86654 77274
rect 86654 77222 86666 77274
rect 86666 77222 86696 77274
rect 86720 77222 86730 77274
rect 86730 77222 86776 77274
rect 86480 77220 86536 77222
rect 86560 77220 86616 77222
rect 86640 77220 86696 77222
rect 86720 77220 86776 77222
rect 87216 76730 87272 76732
rect 87296 76730 87352 76732
rect 87376 76730 87432 76732
rect 87456 76730 87512 76732
rect 85818 76616 85874 76672
rect 87216 76678 87262 76730
rect 87262 76678 87272 76730
rect 87296 76678 87326 76730
rect 87326 76678 87338 76730
rect 87338 76678 87352 76730
rect 87376 76678 87390 76730
rect 87390 76678 87402 76730
rect 87402 76678 87432 76730
rect 87456 76678 87466 76730
rect 87466 76678 87512 76730
rect 87216 76676 87272 76678
rect 87296 76676 87352 76678
rect 87376 76676 87432 76678
rect 87456 76676 87512 76678
rect 88026 76480 88082 76536
rect 86480 76186 86536 76188
rect 86560 76186 86616 76188
rect 86640 76186 86696 76188
rect 86720 76186 86776 76188
rect 86480 76134 86526 76186
rect 86526 76134 86536 76186
rect 86560 76134 86590 76186
rect 86590 76134 86602 76186
rect 86602 76134 86616 76186
rect 86640 76134 86654 76186
rect 86654 76134 86666 76186
rect 86666 76134 86696 76186
rect 86720 76134 86730 76186
rect 86730 76134 86776 76186
rect 86480 76132 86536 76134
rect 86560 76132 86616 76134
rect 86640 76132 86696 76134
rect 86720 76132 86776 76134
rect 88210 75836 88212 75856
rect 88212 75836 88264 75856
rect 88264 75836 88266 75856
rect 88210 75800 88266 75836
rect 87216 75642 87272 75644
rect 87296 75642 87352 75644
rect 87376 75642 87432 75644
rect 87456 75642 87512 75644
rect 85818 75528 85874 75584
rect 87216 75590 87262 75642
rect 87262 75590 87272 75642
rect 87296 75590 87326 75642
rect 87326 75590 87338 75642
rect 87338 75590 87352 75642
rect 87376 75590 87390 75642
rect 87390 75590 87402 75642
rect 87402 75590 87432 75642
rect 87456 75590 87466 75642
rect 87466 75590 87512 75642
rect 87216 75588 87272 75590
rect 87296 75588 87352 75590
rect 87376 75588 87432 75590
rect 87456 75588 87512 75590
rect 86480 75098 86536 75100
rect 86560 75098 86616 75100
rect 86640 75098 86696 75100
rect 86720 75098 86776 75100
rect 86480 75046 86526 75098
rect 86526 75046 86536 75098
rect 86560 75046 86590 75098
rect 86590 75046 86602 75098
rect 86602 75046 86616 75098
rect 86640 75046 86654 75098
rect 86654 75046 86666 75098
rect 86666 75046 86696 75098
rect 86720 75046 86730 75098
rect 86730 75046 86776 75098
rect 86480 75044 86536 75046
rect 86560 75044 86616 75046
rect 86640 75044 86696 75046
rect 86720 75044 86776 75046
rect 87216 74554 87272 74556
rect 87296 74554 87352 74556
rect 87376 74554 87432 74556
rect 87456 74554 87512 74556
rect 84530 74440 84586 74496
rect 87216 74502 87262 74554
rect 87262 74502 87272 74554
rect 87296 74502 87326 74554
rect 87326 74502 87338 74554
rect 87338 74502 87352 74554
rect 87376 74502 87390 74554
rect 87390 74502 87402 74554
rect 87402 74502 87432 74554
rect 87456 74502 87466 74554
rect 87466 74502 87512 74554
rect 87216 74500 87272 74502
rect 87296 74500 87352 74502
rect 87376 74500 87432 74502
rect 87456 74500 87512 74502
rect 88578 74440 88634 74496
rect 86480 74010 86536 74012
rect 86560 74010 86616 74012
rect 86640 74010 86696 74012
rect 86720 74010 86776 74012
rect 86480 73958 86526 74010
rect 86526 73958 86536 74010
rect 86560 73958 86590 74010
rect 86590 73958 86602 74010
rect 86602 73958 86616 74010
rect 86640 73958 86654 74010
rect 86654 73958 86666 74010
rect 86666 73958 86696 74010
rect 86720 73958 86730 74010
rect 86730 73958 86776 74010
rect 86480 73956 86536 73958
rect 86560 73956 86616 73958
rect 86640 73956 86696 73958
rect 86720 73956 86776 73958
rect 87216 73466 87272 73468
rect 87296 73466 87352 73468
rect 87376 73466 87432 73468
rect 87456 73466 87512 73468
rect 84806 73352 84862 73408
rect 87216 73414 87262 73466
rect 87262 73414 87272 73466
rect 87296 73414 87326 73466
rect 87326 73414 87338 73466
rect 87338 73414 87352 73466
rect 87376 73414 87390 73466
rect 87390 73414 87402 73466
rect 87402 73414 87432 73466
rect 87456 73414 87466 73466
rect 87466 73414 87512 73466
rect 87216 73412 87272 73414
rect 87296 73412 87352 73414
rect 87376 73412 87432 73414
rect 87456 73412 87512 73414
rect 88210 73080 88266 73136
rect 86480 72922 86536 72924
rect 86560 72922 86616 72924
rect 86640 72922 86696 72924
rect 86720 72922 86776 72924
rect 86480 72870 86526 72922
rect 86526 72870 86536 72922
rect 86560 72870 86590 72922
rect 86590 72870 86602 72922
rect 86602 72870 86616 72922
rect 86640 72870 86654 72922
rect 86654 72870 86666 72922
rect 86666 72870 86696 72922
rect 86720 72870 86730 72922
rect 86730 72870 86776 72922
rect 86480 72868 86536 72870
rect 86560 72868 86616 72870
rect 86640 72868 86696 72870
rect 86720 72868 86776 72870
rect 87216 72378 87272 72380
rect 87296 72378 87352 72380
rect 87376 72378 87432 72380
rect 87456 72378 87512 72380
rect 87216 72326 87262 72378
rect 87262 72326 87272 72378
rect 87296 72326 87326 72378
rect 87326 72326 87338 72378
rect 87338 72326 87352 72378
rect 87376 72326 87390 72378
rect 87390 72326 87402 72378
rect 87402 72326 87432 72378
rect 87456 72326 87466 72378
rect 87466 72326 87512 72378
rect 87216 72324 87272 72326
rect 87296 72324 87352 72326
rect 87376 72324 87432 72326
rect 87456 72324 87512 72326
rect 88210 72400 88266 72456
rect 87842 72128 87898 72184
rect 86480 71834 86536 71836
rect 86560 71834 86616 71836
rect 86640 71834 86696 71836
rect 86720 71834 86776 71836
rect 86480 71782 86526 71834
rect 86526 71782 86536 71834
rect 86560 71782 86590 71834
rect 86590 71782 86602 71834
rect 86602 71782 86616 71834
rect 86640 71782 86654 71834
rect 86654 71782 86666 71834
rect 86666 71782 86696 71834
rect 86720 71782 86730 71834
rect 86730 71782 86776 71834
rect 86480 71780 86536 71782
rect 86560 71780 86616 71782
rect 86640 71780 86696 71782
rect 86720 71780 86776 71782
rect 87216 71290 87272 71292
rect 87296 71290 87352 71292
rect 87376 71290 87432 71292
rect 87456 71290 87512 71292
rect 85818 71176 85874 71232
rect 87216 71238 87262 71290
rect 87262 71238 87272 71290
rect 87296 71238 87326 71290
rect 87326 71238 87338 71290
rect 87338 71238 87352 71290
rect 87376 71238 87390 71290
rect 87390 71238 87402 71290
rect 87402 71238 87432 71290
rect 87456 71238 87466 71290
rect 87466 71238 87512 71290
rect 87216 71236 87272 71238
rect 87296 71236 87352 71238
rect 87376 71236 87432 71238
rect 87456 71236 87512 71238
rect 88210 71040 88266 71096
rect 86480 70746 86536 70748
rect 86560 70746 86616 70748
rect 86640 70746 86696 70748
rect 86720 70746 86776 70748
rect 86480 70694 86526 70746
rect 86526 70694 86536 70746
rect 86560 70694 86590 70746
rect 86590 70694 86602 70746
rect 86602 70694 86616 70746
rect 86640 70694 86654 70746
rect 86654 70694 86666 70746
rect 86666 70694 86696 70746
rect 86720 70694 86730 70746
rect 86730 70694 86776 70746
rect 86480 70692 86536 70694
rect 86560 70692 86616 70694
rect 86640 70692 86696 70694
rect 86720 70692 86776 70694
rect 88210 70396 88212 70416
rect 88212 70396 88264 70416
rect 88264 70396 88266 70416
rect 88210 70360 88266 70396
rect 87216 70202 87272 70204
rect 87296 70202 87352 70204
rect 87376 70202 87432 70204
rect 87456 70202 87512 70204
rect 85818 70088 85874 70144
rect 87216 70150 87262 70202
rect 87262 70150 87272 70202
rect 87296 70150 87326 70202
rect 87326 70150 87338 70202
rect 87338 70150 87352 70202
rect 87376 70150 87390 70202
rect 87390 70150 87402 70202
rect 87402 70150 87432 70202
rect 87456 70150 87466 70202
rect 87466 70150 87512 70202
rect 87216 70148 87272 70150
rect 87296 70148 87352 70150
rect 87376 70148 87432 70150
rect 87456 70148 87512 70150
rect 86480 69658 86536 69660
rect 86560 69658 86616 69660
rect 86640 69658 86696 69660
rect 86720 69658 86776 69660
rect 86480 69606 86526 69658
rect 86526 69606 86536 69658
rect 86560 69606 86590 69658
rect 86590 69606 86602 69658
rect 86602 69606 86616 69658
rect 86640 69606 86654 69658
rect 86654 69606 86666 69658
rect 86666 69606 86696 69658
rect 86720 69606 86730 69658
rect 86730 69606 86776 69658
rect 86480 69604 86536 69606
rect 86560 69604 86616 69606
rect 86640 69604 86696 69606
rect 86720 69604 86776 69606
rect 87216 69114 87272 69116
rect 87296 69114 87352 69116
rect 87376 69114 87432 69116
rect 87456 69114 87512 69116
rect 84806 69000 84862 69056
rect 87216 69062 87262 69114
rect 87262 69062 87272 69114
rect 87296 69062 87326 69114
rect 87326 69062 87338 69114
rect 87338 69062 87352 69114
rect 87376 69062 87390 69114
rect 87390 69062 87402 69114
rect 87402 69062 87432 69114
rect 87456 69062 87466 69114
rect 87466 69062 87512 69114
rect 87216 69060 87272 69062
rect 87296 69060 87352 69062
rect 87376 69060 87432 69062
rect 87456 69060 87512 69062
rect 88578 69000 88634 69056
rect 86480 68570 86536 68572
rect 86560 68570 86616 68572
rect 86640 68570 86696 68572
rect 86720 68570 86776 68572
rect 86480 68518 86526 68570
rect 86526 68518 86536 68570
rect 86560 68518 86590 68570
rect 86590 68518 86602 68570
rect 86602 68518 86616 68570
rect 86640 68518 86654 68570
rect 86654 68518 86666 68570
rect 86666 68518 86696 68570
rect 86720 68518 86730 68570
rect 86730 68518 86776 68570
rect 86480 68516 86536 68518
rect 86560 68516 86616 68518
rect 86640 68516 86696 68518
rect 86720 68516 86776 68518
rect 87216 68026 87272 68028
rect 87296 68026 87352 68028
rect 87376 68026 87432 68028
rect 87456 68026 87512 68028
rect 85266 67912 85322 67968
rect 87216 67974 87262 68026
rect 87262 67974 87272 68026
rect 87296 67974 87326 68026
rect 87326 67974 87338 68026
rect 87338 67974 87352 68026
rect 87376 67974 87390 68026
rect 87390 67974 87402 68026
rect 87402 67974 87432 68026
rect 87456 67974 87466 68026
rect 87466 67974 87512 68026
rect 87216 67972 87272 67974
rect 87296 67972 87352 67974
rect 87376 67972 87432 67974
rect 87456 67972 87512 67974
rect 88210 67640 88266 67696
rect 86480 67482 86536 67484
rect 86560 67482 86616 67484
rect 86640 67482 86696 67484
rect 86720 67482 86776 67484
rect 86480 67430 86526 67482
rect 86526 67430 86536 67482
rect 86560 67430 86590 67482
rect 86590 67430 86602 67482
rect 86602 67430 86616 67482
rect 86640 67430 86654 67482
rect 86654 67430 86666 67482
rect 86666 67430 86696 67482
rect 86720 67430 86730 67482
rect 86730 67430 86776 67482
rect 86480 67428 86536 67430
rect 86560 67428 86616 67430
rect 86640 67428 86696 67430
rect 86720 67428 86776 67430
rect 88210 66960 88266 67016
rect 87216 66938 87272 66940
rect 87296 66938 87352 66940
rect 87376 66938 87432 66940
rect 87456 66938 87512 66940
rect 85818 66824 85874 66880
rect 87216 66886 87262 66938
rect 87262 66886 87272 66938
rect 87296 66886 87326 66938
rect 87326 66886 87338 66938
rect 87338 66886 87352 66938
rect 87376 66886 87390 66938
rect 87390 66886 87402 66938
rect 87402 66886 87432 66938
rect 87456 66886 87466 66938
rect 87466 66886 87512 66938
rect 87216 66884 87272 66886
rect 87296 66884 87352 66886
rect 87376 66884 87432 66886
rect 87456 66884 87512 66886
rect 86480 66394 86536 66396
rect 86560 66394 86616 66396
rect 86640 66394 86696 66396
rect 86720 66394 86776 66396
rect 86480 66342 86526 66394
rect 86526 66342 86536 66394
rect 86560 66342 86590 66394
rect 86590 66342 86602 66394
rect 86602 66342 86616 66394
rect 86640 66342 86654 66394
rect 86654 66342 86666 66394
rect 86666 66342 86696 66394
rect 86720 66342 86730 66394
rect 86730 66342 86776 66394
rect 86480 66340 86536 66342
rect 86560 66340 86616 66342
rect 86640 66340 86696 66342
rect 86720 66340 86776 66342
rect 87216 65850 87272 65852
rect 87296 65850 87352 65852
rect 87376 65850 87432 65852
rect 87456 65850 87512 65852
rect 85818 65736 85874 65792
rect 87216 65798 87262 65850
rect 87262 65798 87272 65850
rect 87296 65798 87326 65850
rect 87326 65798 87338 65850
rect 87338 65798 87352 65850
rect 87376 65798 87390 65850
rect 87390 65798 87402 65850
rect 87402 65798 87432 65850
rect 87456 65798 87466 65850
rect 87466 65798 87512 65850
rect 87216 65796 87272 65798
rect 87296 65796 87352 65798
rect 87376 65796 87432 65798
rect 87456 65796 87512 65798
rect 88210 65600 88266 65656
rect 86480 65306 86536 65308
rect 86560 65306 86616 65308
rect 86640 65306 86696 65308
rect 86720 65306 86776 65308
rect 86480 65254 86526 65306
rect 86526 65254 86536 65306
rect 86560 65254 86590 65306
rect 86590 65254 86602 65306
rect 86602 65254 86616 65306
rect 86640 65254 86654 65306
rect 86654 65254 86666 65306
rect 86666 65254 86696 65306
rect 86720 65254 86730 65306
rect 86730 65254 86776 65306
rect 86480 65252 86536 65254
rect 86560 65252 86616 65254
rect 86640 65252 86696 65254
rect 86720 65252 86776 65254
rect 88394 64920 88450 64976
rect 87216 64762 87272 64764
rect 87296 64762 87352 64764
rect 87376 64762 87432 64764
rect 87456 64762 87512 64764
rect 85818 64648 85874 64704
rect 87216 64710 87262 64762
rect 87262 64710 87272 64762
rect 87296 64710 87326 64762
rect 87326 64710 87338 64762
rect 87338 64710 87352 64762
rect 87376 64710 87390 64762
rect 87390 64710 87402 64762
rect 87402 64710 87432 64762
rect 87456 64710 87466 64762
rect 87466 64710 87512 64762
rect 87216 64708 87272 64710
rect 87296 64708 87352 64710
rect 87376 64708 87432 64710
rect 87456 64708 87512 64710
rect 86480 64218 86536 64220
rect 86560 64218 86616 64220
rect 86640 64218 86696 64220
rect 86720 64218 86776 64220
rect 86480 64166 86526 64218
rect 86526 64166 86536 64218
rect 86560 64166 86590 64218
rect 86590 64166 86602 64218
rect 86602 64166 86616 64218
rect 86640 64166 86654 64218
rect 86654 64166 86666 64218
rect 86666 64166 86696 64218
rect 86720 64166 86730 64218
rect 86730 64166 86776 64218
rect 86480 64164 86536 64166
rect 86560 64164 86616 64166
rect 86640 64164 86696 64166
rect 86720 64164 86776 64166
rect 87216 63674 87272 63676
rect 87296 63674 87352 63676
rect 87376 63674 87432 63676
rect 87456 63674 87512 63676
rect 84530 63560 84586 63616
rect 87216 63622 87262 63674
rect 87262 63622 87272 63674
rect 87296 63622 87326 63674
rect 87326 63622 87338 63674
rect 87338 63622 87352 63674
rect 87376 63622 87390 63674
rect 87390 63622 87402 63674
rect 87402 63622 87432 63674
rect 87456 63622 87466 63674
rect 87466 63622 87512 63674
rect 87216 63620 87272 63622
rect 87296 63620 87352 63622
rect 87376 63620 87432 63622
rect 87456 63620 87512 63622
rect 88578 63560 88634 63616
rect 86480 63130 86536 63132
rect 86560 63130 86616 63132
rect 86640 63130 86696 63132
rect 86720 63130 86776 63132
rect 86480 63078 86526 63130
rect 86526 63078 86536 63130
rect 86560 63078 86590 63130
rect 86590 63078 86602 63130
rect 86602 63078 86616 63130
rect 86640 63078 86654 63130
rect 86654 63078 86666 63130
rect 86666 63078 86696 63130
rect 86720 63078 86730 63130
rect 86730 63078 86776 63130
rect 86480 63076 86536 63078
rect 86560 63076 86616 63078
rect 86640 63076 86696 63078
rect 86720 63076 86776 63078
rect 87216 62586 87272 62588
rect 87296 62586 87352 62588
rect 87376 62586 87432 62588
rect 87456 62586 87512 62588
rect 84806 62472 84862 62528
rect 87216 62534 87262 62586
rect 87262 62534 87272 62586
rect 87296 62534 87326 62586
rect 87326 62534 87338 62586
rect 87338 62534 87352 62586
rect 87376 62534 87390 62586
rect 87390 62534 87402 62586
rect 87402 62534 87432 62586
rect 87456 62534 87466 62586
rect 87466 62534 87512 62586
rect 87216 62532 87272 62534
rect 87296 62532 87352 62534
rect 87376 62532 87432 62534
rect 87456 62532 87512 62534
rect 88394 62200 88450 62256
rect 86480 62042 86536 62044
rect 86560 62042 86616 62044
rect 86640 62042 86696 62044
rect 86720 62042 86776 62044
rect 86480 61990 86526 62042
rect 86526 61990 86536 62042
rect 86560 61990 86590 62042
rect 86590 61990 86602 62042
rect 86602 61990 86616 62042
rect 86640 61990 86654 62042
rect 86654 61990 86666 62042
rect 86666 61990 86696 62042
rect 86720 61990 86730 62042
rect 86730 61990 86776 62042
rect 86480 61988 86536 61990
rect 86560 61988 86616 61990
rect 86640 61988 86696 61990
rect 86720 61988 86776 61990
rect 88210 61556 88212 61576
rect 88212 61556 88264 61576
rect 88264 61556 88266 61576
rect 88210 61520 88266 61556
rect 87216 61498 87272 61500
rect 87296 61498 87352 61500
rect 87376 61498 87432 61500
rect 87456 61498 87512 61500
rect 85818 61384 85874 61440
rect 87216 61446 87262 61498
rect 87262 61446 87272 61498
rect 87296 61446 87326 61498
rect 87326 61446 87338 61498
rect 87338 61446 87352 61498
rect 87376 61446 87390 61498
rect 87390 61446 87402 61498
rect 87402 61446 87432 61498
rect 87456 61446 87466 61498
rect 87466 61446 87512 61498
rect 87216 61444 87272 61446
rect 87296 61444 87352 61446
rect 87376 61444 87432 61446
rect 87456 61444 87512 61446
rect 86480 60954 86536 60956
rect 86560 60954 86616 60956
rect 86640 60954 86696 60956
rect 86720 60954 86776 60956
rect 86480 60902 86526 60954
rect 86526 60902 86536 60954
rect 86560 60902 86590 60954
rect 86590 60902 86602 60954
rect 86602 60902 86616 60954
rect 86640 60902 86654 60954
rect 86654 60902 86666 60954
rect 86666 60902 86696 60954
rect 86720 60902 86730 60954
rect 86730 60902 86776 60954
rect 86480 60900 86536 60902
rect 86560 60900 86616 60902
rect 86640 60900 86696 60902
rect 86720 60900 86776 60902
rect 87216 60410 87272 60412
rect 87296 60410 87352 60412
rect 87376 60410 87432 60412
rect 87456 60410 87512 60412
rect 85818 60296 85874 60352
rect 87216 60358 87262 60410
rect 87262 60358 87272 60410
rect 87296 60358 87326 60410
rect 87326 60358 87338 60410
rect 87338 60358 87352 60410
rect 87376 60358 87390 60410
rect 87390 60358 87402 60410
rect 87402 60358 87432 60410
rect 87456 60358 87466 60410
rect 87466 60358 87512 60410
rect 87216 60356 87272 60358
rect 87296 60356 87352 60358
rect 87376 60356 87432 60358
rect 87456 60356 87512 60358
rect 88210 60160 88266 60216
rect 86480 59866 86536 59868
rect 86560 59866 86616 59868
rect 86640 59866 86696 59868
rect 86720 59866 86776 59868
rect 86480 59814 86526 59866
rect 86526 59814 86536 59866
rect 86560 59814 86590 59866
rect 86590 59814 86602 59866
rect 86602 59814 86616 59866
rect 86640 59814 86654 59866
rect 86654 59814 86666 59866
rect 86666 59814 86696 59866
rect 86720 59814 86730 59866
rect 86730 59814 86776 59866
rect 86480 59812 86536 59814
rect 86560 59812 86616 59814
rect 86640 59812 86696 59814
rect 86720 59812 86776 59814
rect 87474 59516 87476 59536
rect 87476 59516 87528 59536
rect 87528 59516 87530 59536
rect 87474 59480 87530 59516
rect 88210 59480 88266 59536
rect 87216 59322 87272 59324
rect 87296 59322 87352 59324
rect 87376 59322 87432 59324
rect 87456 59322 87512 59324
rect 87216 59270 87262 59322
rect 87262 59270 87272 59322
rect 87296 59270 87326 59322
rect 87326 59270 87338 59322
rect 87338 59270 87352 59322
rect 87376 59270 87390 59322
rect 87390 59270 87402 59322
rect 87402 59270 87432 59322
rect 87456 59270 87466 59322
rect 87466 59270 87512 59322
rect 87216 59268 87272 59270
rect 87296 59268 87352 59270
rect 87376 59268 87432 59270
rect 87456 59268 87512 59270
rect 86480 58778 86536 58780
rect 86560 58778 86616 58780
rect 86640 58778 86696 58780
rect 86720 58778 86776 58780
rect 86480 58726 86526 58778
rect 86526 58726 86536 58778
rect 86560 58726 86590 58778
rect 86590 58726 86602 58778
rect 86602 58726 86616 58778
rect 86640 58726 86654 58778
rect 86654 58726 86666 58778
rect 86666 58726 86696 58778
rect 86720 58726 86730 58778
rect 86730 58726 86776 58778
rect 86480 58724 86536 58726
rect 86560 58724 86616 58726
rect 86640 58724 86696 58726
rect 86720 58724 86776 58726
rect 87216 58234 87272 58236
rect 87296 58234 87352 58236
rect 87376 58234 87432 58236
rect 87456 58234 87512 58236
rect 85082 58120 85138 58176
rect 87216 58182 87262 58234
rect 87262 58182 87272 58234
rect 87296 58182 87326 58234
rect 87326 58182 87338 58234
rect 87338 58182 87352 58234
rect 87376 58182 87390 58234
rect 87390 58182 87402 58234
rect 87402 58182 87432 58234
rect 87456 58182 87466 58234
rect 87466 58182 87512 58234
rect 87216 58180 87272 58182
rect 87296 58180 87352 58182
rect 87376 58180 87432 58182
rect 87456 58180 87512 58182
rect 88578 58120 88634 58176
rect 86480 57690 86536 57692
rect 86560 57690 86616 57692
rect 86640 57690 86696 57692
rect 86720 57690 86776 57692
rect 86480 57638 86526 57690
rect 86526 57638 86536 57690
rect 86560 57638 86590 57690
rect 86590 57638 86602 57690
rect 86602 57638 86616 57690
rect 86640 57638 86654 57690
rect 86654 57638 86666 57690
rect 86666 57638 86696 57690
rect 86720 57638 86730 57690
rect 86730 57638 86776 57690
rect 86480 57636 86536 57638
rect 86560 57636 86616 57638
rect 86640 57636 86696 57638
rect 86720 57636 86776 57638
rect 87216 57146 87272 57148
rect 87296 57146 87352 57148
rect 87376 57146 87432 57148
rect 87456 57146 87512 57148
rect 87216 57094 87262 57146
rect 87262 57094 87272 57146
rect 87296 57094 87326 57146
rect 87326 57094 87338 57146
rect 87338 57094 87352 57146
rect 87376 57094 87390 57146
rect 87390 57094 87402 57146
rect 87402 57094 87432 57146
rect 87456 57094 87466 57146
rect 87466 57094 87512 57146
rect 87216 57092 87272 57094
rect 87296 57092 87352 57094
rect 87376 57092 87432 57094
rect 87456 57092 87512 57094
rect 87566 56916 87622 56952
rect 87566 56896 87568 56916
rect 87568 56896 87620 56916
rect 87620 56896 87622 56916
rect 88578 56760 88634 56816
rect 86480 56602 86536 56604
rect 86560 56602 86616 56604
rect 86640 56602 86696 56604
rect 86720 56602 86776 56604
rect 86480 56550 86526 56602
rect 86526 56550 86536 56602
rect 86560 56550 86590 56602
rect 86590 56550 86602 56602
rect 86602 56550 86616 56602
rect 86640 56550 86654 56602
rect 86654 56550 86666 56602
rect 86666 56550 86696 56602
rect 86720 56550 86730 56602
rect 86730 56550 86776 56602
rect 86480 56548 86536 56550
rect 86560 56548 86616 56550
rect 86640 56548 86696 56550
rect 86720 56548 86776 56550
rect 88210 56116 88212 56136
rect 88212 56116 88264 56136
rect 88264 56116 88266 56136
rect 88210 56080 88266 56116
rect 87216 56058 87272 56060
rect 87296 56058 87352 56060
rect 87376 56058 87432 56060
rect 87456 56058 87512 56060
rect 85818 55944 85874 56000
rect 87216 56006 87262 56058
rect 87262 56006 87272 56058
rect 87296 56006 87326 56058
rect 87326 56006 87338 56058
rect 87338 56006 87352 56058
rect 87376 56006 87390 56058
rect 87390 56006 87402 56058
rect 87402 56006 87432 56058
rect 87456 56006 87466 56058
rect 87466 56006 87512 56058
rect 87216 56004 87272 56006
rect 87296 56004 87352 56006
rect 87376 56004 87432 56006
rect 87456 56004 87512 56006
rect 86480 55514 86536 55516
rect 86560 55514 86616 55516
rect 86640 55514 86696 55516
rect 86720 55514 86776 55516
rect 86480 55462 86526 55514
rect 86526 55462 86536 55514
rect 86560 55462 86590 55514
rect 86590 55462 86602 55514
rect 86602 55462 86616 55514
rect 86640 55462 86654 55514
rect 86654 55462 86666 55514
rect 86666 55462 86696 55514
rect 86720 55462 86730 55514
rect 86730 55462 86776 55514
rect 86480 55460 86536 55462
rect 86560 55460 86616 55462
rect 86640 55460 86696 55462
rect 86720 55460 86776 55462
rect 87216 54970 87272 54972
rect 87296 54970 87352 54972
rect 87376 54970 87432 54972
rect 87456 54970 87512 54972
rect 85818 54856 85874 54912
rect 87216 54918 87262 54970
rect 87262 54918 87272 54970
rect 87296 54918 87326 54970
rect 87326 54918 87338 54970
rect 87338 54918 87352 54970
rect 87376 54918 87390 54970
rect 87390 54918 87402 54970
rect 87402 54918 87432 54970
rect 87456 54918 87466 54970
rect 87466 54918 87512 54970
rect 87216 54916 87272 54918
rect 87296 54916 87352 54918
rect 87376 54916 87432 54918
rect 87456 54916 87512 54918
rect 88210 54720 88266 54776
rect 86480 54426 86536 54428
rect 86560 54426 86616 54428
rect 86640 54426 86696 54428
rect 86720 54426 86776 54428
rect 86480 54374 86526 54426
rect 86526 54374 86536 54426
rect 86560 54374 86590 54426
rect 86590 54374 86602 54426
rect 86602 54374 86616 54426
rect 86640 54374 86654 54426
rect 86654 54374 86666 54426
rect 86666 54374 86696 54426
rect 86720 54374 86730 54426
rect 86730 54374 86776 54426
rect 86480 54372 86536 54374
rect 86560 54372 86616 54374
rect 86640 54372 86696 54374
rect 86720 54372 86776 54374
rect 88210 54076 88212 54096
rect 88212 54076 88264 54096
rect 88264 54076 88266 54096
rect 88210 54040 88266 54076
rect 87216 53882 87272 53884
rect 87296 53882 87352 53884
rect 87376 53882 87432 53884
rect 87456 53882 87512 53884
rect 84530 53768 84586 53824
rect 87216 53830 87262 53882
rect 87262 53830 87272 53882
rect 87296 53830 87326 53882
rect 87326 53830 87338 53882
rect 87338 53830 87352 53882
rect 87376 53830 87390 53882
rect 87390 53830 87402 53882
rect 87402 53830 87432 53882
rect 87456 53830 87466 53882
rect 87466 53830 87512 53882
rect 87216 53828 87272 53830
rect 87296 53828 87352 53830
rect 87376 53828 87432 53830
rect 87456 53828 87512 53830
rect 86480 53338 86536 53340
rect 86560 53338 86616 53340
rect 86640 53338 86696 53340
rect 86720 53338 86776 53340
rect 86480 53286 86526 53338
rect 86526 53286 86536 53338
rect 86560 53286 86590 53338
rect 86590 53286 86602 53338
rect 86602 53286 86616 53338
rect 86640 53286 86654 53338
rect 86654 53286 86666 53338
rect 86666 53286 86696 53338
rect 86720 53286 86730 53338
rect 86730 53286 86776 53338
rect 86480 53284 86536 53286
rect 86560 53284 86616 53286
rect 86640 53284 86696 53286
rect 86720 53284 86776 53286
rect 87566 52988 87568 53008
rect 87568 52988 87620 53008
rect 87620 52988 87622 53008
rect 87566 52952 87622 52988
rect 87216 52794 87272 52796
rect 87296 52794 87352 52796
rect 87376 52794 87432 52796
rect 87456 52794 87512 52796
rect 87216 52742 87262 52794
rect 87262 52742 87272 52794
rect 87296 52742 87326 52794
rect 87326 52742 87338 52794
rect 87338 52742 87352 52794
rect 87376 52742 87390 52794
rect 87390 52742 87402 52794
rect 87402 52742 87432 52794
rect 87456 52742 87466 52794
rect 87466 52742 87512 52794
rect 87216 52740 87272 52742
rect 87296 52740 87352 52742
rect 87376 52740 87432 52742
rect 87456 52740 87512 52742
rect 88210 52680 88266 52736
rect 86480 52250 86536 52252
rect 86560 52250 86616 52252
rect 86640 52250 86696 52252
rect 86720 52250 86776 52252
rect 86480 52198 86526 52250
rect 86526 52198 86536 52250
rect 86560 52198 86590 52250
rect 86590 52198 86602 52250
rect 86602 52198 86616 52250
rect 86640 52198 86654 52250
rect 86654 52198 86666 52250
rect 86666 52198 86696 52250
rect 86720 52198 86730 52250
rect 86730 52198 86776 52250
rect 86480 52196 86536 52198
rect 86560 52196 86616 52198
rect 86640 52196 86696 52198
rect 86720 52196 86776 52198
rect 87216 51706 87272 51708
rect 87296 51706 87352 51708
rect 87376 51706 87432 51708
rect 87456 51706 87512 51708
rect 87216 51654 87262 51706
rect 87262 51654 87272 51706
rect 87296 51654 87326 51706
rect 87326 51654 87338 51706
rect 87338 51654 87352 51706
rect 87376 51654 87390 51706
rect 87390 51654 87402 51706
rect 87402 51654 87432 51706
rect 87456 51654 87466 51706
rect 87466 51654 87512 51706
rect 87216 51652 87272 51654
rect 87296 51652 87352 51654
rect 87376 51652 87432 51654
rect 87456 51652 87512 51654
rect 87566 51476 87622 51512
rect 87566 51456 87568 51476
rect 87568 51456 87620 51476
rect 87620 51456 87622 51476
rect 88210 51340 88266 51376
rect 88210 51320 88212 51340
rect 88212 51320 88264 51340
rect 88264 51320 88266 51340
rect 86480 51162 86536 51164
rect 86560 51162 86616 51164
rect 86640 51162 86696 51164
rect 86720 51162 86776 51164
rect 86480 51110 86526 51162
rect 86526 51110 86536 51162
rect 86560 51110 86590 51162
rect 86590 51110 86602 51162
rect 86602 51110 86616 51162
rect 86640 51110 86654 51162
rect 86654 51110 86666 51162
rect 86666 51110 86696 51162
rect 86720 51110 86730 51162
rect 86730 51110 86776 51162
rect 86480 51108 86536 51110
rect 86560 51108 86616 51110
rect 86640 51108 86696 51110
rect 86720 51108 86776 51110
rect 87216 50618 87272 50620
rect 87296 50618 87352 50620
rect 87376 50618 87432 50620
rect 87456 50618 87512 50620
rect 85450 50504 85506 50560
rect 85634 50504 85690 50560
rect 87216 50566 87262 50618
rect 87262 50566 87272 50618
rect 87296 50566 87326 50618
rect 87326 50566 87338 50618
rect 87338 50566 87352 50618
rect 87376 50566 87390 50618
rect 87390 50566 87402 50618
rect 87402 50566 87432 50618
rect 87456 50566 87466 50618
rect 87466 50566 87512 50618
rect 87216 50564 87272 50566
rect 87296 50564 87352 50566
rect 87376 50564 87432 50566
rect 87456 50564 87512 50566
rect 85358 48328 85414 48384
rect 83610 44588 83666 44644
rect 84806 35952 84862 36008
rect 84806 30512 84862 30568
rect 84806 24936 84862 24992
rect 84806 20720 84862 20776
rect 84806 15280 84862 15336
rect 83426 14124 83482 14180
rect 46442 10928 46498 10984
rect 83334 10860 83390 10916
rect 46442 10112 46498 10168
rect 54528 7642 54584 7644
rect 54608 7642 54664 7644
rect 54688 7642 54744 7644
rect 54768 7642 54824 7644
rect 54528 7590 54574 7642
rect 54574 7590 54584 7642
rect 54608 7590 54638 7642
rect 54638 7590 54650 7642
rect 54650 7590 54664 7642
rect 54688 7590 54702 7642
rect 54702 7590 54714 7642
rect 54714 7590 54744 7642
rect 54768 7590 54778 7642
rect 54778 7590 54824 7642
rect 54528 7588 54584 7590
rect 54608 7588 54664 7590
rect 54688 7588 54744 7590
rect 54768 7588 54824 7590
rect 55188 7098 55244 7100
rect 55268 7098 55324 7100
rect 55348 7098 55404 7100
rect 55428 7098 55484 7100
rect 55188 7046 55234 7098
rect 55234 7046 55244 7098
rect 55268 7046 55298 7098
rect 55298 7046 55310 7098
rect 55310 7046 55324 7098
rect 55348 7046 55362 7098
rect 55362 7046 55374 7098
rect 55374 7046 55404 7098
rect 55428 7046 55438 7098
rect 55438 7046 55484 7098
rect 55188 7044 55244 7046
rect 55268 7044 55324 7046
rect 55348 7044 55404 7046
rect 55428 7044 55484 7046
rect 54528 6554 54584 6556
rect 54608 6554 54664 6556
rect 54688 6554 54744 6556
rect 54768 6554 54824 6556
rect 54528 6502 54574 6554
rect 54574 6502 54584 6554
rect 54608 6502 54638 6554
rect 54638 6502 54650 6554
rect 54650 6502 54664 6554
rect 54688 6502 54702 6554
rect 54702 6502 54714 6554
rect 54714 6502 54744 6554
rect 54768 6502 54778 6554
rect 54778 6502 54824 6554
rect 54528 6500 54584 6502
rect 54608 6500 54664 6502
rect 54688 6500 54744 6502
rect 54768 6500 54824 6502
rect 55188 6010 55244 6012
rect 55268 6010 55324 6012
rect 55348 6010 55404 6012
rect 55428 6010 55484 6012
rect 55188 5958 55234 6010
rect 55234 5958 55244 6010
rect 55268 5958 55298 6010
rect 55298 5958 55310 6010
rect 55310 5958 55324 6010
rect 55348 5958 55362 6010
rect 55362 5958 55374 6010
rect 55374 5958 55404 6010
rect 55428 5958 55438 6010
rect 55438 5958 55484 6010
rect 55188 5956 55244 5958
rect 55268 5956 55324 5958
rect 55348 5956 55404 5958
rect 55428 5956 55484 5958
rect 54528 5466 54584 5468
rect 54608 5466 54664 5468
rect 54688 5466 54744 5468
rect 54768 5466 54824 5468
rect 54528 5414 54574 5466
rect 54574 5414 54584 5466
rect 54608 5414 54638 5466
rect 54638 5414 54650 5466
rect 54650 5414 54664 5466
rect 54688 5414 54702 5466
rect 54702 5414 54714 5466
rect 54714 5414 54744 5466
rect 54768 5414 54778 5466
rect 54778 5414 54824 5466
rect 54528 5412 54584 5414
rect 54608 5412 54664 5414
rect 54688 5412 54744 5414
rect 54768 5412 54824 5414
rect 72928 7642 72984 7644
rect 73008 7642 73064 7644
rect 73088 7642 73144 7644
rect 73168 7642 73224 7644
rect 72928 7590 72974 7642
rect 72974 7590 72984 7642
rect 73008 7590 73038 7642
rect 73038 7590 73050 7642
rect 73050 7590 73064 7642
rect 73088 7590 73102 7642
rect 73102 7590 73114 7642
rect 73114 7590 73144 7642
rect 73168 7590 73178 7642
rect 73178 7590 73224 7642
rect 72928 7588 72984 7590
rect 73008 7588 73064 7590
rect 73088 7588 73144 7590
rect 73168 7588 73224 7590
rect 72928 6554 72984 6556
rect 73008 6554 73064 6556
rect 73088 6554 73144 6556
rect 73168 6554 73224 6556
rect 72928 6502 72974 6554
rect 72974 6502 72984 6554
rect 73008 6502 73038 6554
rect 73038 6502 73050 6554
rect 73050 6502 73064 6554
rect 73088 6502 73102 6554
rect 73102 6502 73114 6554
rect 73114 6502 73144 6554
rect 73168 6502 73178 6554
rect 73178 6502 73224 6554
rect 72928 6500 72984 6502
rect 73008 6500 73064 6502
rect 73088 6500 73144 6502
rect 73168 6500 73224 6502
rect 72928 5466 72984 5468
rect 73008 5466 73064 5468
rect 73088 5466 73144 5468
rect 73168 5466 73224 5468
rect 72928 5414 72974 5466
rect 72974 5414 72984 5466
rect 73008 5414 73038 5466
rect 73038 5414 73050 5466
rect 73050 5414 73064 5466
rect 73088 5414 73102 5466
rect 73102 5414 73114 5466
rect 73114 5414 73144 5466
rect 73168 5414 73178 5466
rect 73178 5414 73224 5466
rect 72928 5412 72984 5414
rect 73008 5412 73064 5414
rect 73088 5412 73144 5414
rect 73168 5412 73224 5414
rect 73588 7098 73644 7100
rect 73668 7098 73724 7100
rect 73748 7098 73804 7100
rect 73828 7098 73884 7100
rect 73588 7046 73634 7098
rect 73634 7046 73644 7098
rect 73668 7046 73698 7098
rect 73698 7046 73710 7098
rect 73710 7046 73724 7098
rect 73748 7046 73762 7098
rect 73762 7046 73774 7098
rect 73774 7046 73804 7098
rect 73828 7046 73838 7098
rect 73838 7046 73884 7098
rect 73588 7044 73644 7046
rect 73668 7044 73724 7046
rect 73748 7044 73804 7046
rect 73828 7044 73884 7046
rect 73588 6010 73644 6012
rect 73668 6010 73724 6012
rect 73748 6010 73804 6012
rect 73828 6010 73884 6012
rect 73588 5958 73634 6010
rect 73634 5958 73644 6010
rect 73668 5958 73698 6010
rect 73698 5958 73710 6010
rect 73710 5958 73724 6010
rect 73748 5958 73762 6010
rect 73762 5958 73774 6010
rect 73774 5958 73804 6010
rect 73828 5958 73838 6010
rect 73838 5958 73884 6010
rect 73588 5956 73644 5958
rect 73668 5956 73724 5958
rect 73748 5956 73804 5958
rect 73828 5956 73884 5958
rect 83610 13036 83666 13092
rect 86480 50074 86536 50076
rect 86560 50074 86616 50076
rect 86640 50074 86696 50076
rect 86720 50074 86776 50076
rect 86480 50022 86526 50074
rect 86526 50022 86536 50074
rect 86560 50022 86590 50074
rect 86590 50022 86602 50074
rect 86602 50022 86616 50074
rect 86640 50022 86654 50074
rect 86654 50022 86666 50074
rect 86666 50022 86696 50074
rect 86720 50022 86730 50074
rect 86730 50022 86776 50074
rect 86480 50020 86536 50022
rect 86560 50020 86616 50022
rect 86640 50020 86696 50022
rect 86720 50020 86776 50022
rect 87216 49530 87272 49532
rect 87296 49530 87352 49532
rect 87376 49530 87432 49532
rect 87456 49530 87512 49532
rect 85634 49416 85690 49472
rect 87216 49478 87262 49530
rect 87262 49478 87272 49530
rect 87296 49478 87326 49530
rect 87326 49478 87338 49530
rect 87338 49478 87352 49530
rect 87376 49478 87390 49530
rect 87390 49478 87402 49530
rect 87402 49478 87432 49530
rect 87456 49478 87466 49530
rect 87466 49478 87512 49530
rect 87216 49476 87272 49478
rect 87296 49476 87352 49478
rect 87376 49476 87432 49478
rect 87456 49476 87512 49478
rect 86480 48986 86536 48988
rect 86560 48986 86616 48988
rect 86640 48986 86696 48988
rect 86720 48986 86776 48988
rect 86480 48934 86526 48986
rect 86526 48934 86536 48986
rect 86560 48934 86590 48986
rect 86590 48934 86602 48986
rect 86602 48934 86616 48986
rect 86640 48934 86654 48986
rect 86654 48934 86666 48986
rect 86666 48934 86696 48986
rect 86720 48934 86730 48986
rect 86730 48934 86776 48986
rect 86480 48932 86536 48934
rect 86560 48932 86616 48934
rect 86640 48932 86696 48934
rect 86720 48932 86776 48934
rect 88210 48636 88212 48656
rect 88212 48636 88264 48656
rect 88264 48636 88266 48656
rect 88210 48600 88266 48636
rect 87216 48442 87272 48444
rect 87296 48442 87352 48444
rect 87376 48442 87432 48444
rect 87456 48442 87512 48444
rect 87216 48390 87262 48442
rect 87262 48390 87272 48442
rect 87296 48390 87326 48442
rect 87326 48390 87338 48442
rect 87338 48390 87352 48442
rect 87376 48390 87390 48442
rect 87390 48390 87402 48442
rect 87402 48390 87432 48442
rect 87456 48390 87466 48442
rect 87466 48390 87512 48442
rect 87216 48388 87272 48390
rect 87296 48388 87352 48390
rect 87376 48388 87432 48390
rect 87456 48388 87512 48390
rect 88210 47956 88212 47976
rect 88212 47956 88264 47976
rect 88264 47956 88266 47976
rect 88210 47920 88266 47956
rect 86480 47898 86536 47900
rect 86560 47898 86616 47900
rect 86640 47898 86696 47900
rect 86720 47898 86776 47900
rect 86480 47846 86526 47898
rect 86526 47846 86536 47898
rect 86560 47846 86590 47898
rect 86590 47846 86602 47898
rect 86602 47846 86616 47898
rect 86640 47846 86654 47898
rect 86654 47846 86666 47898
rect 86666 47846 86696 47898
rect 86720 47846 86730 47898
rect 86730 47846 86776 47898
rect 86480 47844 86536 47846
rect 86560 47844 86616 47846
rect 86640 47844 86696 47846
rect 86720 47844 86776 47846
rect 87216 47354 87272 47356
rect 87296 47354 87352 47356
rect 87376 47354 87432 47356
rect 87456 47354 87512 47356
rect 85818 47240 85874 47296
rect 87216 47302 87262 47354
rect 87262 47302 87272 47354
rect 87296 47302 87326 47354
rect 87326 47302 87338 47354
rect 87338 47302 87352 47354
rect 87376 47302 87390 47354
rect 87390 47302 87402 47354
rect 87402 47302 87432 47354
rect 87456 47302 87466 47354
rect 87466 47302 87512 47354
rect 87216 47300 87272 47302
rect 87296 47300 87352 47302
rect 87376 47300 87432 47302
rect 87456 47300 87512 47302
rect 88210 47240 88266 47296
rect 86480 46810 86536 46812
rect 86560 46810 86616 46812
rect 86640 46810 86696 46812
rect 86720 46810 86776 46812
rect 86480 46758 86526 46810
rect 86526 46758 86536 46810
rect 86560 46758 86590 46810
rect 86590 46758 86602 46810
rect 86602 46758 86616 46810
rect 86640 46758 86654 46810
rect 86654 46758 86666 46810
rect 86666 46758 86696 46810
rect 86720 46758 86730 46810
rect 86730 46758 86776 46810
rect 86480 46756 86536 46758
rect 86560 46756 86616 46758
rect 86640 46756 86696 46758
rect 86720 46756 86776 46758
rect 88210 46560 88266 46616
rect 87216 46266 87272 46268
rect 87296 46266 87352 46268
rect 87376 46266 87432 46268
rect 87456 46266 87512 46268
rect 87216 46214 87262 46266
rect 87262 46214 87272 46266
rect 87296 46214 87326 46266
rect 87326 46214 87338 46266
rect 87338 46214 87352 46266
rect 87376 46214 87390 46266
rect 87390 46214 87402 46266
rect 87402 46214 87432 46266
rect 87456 46214 87466 46266
rect 87466 46214 87512 46266
rect 87216 46212 87272 46214
rect 87296 46212 87352 46214
rect 87376 46212 87432 46214
rect 87456 46212 87512 46214
rect 86480 45722 86536 45724
rect 86560 45722 86616 45724
rect 86640 45722 86696 45724
rect 86720 45722 86776 45724
rect 86480 45670 86526 45722
rect 86526 45670 86536 45722
rect 86560 45670 86590 45722
rect 86590 45670 86602 45722
rect 86602 45670 86616 45722
rect 86640 45670 86654 45722
rect 86654 45670 86666 45722
rect 86666 45670 86696 45722
rect 86720 45670 86730 45722
rect 86730 45670 86776 45722
rect 86480 45668 86536 45670
rect 86560 45668 86616 45670
rect 86640 45668 86696 45670
rect 86720 45668 86776 45670
rect 86002 45372 86004 45392
rect 86004 45372 86056 45392
rect 86056 45372 86058 45392
rect 86002 45336 86058 45372
rect 86186 45236 86188 45256
rect 86188 45236 86240 45256
rect 86240 45236 86242 45256
rect 86186 45200 86242 45236
rect 88210 45200 88266 45256
rect 87216 45178 87272 45180
rect 87296 45178 87352 45180
rect 87376 45178 87432 45180
rect 87456 45178 87512 45180
rect 85634 45064 85690 45120
rect 87216 45126 87262 45178
rect 87262 45126 87272 45178
rect 87296 45126 87326 45178
rect 87326 45126 87338 45178
rect 87338 45126 87352 45178
rect 87376 45126 87390 45178
rect 87390 45126 87402 45178
rect 87402 45126 87432 45178
rect 87456 45126 87466 45178
rect 87466 45126 87512 45178
rect 87216 45124 87272 45126
rect 87296 45124 87352 45126
rect 87376 45124 87432 45126
rect 87456 45124 87512 45126
rect 86480 44634 86536 44636
rect 86560 44634 86616 44636
rect 86640 44634 86696 44636
rect 86720 44634 86776 44636
rect 86480 44582 86526 44634
rect 86526 44582 86536 44634
rect 86560 44582 86590 44634
rect 86590 44582 86602 44634
rect 86602 44582 86616 44634
rect 86640 44582 86654 44634
rect 86654 44582 86666 44634
rect 86666 44582 86696 44634
rect 86720 44582 86730 44634
rect 86730 44582 86776 44634
rect 86480 44580 86536 44582
rect 86560 44580 86616 44582
rect 86640 44580 86696 44582
rect 86720 44580 86776 44582
rect 88210 44520 88266 44576
rect 87216 44090 87272 44092
rect 87296 44090 87352 44092
rect 87376 44090 87432 44092
rect 87456 44090 87512 44092
rect 87216 44038 87262 44090
rect 87262 44038 87272 44090
rect 87296 44038 87326 44090
rect 87326 44038 87338 44090
rect 87338 44038 87352 44090
rect 87376 44038 87390 44090
rect 87390 44038 87402 44090
rect 87402 44038 87432 44090
rect 87456 44038 87466 44090
rect 87466 44038 87512 44090
rect 87216 44036 87272 44038
rect 87296 44036 87352 44038
rect 87376 44036 87432 44038
rect 87456 44036 87512 44038
rect 88210 43840 88266 43896
rect 86480 43546 86536 43548
rect 86560 43546 86616 43548
rect 86640 43546 86696 43548
rect 86720 43546 86776 43548
rect 85818 43432 85874 43488
rect 86480 43494 86526 43546
rect 86526 43494 86536 43546
rect 86560 43494 86590 43546
rect 86590 43494 86602 43546
rect 86602 43494 86616 43546
rect 86640 43494 86654 43546
rect 86654 43494 86666 43546
rect 86666 43494 86696 43546
rect 86720 43494 86730 43546
rect 86730 43494 86776 43546
rect 86480 43492 86536 43494
rect 86560 43492 86616 43494
rect 86640 43492 86696 43494
rect 86720 43492 86776 43494
rect 88210 43196 88212 43216
rect 88212 43196 88264 43216
rect 88264 43196 88266 43216
rect 88210 43160 88266 43196
rect 87216 43002 87272 43004
rect 87296 43002 87352 43004
rect 87376 43002 87432 43004
rect 87456 43002 87512 43004
rect 87216 42950 87262 43002
rect 87262 42950 87272 43002
rect 87296 42950 87326 43002
rect 87326 42950 87338 43002
rect 87338 42950 87352 43002
rect 87376 42950 87390 43002
rect 87390 42950 87402 43002
rect 87402 42950 87432 43002
rect 87456 42950 87466 43002
rect 87466 42950 87512 43002
rect 87216 42948 87272 42950
rect 87296 42948 87352 42950
rect 87376 42948 87432 42950
rect 87456 42948 87512 42950
rect 85818 42480 85874 42536
rect 88210 42480 88266 42536
rect 86480 42458 86536 42460
rect 86560 42458 86616 42460
rect 86640 42458 86696 42460
rect 86720 42458 86776 42460
rect 86480 42406 86526 42458
rect 86526 42406 86536 42458
rect 86560 42406 86590 42458
rect 86590 42406 86602 42458
rect 86602 42406 86616 42458
rect 86640 42406 86654 42458
rect 86654 42406 86666 42458
rect 86666 42406 86696 42458
rect 86720 42406 86730 42458
rect 86730 42406 86776 42458
rect 86480 42404 86536 42406
rect 86560 42404 86616 42406
rect 86640 42404 86696 42406
rect 86720 42404 86776 42406
rect 87216 41914 87272 41916
rect 87296 41914 87352 41916
rect 87376 41914 87432 41916
rect 87456 41914 87512 41916
rect 87216 41862 87262 41914
rect 87262 41862 87272 41914
rect 87296 41862 87326 41914
rect 87326 41862 87338 41914
rect 87338 41862 87352 41914
rect 87376 41862 87390 41914
rect 87390 41862 87402 41914
rect 87402 41862 87432 41914
rect 87456 41862 87466 41914
rect 87466 41862 87512 41914
rect 87216 41860 87272 41862
rect 87296 41860 87352 41862
rect 87376 41860 87432 41862
rect 87456 41860 87512 41862
rect 87566 41528 87622 41584
rect 86480 41370 86536 41372
rect 86560 41370 86616 41372
rect 86640 41370 86696 41372
rect 86720 41370 86776 41372
rect 86480 41318 86526 41370
rect 86526 41318 86536 41370
rect 86560 41318 86590 41370
rect 86590 41318 86602 41370
rect 86602 41318 86616 41370
rect 86640 41318 86654 41370
rect 86654 41318 86666 41370
rect 86666 41318 86696 41370
rect 86720 41318 86730 41370
rect 86730 41318 86776 41370
rect 86480 41316 86536 41318
rect 86560 41316 86616 41318
rect 86640 41316 86696 41318
rect 86720 41316 86776 41318
rect 88210 41120 88266 41176
rect 87216 40826 87272 40828
rect 87296 40826 87352 40828
rect 87376 40826 87432 40828
rect 87456 40826 87512 40828
rect 87216 40774 87262 40826
rect 87262 40774 87272 40826
rect 87296 40774 87326 40826
rect 87326 40774 87338 40826
rect 87338 40774 87352 40826
rect 87376 40774 87390 40826
rect 87390 40774 87402 40826
rect 87402 40774 87432 40826
rect 87456 40774 87466 40826
rect 87466 40774 87512 40826
rect 87216 40772 87272 40774
rect 87296 40772 87352 40774
rect 87376 40772 87432 40774
rect 87456 40772 87512 40774
rect 87934 40476 87936 40496
rect 87936 40476 87988 40496
rect 87988 40476 87990 40496
rect 87934 40440 87990 40476
rect 88210 40476 88212 40496
rect 88212 40476 88264 40496
rect 88264 40476 88266 40496
rect 88210 40440 88266 40476
rect 86480 40282 86536 40284
rect 86560 40282 86616 40284
rect 86640 40282 86696 40284
rect 86720 40282 86776 40284
rect 86480 40230 86526 40282
rect 86526 40230 86536 40282
rect 86560 40230 86590 40282
rect 86590 40230 86602 40282
rect 86602 40230 86616 40282
rect 86640 40230 86654 40282
rect 86654 40230 86666 40282
rect 86666 40230 86696 40282
rect 86720 40230 86730 40282
rect 86730 40230 86776 40282
rect 86480 40228 86536 40230
rect 86560 40228 86616 40230
rect 86640 40228 86696 40230
rect 86720 40228 86776 40230
rect 87216 39738 87272 39740
rect 87296 39738 87352 39740
rect 87376 39738 87432 39740
rect 87456 39738 87512 39740
rect 87216 39686 87262 39738
rect 87262 39686 87272 39738
rect 87296 39686 87326 39738
rect 87326 39686 87338 39738
rect 87338 39686 87352 39738
rect 87376 39686 87390 39738
rect 87390 39686 87402 39738
rect 87402 39686 87432 39738
rect 87456 39686 87466 39738
rect 87466 39686 87512 39738
rect 87216 39684 87272 39686
rect 87296 39684 87352 39686
rect 87376 39684 87432 39686
rect 87456 39684 87512 39686
rect 87566 39372 87622 39408
rect 87566 39352 87568 39372
rect 87568 39352 87620 39372
rect 87620 39352 87622 39372
rect 86480 39194 86536 39196
rect 86560 39194 86616 39196
rect 86640 39194 86696 39196
rect 86720 39194 86776 39196
rect 86480 39142 86526 39194
rect 86526 39142 86536 39194
rect 86560 39142 86590 39194
rect 86590 39142 86602 39194
rect 86602 39142 86616 39194
rect 86640 39142 86654 39194
rect 86654 39142 86666 39194
rect 86666 39142 86696 39194
rect 86720 39142 86730 39194
rect 86730 39142 86776 39194
rect 86480 39140 86536 39142
rect 86560 39140 86616 39142
rect 86640 39140 86696 39142
rect 86720 39140 86776 39142
rect 88210 39080 88266 39136
rect 87216 38650 87272 38652
rect 87296 38650 87352 38652
rect 87376 38650 87432 38652
rect 87456 38650 87512 38652
rect 87216 38598 87262 38650
rect 87262 38598 87272 38650
rect 87296 38598 87326 38650
rect 87326 38598 87338 38650
rect 87338 38598 87352 38650
rect 87376 38598 87390 38650
rect 87390 38598 87402 38650
rect 87402 38598 87432 38650
rect 87456 38598 87466 38650
rect 87466 38598 87512 38650
rect 87216 38596 87272 38598
rect 87296 38596 87352 38598
rect 87376 38596 87432 38598
rect 87456 38596 87512 38598
rect 86480 38106 86536 38108
rect 86560 38106 86616 38108
rect 86640 38106 86696 38108
rect 86720 38106 86776 38108
rect 85818 37992 85874 38048
rect 86480 38054 86526 38106
rect 86526 38054 86536 38106
rect 86560 38054 86590 38106
rect 86590 38054 86602 38106
rect 86602 38054 86616 38106
rect 86640 38054 86654 38106
rect 86654 38054 86666 38106
rect 86666 38054 86696 38106
rect 86720 38054 86730 38106
rect 86730 38054 86776 38106
rect 86480 38052 86536 38054
rect 86560 38052 86616 38054
rect 86640 38052 86696 38054
rect 86720 38052 86776 38054
rect 88210 37756 88212 37776
rect 88212 37756 88264 37776
rect 88264 37756 88266 37776
rect 88210 37720 88266 37756
rect 87216 37562 87272 37564
rect 87296 37562 87352 37564
rect 87376 37562 87432 37564
rect 87456 37562 87512 37564
rect 87216 37510 87262 37562
rect 87262 37510 87272 37562
rect 87296 37510 87326 37562
rect 87326 37510 87338 37562
rect 87338 37510 87352 37562
rect 87376 37510 87390 37562
rect 87390 37510 87402 37562
rect 87402 37510 87432 37562
rect 87456 37510 87466 37562
rect 87466 37510 87512 37562
rect 87216 37508 87272 37510
rect 87296 37508 87352 37510
rect 87376 37508 87432 37510
rect 87456 37508 87512 37510
rect 85818 37040 85874 37096
rect 88210 37040 88266 37096
rect 86480 37018 86536 37020
rect 86560 37018 86616 37020
rect 86640 37018 86696 37020
rect 86720 37018 86776 37020
rect 86480 36966 86526 37018
rect 86526 36966 86536 37018
rect 86560 36966 86590 37018
rect 86590 36966 86602 37018
rect 86602 36966 86616 37018
rect 86640 36966 86654 37018
rect 86654 36966 86666 37018
rect 86666 36966 86696 37018
rect 86720 36966 86730 37018
rect 86730 36966 86776 37018
rect 86480 36964 86536 36966
rect 86560 36964 86616 36966
rect 86640 36964 86696 36966
rect 86720 36964 86776 36966
rect 87216 36474 87272 36476
rect 87296 36474 87352 36476
rect 87376 36474 87432 36476
rect 87456 36474 87512 36476
rect 87216 36422 87262 36474
rect 87262 36422 87272 36474
rect 87296 36422 87326 36474
rect 87326 36422 87338 36474
rect 87338 36422 87352 36474
rect 87376 36422 87390 36474
rect 87390 36422 87402 36474
rect 87402 36422 87432 36474
rect 87456 36422 87466 36474
rect 87466 36422 87512 36474
rect 87216 36420 87272 36422
rect 87296 36420 87352 36422
rect 87376 36420 87432 36422
rect 87456 36420 87512 36422
rect 86480 35930 86536 35932
rect 86560 35930 86616 35932
rect 86640 35930 86696 35932
rect 86720 35930 86776 35932
rect 86480 35878 86526 35930
rect 86526 35878 86536 35930
rect 86560 35878 86590 35930
rect 86590 35878 86602 35930
rect 86602 35878 86616 35930
rect 86640 35878 86654 35930
rect 86654 35878 86666 35930
rect 86666 35878 86696 35930
rect 86720 35878 86730 35930
rect 86730 35878 86776 35930
rect 86480 35876 86536 35878
rect 86560 35876 86616 35878
rect 86640 35876 86696 35878
rect 86720 35876 86776 35878
rect 88578 35680 88634 35736
rect 87216 35386 87272 35388
rect 87296 35386 87352 35388
rect 87376 35386 87432 35388
rect 87456 35386 87512 35388
rect 87216 35334 87262 35386
rect 87262 35334 87272 35386
rect 87296 35334 87326 35386
rect 87326 35334 87338 35386
rect 87338 35334 87352 35386
rect 87376 35334 87390 35386
rect 87390 35334 87402 35386
rect 87402 35334 87432 35386
rect 87456 35334 87466 35386
rect 87466 35334 87512 35386
rect 87216 35332 87272 35334
rect 87296 35332 87352 35334
rect 87376 35332 87432 35334
rect 87456 35332 87512 35334
rect 88210 35000 88266 35056
rect 85818 34864 85874 34920
rect 86480 34842 86536 34844
rect 86560 34842 86616 34844
rect 86640 34842 86696 34844
rect 86720 34842 86776 34844
rect 86480 34790 86526 34842
rect 86526 34790 86536 34842
rect 86560 34790 86590 34842
rect 86590 34790 86602 34842
rect 86602 34790 86616 34842
rect 86640 34790 86654 34842
rect 86654 34790 86666 34842
rect 86666 34790 86696 34842
rect 86720 34790 86730 34842
rect 86730 34790 86776 34842
rect 86480 34788 86536 34790
rect 86560 34788 86616 34790
rect 86640 34788 86696 34790
rect 86720 34788 86776 34790
rect 87216 34298 87272 34300
rect 87296 34298 87352 34300
rect 87376 34298 87432 34300
rect 87456 34298 87512 34300
rect 87216 34246 87262 34298
rect 87262 34246 87272 34298
rect 87296 34246 87326 34298
rect 87326 34246 87338 34298
rect 87338 34246 87352 34298
rect 87376 34246 87390 34298
rect 87390 34246 87402 34298
rect 87402 34246 87432 34298
rect 87456 34246 87466 34298
rect 87466 34246 87512 34298
rect 87216 34244 87272 34246
rect 87296 34244 87352 34246
rect 87376 34244 87432 34246
rect 87456 34244 87512 34246
rect 85818 33776 85874 33832
rect 86480 33754 86536 33756
rect 86560 33754 86616 33756
rect 86640 33754 86696 33756
rect 86720 33754 86776 33756
rect 86480 33702 86526 33754
rect 86526 33702 86536 33754
rect 86560 33702 86590 33754
rect 86590 33702 86602 33754
rect 86602 33702 86616 33754
rect 86640 33702 86654 33754
rect 86654 33702 86666 33754
rect 86666 33702 86696 33754
rect 86720 33702 86730 33754
rect 86730 33702 86776 33754
rect 86480 33700 86536 33702
rect 86560 33700 86616 33702
rect 86640 33700 86696 33702
rect 86720 33700 86776 33702
rect 88210 33640 88266 33696
rect 87216 33210 87272 33212
rect 87296 33210 87352 33212
rect 87376 33210 87432 33212
rect 87456 33210 87512 33212
rect 87216 33158 87262 33210
rect 87262 33158 87272 33210
rect 87296 33158 87326 33210
rect 87326 33158 87338 33210
rect 87338 33158 87352 33210
rect 87376 33158 87390 33210
rect 87390 33158 87402 33210
rect 87402 33158 87432 33210
rect 87456 33158 87466 33210
rect 87466 33158 87512 33210
rect 87216 33156 87272 33158
rect 87296 33156 87352 33158
rect 87376 33156 87432 33158
rect 87456 33156 87512 33158
rect 86480 32666 86536 32668
rect 86560 32666 86616 32668
rect 86640 32666 86696 32668
rect 86720 32666 86776 32668
rect 85818 32552 85874 32608
rect 86480 32614 86526 32666
rect 86526 32614 86536 32666
rect 86560 32614 86590 32666
rect 86590 32614 86602 32666
rect 86602 32614 86616 32666
rect 86640 32614 86654 32666
rect 86654 32614 86666 32666
rect 86666 32614 86696 32666
rect 86720 32614 86730 32666
rect 86730 32614 86776 32666
rect 86480 32612 86536 32614
rect 86560 32612 86616 32614
rect 86640 32612 86696 32614
rect 86720 32612 86776 32614
rect 88210 32316 88212 32336
rect 88212 32316 88264 32336
rect 88264 32316 88266 32336
rect 88210 32280 88266 32316
rect 87216 32122 87272 32124
rect 87296 32122 87352 32124
rect 87376 32122 87432 32124
rect 87456 32122 87512 32124
rect 87216 32070 87262 32122
rect 87262 32070 87272 32122
rect 87296 32070 87326 32122
rect 87326 32070 87338 32122
rect 87338 32070 87352 32122
rect 87376 32070 87390 32122
rect 87390 32070 87402 32122
rect 87402 32070 87432 32122
rect 87456 32070 87466 32122
rect 87466 32070 87512 32122
rect 87216 32068 87272 32070
rect 87296 32068 87352 32070
rect 87376 32068 87432 32070
rect 87456 32068 87512 32070
rect 85818 31600 85874 31656
rect 88210 31600 88266 31656
rect 86480 31578 86536 31580
rect 86560 31578 86616 31580
rect 86640 31578 86696 31580
rect 86720 31578 86776 31580
rect 86480 31526 86526 31578
rect 86526 31526 86536 31578
rect 86560 31526 86590 31578
rect 86590 31526 86602 31578
rect 86602 31526 86616 31578
rect 86640 31526 86654 31578
rect 86654 31526 86666 31578
rect 86666 31526 86696 31578
rect 86720 31526 86730 31578
rect 86730 31526 86776 31578
rect 86480 31524 86536 31526
rect 86560 31524 86616 31526
rect 86640 31524 86696 31526
rect 86720 31524 86776 31526
rect 87216 31034 87272 31036
rect 87296 31034 87352 31036
rect 87376 31034 87432 31036
rect 87456 31034 87512 31036
rect 87216 30982 87262 31034
rect 87262 30982 87272 31034
rect 87296 30982 87326 31034
rect 87326 30982 87338 31034
rect 87338 30982 87352 31034
rect 87376 30982 87390 31034
rect 87390 30982 87402 31034
rect 87402 30982 87432 31034
rect 87456 30982 87466 31034
rect 87466 30982 87512 31034
rect 87216 30980 87272 30982
rect 87296 30980 87352 30982
rect 87376 30980 87432 30982
rect 87456 30980 87512 30982
rect 86480 30490 86536 30492
rect 86560 30490 86616 30492
rect 86640 30490 86696 30492
rect 86720 30490 86776 30492
rect 86480 30438 86526 30490
rect 86526 30438 86536 30490
rect 86560 30438 86590 30490
rect 86590 30438 86602 30490
rect 86602 30438 86616 30490
rect 86640 30438 86654 30490
rect 86654 30438 86666 30490
rect 86666 30438 86696 30490
rect 86720 30438 86730 30490
rect 86730 30438 86776 30490
rect 86480 30436 86536 30438
rect 86560 30436 86616 30438
rect 86640 30436 86696 30438
rect 86720 30436 86776 30438
rect 88578 30240 88634 30296
rect 87216 29946 87272 29948
rect 87296 29946 87352 29948
rect 87376 29946 87432 29948
rect 87456 29946 87512 29948
rect 87216 29894 87262 29946
rect 87262 29894 87272 29946
rect 87296 29894 87326 29946
rect 87326 29894 87338 29946
rect 87338 29894 87352 29946
rect 87376 29894 87390 29946
rect 87390 29894 87402 29946
rect 87402 29894 87432 29946
rect 87456 29894 87466 29946
rect 87466 29894 87512 29946
rect 87216 29892 87272 29894
rect 87296 29892 87352 29894
rect 87376 29892 87432 29894
rect 87456 29892 87512 29894
rect 88394 29560 88450 29616
rect 85818 29424 85874 29480
rect 86480 29402 86536 29404
rect 86560 29402 86616 29404
rect 86640 29402 86696 29404
rect 86720 29402 86776 29404
rect 86480 29350 86526 29402
rect 86526 29350 86536 29402
rect 86560 29350 86590 29402
rect 86590 29350 86602 29402
rect 86602 29350 86616 29402
rect 86640 29350 86654 29402
rect 86654 29350 86666 29402
rect 86666 29350 86696 29402
rect 86720 29350 86730 29402
rect 86730 29350 86776 29402
rect 86480 29348 86536 29350
rect 86560 29348 86616 29350
rect 86640 29348 86696 29350
rect 86720 29348 86776 29350
rect 87216 28858 87272 28860
rect 87296 28858 87352 28860
rect 87376 28858 87432 28860
rect 87456 28858 87512 28860
rect 87216 28806 87262 28858
rect 87262 28806 87272 28858
rect 87296 28806 87326 28858
rect 87326 28806 87338 28858
rect 87338 28806 87352 28858
rect 87376 28806 87390 28858
rect 87390 28806 87402 28858
rect 87402 28806 87432 28858
rect 87456 28806 87466 28858
rect 87466 28806 87512 28858
rect 87216 28804 87272 28806
rect 87296 28804 87352 28806
rect 87376 28804 87432 28806
rect 87456 28804 87512 28806
rect 85818 28336 85874 28392
rect 86480 28314 86536 28316
rect 86560 28314 86616 28316
rect 86640 28314 86696 28316
rect 86720 28314 86776 28316
rect 86480 28262 86526 28314
rect 86526 28262 86536 28314
rect 86560 28262 86590 28314
rect 86590 28262 86602 28314
rect 86602 28262 86616 28314
rect 86640 28262 86654 28314
rect 86654 28262 86666 28314
rect 86666 28262 86696 28314
rect 86720 28262 86730 28314
rect 86730 28262 86776 28314
rect 86480 28260 86536 28262
rect 86560 28260 86616 28262
rect 86640 28260 86696 28262
rect 86720 28260 86776 28262
rect 88210 28200 88266 28256
rect 87216 27770 87272 27772
rect 87296 27770 87352 27772
rect 87376 27770 87432 27772
rect 87456 27770 87512 27772
rect 87216 27718 87262 27770
rect 87262 27718 87272 27770
rect 87296 27718 87326 27770
rect 87326 27718 87338 27770
rect 87338 27718 87352 27770
rect 87376 27718 87390 27770
rect 87390 27718 87402 27770
rect 87402 27718 87432 27770
rect 87456 27718 87466 27770
rect 87466 27718 87512 27770
rect 87216 27716 87272 27718
rect 87296 27716 87352 27718
rect 87376 27716 87432 27718
rect 87456 27716 87512 27718
rect 86480 27226 86536 27228
rect 86560 27226 86616 27228
rect 86640 27226 86696 27228
rect 86720 27226 86776 27228
rect 85818 27112 85874 27168
rect 86480 27174 86526 27226
rect 86526 27174 86536 27226
rect 86560 27174 86590 27226
rect 86590 27174 86602 27226
rect 86602 27174 86616 27226
rect 86640 27174 86654 27226
rect 86654 27174 86666 27226
rect 86666 27174 86696 27226
rect 86720 27174 86730 27226
rect 86730 27174 86776 27226
rect 86480 27172 86536 27174
rect 86560 27172 86616 27174
rect 86640 27172 86696 27174
rect 86720 27172 86776 27174
rect 88394 26840 88450 26896
rect 87216 26682 87272 26684
rect 87296 26682 87352 26684
rect 87376 26682 87432 26684
rect 87456 26682 87512 26684
rect 87216 26630 87262 26682
rect 87262 26630 87272 26682
rect 87296 26630 87326 26682
rect 87326 26630 87338 26682
rect 87338 26630 87352 26682
rect 87376 26630 87390 26682
rect 87390 26630 87402 26682
rect 87402 26630 87432 26682
rect 87456 26630 87466 26682
rect 87466 26630 87512 26682
rect 87216 26628 87272 26630
rect 87296 26628 87352 26630
rect 87376 26628 87432 26630
rect 87456 26628 87512 26630
rect 87566 26296 87622 26352
rect 88210 26196 88212 26216
rect 88212 26196 88264 26216
rect 88264 26196 88266 26216
rect 88210 26160 88266 26196
rect 86480 26138 86536 26140
rect 86560 26138 86616 26140
rect 86640 26138 86696 26140
rect 86720 26138 86776 26140
rect 86480 26086 86526 26138
rect 86526 26086 86536 26138
rect 86560 26086 86590 26138
rect 86590 26086 86602 26138
rect 86602 26086 86616 26138
rect 86640 26086 86654 26138
rect 86654 26086 86666 26138
rect 86666 26086 86696 26138
rect 86720 26086 86730 26138
rect 86730 26086 86776 26138
rect 86480 26084 86536 26086
rect 86560 26084 86616 26086
rect 86640 26084 86696 26086
rect 86720 26084 86776 26086
rect 87216 25594 87272 25596
rect 87296 25594 87352 25596
rect 87376 25594 87432 25596
rect 87456 25594 87512 25596
rect 87216 25542 87262 25594
rect 87262 25542 87272 25594
rect 87296 25542 87326 25594
rect 87326 25542 87338 25594
rect 87338 25542 87352 25594
rect 87376 25542 87390 25594
rect 87390 25542 87402 25594
rect 87402 25542 87432 25594
rect 87456 25542 87466 25594
rect 87466 25542 87512 25594
rect 87216 25540 87272 25542
rect 87296 25540 87352 25542
rect 87376 25540 87432 25542
rect 87456 25540 87512 25542
rect 86480 25050 86536 25052
rect 86560 25050 86616 25052
rect 86640 25050 86696 25052
rect 86720 25050 86776 25052
rect 86480 24998 86526 25050
rect 86526 24998 86536 25050
rect 86560 24998 86590 25050
rect 86590 24998 86602 25050
rect 86602 24998 86616 25050
rect 86640 24998 86654 25050
rect 86654 24998 86666 25050
rect 86666 24998 86696 25050
rect 86720 24998 86730 25050
rect 86730 24998 86776 25050
rect 86480 24996 86536 24998
rect 86560 24996 86616 24998
rect 86640 24996 86696 24998
rect 86720 24996 86776 24998
rect 88578 24800 88634 24856
rect 87216 24506 87272 24508
rect 87296 24506 87352 24508
rect 87376 24506 87432 24508
rect 87456 24506 87512 24508
rect 87216 24454 87262 24506
rect 87262 24454 87272 24506
rect 87296 24454 87326 24506
rect 87326 24454 87338 24506
rect 87338 24454 87352 24506
rect 87376 24454 87390 24506
rect 87390 24454 87402 24506
rect 87402 24454 87432 24506
rect 87456 24454 87466 24506
rect 87466 24454 87512 24506
rect 87216 24452 87272 24454
rect 87296 24452 87352 24454
rect 87376 24452 87432 24454
rect 87456 24452 87512 24454
rect 87566 24120 87622 24176
rect 88486 24140 88542 24176
rect 88486 24120 88488 24140
rect 88488 24120 88540 24140
rect 88540 24120 88542 24140
rect 86480 23962 86536 23964
rect 86560 23962 86616 23964
rect 86640 23962 86696 23964
rect 86720 23962 86776 23964
rect 86480 23910 86526 23962
rect 86526 23910 86536 23962
rect 86560 23910 86590 23962
rect 86590 23910 86602 23962
rect 86602 23910 86616 23962
rect 86640 23910 86654 23962
rect 86654 23910 86666 23962
rect 86666 23910 86696 23962
rect 86720 23910 86730 23962
rect 86730 23910 86776 23962
rect 86480 23908 86536 23910
rect 86560 23908 86616 23910
rect 86640 23908 86696 23910
rect 86720 23908 86776 23910
rect 87216 23418 87272 23420
rect 87296 23418 87352 23420
rect 87376 23418 87432 23420
rect 87456 23418 87512 23420
rect 87216 23366 87262 23418
rect 87262 23366 87272 23418
rect 87296 23366 87326 23418
rect 87326 23366 87338 23418
rect 87338 23366 87352 23418
rect 87376 23366 87390 23418
rect 87390 23366 87402 23418
rect 87402 23366 87432 23418
rect 87456 23366 87466 23418
rect 87466 23366 87512 23418
rect 87216 23364 87272 23366
rect 87296 23364 87352 23366
rect 87376 23364 87432 23366
rect 87456 23364 87512 23366
rect 85818 22896 85874 22952
rect 86480 22874 86536 22876
rect 86560 22874 86616 22876
rect 86640 22874 86696 22876
rect 86720 22874 86776 22876
rect 86480 22822 86526 22874
rect 86526 22822 86536 22874
rect 86560 22822 86590 22874
rect 86590 22822 86602 22874
rect 86602 22822 86616 22874
rect 86640 22822 86654 22874
rect 86654 22822 86666 22874
rect 86666 22822 86696 22874
rect 86720 22822 86730 22874
rect 86730 22822 86776 22874
rect 86480 22820 86536 22822
rect 86560 22820 86616 22822
rect 86640 22820 86696 22822
rect 86720 22820 86776 22822
rect 88210 22760 88266 22816
rect 87216 22330 87272 22332
rect 87296 22330 87352 22332
rect 87376 22330 87432 22332
rect 87456 22330 87512 22332
rect 87216 22278 87262 22330
rect 87262 22278 87272 22330
rect 87296 22278 87326 22330
rect 87326 22278 87338 22330
rect 87338 22278 87352 22330
rect 87376 22278 87390 22330
rect 87390 22278 87402 22330
rect 87402 22278 87432 22330
rect 87456 22278 87466 22330
rect 87466 22278 87512 22330
rect 87216 22276 87272 22278
rect 87296 22276 87352 22278
rect 87376 22276 87432 22278
rect 87456 22276 87512 22278
rect 86480 21786 86536 21788
rect 86560 21786 86616 21788
rect 86640 21786 86696 21788
rect 86720 21786 86776 21788
rect 85818 21672 85874 21728
rect 86480 21734 86526 21786
rect 86526 21734 86536 21786
rect 86560 21734 86590 21786
rect 86590 21734 86602 21786
rect 86602 21734 86616 21786
rect 86640 21734 86654 21786
rect 86654 21734 86666 21786
rect 86666 21734 86696 21786
rect 86720 21734 86730 21786
rect 86730 21734 86776 21786
rect 86480 21732 86536 21734
rect 86560 21732 86616 21734
rect 86640 21732 86696 21734
rect 86720 21732 86776 21734
rect 88394 21400 88450 21456
rect 87216 21242 87272 21244
rect 87296 21242 87352 21244
rect 87376 21242 87432 21244
rect 87456 21242 87512 21244
rect 87216 21190 87262 21242
rect 87262 21190 87272 21242
rect 87296 21190 87326 21242
rect 87326 21190 87338 21242
rect 87338 21190 87352 21242
rect 87376 21190 87390 21242
rect 87390 21190 87402 21242
rect 87402 21190 87432 21242
rect 87456 21190 87466 21242
rect 87466 21190 87512 21242
rect 87216 21188 87272 21190
rect 87296 21188 87352 21190
rect 87376 21188 87432 21190
rect 87456 21188 87512 21190
rect 88578 20720 88634 20776
rect 86480 20698 86536 20700
rect 86560 20698 86616 20700
rect 86640 20698 86696 20700
rect 86720 20698 86776 20700
rect 86480 20646 86526 20698
rect 86526 20646 86536 20698
rect 86560 20646 86590 20698
rect 86590 20646 86602 20698
rect 86602 20646 86616 20698
rect 86640 20646 86654 20698
rect 86654 20646 86666 20698
rect 86666 20646 86696 20698
rect 86720 20646 86730 20698
rect 86730 20646 86776 20698
rect 86480 20644 86536 20646
rect 86560 20644 86616 20646
rect 86640 20644 86696 20646
rect 86720 20644 86776 20646
rect 87216 20154 87272 20156
rect 87296 20154 87352 20156
rect 87376 20154 87432 20156
rect 87456 20154 87512 20156
rect 87216 20102 87262 20154
rect 87262 20102 87272 20154
rect 87296 20102 87326 20154
rect 87326 20102 87338 20154
rect 87338 20102 87352 20154
rect 87376 20102 87390 20154
rect 87390 20102 87402 20154
rect 87402 20102 87432 20154
rect 87456 20102 87466 20154
rect 87466 20102 87512 20154
rect 87216 20100 87272 20102
rect 87296 20100 87352 20102
rect 87376 20100 87432 20102
rect 87456 20100 87512 20102
rect 87566 19768 87622 19824
rect 86480 19610 86536 19612
rect 86560 19610 86616 19612
rect 86640 19610 86696 19612
rect 86720 19610 86776 19612
rect 86480 19558 86526 19610
rect 86526 19558 86536 19610
rect 86560 19558 86590 19610
rect 86590 19558 86602 19610
rect 86602 19558 86616 19610
rect 86640 19558 86654 19610
rect 86654 19558 86666 19610
rect 86666 19558 86696 19610
rect 86720 19558 86730 19610
rect 86730 19558 86776 19610
rect 86480 19556 86536 19558
rect 86560 19556 86616 19558
rect 86640 19556 86696 19558
rect 86720 19556 86776 19558
rect 88670 19360 88726 19416
rect 87216 19066 87272 19068
rect 87296 19066 87352 19068
rect 87376 19066 87432 19068
rect 87456 19066 87512 19068
rect 87216 19014 87262 19066
rect 87262 19014 87272 19066
rect 87296 19014 87326 19066
rect 87326 19014 87338 19066
rect 87338 19014 87352 19066
rect 87376 19014 87390 19066
rect 87390 19014 87402 19066
rect 87402 19014 87432 19066
rect 87456 19014 87466 19066
rect 87466 19014 87512 19066
rect 87216 19012 87272 19014
rect 87296 19012 87352 19014
rect 87376 19012 87432 19014
rect 87456 19012 87512 19014
rect 87290 18680 87346 18736
rect 88210 18700 88266 18736
rect 88210 18680 88212 18700
rect 88212 18680 88264 18700
rect 88264 18680 88266 18700
rect 86480 18522 86536 18524
rect 86560 18522 86616 18524
rect 86640 18522 86696 18524
rect 86720 18522 86776 18524
rect 86480 18470 86526 18522
rect 86526 18470 86536 18522
rect 86560 18470 86590 18522
rect 86590 18470 86602 18522
rect 86602 18470 86616 18522
rect 86640 18470 86654 18522
rect 86654 18470 86666 18522
rect 86666 18470 86696 18522
rect 86720 18470 86730 18522
rect 86730 18470 86776 18522
rect 86480 18468 86536 18470
rect 86560 18468 86616 18470
rect 86640 18468 86696 18470
rect 86720 18468 86776 18470
rect 87216 17978 87272 17980
rect 87296 17978 87352 17980
rect 87376 17978 87432 17980
rect 87456 17978 87512 17980
rect 87216 17926 87262 17978
rect 87262 17926 87272 17978
rect 87296 17926 87326 17978
rect 87326 17926 87338 17978
rect 87338 17926 87352 17978
rect 87376 17926 87390 17978
rect 87390 17926 87402 17978
rect 87402 17926 87432 17978
rect 87456 17926 87466 17978
rect 87466 17926 87512 17978
rect 87216 17924 87272 17926
rect 87296 17924 87352 17926
rect 87376 17924 87432 17926
rect 87456 17924 87512 17926
rect 85818 17456 85874 17512
rect 86480 17434 86536 17436
rect 86560 17434 86616 17436
rect 86640 17434 86696 17436
rect 86720 17434 86776 17436
rect 86480 17382 86526 17434
rect 86526 17382 86536 17434
rect 86560 17382 86590 17434
rect 86590 17382 86602 17434
rect 86602 17382 86616 17434
rect 86640 17382 86654 17434
rect 86654 17382 86666 17434
rect 86666 17382 86696 17434
rect 86720 17382 86730 17434
rect 86730 17382 86776 17434
rect 86480 17380 86536 17382
rect 86560 17380 86616 17382
rect 86640 17380 86696 17382
rect 86720 17380 86776 17382
rect 88210 17320 88266 17376
rect 87216 16890 87272 16892
rect 87296 16890 87352 16892
rect 87376 16890 87432 16892
rect 87456 16890 87512 16892
rect 87216 16838 87262 16890
rect 87262 16838 87272 16890
rect 87296 16838 87326 16890
rect 87326 16838 87338 16890
rect 87338 16838 87352 16890
rect 87376 16838 87390 16890
rect 87390 16838 87402 16890
rect 87402 16838 87432 16890
rect 87456 16838 87466 16890
rect 87466 16838 87512 16890
rect 87216 16836 87272 16838
rect 87296 16836 87352 16838
rect 87376 16836 87432 16838
rect 87456 16836 87512 16838
rect 86480 16346 86536 16348
rect 86560 16346 86616 16348
rect 86640 16346 86696 16348
rect 86720 16346 86776 16348
rect 85818 16232 85874 16288
rect 86480 16294 86526 16346
rect 86526 16294 86536 16346
rect 86560 16294 86590 16346
rect 86590 16294 86602 16346
rect 86602 16294 86616 16346
rect 86640 16294 86654 16346
rect 86654 16294 86666 16346
rect 86666 16294 86696 16346
rect 86720 16294 86730 16346
rect 86730 16294 86776 16346
rect 86480 16292 86536 16294
rect 86560 16292 86616 16294
rect 86640 16292 86696 16294
rect 86720 16292 86776 16294
rect 88210 15960 88266 16016
rect 87216 15802 87272 15804
rect 87296 15802 87352 15804
rect 87376 15802 87432 15804
rect 87456 15802 87512 15804
rect 87216 15750 87262 15802
rect 87262 15750 87272 15802
rect 87296 15750 87326 15802
rect 87326 15750 87338 15802
rect 87338 15750 87352 15802
rect 87376 15750 87390 15802
rect 87390 15750 87402 15802
rect 87402 15750 87432 15802
rect 87456 15750 87466 15802
rect 87466 15750 87512 15802
rect 87216 15748 87272 15750
rect 87296 15748 87352 15750
rect 87376 15748 87432 15750
rect 87456 15748 87512 15750
rect 88578 15280 88634 15336
rect 86480 15258 86536 15260
rect 86560 15258 86616 15260
rect 86640 15258 86696 15260
rect 86720 15258 86776 15260
rect 86480 15206 86526 15258
rect 86526 15206 86536 15258
rect 86560 15206 86590 15258
rect 86590 15206 86602 15258
rect 86602 15206 86616 15258
rect 86640 15206 86654 15258
rect 86654 15206 86666 15258
rect 86666 15206 86696 15258
rect 86720 15206 86730 15258
rect 86730 15206 86776 15258
rect 86480 15204 86536 15206
rect 86560 15204 86616 15206
rect 86640 15204 86696 15206
rect 86720 15204 86776 15206
rect 87216 14714 87272 14716
rect 87296 14714 87352 14716
rect 87376 14714 87432 14716
rect 87456 14714 87512 14716
rect 87216 14662 87262 14714
rect 87262 14662 87272 14714
rect 87296 14662 87326 14714
rect 87326 14662 87338 14714
rect 87338 14662 87352 14714
rect 87376 14662 87390 14714
rect 87390 14662 87402 14714
rect 87402 14662 87432 14714
rect 87456 14662 87466 14714
rect 87466 14662 87512 14714
rect 87216 14660 87272 14662
rect 87296 14660 87352 14662
rect 87376 14660 87432 14662
rect 87456 14660 87512 14662
rect 88026 14600 88082 14656
rect 86480 14170 86536 14172
rect 86560 14170 86616 14172
rect 86640 14170 86696 14172
rect 86720 14170 86776 14172
rect 86480 14118 86526 14170
rect 86526 14118 86536 14170
rect 86560 14118 86590 14170
rect 86590 14118 86602 14170
rect 86602 14118 86616 14170
rect 86640 14118 86654 14170
rect 86654 14118 86666 14170
rect 86666 14118 86696 14170
rect 86720 14118 86730 14170
rect 86730 14118 86776 14170
rect 86480 14116 86536 14118
rect 86560 14116 86616 14118
rect 86640 14116 86696 14118
rect 86720 14116 86776 14118
rect 87216 13626 87272 13628
rect 87296 13626 87352 13628
rect 87376 13626 87432 13628
rect 87456 13626 87512 13628
rect 87216 13574 87262 13626
rect 87262 13574 87272 13626
rect 87296 13574 87326 13626
rect 87326 13574 87338 13626
rect 87338 13574 87352 13626
rect 87376 13574 87390 13626
rect 87390 13574 87402 13626
rect 87402 13574 87432 13626
rect 87456 13574 87466 13626
rect 87466 13574 87512 13626
rect 87216 13572 87272 13574
rect 87296 13572 87352 13574
rect 87376 13572 87432 13574
rect 87456 13572 87512 13574
rect 86480 13082 86536 13084
rect 86560 13082 86616 13084
rect 86640 13082 86696 13084
rect 86720 13082 86776 13084
rect 86480 13030 86526 13082
rect 86526 13030 86536 13082
rect 86560 13030 86590 13082
rect 86590 13030 86602 13082
rect 86602 13030 86616 13082
rect 86640 13030 86654 13082
rect 86654 13030 86666 13082
rect 86666 13030 86696 13082
rect 86720 13030 86730 13082
rect 86730 13030 86776 13082
rect 86480 13028 86536 13030
rect 86560 13028 86616 13030
rect 86640 13028 86696 13030
rect 86720 13028 86776 13030
rect 88210 13240 88266 13296
rect 87216 12538 87272 12540
rect 87296 12538 87352 12540
rect 87376 12538 87432 12540
rect 87456 12538 87512 12540
rect 87216 12486 87262 12538
rect 87262 12486 87272 12538
rect 87296 12486 87326 12538
rect 87326 12486 87338 12538
rect 87338 12486 87352 12538
rect 87376 12486 87390 12538
rect 87390 12486 87402 12538
rect 87402 12486 87432 12538
rect 87456 12486 87466 12538
rect 87466 12486 87512 12538
rect 87216 12484 87272 12486
rect 87296 12484 87352 12486
rect 87376 12484 87432 12486
rect 87456 12484 87512 12486
rect 88578 12560 88634 12616
rect 83610 11948 83666 12004
rect 86480 11994 86536 11996
rect 86560 11994 86616 11996
rect 86640 11994 86696 11996
rect 86720 11994 86776 11996
rect 86480 11942 86526 11994
rect 86526 11942 86536 11994
rect 86560 11942 86590 11994
rect 86590 11942 86602 11994
rect 86602 11942 86616 11994
rect 86640 11942 86654 11994
rect 86654 11942 86666 11994
rect 86666 11942 86696 11994
rect 86720 11942 86730 11994
rect 86730 11942 86776 11994
rect 86480 11940 86536 11942
rect 86560 11940 86616 11942
rect 86640 11940 86696 11942
rect 86720 11940 86776 11942
rect 87216 11450 87272 11452
rect 87296 11450 87352 11452
rect 87376 11450 87432 11452
rect 87456 11450 87512 11452
rect 87216 11398 87262 11450
rect 87262 11398 87272 11450
rect 87296 11398 87326 11450
rect 87326 11398 87338 11450
rect 87338 11398 87352 11450
rect 87376 11398 87390 11450
rect 87390 11398 87402 11450
rect 87402 11398 87432 11450
rect 87456 11398 87466 11450
rect 87466 11398 87512 11450
rect 87216 11396 87272 11398
rect 87296 11396 87352 11398
rect 87376 11396 87432 11398
rect 87456 11396 87512 11398
rect 86480 10906 86536 10908
rect 86560 10906 86616 10908
rect 86640 10906 86696 10908
rect 86720 10906 86776 10908
rect 86480 10854 86526 10906
rect 86526 10854 86536 10906
rect 86560 10854 86590 10906
rect 86590 10854 86602 10906
rect 86602 10854 86616 10906
rect 86640 10854 86654 10906
rect 86654 10854 86666 10906
rect 86666 10854 86696 10906
rect 86720 10854 86730 10906
rect 86730 10854 86776 10906
rect 86480 10852 86536 10854
rect 86560 10852 86616 10854
rect 86640 10852 86696 10854
rect 86720 10852 86776 10854
rect 88210 10556 88212 10576
rect 88212 10556 88264 10576
rect 88264 10556 88266 10576
rect 88210 10520 88266 10556
rect 87216 10362 87272 10364
rect 87296 10362 87352 10364
rect 87376 10362 87432 10364
rect 87456 10362 87512 10364
rect 87216 10310 87262 10362
rect 87262 10310 87272 10362
rect 87296 10310 87326 10362
rect 87326 10310 87338 10362
rect 87338 10310 87352 10362
rect 87376 10310 87390 10362
rect 87390 10310 87402 10362
rect 87402 10310 87432 10362
rect 87456 10310 87466 10362
rect 87466 10310 87512 10362
rect 87216 10308 87272 10310
rect 87296 10308 87352 10310
rect 87376 10308 87432 10310
rect 87456 10308 87512 10310
rect 86480 9818 86536 9820
rect 86560 9818 86616 9820
rect 86640 9818 86696 9820
rect 86720 9818 86776 9820
rect 86480 9766 86526 9818
rect 86526 9766 86536 9818
rect 86560 9766 86590 9818
rect 86590 9766 86602 9818
rect 86602 9766 86616 9818
rect 86640 9766 86654 9818
rect 86654 9766 86666 9818
rect 86666 9766 86696 9818
rect 86720 9766 86730 9818
rect 86730 9766 86776 9818
rect 86480 9764 86536 9766
rect 86560 9764 86616 9766
rect 86640 9764 86696 9766
rect 86720 9764 86776 9766
rect 87216 9274 87272 9276
rect 87296 9274 87352 9276
rect 87376 9274 87432 9276
rect 87456 9274 87512 9276
rect 87216 9222 87262 9274
rect 87262 9222 87272 9274
rect 87296 9222 87326 9274
rect 87326 9222 87338 9274
rect 87338 9222 87352 9274
rect 87376 9222 87390 9274
rect 87390 9222 87402 9274
rect 87402 9222 87432 9274
rect 87456 9222 87466 9274
rect 87466 9222 87512 9274
rect 87216 9220 87272 9222
rect 87296 9220 87352 9222
rect 87376 9220 87432 9222
rect 87456 9220 87512 9222
rect 86480 8730 86536 8732
rect 86560 8730 86616 8732
rect 86640 8730 86696 8732
rect 86720 8730 86776 8732
rect 86480 8678 86526 8730
rect 86526 8678 86536 8730
rect 86560 8678 86590 8730
rect 86590 8678 86602 8730
rect 86602 8678 86616 8730
rect 86640 8678 86654 8730
rect 86654 8678 86666 8730
rect 86666 8678 86696 8730
rect 86720 8678 86730 8730
rect 86730 8678 86776 8730
rect 86480 8676 86536 8678
rect 86560 8676 86616 8678
rect 86640 8676 86696 8678
rect 86720 8676 86776 8678
rect 87216 8186 87272 8188
rect 87296 8186 87352 8188
rect 87376 8186 87432 8188
rect 87456 8186 87512 8188
rect 87216 8134 87262 8186
rect 87262 8134 87272 8186
rect 87296 8134 87326 8186
rect 87326 8134 87338 8186
rect 87338 8134 87352 8186
rect 87376 8134 87390 8186
rect 87390 8134 87402 8186
rect 87402 8134 87432 8186
rect 87456 8134 87466 8186
rect 87466 8134 87512 8186
rect 87216 8132 87272 8134
rect 87296 8132 87352 8134
rect 87376 8132 87432 8134
rect 87456 8132 87512 8134
rect 86480 7642 86536 7644
rect 86560 7642 86616 7644
rect 86640 7642 86696 7644
rect 86720 7642 86776 7644
rect 86480 7590 86526 7642
rect 86526 7590 86536 7642
rect 86560 7590 86590 7642
rect 86590 7590 86602 7642
rect 86602 7590 86616 7642
rect 86640 7590 86654 7642
rect 86654 7590 86666 7642
rect 86666 7590 86696 7642
rect 86720 7590 86730 7642
rect 86730 7590 86776 7642
rect 86480 7588 86536 7590
rect 86560 7588 86616 7590
rect 86640 7588 86696 7590
rect 86720 7588 86776 7590
rect 87216 7098 87272 7100
rect 87296 7098 87352 7100
rect 87376 7098 87432 7100
rect 87456 7098 87512 7100
rect 87216 7046 87262 7098
rect 87262 7046 87272 7098
rect 87296 7046 87326 7098
rect 87326 7046 87338 7098
rect 87338 7046 87352 7098
rect 87376 7046 87390 7098
rect 87390 7046 87402 7098
rect 87402 7046 87432 7098
rect 87456 7046 87466 7098
rect 87466 7046 87512 7098
rect 87216 7044 87272 7046
rect 87296 7044 87352 7046
rect 87376 7044 87432 7046
rect 87456 7044 87512 7046
rect 18388 4922 18444 4924
rect 18468 4922 18524 4924
rect 18548 4922 18604 4924
rect 18628 4922 18684 4924
rect 18388 4870 18434 4922
rect 18434 4870 18444 4922
rect 18468 4870 18498 4922
rect 18498 4870 18510 4922
rect 18510 4870 18524 4922
rect 18548 4870 18562 4922
rect 18562 4870 18574 4922
rect 18574 4870 18604 4922
rect 18628 4870 18638 4922
rect 18638 4870 18684 4922
rect 18388 4868 18444 4870
rect 18468 4868 18524 4870
rect 18548 4868 18604 4870
rect 18628 4868 18684 4870
rect 36788 4922 36844 4924
rect 36868 4922 36924 4924
rect 36948 4922 37004 4924
rect 37028 4922 37084 4924
rect 36788 4870 36834 4922
rect 36834 4870 36844 4922
rect 36868 4870 36898 4922
rect 36898 4870 36910 4922
rect 36910 4870 36924 4922
rect 36948 4870 36962 4922
rect 36962 4870 36974 4922
rect 36974 4870 37004 4922
rect 37028 4870 37038 4922
rect 37038 4870 37084 4922
rect 36788 4868 36844 4870
rect 36868 4868 36924 4870
rect 36948 4868 37004 4870
rect 37028 4868 37084 4870
rect 55188 4922 55244 4924
rect 55268 4922 55324 4924
rect 55348 4922 55404 4924
rect 55428 4922 55484 4924
rect 55188 4870 55234 4922
rect 55234 4870 55244 4922
rect 55268 4870 55298 4922
rect 55298 4870 55310 4922
rect 55310 4870 55324 4922
rect 55348 4870 55362 4922
rect 55362 4870 55374 4922
rect 55374 4870 55404 4922
rect 55428 4870 55438 4922
rect 55438 4870 55484 4922
rect 55188 4868 55244 4870
rect 55268 4868 55324 4870
rect 55348 4868 55404 4870
rect 55428 4868 55484 4870
rect 73588 4922 73644 4924
rect 73668 4922 73724 4924
rect 73748 4922 73804 4924
rect 73828 4922 73884 4924
rect 73588 4870 73634 4922
rect 73634 4870 73644 4922
rect 73668 4870 73698 4922
rect 73698 4870 73710 4922
rect 73710 4870 73724 4922
rect 73748 4870 73762 4922
rect 73762 4870 73774 4922
rect 73774 4870 73804 4922
rect 73828 4870 73838 4922
rect 73838 4870 73884 4922
rect 73588 4868 73644 4870
rect 73668 4868 73724 4870
rect 73748 4868 73804 4870
rect 73828 4868 73884 4870
<< metal3 >>
rect 18378 87616 18694 87617
rect 18378 87552 18384 87616
rect 18448 87552 18464 87616
rect 18528 87552 18544 87616
rect 18608 87552 18624 87616
rect 18688 87552 18694 87616
rect 18378 87551 18694 87552
rect 36778 87616 37094 87617
rect 36778 87552 36784 87616
rect 36848 87552 36864 87616
rect 36928 87552 36944 87616
rect 37008 87552 37024 87616
rect 37088 87552 37094 87616
rect 36778 87551 37094 87552
rect 55178 87616 55494 87617
rect 55178 87552 55184 87616
rect 55248 87552 55264 87616
rect 55328 87552 55344 87616
rect 55408 87552 55424 87616
rect 55488 87552 55494 87616
rect 55178 87551 55494 87552
rect 73578 87616 73894 87617
rect 73578 87552 73584 87616
rect 73648 87552 73664 87616
rect 73728 87552 73744 87616
rect 73808 87552 73824 87616
rect 73888 87552 73894 87616
rect 73578 87551 73894 87552
rect 17718 87072 18034 87073
rect 17718 87008 17724 87072
rect 17788 87008 17804 87072
rect 17868 87008 17884 87072
rect 17948 87008 17964 87072
rect 18028 87008 18034 87072
rect 17718 87007 18034 87008
rect 36118 87072 36434 87073
rect 36118 87008 36124 87072
rect 36188 87008 36204 87072
rect 36268 87008 36284 87072
rect 36348 87008 36364 87072
rect 36428 87008 36434 87072
rect 36118 87007 36434 87008
rect 54518 87072 54834 87073
rect 54518 87008 54524 87072
rect 54588 87008 54604 87072
rect 54668 87008 54684 87072
rect 54748 87008 54764 87072
rect 54828 87008 54834 87072
rect 54518 87007 54834 87008
rect 72918 87072 73234 87073
rect 72918 87008 72924 87072
rect 72988 87008 73004 87072
rect 73068 87008 73084 87072
rect 73148 87008 73164 87072
rect 73228 87008 73234 87072
rect 72918 87007 73234 87008
rect 18378 86528 18694 86529
rect 18378 86464 18384 86528
rect 18448 86464 18464 86528
rect 18528 86464 18544 86528
rect 18608 86464 18624 86528
rect 18688 86464 18694 86528
rect 18378 86463 18694 86464
rect 36778 86528 37094 86529
rect 36778 86464 36784 86528
rect 36848 86464 36864 86528
rect 36928 86464 36944 86528
rect 37008 86464 37024 86528
rect 37088 86464 37094 86528
rect 36778 86463 37094 86464
rect 55178 86528 55494 86529
rect 55178 86464 55184 86528
rect 55248 86464 55264 86528
rect 55328 86464 55344 86528
rect 55408 86464 55424 86528
rect 55488 86464 55494 86528
rect 55178 86463 55494 86464
rect 73578 86528 73894 86529
rect 73578 86464 73584 86528
rect 73648 86464 73664 86528
rect 73728 86464 73744 86528
rect 73808 86464 73824 86528
rect 73888 86464 73894 86528
rect 73578 86463 73894 86464
rect 17718 85984 18034 85985
rect 17718 85920 17724 85984
rect 17788 85920 17804 85984
rect 17868 85920 17884 85984
rect 17948 85920 17964 85984
rect 18028 85920 18034 85984
rect 17718 85919 18034 85920
rect 36118 85984 36434 85985
rect 36118 85920 36124 85984
rect 36188 85920 36204 85984
rect 36268 85920 36284 85984
rect 36348 85920 36364 85984
rect 36428 85920 36434 85984
rect 36118 85919 36434 85920
rect 54518 85984 54834 85985
rect 54518 85920 54524 85984
rect 54588 85920 54604 85984
rect 54668 85920 54684 85984
rect 54748 85920 54764 85984
rect 54828 85920 54834 85984
rect 54518 85919 54834 85920
rect 72918 85984 73234 85985
rect 72918 85920 72924 85984
rect 72988 85920 73004 85984
rect 73068 85920 73084 85984
rect 73148 85920 73164 85984
rect 73228 85920 73234 85984
rect 72918 85919 73234 85920
rect 18378 85440 18694 85441
rect 18378 85376 18384 85440
rect 18448 85376 18464 85440
rect 18528 85376 18544 85440
rect 18608 85376 18624 85440
rect 18688 85376 18694 85440
rect 18378 85375 18694 85376
rect 36778 85440 37094 85441
rect 36778 85376 36784 85440
rect 36848 85376 36864 85440
rect 36928 85376 36944 85440
rect 37008 85376 37024 85440
rect 37088 85376 37094 85440
rect 36778 85375 37094 85376
rect 55178 85440 55494 85441
rect 55178 85376 55184 85440
rect 55248 85376 55264 85440
rect 55328 85376 55344 85440
rect 55408 85376 55424 85440
rect 55488 85376 55494 85440
rect 55178 85375 55494 85376
rect 73578 85440 73894 85441
rect 73578 85376 73584 85440
rect 73648 85376 73664 85440
rect 73728 85376 73744 85440
rect 73808 85376 73824 85440
rect 73888 85376 73894 85440
rect 73578 85375 73894 85376
rect 5878 84896 6194 84897
rect 5878 84832 5884 84896
rect 5948 84832 5964 84896
rect 6028 84832 6044 84896
rect 6108 84832 6124 84896
rect 6188 84832 6194 84896
rect 5878 84831 6194 84832
rect 17718 84896 18034 84897
rect 17718 84832 17724 84896
rect 17788 84832 17804 84896
rect 17868 84832 17884 84896
rect 17948 84832 17964 84896
rect 18028 84832 18034 84896
rect 17718 84831 18034 84832
rect 36118 84896 36434 84897
rect 36118 84832 36124 84896
rect 36188 84832 36204 84896
rect 36268 84832 36284 84896
rect 36348 84832 36364 84896
rect 36428 84832 36434 84896
rect 36118 84831 36434 84832
rect 54518 84896 54834 84897
rect 54518 84832 54524 84896
rect 54588 84832 54604 84896
rect 54668 84832 54684 84896
rect 54748 84832 54764 84896
rect 54828 84832 54834 84896
rect 54518 84831 54834 84832
rect 72918 84896 73234 84897
rect 72918 84832 72924 84896
rect 72988 84832 73004 84896
rect 73068 84832 73084 84896
rect 73148 84832 73164 84896
rect 73228 84832 73234 84896
rect 72918 84831 73234 84832
rect 86470 84896 86786 84897
rect 86470 84832 86476 84896
rect 86540 84832 86556 84896
rect 86620 84832 86636 84896
rect 86700 84832 86716 84896
rect 86780 84832 86786 84896
rect 86470 84831 86786 84832
rect 6614 84352 6930 84353
rect 6614 84288 6620 84352
rect 6684 84288 6700 84352
rect 6764 84288 6780 84352
rect 6844 84288 6860 84352
rect 6924 84288 6930 84352
rect 6614 84287 6930 84288
rect 18378 84352 18694 84353
rect 18378 84288 18384 84352
rect 18448 84288 18464 84352
rect 18528 84288 18544 84352
rect 18608 84288 18624 84352
rect 18688 84288 18694 84352
rect 18378 84287 18694 84288
rect 36778 84352 37094 84353
rect 36778 84288 36784 84352
rect 36848 84288 36864 84352
rect 36928 84288 36944 84352
rect 37008 84288 37024 84352
rect 37088 84288 37094 84352
rect 36778 84287 37094 84288
rect 55178 84352 55494 84353
rect 55178 84288 55184 84352
rect 55248 84288 55264 84352
rect 55328 84288 55344 84352
rect 55408 84288 55424 84352
rect 55488 84288 55494 84352
rect 55178 84287 55494 84288
rect 73578 84352 73894 84353
rect 73578 84288 73584 84352
rect 73648 84288 73664 84352
rect 73728 84288 73744 84352
rect 73808 84288 73824 84352
rect 73888 84288 73894 84352
rect 73578 84287 73894 84288
rect 87206 84352 87522 84353
rect 87206 84288 87212 84352
rect 87276 84288 87292 84352
rect 87356 84288 87372 84352
rect 87436 84288 87452 84352
rect 87516 84288 87522 84352
rect 87206 84287 87522 84288
rect 5878 83808 6194 83809
rect 5878 83744 5884 83808
rect 5948 83744 5964 83808
rect 6028 83744 6044 83808
rect 6108 83744 6124 83808
rect 6188 83744 6194 83808
rect 5878 83743 6194 83744
rect 86470 83808 86786 83809
rect 86470 83744 86476 83808
rect 86540 83744 86556 83808
rect 86620 83744 86636 83808
rect 86700 83744 86716 83808
rect 86780 83744 86786 83808
rect 86470 83743 86786 83744
rect 6614 83264 6930 83265
rect 6614 83200 6620 83264
rect 6684 83200 6700 83264
rect 6764 83200 6780 83264
rect 6844 83200 6860 83264
rect 6924 83200 6930 83264
rect 6614 83199 6930 83200
rect 87206 83264 87522 83265
rect 87206 83200 87212 83264
rect 87276 83200 87292 83264
rect 87356 83200 87372 83264
rect 87436 83200 87452 83264
rect 87516 83200 87522 83264
rect 87206 83199 87522 83200
rect 5878 82720 6194 82721
rect 5878 82656 5884 82720
rect 5948 82656 5964 82720
rect 6028 82656 6044 82720
rect 6108 82656 6124 82720
rect 6188 82656 6194 82720
rect 5878 82655 6194 82656
rect 86470 82720 86786 82721
rect 86470 82656 86476 82720
rect 86540 82656 86556 82720
rect 86620 82656 86636 82720
rect 86700 82656 86716 82720
rect 86780 82656 86786 82720
rect 86470 82655 86786 82656
rect 6614 82176 6930 82177
rect 6614 82112 6620 82176
rect 6684 82112 6700 82176
rect 6764 82112 6780 82176
rect 6844 82112 6860 82176
rect 6924 82112 6930 82176
rect 6614 82111 6930 82112
rect 87206 82176 87522 82177
rect 87206 82112 87212 82176
rect 87276 82112 87292 82176
rect 87356 82112 87372 82176
rect 87436 82112 87452 82176
rect 87516 82112 87522 82176
rect 87206 82111 87522 82112
rect 47081 81706 47147 81709
rect 47955 81706 48021 81709
rect 47081 81704 48021 81706
rect 47081 81648 47086 81704
rect 47142 81648 47960 81704
rect 48016 81648 48021 81704
rect 47081 81646 48021 81648
rect 47081 81643 47147 81646
rect 47955 81643 48021 81646
rect 5878 81632 6194 81633
rect 5878 81568 5884 81632
rect 5948 81568 5964 81632
rect 6028 81568 6044 81632
rect 6108 81568 6124 81632
rect 6188 81568 6194 81632
rect 5878 81567 6194 81568
rect 86470 81632 86786 81633
rect 86470 81568 86476 81632
rect 86540 81568 86556 81632
rect 86620 81568 86636 81632
rect 86700 81568 86716 81632
rect 86780 81568 86786 81632
rect 86470 81567 86786 81568
rect 3000 81298 3800 81328
rect 4117 81298 4183 81301
rect 3000 81296 4183 81298
rect 3000 81240 4122 81296
rect 4178 81240 4183 81296
rect 3000 81238 4183 81240
rect 3000 81208 3800 81238
rect 4117 81235 4183 81238
rect 88205 81298 88271 81301
rect 89200 81298 90000 81328
rect 88205 81296 90000 81298
rect 88205 81240 88210 81296
rect 88266 81240 90000 81296
rect 88205 81238 90000 81240
rect 88205 81235 88271 81238
rect 89200 81208 90000 81238
rect 6614 81088 6930 81089
rect 6614 81024 6620 81088
rect 6684 81024 6700 81088
rect 6764 81024 6780 81088
rect 6844 81024 6860 81088
rect 6924 81024 6930 81088
rect 87206 81088 87522 81089
rect 6614 81023 6930 81024
rect 8533 81026 8599 81029
rect 84341 81026 84407 81029
rect 8533 81024 10084 81026
rect 8533 80968 8538 81024
rect 8594 80968 10084 81024
rect 8533 80966 10084 80968
rect 45596 80966 47436 81026
rect 83132 81024 84407 81026
rect 83132 80968 84346 81024
rect 84402 80968 84407 81024
rect 87206 81024 87212 81088
rect 87276 81024 87292 81088
rect 87356 81024 87372 81088
rect 87436 81024 87452 81088
rect 87516 81024 87522 81088
rect 87206 81023 87522 81024
rect 83132 80966 84407 80968
rect 8533 80963 8599 80966
rect 84341 80963 84407 80966
rect 5878 80544 6194 80545
rect 5878 80480 5884 80544
rect 5948 80480 5964 80544
rect 6028 80480 6044 80544
rect 6108 80480 6124 80544
rect 6188 80480 6194 80544
rect 5878 80479 6194 80480
rect 86470 80544 86786 80545
rect 86470 80480 86476 80544
rect 86540 80480 86556 80544
rect 86620 80480 86636 80544
rect 86700 80480 86716 80544
rect 86780 80480 86786 80544
rect 86470 80479 86786 80480
rect 6614 80000 6930 80001
rect 3000 79938 3800 79968
rect 4117 79938 4183 79941
rect 3000 79936 4183 79938
rect 3000 79880 4122 79936
rect 4178 79880 4183 79936
rect 6614 79936 6620 80000
rect 6684 79936 6700 80000
rect 6764 79936 6780 80000
rect 6844 79936 6860 80000
rect 6924 79936 6930 80000
rect 87206 80000 87522 80001
rect 6614 79935 6930 79936
rect 8533 79938 8599 79941
rect 85813 79938 85879 79941
rect 8533 79936 10084 79938
rect 3000 79878 4183 79880
rect 3000 79848 3800 79878
rect 4117 79875 4183 79878
rect 8533 79880 8538 79936
rect 8594 79880 10084 79936
rect 8533 79878 10084 79880
rect 45596 79878 47436 79938
rect 83132 79936 85879 79938
rect 83132 79880 85818 79936
rect 85874 79880 85879 79936
rect 87206 79936 87212 80000
rect 87276 79936 87292 80000
rect 87356 79936 87372 80000
rect 87436 79936 87452 80000
rect 87516 79936 87522 80000
rect 87206 79935 87522 79936
rect 88205 79938 88271 79941
rect 89200 79938 90000 79968
rect 88205 79936 90000 79938
rect 83132 79878 85879 79880
rect 8533 79875 8599 79878
rect 85813 79875 85879 79878
rect 88205 79880 88210 79936
rect 88266 79880 90000 79936
rect 88205 79878 90000 79880
rect 88205 79875 88271 79878
rect 89200 79848 90000 79878
rect 5878 79456 6194 79457
rect 5878 79392 5884 79456
rect 5948 79392 5964 79456
rect 6028 79392 6044 79456
rect 6108 79392 6124 79456
rect 6188 79392 6194 79456
rect 5878 79391 6194 79392
rect 86470 79456 86786 79457
rect 86470 79392 86476 79456
rect 86540 79392 86556 79456
rect 86620 79392 86636 79456
rect 86700 79392 86716 79456
rect 86780 79392 86786 79456
rect 86470 79391 86786 79392
rect 6614 78912 6930 78913
rect 6614 78848 6620 78912
rect 6684 78848 6700 78912
rect 6764 78848 6780 78912
rect 6844 78848 6860 78912
rect 6924 78848 6930 78912
rect 87206 78912 87522 78913
rect 6614 78847 6930 78848
rect 8533 78850 8599 78853
rect 85813 78850 85879 78853
rect 8533 78848 10084 78850
rect 8533 78792 8538 78848
rect 8594 78792 10084 78848
rect 8533 78790 10084 78792
rect 45596 78790 47436 78850
rect 83132 78848 85879 78850
rect 83132 78792 85818 78848
rect 85874 78792 85879 78848
rect 87206 78848 87212 78912
rect 87276 78848 87292 78912
rect 87356 78848 87372 78912
rect 87436 78848 87452 78912
rect 87516 78848 87522 78912
rect 87206 78847 87522 78848
rect 83132 78790 85879 78792
rect 8533 78787 8599 78790
rect 85813 78787 85879 78790
rect 3000 78578 3800 78608
rect 4117 78578 4183 78581
rect 3000 78576 4183 78578
rect 3000 78520 4122 78576
rect 4178 78520 4183 78576
rect 3000 78518 4183 78520
rect 3000 78488 3800 78518
rect 4117 78515 4183 78518
rect 88205 78578 88271 78581
rect 89200 78578 90000 78608
rect 88205 78576 90000 78578
rect 88205 78520 88210 78576
rect 88266 78520 90000 78576
rect 88205 78518 90000 78520
rect 88205 78515 88271 78518
rect 89200 78488 90000 78518
rect 5878 78368 6194 78369
rect 5878 78304 5884 78368
rect 5948 78304 5964 78368
rect 6028 78304 6044 78368
rect 6108 78304 6124 78368
rect 6188 78304 6194 78368
rect 5878 78303 6194 78304
rect 86470 78368 86786 78369
rect 86470 78304 86476 78368
rect 86540 78304 86556 78368
rect 86620 78304 86636 78368
rect 86700 78304 86716 78368
rect 86780 78304 86786 78368
rect 86470 78303 86786 78304
rect 3000 77898 3800 77928
rect 4117 77898 4183 77901
rect 3000 77896 4183 77898
rect 3000 77840 4122 77896
rect 4178 77840 4183 77896
rect 3000 77838 4183 77840
rect 3000 77808 3800 77838
rect 4117 77835 4183 77838
rect 88205 77898 88271 77901
rect 89200 77898 90000 77928
rect 88205 77896 90000 77898
rect 88205 77840 88210 77896
rect 88266 77840 90000 77896
rect 88205 77838 90000 77840
rect 88205 77835 88271 77838
rect 6614 77824 6930 77825
rect 6614 77760 6620 77824
rect 6684 77760 6700 77824
rect 6764 77760 6780 77824
rect 6844 77760 6860 77824
rect 6924 77760 6930 77824
rect 87206 77824 87522 77825
rect 6614 77759 6930 77760
rect 8533 77762 8599 77765
rect 85813 77762 85879 77765
rect 8533 77760 10084 77762
rect 8533 77704 8538 77760
rect 8594 77704 10084 77760
rect 8533 77702 10084 77704
rect 45596 77702 47436 77762
rect 83132 77760 85879 77762
rect 83132 77704 85818 77760
rect 85874 77704 85879 77760
rect 87206 77760 87212 77824
rect 87276 77760 87292 77824
rect 87356 77760 87372 77824
rect 87436 77760 87452 77824
rect 87516 77760 87522 77824
rect 89200 77808 90000 77838
rect 87206 77759 87522 77760
rect 83132 77702 85879 77704
rect 8533 77699 8599 77702
rect 85813 77699 85879 77702
rect 5878 77280 6194 77281
rect 5878 77216 5884 77280
rect 5948 77216 5964 77280
rect 6028 77216 6044 77280
rect 6108 77216 6124 77280
rect 6188 77216 6194 77280
rect 5878 77215 6194 77216
rect 86470 77280 86786 77281
rect 86470 77216 86476 77280
rect 86540 77216 86556 77280
rect 86620 77216 86636 77280
rect 86700 77216 86716 77280
rect 86780 77216 86786 77280
rect 86470 77215 86786 77216
rect 6614 76736 6930 76737
rect 6614 76672 6620 76736
rect 6684 76672 6700 76736
rect 6764 76672 6780 76736
rect 6844 76672 6860 76736
rect 6924 76672 6930 76736
rect 87206 76736 87522 76737
rect 6614 76671 6930 76672
rect 8533 76674 8599 76677
rect 85813 76674 85879 76677
rect 8533 76672 10084 76674
rect 8533 76616 8538 76672
rect 8594 76616 10084 76672
rect 8533 76614 10084 76616
rect 45596 76614 47436 76674
rect 83132 76672 85879 76674
rect 83132 76616 85818 76672
rect 85874 76616 85879 76672
rect 87206 76672 87212 76736
rect 87276 76672 87292 76736
rect 87356 76672 87372 76736
rect 87436 76672 87452 76736
rect 87516 76672 87522 76736
rect 87206 76671 87522 76672
rect 83132 76614 85879 76616
rect 8533 76611 8599 76614
rect 85813 76611 85879 76614
rect 3000 76538 3800 76568
rect 4209 76538 4275 76541
rect 3000 76536 4275 76538
rect 3000 76480 4214 76536
rect 4270 76480 4275 76536
rect 3000 76478 4275 76480
rect 3000 76448 3800 76478
rect 4209 76475 4275 76478
rect 88021 76538 88087 76541
rect 89200 76538 90000 76568
rect 88021 76536 90000 76538
rect 88021 76480 88026 76536
rect 88082 76480 90000 76536
rect 88021 76478 90000 76480
rect 88021 76475 88087 76478
rect 89200 76448 90000 76478
rect 5878 76192 6194 76193
rect 5878 76128 5884 76192
rect 5948 76128 5964 76192
rect 6028 76128 6044 76192
rect 6108 76128 6124 76192
rect 6188 76128 6194 76192
rect 5878 76127 6194 76128
rect 86470 76192 86786 76193
rect 86470 76128 86476 76192
rect 86540 76128 86556 76192
rect 86620 76128 86636 76192
rect 86700 76128 86716 76192
rect 86780 76128 86786 76192
rect 86470 76127 86786 76128
rect 3000 75858 3800 75888
rect 4117 75858 4183 75861
rect 3000 75856 4183 75858
rect 3000 75800 4122 75856
rect 4178 75800 4183 75856
rect 3000 75798 4183 75800
rect 3000 75768 3800 75798
rect 4117 75795 4183 75798
rect 88205 75858 88271 75861
rect 89200 75858 90000 75888
rect 88205 75856 90000 75858
rect 88205 75800 88210 75856
rect 88266 75800 90000 75856
rect 88205 75798 90000 75800
rect 88205 75795 88271 75798
rect 89200 75768 90000 75798
rect 6614 75648 6930 75649
rect 6614 75584 6620 75648
rect 6684 75584 6700 75648
rect 6764 75584 6780 75648
rect 6844 75584 6860 75648
rect 6924 75584 6930 75648
rect 87206 75648 87522 75649
rect 6614 75583 6930 75584
rect 8533 75586 8599 75589
rect 85813 75586 85879 75589
rect 8533 75584 10084 75586
rect 8533 75528 8538 75584
rect 8594 75528 10084 75584
rect 8533 75526 10084 75528
rect 45596 75526 47436 75586
rect 83132 75584 85879 75586
rect 83132 75528 85818 75584
rect 85874 75528 85879 75584
rect 87206 75584 87212 75648
rect 87276 75584 87292 75648
rect 87356 75584 87372 75648
rect 87436 75584 87452 75648
rect 87516 75584 87522 75648
rect 87206 75583 87522 75584
rect 83132 75526 85879 75528
rect 8533 75523 8599 75526
rect 85813 75523 85879 75526
rect 5878 75104 6194 75105
rect 5878 75040 5884 75104
rect 5948 75040 5964 75104
rect 6028 75040 6044 75104
rect 6108 75040 6124 75104
rect 6188 75040 6194 75104
rect 5878 75039 6194 75040
rect 86470 75104 86786 75105
rect 86470 75040 86476 75104
rect 86540 75040 86556 75104
rect 86620 75040 86636 75104
rect 86700 75040 86716 75104
rect 86780 75040 86786 75104
rect 86470 75039 86786 75040
rect 5405 74770 5471 74773
rect 5405 74768 10114 74770
rect 5405 74712 5410 74768
rect 5466 74712 10114 74768
rect 5405 74710 10114 74712
rect 5405 74707 5471 74710
rect 6614 74560 6930 74561
rect 3000 74498 3800 74528
rect 4117 74498 4183 74501
rect 3000 74496 4183 74498
rect 3000 74440 4122 74496
rect 4178 74440 4183 74496
rect 6614 74496 6620 74560
rect 6684 74496 6700 74560
rect 6764 74496 6780 74560
rect 6844 74496 6860 74560
rect 6924 74496 6930 74560
rect 6614 74495 6930 74496
rect 10054 74468 10114 74710
rect 87206 74560 87522 74561
rect 84525 74498 84591 74501
rect 3000 74438 4183 74440
rect 45596 74438 47436 74498
rect 83132 74496 84591 74498
rect 83132 74440 84530 74496
rect 84586 74440 84591 74496
rect 87206 74496 87212 74560
rect 87276 74496 87292 74560
rect 87356 74496 87372 74560
rect 87436 74496 87452 74560
rect 87516 74496 87522 74560
rect 87206 74495 87522 74496
rect 88573 74498 88639 74501
rect 89200 74498 90000 74528
rect 88573 74496 90000 74498
rect 83132 74438 84591 74440
rect 3000 74408 3800 74438
rect 4117 74435 4183 74438
rect 84525 74435 84591 74438
rect 88573 74440 88578 74496
rect 88634 74440 90000 74496
rect 88573 74438 90000 74440
rect 88573 74435 88639 74438
rect 89200 74408 90000 74438
rect 5878 74016 6194 74017
rect 5878 73952 5884 74016
rect 5948 73952 5964 74016
rect 6028 73952 6044 74016
rect 6108 73952 6124 74016
rect 6188 73952 6194 74016
rect 5878 73951 6194 73952
rect 86470 74016 86786 74017
rect 86470 73952 86476 74016
rect 86540 73952 86556 74016
rect 86620 73952 86636 74016
rect 86700 73952 86716 74016
rect 86780 73952 86786 74016
rect 86470 73951 86786 73952
rect 5405 73682 5471 73685
rect 5405 73680 10114 73682
rect 5405 73624 5410 73680
rect 5466 73624 10114 73680
rect 5405 73622 10114 73624
rect 5405 73619 5471 73622
rect 6614 73472 6930 73473
rect 6614 73408 6620 73472
rect 6684 73408 6700 73472
rect 6764 73408 6780 73472
rect 6844 73408 6860 73472
rect 6924 73408 6930 73472
rect 6614 73407 6930 73408
rect 10054 73380 10114 73622
rect 87206 73472 87522 73473
rect 84801 73410 84867 73413
rect 45596 73350 47436 73410
rect 83132 73408 84867 73410
rect 83132 73352 84806 73408
rect 84862 73352 84867 73408
rect 87206 73408 87212 73472
rect 87276 73408 87292 73472
rect 87356 73408 87372 73472
rect 87436 73408 87452 73472
rect 87516 73408 87522 73472
rect 87206 73407 87522 73408
rect 83132 73350 84867 73352
rect 84801 73347 84867 73350
rect 3000 73138 3800 73168
rect 4117 73138 4183 73141
rect 3000 73136 4183 73138
rect 3000 73080 4122 73136
rect 4178 73080 4183 73136
rect 3000 73078 4183 73080
rect 3000 73048 3800 73078
rect 4117 73075 4183 73078
rect 88205 73138 88271 73141
rect 89200 73138 90000 73168
rect 88205 73136 90000 73138
rect 88205 73080 88210 73136
rect 88266 73080 90000 73136
rect 88205 73078 90000 73080
rect 88205 73075 88271 73078
rect 89200 73048 90000 73078
rect 5878 72928 6194 72929
rect 5878 72864 5884 72928
rect 5948 72864 5964 72928
rect 6028 72864 6044 72928
rect 6108 72864 6124 72928
rect 6188 72864 6194 72928
rect 5878 72863 6194 72864
rect 86470 72928 86786 72929
rect 86470 72864 86476 72928
rect 86540 72864 86556 72928
rect 86620 72864 86636 72928
rect 86700 72864 86716 72928
rect 86780 72864 86786 72928
rect 86470 72863 86786 72864
rect 3000 72458 3800 72488
rect 4117 72458 4183 72461
rect 3000 72456 4183 72458
rect 3000 72400 4122 72456
rect 4178 72400 4183 72456
rect 3000 72398 4183 72400
rect 3000 72368 3800 72398
rect 4117 72395 4183 72398
rect 88205 72458 88271 72461
rect 89200 72458 90000 72488
rect 88205 72456 90000 72458
rect 88205 72400 88210 72456
rect 88266 72400 90000 72456
rect 88205 72398 90000 72400
rect 88205 72395 88271 72398
rect 6614 72384 6930 72385
rect 6614 72320 6620 72384
rect 6684 72320 6700 72384
rect 6764 72320 6780 72384
rect 6844 72320 6860 72384
rect 6924 72320 6930 72384
rect 87206 72384 87522 72385
rect 6614 72319 6930 72320
rect 8533 72322 8599 72325
rect 8533 72320 10084 72322
rect 8533 72264 8538 72320
rect 8594 72264 10084 72320
rect 8533 72262 10084 72264
rect 45596 72262 47436 72322
rect 83132 72262 84634 72322
rect 87206 72320 87212 72384
rect 87276 72320 87292 72384
rect 87356 72320 87372 72384
rect 87436 72320 87452 72384
rect 87516 72320 87522 72384
rect 89200 72368 90000 72398
rect 87206 72319 87522 72320
rect 8533 72259 8599 72262
rect 84574 72186 84634 72262
rect 87837 72186 87903 72189
rect 84574 72184 87903 72186
rect 84574 72128 87842 72184
rect 87898 72128 87903 72184
rect 84574 72126 87903 72128
rect 87837 72123 87903 72126
rect 5878 71840 6194 71841
rect 5878 71776 5884 71840
rect 5948 71776 5964 71840
rect 6028 71776 6044 71840
rect 6108 71776 6124 71840
rect 6188 71776 6194 71840
rect 5878 71775 6194 71776
rect 86470 71840 86786 71841
rect 86470 71776 86476 71840
rect 86540 71776 86556 71840
rect 86620 71776 86636 71840
rect 86700 71776 86716 71840
rect 86780 71776 86786 71840
rect 86470 71775 86786 71776
rect 6614 71296 6930 71297
rect 6614 71232 6620 71296
rect 6684 71232 6700 71296
rect 6764 71232 6780 71296
rect 6844 71232 6860 71296
rect 6924 71232 6930 71296
rect 87206 71296 87522 71297
rect 6614 71231 6930 71232
rect 8533 71234 8599 71237
rect 85813 71234 85879 71237
rect 8533 71232 10084 71234
rect 8533 71176 8538 71232
rect 8594 71176 10084 71232
rect 8533 71174 10084 71176
rect 45596 71174 47436 71234
rect 83132 71232 85879 71234
rect 83132 71176 85818 71232
rect 85874 71176 85879 71232
rect 87206 71232 87212 71296
rect 87276 71232 87292 71296
rect 87356 71232 87372 71296
rect 87436 71232 87452 71296
rect 87516 71232 87522 71296
rect 87206 71231 87522 71232
rect 83132 71174 85879 71176
rect 8533 71171 8599 71174
rect 85813 71171 85879 71174
rect 3000 71098 3800 71128
rect 4209 71098 4275 71101
rect 3000 71096 4275 71098
rect 3000 71040 4214 71096
rect 4270 71040 4275 71096
rect 3000 71038 4275 71040
rect 3000 71008 3800 71038
rect 4209 71035 4275 71038
rect 88205 71098 88271 71101
rect 89200 71098 90000 71128
rect 88205 71096 90000 71098
rect 88205 71040 88210 71096
rect 88266 71040 90000 71096
rect 88205 71038 90000 71040
rect 88205 71035 88271 71038
rect 89200 71008 90000 71038
rect 5878 70752 6194 70753
rect 5878 70688 5884 70752
rect 5948 70688 5964 70752
rect 6028 70688 6044 70752
rect 6108 70688 6124 70752
rect 6188 70688 6194 70752
rect 5878 70687 6194 70688
rect 86470 70752 86786 70753
rect 86470 70688 86476 70752
rect 86540 70688 86556 70752
rect 86620 70688 86636 70752
rect 86700 70688 86716 70752
rect 86780 70688 86786 70752
rect 86470 70687 86786 70688
rect 3000 70418 3800 70448
rect 4117 70418 4183 70421
rect 3000 70416 4183 70418
rect 3000 70360 4122 70416
rect 4178 70360 4183 70416
rect 3000 70358 4183 70360
rect 3000 70328 3800 70358
rect 4117 70355 4183 70358
rect 88205 70418 88271 70421
rect 89200 70418 90000 70448
rect 88205 70416 90000 70418
rect 88205 70360 88210 70416
rect 88266 70360 90000 70416
rect 88205 70358 90000 70360
rect 88205 70355 88271 70358
rect 89200 70328 90000 70358
rect 6614 70208 6930 70209
rect 6614 70144 6620 70208
rect 6684 70144 6700 70208
rect 6764 70144 6780 70208
rect 6844 70144 6860 70208
rect 6924 70144 6930 70208
rect 87206 70208 87522 70209
rect 6614 70143 6930 70144
rect 8533 70146 8599 70149
rect 85813 70146 85879 70149
rect 8533 70144 10084 70146
rect 8533 70088 8538 70144
rect 8594 70088 10084 70144
rect 8533 70086 10084 70088
rect 45596 70086 47436 70146
rect 83132 70144 85879 70146
rect 83132 70088 85818 70144
rect 85874 70088 85879 70144
rect 87206 70144 87212 70208
rect 87276 70144 87292 70208
rect 87356 70144 87372 70208
rect 87436 70144 87452 70208
rect 87516 70144 87522 70208
rect 87206 70143 87522 70144
rect 83132 70086 85879 70088
rect 8533 70083 8599 70086
rect 85813 70083 85879 70086
rect 5878 69664 6194 69665
rect 5878 69600 5884 69664
rect 5948 69600 5964 69664
rect 6028 69600 6044 69664
rect 6108 69600 6124 69664
rect 6188 69600 6194 69664
rect 5878 69599 6194 69600
rect 86470 69664 86786 69665
rect 86470 69600 86476 69664
rect 86540 69600 86556 69664
rect 86620 69600 86636 69664
rect 86700 69600 86716 69664
rect 86780 69600 86786 69664
rect 86470 69599 86786 69600
rect 6614 69120 6930 69121
rect 3000 69058 3800 69088
rect 4117 69058 4183 69061
rect 3000 69056 4183 69058
rect 3000 69000 4122 69056
rect 4178 69000 4183 69056
rect 6614 69056 6620 69120
rect 6684 69056 6700 69120
rect 6764 69056 6780 69120
rect 6844 69056 6860 69120
rect 6924 69056 6930 69120
rect 87206 69120 87522 69121
rect 84801 69058 84867 69061
rect 6614 69055 6930 69056
rect 3000 68998 4183 69000
rect 3000 68968 3800 68998
rect 4117 68995 4183 68998
rect 5405 68922 5471 68925
rect 10054 68922 10114 69028
rect 45596 68998 47436 69058
rect 83132 69056 84867 69058
rect 83132 69000 84806 69056
rect 84862 69000 84867 69056
rect 87206 69056 87212 69120
rect 87276 69056 87292 69120
rect 87356 69056 87372 69120
rect 87436 69056 87452 69120
rect 87516 69056 87522 69120
rect 87206 69055 87522 69056
rect 88573 69058 88639 69061
rect 89200 69058 90000 69088
rect 88573 69056 90000 69058
rect 83132 68998 84867 69000
rect 84801 68995 84867 68998
rect 88573 69000 88578 69056
rect 88634 69000 90000 69056
rect 88573 68998 90000 69000
rect 88573 68995 88639 68998
rect 89200 68968 90000 68998
rect 5405 68920 10114 68922
rect 5405 68864 5410 68920
rect 5466 68864 10114 68920
rect 5405 68862 10114 68864
rect 5405 68859 5471 68862
rect 5878 68576 6194 68577
rect 5878 68512 5884 68576
rect 5948 68512 5964 68576
rect 6028 68512 6044 68576
rect 6108 68512 6124 68576
rect 6188 68512 6194 68576
rect 5878 68511 6194 68512
rect 86470 68576 86786 68577
rect 86470 68512 86476 68576
rect 86540 68512 86556 68576
rect 86620 68512 86636 68576
rect 86700 68512 86716 68576
rect 86780 68512 86786 68576
rect 86470 68511 86786 68512
rect 5405 68242 5471 68245
rect 5405 68240 10114 68242
rect 5405 68184 5410 68240
rect 5466 68184 10114 68240
rect 5405 68182 10114 68184
rect 5405 68179 5471 68182
rect 6614 68032 6930 68033
rect 6614 67968 6620 68032
rect 6684 67968 6700 68032
rect 6764 67968 6780 68032
rect 6844 67968 6860 68032
rect 6924 67968 6930 68032
rect 6614 67967 6930 67968
rect 10054 67940 10114 68182
rect 87206 68032 87522 68033
rect 85261 67970 85327 67973
rect 45596 67910 47436 67970
rect 83132 67968 85327 67970
rect 83132 67912 85266 67968
rect 85322 67912 85327 67968
rect 87206 67968 87212 68032
rect 87276 67968 87292 68032
rect 87356 67968 87372 68032
rect 87436 67968 87452 68032
rect 87516 67968 87522 68032
rect 87206 67967 87522 67968
rect 83132 67910 85327 67912
rect 85261 67907 85327 67910
rect 3000 67698 3800 67728
rect 4025 67698 4091 67701
rect 3000 67696 4091 67698
rect 3000 67640 4030 67696
rect 4086 67640 4091 67696
rect 3000 67638 4091 67640
rect 3000 67608 3800 67638
rect 4025 67635 4091 67638
rect 88205 67698 88271 67701
rect 89200 67698 90000 67728
rect 88205 67696 90000 67698
rect 88205 67640 88210 67696
rect 88266 67640 90000 67696
rect 88205 67638 90000 67640
rect 88205 67635 88271 67638
rect 89200 67608 90000 67638
rect 5878 67488 6194 67489
rect 5878 67424 5884 67488
rect 5948 67424 5964 67488
rect 6028 67424 6044 67488
rect 6108 67424 6124 67488
rect 6188 67424 6194 67488
rect 5878 67423 6194 67424
rect 86470 67488 86786 67489
rect 86470 67424 86476 67488
rect 86540 67424 86556 67488
rect 86620 67424 86636 67488
rect 86700 67424 86716 67488
rect 86780 67424 86786 67488
rect 86470 67423 86786 67424
rect 3000 67018 3800 67048
rect 4117 67018 4183 67021
rect 3000 67016 4183 67018
rect 3000 66960 4122 67016
rect 4178 66960 4183 67016
rect 3000 66958 4183 66960
rect 3000 66928 3800 66958
rect 4117 66955 4183 66958
rect 88205 67018 88271 67021
rect 89200 67018 90000 67048
rect 88205 67016 90000 67018
rect 88205 66960 88210 67016
rect 88266 66960 90000 67016
rect 88205 66958 90000 66960
rect 88205 66955 88271 66958
rect 6614 66944 6930 66945
rect 6614 66880 6620 66944
rect 6684 66880 6700 66944
rect 6764 66880 6780 66944
rect 6844 66880 6860 66944
rect 6924 66880 6930 66944
rect 87206 66944 87522 66945
rect 6614 66879 6930 66880
rect 8533 66882 8599 66885
rect 85813 66882 85879 66885
rect 8533 66880 10084 66882
rect 8533 66824 8538 66880
rect 8594 66824 10084 66880
rect 8533 66822 10084 66824
rect 45596 66822 47436 66882
rect 83132 66880 85879 66882
rect 83132 66824 85818 66880
rect 85874 66824 85879 66880
rect 87206 66880 87212 66944
rect 87276 66880 87292 66944
rect 87356 66880 87372 66944
rect 87436 66880 87452 66944
rect 87516 66880 87522 66944
rect 89200 66928 90000 66958
rect 87206 66879 87522 66880
rect 83132 66822 85879 66824
rect 8533 66819 8599 66822
rect 85813 66819 85879 66822
rect 5878 66400 6194 66401
rect 5878 66336 5884 66400
rect 5948 66336 5964 66400
rect 6028 66336 6044 66400
rect 6108 66336 6124 66400
rect 6188 66336 6194 66400
rect 5878 66335 6194 66336
rect 86470 66400 86786 66401
rect 86470 66336 86476 66400
rect 86540 66336 86556 66400
rect 86620 66336 86636 66400
rect 86700 66336 86716 66400
rect 86780 66336 86786 66400
rect 86470 66335 86786 66336
rect 6614 65856 6930 65857
rect 6614 65792 6620 65856
rect 6684 65792 6700 65856
rect 6764 65792 6780 65856
rect 6844 65792 6860 65856
rect 6924 65792 6930 65856
rect 87206 65856 87522 65857
rect 6614 65791 6930 65792
rect 8533 65794 8599 65797
rect 85813 65794 85879 65797
rect 8533 65792 10084 65794
rect 8533 65736 8538 65792
rect 8594 65736 10084 65792
rect 8533 65734 10084 65736
rect 45596 65734 47436 65794
rect 83132 65792 85879 65794
rect 83132 65736 85818 65792
rect 85874 65736 85879 65792
rect 87206 65792 87212 65856
rect 87276 65792 87292 65856
rect 87356 65792 87372 65856
rect 87436 65792 87452 65856
rect 87516 65792 87522 65856
rect 87206 65791 87522 65792
rect 83132 65734 85879 65736
rect 8533 65731 8599 65734
rect 85813 65731 85879 65734
rect 3000 65658 3800 65688
rect 4301 65658 4367 65661
rect 3000 65656 4367 65658
rect 3000 65600 4306 65656
rect 4362 65600 4367 65656
rect 3000 65598 4367 65600
rect 3000 65568 3800 65598
rect 4301 65595 4367 65598
rect 88205 65658 88271 65661
rect 89200 65658 90000 65688
rect 88205 65656 90000 65658
rect 88205 65600 88210 65656
rect 88266 65600 90000 65656
rect 88205 65598 90000 65600
rect 88205 65595 88271 65598
rect 89200 65568 90000 65598
rect 5878 65312 6194 65313
rect 5878 65248 5884 65312
rect 5948 65248 5964 65312
rect 6028 65248 6044 65312
rect 6108 65248 6124 65312
rect 6188 65248 6194 65312
rect 5878 65247 6194 65248
rect 86470 65312 86786 65313
rect 86470 65248 86476 65312
rect 86540 65248 86556 65312
rect 86620 65248 86636 65312
rect 86700 65248 86716 65312
rect 86780 65248 86786 65312
rect 86470 65247 86786 65248
rect 3000 64978 3800 65008
rect 4301 64978 4367 64981
rect 3000 64976 4367 64978
rect 3000 64920 4306 64976
rect 4362 64920 4367 64976
rect 3000 64918 4367 64920
rect 3000 64888 3800 64918
rect 4301 64915 4367 64918
rect 88389 64978 88455 64981
rect 89200 64978 90000 65008
rect 88389 64976 90000 64978
rect 88389 64920 88394 64976
rect 88450 64920 90000 64976
rect 88389 64918 90000 64920
rect 88389 64915 88455 64918
rect 89200 64888 90000 64918
rect 6614 64768 6930 64769
rect 6614 64704 6620 64768
rect 6684 64704 6700 64768
rect 6764 64704 6780 64768
rect 6844 64704 6860 64768
rect 6924 64704 6930 64768
rect 87206 64768 87522 64769
rect 6614 64703 6930 64704
rect 8533 64706 8599 64709
rect 85813 64706 85879 64709
rect 8533 64704 10084 64706
rect 8533 64648 8538 64704
rect 8594 64648 10084 64704
rect 8533 64646 10084 64648
rect 45596 64646 47436 64706
rect 83132 64704 85879 64706
rect 83132 64648 85818 64704
rect 85874 64648 85879 64704
rect 87206 64704 87212 64768
rect 87276 64704 87292 64768
rect 87356 64704 87372 64768
rect 87436 64704 87452 64768
rect 87516 64704 87522 64768
rect 87206 64703 87522 64704
rect 83132 64646 85879 64648
rect 8533 64643 8599 64646
rect 85813 64643 85879 64646
rect 5878 64224 6194 64225
rect 5878 64160 5884 64224
rect 5948 64160 5964 64224
rect 6028 64160 6044 64224
rect 6108 64160 6124 64224
rect 6188 64160 6194 64224
rect 5878 64159 6194 64160
rect 86470 64224 86786 64225
rect 86470 64160 86476 64224
rect 86540 64160 86556 64224
rect 86620 64160 86636 64224
rect 86700 64160 86716 64224
rect 86780 64160 86786 64224
rect 86470 64159 86786 64160
rect 6614 63680 6930 63681
rect 3000 63618 3800 63648
rect 4301 63618 4367 63621
rect 3000 63616 4367 63618
rect 3000 63560 4306 63616
rect 4362 63560 4367 63616
rect 6614 63616 6620 63680
rect 6684 63616 6700 63680
rect 6764 63616 6780 63680
rect 6844 63616 6860 63680
rect 6924 63616 6930 63680
rect 87206 63680 87522 63681
rect 84525 63618 84591 63621
rect 6614 63615 6930 63616
rect 3000 63558 4367 63560
rect 3000 63528 3800 63558
rect 4301 63555 4367 63558
rect 5681 63482 5747 63485
rect 10054 63482 10114 63588
rect 45596 63558 47436 63618
rect 83132 63616 84591 63618
rect 83132 63560 84530 63616
rect 84586 63560 84591 63616
rect 87206 63616 87212 63680
rect 87276 63616 87292 63680
rect 87356 63616 87372 63680
rect 87436 63616 87452 63680
rect 87516 63616 87522 63680
rect 87206 63615 87522 63616
rect 88573 63618 88639 63621
rect 89200 63618 90000 63648
rect 88573 63616 90000 63618
rect 83132 63558 84591 63560
rect 84525 63555 84591 63558
rect 88573 63560 88578 63616
rect 88634 63560 90000 63616
rect 88573 63558 90000 63560
rect 88573 63555 88639 63558
rect 89200 63528 90000 63558
rect 5681 63480 10114 63482
rect 5681 63424 5686 63480
rect 5742 63424 10114 63480
rect 5681 63422 10114 63424
rect 5681 63419 5747 63422
rect 5878 63136 6194 63137
rect 5878 63072 5884 63136
rect 5948 63072 5964 63136
rect 6028 63072 6044 63136
rect 6108 63072 6124 63136
rect 6188 63072 6194 63136
rect 5878 63071 6194 63072
rect 86470 63136 86786 63137
rect 86470 63072 86476 63136
rect 86540 63072 86556 63136
rect 86620 63072 86636 63136
rect 86700 63072 86716 63136
rect 86780 63072 86786 63136
rect 86470 63071 86786 63072
rect 6614 62592 6930 62593
rect 6614 62528 6620 62592
rect 6684 62528 6700 62592
rect 6764 62528 6780 62592
rect 6844 62528 6860 62592
rect 6924 62528 6930 62592
rect 87206 62592 87522 62593
rect 84801 62530 84867 62533
rect 6614 62527 6930 62528
rect 5681 62394 5747 62397
rect 10054 62394 10114 62500
rect 45596 62470 47436 62530
rect 83132 62528 84867 62530
rect 83132 62472 84806 62528
rect 84862 62472 84867 62528
rect 87206 62528 87212 62592
rect 87276 62528 87292 62592
rect 87356 62528 87372 62592
rect 87436 62528 87452 62592
rect 87516 62528 87522 62592
rect 87206 62527 87522 62528
rect 83132 62470 84867 62472
rect 84801 62467 84867 62470
rect 5681 62392 10114 62394
rect 5681 62336 5686 62392
rect 5742 62336 10114 62392
rect 5681 62334 10114 62336
rect 5681 62331 5747 62334
rect 3000 62258 3800 62288
rect 4301 62258 4367 62261
rect 3000 62256 4367 62258
rect 3000 62200 4306 62256
rect 4362 62200 4367 62256
rect 3000 62198 4367 62200
rect 3000 62168 3800 62198
rect 4301 62195 4367 62198
rect 88389 62258 88455 62261
rect 89200 62258 90000 62288
rect 88389 62256 90000 62258
rect 88389 62200 88394 62256
rect 88450 62200 90000 62256
rect 88389 62198 90000 62200
rect 88389 62195 88455 62198
rect 89200 62168 90000 62198
rect 5878 62048 6194 62049
rect 5878 61984 5884 62048
rect 5948 61984 5964 62048
rect 6028 61984 6044 62048
rect 6108 61984 6124 62048
rect 6188 61984 6194 62048
rect 5878 61983 6194 61984
rect 86470 62048 86786 62049
rect 86470 61984 86476 62048
rect 86540 61984 86556 62048
rect 86620 61984 86636 62048
rect 86700 61984 86716 62048
rect 86780 61984 86786 62048
rect 86470 61983 86786 61984
rect 3000 61578 3800 61608
rect 4301 61578 4367 61581
rect 3000 61576 4367 61578
rect 3000 61520 4306 61576
rect 4362 61520 4367 61576
rect 3000 61518 4367 61520
rect 3000 61488 3800 61518
rect 4301 61515 4367 61518
rect 88205 61578 88271 61581
rect 89200 61578 90000 61608
rect 88205 61576 90000 61578
rect 88205 61520 88210 61576
rect 88266 61520 90000 61576
rect 88205 61518 90000 61520
rect 88205 61515 88271 61518
rect 6614 61504 6930 61505
rect 6614 61440 6620 61504
rect 6684 61440 6700 61504
rect 6764 61440 6780 61504
rect 6844 61440 6860 61504
rect 6924 61440 6930 61504
rect 87206 61504 87522 61505
rect 6614 61439 6930 61440
rect 8533 61442 8599 61445
rect 85813 61442 85879 61445
rect 8533 61440 10084 61442
rect 8533 61384 8538 61440
rect 8594 61384 10084 61440
rect 8533 61382 10084 61384
rect 45596 61382 47436 61442
rect 83132 61440 85879 61442
rect 83132 61384 85818 61440
rect 85874 61384 85879 61440
rect 87206 61440 87212 61504
rect 87276 61440 87292 61504
rect 87356 61440 87372 61504
rect 87436 61440 87452 61504
rect 87516 61440 87522 61504
rect 89200 61488 90000 61518
rect 87206 61439 87522 61440
rect 83132 61382 85879 61384
rect 8533 61379 8599 61382
rect 85813 61379 85879 61382
rect 5878 60960 6194 60961
rect 5878 60896 5884 60960
rect 5948 60896 5964 60960
rect 6028 60896 6044 60960
rect 6108 60896 6124 60960
rect 6188 60896 6194 60960
rect 5878 60895 6194 60896
rect 86470 60960 86786 60961
rect 86470 60896 86476 60960
rect 86540 60896 86556 60960
rect 86620 60896 86636 60960
rect 86700 60896 86716 60960
rect 86780 60896 86786 60960
rect 86470 60895 86786 60896
rect 6614 60416 6930 60417
rect 6614 60352 6620 60416
rect 6684 60352 6700 60416
rect 6764 60352 6780 60416
rect 6844 60352 6860 60416
rect 6924 60352 6930 60416
rect 87206 60416 87522 60417
rect 6614 60351 6930 60352
rect 8533 60354 8599 60357
rect 85813 60354 85879 60357
rect 8533 60352 10084 60354
rect 8533 60296 8538 60352
rect 8594 60296 10084 60352
rect 8533 60294 10084 60296
rect 45596 60294 47436 60354
rect 83132 60352 85879 60354
rect 83132 60296 85818 60352
rect 85874 60296 85879 60352
rect 87206 60352 87212 60416
rect 87276 60352 87292 60416
rect 87356 60352 87372 60416
rect 87436 60352 87452 60416
rect 87516 60352 87522 60416
rect 87206 60351 87522 60352
rect 83132 60294 85879 60296
rect 8533 60291 8599 60294
rect 85813 60291 85879 60294
rect 3000 60218 3800 60248
rect 4301 60218 4367 60221
rect 3000 60216 4367 60218
rect 3000 60160 4306 60216
rect 4362 60160 4367 60216
rect 3000 60158 4367 60160
rect 3000 60128 3800 60158
rect 4301 60155 4367 60158
rect 88205 60218 88271 60221
rect 89200 60218 90000 60248
rect 88205 60216 90000 60218
rect 88205 60160 88210 60216
rect 88266 60160 90000 60216
rect 88205 60158 90000 60160
rect 88205 60155 88271 60158
rect 89200 60128 90000 60158
rect 5878 59872 6194 59873
rect 5878 59808 5884 59872
rect 5948 59808 5964 59872
rect 6028 59808 6044 59872
rect 6108 59808 6124 59872
rect 6188 59808 6194 59872
rect 5878 59807 6194 59808
rect 86470 59872 86786 59873
rect 86470 59808 86476 59872
rect 86540 59808 86556 59872
rect 86620 59808 86636 59872
rect 86700 59808 86716 59872
rect 86780 59808 86786 59872
rect 86470 59807 86786 59808
rect 3000 59538 3800 59568
rect 4301 59538 4367 59541
rect 87469 59538 87535 59541
rect 3000 59536 4367 59538
rect 3000 59480 4306 59536
rect 4362 59480 4367 59536
rect 3000 59478 4367 59480
rect 3000 59448 3800 59478
rect 4301 59475 4367 59478
rect 84758 59536 87535 59538
rect 84758 59480 87474 59536
rect 87530 59480 87535 59536
rect 84758 59478 87535 59480
rect 6614 59328 6930 59329
rect 6614 59264 6620 59328
rect 6684 59264 6700 59328
rect 6764 59264 6780 59328
rect 6844 59264 6860 59328
rect 6924 59264 6930 59328
rect 6614 59263 6930 59264
rect 8533 59266 8599 59269
rect 84758 59266 84818 59478
rect 87469 59475 87535 59478
rect 88205 59538 88271 59541
rect 89200 59538 90000 59568
rect 88205 59536 90000 59538
rect 88205 59480 88210 59536
rect 88266 59480 90000 59536
rect 88205 59478 90000 59480
rect 88205 59475 88271 59478
rect 89200 59448 90000 59478
rect 8533 59264 10084 59266
rect 8533 59208 8538 59264
rect 8594 59208 10084 59264
rect 8533 59206 10084 59208
rect 45596 59206 47436 59266
rect 83132 59206 84818 59266
rect 87206 59328 87522 59329
rect 87206 59264 87212 59328
rect 87276 59264 87292 59328
rect 87356 59264 87372 59328
rect 87436 59264 87452 59328
rect 87516 59264 87522 59328
rect 87206 59263 87522 59264
rect 8533 59203 8599 59206
rect 5878 58784 6194 58785
rect 5878 58720 5884 58784
rect 5948 58720 5964 58784
rect 6028 58720 6044 58784
rect 6108 58720 6124 58784
rect 6188 58720 6194 58784
rect 5878 58719 6194 58720
rect 86470 58784 86786 58785
rect 86470 58720 86476 58784
rect 86540 58720 86556 58784
rect 86620 58720 86636 58784
rect 86700 58720 86716 58784
rect 86780 58720 86786 58784
rect 86470 58719 86786 58720
rect 6614 58240 6930 58241
rect 3000 58178 3800 58208
rect 4301 58178 4367 58181
rect 3000 58176 4367 58178
rect 3000 58120 4306 58176
rect 4362 58120 4367 58176
rect 6614 58176 6620 58240
rect 6684 58176 6700 58240
rect 6764 58176 6780 58240
rect 6844 58176 6860 58240
rect 6924 58176 6930 58240
rect 87206 58240 87522 58241
rect 85077 58178 85143 58181
rect 6614 58175 6930 58176
rect 3000 58118 4367 58120
rect 3000 58088 3800 58118
rect 4301 58115 4367 58118
rect 5405 58042 5471 58045
rect 10054 58042 10114 58148
rect 45596 58118 47436 58178
rect 83132 58176 85143 58178
rect 83132 58120 85082 58176
rect 85138 58120 85143 58176
rect 87206 58176 87212 58240
rect 87276 58176 87292 58240
rect 87356 58176 87372 58240
rect 87436 58176 87452 58240
rect 87516 58176 87522 58240
rect 87206 58175 87522 58176
rect 88573 58178 88639 58181
rect 89200 58178 90000 58208
rect 88573 58176 90000 58178
rect 83132 58118 85143 58120
rect 85077 58115 85143 58118
rect 88573 58120 88578 58176
rect 88634 58120 90000 58176
rect 88573 58118 90000 58120
rect 88573 58115 88639 58118
rect 89200 58088 90000 58118
rect 5405 58040 10114 58042
rect 5405 57984 5410 58040
rect 5466 57984 10114 58040
rect 5405 57982 10114 57984
rect 5405 57979 5471 57982
rect 5878 57696 6194 57697
rect 5878 57632 5884 57696
rect 5948 57632 5964 57696
rect 6028 57632 6044 57696
rect 6108 57632 6124 57696
rect 6188 57632 6194 57696
rect 5878 57631 6194 57632
rect 86470 57696 86786 57697
rect 86470 57632 86476 57696
rect 86540 57632 86556 57696
rect 86620 57632 86636 57696
rect 86700 57632 86716 57696
rect 86780 57632 86786 57696
rect 86470 57631 86786 57632
rect 6614 57152 6930 57153
rect 6614 57088 6620 57152
rect 6684 57088 6700 57152
rect 6764 57088 6780 57152
rect 6844 57088 6860 57152
rect 6924 57088 6930 57152
rect 87206 57152 87522 57153
rect 6614 57087 6930 57088
rect 9913 56954 9979 56957
rect 10054 56954 10114 57060
rect 45596 57030 47436 57090
rect 83132 57030 84082 57090
rect 87206 57088 87212 57152
rect 87276 57088 87292 57152
rect 87356 57088 87372 57152
rect 87436 57088 87452 57152
rect 87516 57088 87522 57152
rect 87206 57087 87522 57088
rect 9913 56952 10114 56954
rect 9913 56896 9918 56952
rect 9974 56896 10114 56952
rect 9913 56894 10114 56896
rect 84022 56954 84082 57030
rect 87561 56954 87627 56957
rect 84022 56952 87627 56954
rect 84022 56896 87566 56952
rect 87622 56896 87627 56952
rect 84022 56894 87627 56896
rect 9913 56891 9979 56894
rect 87561 56891 87627 56894
rect 3000 56818 3800 56848
rect 4301 56818 4367 56821
rect 3000 56816 4367 56818
rect 3000 56760 4306 56816
rect 4362 56760 4367 56816
rect 3000 56758 4367 56760
rect 3000 56728 3800 56758
rect 4301 56755 4367 56758
rect 88573 56818 88639 56821
rect 89200 56818 90000 56848
rect 88573 56816 90000 56818
rect 88573 56760 88578 56816
rect 88634 56760 90000 56816
rect 88573 56758 90000 56760
rect 88573 56755 88639 56758
rect 89200 56728 90000 56758
rect 5878 56608 6194 56609
rect 5878 56544 5884 56608
rect 5948 56544 5964 56608
rect 6028 56544 6044 56608
rect 6108 56544 6124 56608
rect 6188 56544 6194 56608
rect 5878 56543 6194 56544
rect 86470 56608 86786 56609
rect 86470 56544 86476 56608
rect 86540 56544 86556 56608
rect 86620 56544 86636 56608
rect 86700 56544 86716 56608
rect 86780 56544 86786 56608
rect 86470 56543 86786 56544
rect 9913 56274 9979 56277
rect 9913 56272 10114 56274
rect 9913 56216 9918 56272
rect 9974 56216 10114 56272
rect 9913 56214 10114 56216
rect 9913 56211 9979 56214
rect 3000 56138 3800 56168
rect 4301 56138 4367 56141
rect 3000 56136 4367 56138
rect 3000 56080 4306 56136
rect 4362 56080 4367 56136
rect 3000 56078 4367 56080
rect 3000 56048 3800 56078
rect 4301 56075 4367 56078
rect 6614 56064 6930 56065
rect 6614 56000 6620 56064
rect 6684 56000 6700 56064
rect 6764 56000 6780 56064
rect 6844 56000 6860 56064
rect 6924 56000 6930 56064
rect 6614 55999 6930 56000
rect 10054 55972 10114 56214
rect 88205 56138 88271 56141
rect 89200 56138 90000 56168
rect 88205 56136 90000 56138
rect 88205 56080 88210 56136
rect 88266 56080 90000 56136
rect 88205 56078 90000 56080
rect 88205 56075 88271 56078
rect 87206 56064 87522 56065
rect 85813 56002 85879 56005
rect 45596 55942 47436 56002
rect 83132 56000 85879 56002
rect 83132 55944 85818 56000
rect 85874 55944 85879 56000
rect 87206 56000 87212 56064
rect 87276 56000 87292 56064
rect 87356 56000 87372 56064
rect 87436 56000 87452 56064
rect 87516 56000 87522 56064
rect 89200 56048 90000 56078
rect 87206 55999 87522 56000
rect 83132 55942 85879 55944
rect 85813 55939 85879 55942
rect 5878 55520 6194 55521
rect 5878 55456 5884 55520
rect 5948 55456 5964 55520
rect 6028 55456 6044 55520
rect 6108 55456 6124 55520
rect 6188 55456 6194 55520
rect 5878 55455 6194 55456
rect 86470 55520 86786 55521
rect 86470 55456 86476 55520
rect 86540 55456 86556 55520
rect 86620 55456 86636 55520
rect 86700 55456 86716 55520
rect 86780 55456 86786 55520
rect 86470 55455 86786 55456
rect 6614 54976 6930 54977
rect 6614 54912 6620 54976
rect 6684 54912 6700 54976
rect 6764 54912 6780 54976
rect 6844 54912 6860 54976
rect 6924 54912 6930 54976
rect 87206 54976 87522 54977
rect 6614 54911 6930 54912
rect 8533 54914 8599 54917
rect 85813 54914 85879 54917
rect 8533 54912 10084 54914
rect 8533 54856 8538 54912
rect 8594 54856 10084 54912
rect 8533 54854 10084 54856
rect 45596 54854 47436 54914
rect 83132 54912 85879 54914
rect 83132 54856 85818 54912
rect 85874 54856 85879 54912
rect 87206 54912 87212 54976
rect 87276 54912 87292 54976
rect 87356 54912 87372 54976
rect 87436 54912 87452 54976
rect 87516 54912 87522 54976
rect 87206 54911 87522 54912
rect 83132 54854 85879 54856
rect 8533 54851 8599 54854
rect 85813 54851 85879 54854
rect 3000 54778 3800 54808
rect 4301 54778 4367 54781
rect 3000 54776 4367 54778
rect 3000 54720 4306 54776
rect 4362 54720 4367 54776
rect 3000 54718 4367 54720
rect 3000 54688 3800 54718
rect 4301 54715 4367 54718
rect 88205 54778 88271 54781
rect 89200 54778 90000 54808
rect 88205 54776 90000 54778
rect 88205 54720 88210 54776
rect 88266 54720 90000 54776
rect 88205 54718 90000 54720
rect 88205 54715 88271 54718
rect 89200 54688 90000 54718
rect 5878 54432 6194 54433
rect 5878 54368 5884 54432
rect 5948 54368 5964 54432
rect 6028 54368 6044 54432
rect 6108 54368 6124 54432
rect 6188 54368 6194 54432
rect 5878 54367 6194 54368
rect 86470 54432 86786 54433
rect 86470 54368 86476 54432
rect 86540 54368 86556 54432
rect 86620 54368 86636 54432
rect 86700 54368 86716 54432
rect 86780 54368 86786 54432
rect 86470 54367 86786 54368
rect 3000 54098 3800 54128
rect 4301 54098 4367 54101
rect 3000 54096 4367 54098
rect 3000 54040 4306 54096
rect 4362 54040 4367 54096
rect 3000 54038 4367 54040
rect 3000 54008 3800 54038
rect 4301 54035 4367 54038
rect 88205 54098 88271 54101
rect 89200 54098 90000 54128
rect 88205 54096 90000 54098
rect 88205 54040 88210 54096
rect 88266 54040 90000 54096
rect 88205 54038 90000 54040
rect 88205 54035 88271 54038
rect 89200 54008 90000 54038
rect 6614 53888 6930 53889
rect 6614 53824 6620 53888
rect 6684 53824 6700 53888
rect 6764 53824 6780 53888
rect 6844 53824 6860 53888
rect 6924 53824 6930 53888
rect 87206 53888 87522 53889
rect 84525 53826 84591 53829
rect 6614 53823 6930 53824
rect 5681 53690 5747 53693
rect 10054 53690 10114 53796
rect 45596 53766 47436 53826
rect 83132 53824 84591 53826
rect 83132 53768 84530 53824
rect 84586 53768 84591 53824
rect 87206 53824 87212 53888
rect 87276 53824 87292 53888
rect 87356 53824 87372 53888
rect 87436 53824 87452 53888
rect 87516 53824 87522 53888
rect 87206 53823 87522 53824
rect 83132 53766 84591 53768
rect 84525 53763 84591 53766
rect 5681 53688 10114 53690
rect 5681 53632 5686 53688
rect 5742 53632 10114 53688
rect 5681 53630 10114 53632
rect 5681 53627 5747 53630
rect 5878 53344 6194 53345
rect 5878 53280 5884 53344
rect 5948 53280 5964 53344
rect 6028 53280 6044 53344
rect 6108 53280 6124 53344
rect 6188 53280 6194 53344
rect 5878 53279 6194 53280
rect 86470 53344 86786 53345
rect 86470 53280 86476 53344
rect 86540 53280 86556 53344
rect 86620 53280 86636 53344
rect 86700 53280 86716 53344
rect 86780 53280 86786 53344
rect 86470 53279 86786 53280
rect 87561 53010 87627 53013
rect 84206 53008 87627 53010
rect 84206 52952 87566 53008
rect 87622 52952 87627 53008
rect 84206 52950 87627 52952
rect 6614 52800 6930 52801
rect 3000 52738 3800 52768
rect 4301 52738 4367 52741
rect 3000 52736 4367 52738
rect 3000 52680 4306 52736
rect 4362 52680 4367 52736
rect 6614 52736 6620 52800
rect 6684 52736 6700 52800
rect 6764 52736 6780 52800
rect 6844 52736 6860 52800
rect 6924 52736 6930 52800
rect 6614 52735 6930 52736
rect 8533 52738 8599 52741
rect 84206 52738 84266 52950
rect 87561 52947 87627 52950
rect 8533 52736 10084 52738
rect 3000 52678 4367 52680
rect 3000 52648 3800 52678
rect 4301 52675 4367 52678
rect 8533 52680 8538 52736
rect 8594 52680 10084 52736
rect 8533 52678 10084 52680
rect 45596 52678 47436 52738
rect 83132 52678 84266 52738
rect 87206 52800 87522 52801
rect 87206 52736 87212 52800
rect 87276 52736 87292 52800
rect 87356 52736 87372 52800
rect 87436 52736 87452 52800
rect 87516 52736 87522 52800
rect 87206 52735 87522 52736
rect 88205 52738 88271 52741
rect 89200 52738 90000 52768
rect 88205 52736 90000 52738
rect 88205 52680 88210 52736
rect 88266 52680 90000 52736
rect 88205 52678 90000 52680
rect 8533 52675 8599 52678
rect 88205 52675 88271 52678
rect 89200 52648 90000 52678
rect 5878 52256 6194 52257
rect 5878 52192 5884 52256
rect 5948 52192 5964 52256
rect 6028 52192 6044 52256
rect 6108 52192 6124 52256
rect 6188 52192 6194 52256
rect 5878 52191 6194 52192
rect 86470 52256 86786 52257
rect 86470 52192 86476 52256
rect 86540 52192 86556 52256
rect 86620 52192 86636 52256
rect 86700 52192 86716 52256
rect 86780 52192 86786 52256
rect 86470 52191 86786 52192
rect 6614 51712 6930 51713
rect 6614 51648 6620 51712
rect 6684 51648 6700 51712
rect 6764 51648 6780 51712
rect 6844 51648 6860 51712
rect 6924 51648 6930 51712
rect 87206 51712 87522 51713
rect 6614 51647 6930 51648
rect 8533 51650 8599 51653
rect 8533 51648 10084 51650
rect 8533 51592 8538 51648
rect 8594 51592 10084 51648
rect 8533 51590 10084 51592
rect 45596 51590 47436 51650
rect 83132 51590 84082 51650
rect 87206 51648 87212 51712
rect 87276 51648 87292 51712
rect 87356 51648 87372 51712
rect 87436 51648 87452 51712
rect 87516 51648 87522 51712
rect 87206 51647 87522 51648
rect 8533 51587 8599 51590
rect 84022 51514 84082 51590
rect 87561 51514 87627 51517
rect 84022 51512 87627 51514
rect 84022 51456 87566 51512
rect 87622 51456 87627 51512
rect 84022 51454 87627 51456
rect 87561 51451 87627 51454
rect 3000 51378 3800 51408
rect 4301 51378 4367 51381
rect 3000 51376 4367 51378
rect 3000 51320 4306 51376
rect 4362 51320 4367 51376
rect 3000 51318 4367 51320
rect 3000 51288 3800 51318
rect 4301 51315 4367 51318
rect 88205 51378 88271 51381
rect 89200 51378 90000 51408
rect 88205 51376 90000 51378
rect 88205 51320 88210 51376
rect 88266 51320 90000 51376
rect 88205 51318 90000 51320
rect 88205 51315 88271 51318
rect 89200 51288 90000 51318
rect 5878 51168 6194 51169
rect 5878 51104 5884 51168
rect 5948 51104 5964 51168
rect 6028 51104 6044 51168
rect 6108 51104 6124 51168
rect 6188 51104 6194 51168
rect 5878 51103 6194 51104
rect 86470 51168 86786 51169
rect 86470 51104 86476 51168
rect 86540 51104 86556 51168
rect 86620 51104 86636 51168
rect 86700 51104 86716 51168
rect 86780 51104 86786 51168
rect 86470 51103 86786 51104
rect 6614 50624 6930 50625
rect 6614 50560 6620 50624
rect 6684 50560 6700 50624
rect 6764 50560 6780 50624
rect 6844 50560 6860 50624
rect 6924 50560 6930 50624
rect 87206 50624 87522 50625
rect 45977 50562 46043 50565
rect 85445 50562 85511 50565
rect 85629 50562 85695 50565
rect 6614 50559 6930 50560
rect 45596 50560 46043 50562
rect 45596 50504 45982 50560
rect 46038 50504 46043 50560
rect 45596 50502 46043 50504
rect 83132 50560 85695 50562
rect 83132 50504 85450 50560
rect 85506 50504 85634 50560
rect 85690 50504 85695 50560
rect 87206 50560 87212 50624
rect 87276 50560 87292 50624
rect 87356 50560 87372 50624
rect 87436 50560 87452 50624
rect 87516 50560 87522 50624
rect 87206 50559 87522 50560
rect 83132 50502 85695 50504
rect 45977 50499 46043 50502
rect 85445 50499 85511 50502
rect 85629 50499 85695 50502
rect 5878 50080 6194 50081
rect 5878 50016 5884 50080
rect 5948 50016 5964 50080
rect 6028 50016 6044 50080
rect 6108 50016 6124 50080
rect 6188 50016 6194 50080
rect 5878 50015 6194 50016
rect 86470 50080 86786 50081
rect 86470 50016 86476 50080
rect 86540 50016 86556 50080
rect 86620 50016 86636 50080
rect 86700 50016 86716 50080
rect 86780 50016 86786 50080
rect 86470 50015 86786 50016
rect 6614 49536 6930 49537
rect 6614 49472 6620 49536
rect 6684 49472 6700 49536
rect 6764 49472 6780 49536
rect 6844 49472 6860 49536
rect 6924 49472 6930 49536
rect 87206 49536 87522 49537
rect 45885 49474 45951 49477
rect 85629 49474 85695 49477
rect 6614 49471 6930 49472
rect 45596 49472 45951 49474
rect 45596 49416 45890 49472
rect 45946 49416 45951 49472
rect 45596 49414 45951 49416
rect 83132 49472 85695 49474
rect 83132 49416 85634 49472
rect 85690 49416 85695 49472
rect 87206 49472 87212 49536
rect 87276 49472 87292 49536
rect 87356 49472 87372 49536
rect 87436 49472 87452 49536
rect 87516 49472 87522 49536
rect 87206 49471 87522 49472
rect 83132 49414 85695 49416
rect 45885 49411 45951 49414
rect 85629 49411 85695 49414
rect 5878 48992 6194 48993
rect 5878 48928 5884 48992
rect 5948 48928 5964 48992
rect 6028 48928 6044 48992
rect 6108 48928 6124 48992
rect 6188 48928 6194 48992
rect 5878 48927 6194 48928
rect 86470 48992 86786 48993
rect 86470 48928 86476 48992
rect 86540 48928 86556 48992
rect 86620 48928 86636 48992
rect 86700 48928 86716 48992
rect 86780 48928 86786 48992
rect 86470 48927 86786 48928
rect 88205 48658 88271 48661
rect 89200 48658 90000 48688
rect 88205 48656 90000 48658
rect 88205 48600 88210 48656
rect 88266 48600 90000 48656
rect 88205 48598 90000 48600
rect 88205 48595 88271 48598
rect 89200 48568 90000 48598
rect 6614 48448 6930 48449
rect 6614 48384 6620 48448
rect 6684 48384 6700 48448
rect 6764 48384 6780 48448
rect 6844 48384 6860 48448
rect 6924 48384 6930 48448
rect 87206 48448 87522 48449
rect 46069 48386 46135 48389
rect 85353 48386 85419 48389
rect 6614 48383 6930 48384
rect 45596 48384 46135 48386
rect 45596 48328 46074 48384
rect 46130 48328 46135 48384
rect 45596 48326 46135 48328
rect 83132 48384 85419 48386
rect 83132 48328 85358 48384
rect 85414 48328 85419 48384
rect 87206 48384 87212 48448
rect 87276 48384 87292 48448
rect 87356 48384 87372 48448
rect 87436 48384 87452 48448
rect 87516 48384 87522 48448
rect 87206 48383 87522 48384
rect 83132 48326 85419 48328
rect 46069 48323 46135 48326
rect 85353 48323 85419 48326
rect 88205 47978 88271 47981
rect 89200 47978 90000 48008
rect 88205 47976 90000 47978
rect 88205 47920 88210 47976
rect 88266 47920 90000 47976
rect 88205 47918 90000 47920
rect 88205 47915 88271 47918
rect 5878 47904 6194 47905
rect 5878 47840 5884 47904
rect 5948 47840 5964 47904
rect 6028 47840 6044 47904
rect 6108 47840 6124 47904
rect 6188 47840 6194 47904
rect 5878 47839 6194 47840
rect 86470 47904 86786 47905
rect 86470 47840 86476 47904
rect 86540 47840 86556 47904
rect 86620 47840 86636 47904
rect 86700 47840 86716 47904
rect 86780 47840 86786 47904
rect 89200 47888 90000 47918
rect 86470 47839 86786 47840
rect 6614 47360 6930 47361
rect 6614 47296 6620 47360
rect 6684 47296 6700 47360
rect 6764 47296 6780 47360
rect 6844 47296 6860 47360
rect 6924 47296 6930 47360
rect 87206 47360 87522 47361
rect 46161 47298 46227 47301
rect 85813 47298 85879 47301
rect 6614 47295 6930 47296
rect 45596 47296 46227 47298
rect 45596 47240 46166 47296
rect 46222 47240 46227 47296
rect 45596 47238 46227 47240
rect 83132 47296 85879 47298
rect 83132 47240 85818 47296
rect 85874 47240 85879 47296
rect 87206 47296 87212 47360
rect 87276 47296 87292 47360
rect 87356 47296 87372 47360
rect 87436 47296 87452 47360
rect 87516 47296 87522 47360
rect 87206 47295 87522 47296
rect 88205 47298 88271 47301
rect 89200 47298 90000 47328
rect 88205 47296 90000 47298
rect 83132 47238 85879 47240
rect 46161 47235 46227 47238
rect 85813 47235 85879 47238
rect 88205 47240 88210 47296
rect 88266 47240 90000 47296
rect 88205 47238 90000 47240
rect 88205 47235 88271 47238
rect 89200 47208 90000 47238
rect 5878 46816 6194 46817
rect 5878 46752 5884 46816
rect 5948 46752 5964 46816
rect 6028 46752 6044 46816
rect 6108 46752 6124 46816
rect 6188 46752 6194 46816
rect 5878 46751 6194 46752
rect 86470 46816 86786 46817
rect 86470 46752 86476 46816
rect 86540 46752 86556 46816
rect 86620 46752 86636 46816
rect 86700 46752 86716 46816
rect 86780 46752 86786 46816
rect 86470 46751 86786 46752
rect 88205 46618 88271 46621
rect 89200 46618 90000 46648
rect 88205 46616 90000 46618
rect 88205 46560 88210 46616
rect 88266 46560 90000 46616
rect 88205 46558 90000 46560
rect 88205 46555 88271 46558
rect 89200 46528 90000 46558
rect 6614 46272 6930 46273
rect 6614 46208 6620 46272
rect 6684 46208 6700 46272
rect 6764 46208 6780 46272
rect 6844 46208 6860 46272
rect 6924 46208 6930 46272
rect 6614 46207 6930 46208
rect 87206 46272 87522 46273
rect 87206 46208 87212 46272
rect 87276 46208 87292 46272
rect 87356 46208 87372 46272
rect 87436 46208 87452 46272
rect 87516 46208 87522 46272
rect 87206 46207 87522 46208
rect 11661 45938 11727 45941
rect 12765 45938 12831 45941
rect 13869 45938 13935 45941
rect 11661 45936 11770 45938
rect 11661 45880 11666 45936
rect 11722 45880 11770 45936
rect 11661 45875 11770 45880
rect 7613 45802 7679 45805
rect 11710 45804 11770 45875
rect 12630 45936 12831 45938
rect 12630 45880 12770 45936
rect 12826 45880 12831 45936
rect 12630 45878 12831 45880
rect 11702 45802 11708 45804
rect 7613 45800 11708 45802
rect 7613 45744 7618 45800
rect 7674 45744 11708 45800
rect 7613 45742 11708 45744
rect 7613 45739 7679 45742
rect 11702 45740 11708 45742
rect 11772 45740 11778 45804
rect 5878 45728 6194 45729
rect 5878 45664 5884 45728
rect 5948 45664 5964 45728
rect 6028 45664 6044 45728
rect 6108 45664 6124 45728
rect 6188 45664 6194 45728
rect 5878 45663 6194 45664
rect 8993 45530 9059 45533
rect 9821 45530 9887 45533
rect 12630 45530 12690 45878
rect 12765 45875 12831 45878
rect 13734 45936 13935 45938
rect 13734 45880 13874 45936
rect 13930 45880 13935 45936
rect 13734 45878 13935 45880
rect 8993 45528 12690 45530
rect 8993 45472 8998 45528
rect 9054 45472 9826 45528
rect 9882 45472 12690 45528
rect 8993 45470 12690 45472
rect 8993 45467 9059 45470
rect 9821 45467 9887 45470
rect 5681 45394 5747 45397
rect 13734 45394 13794 45878
rect 13869 45875 13935 45878
rect 49059 45936 49125 45941
rect 49059 45880 49064 45936
rect 49120 45880 49125 45936
rect 49059 45875 49125 45880
rect 51129 45938 51195 45941
rect 51129 45936 52066 45938
rect 51129 45880 51134 45936
rect 51190 45880 52066 45936
rect 51129 45878 52066 45880
rect 51129 45875 51195 45878
rect 49062 45802 49122 45875
rect 52006 45802 52066 45878
rect 5681 45392 13794 45394
rect 5681 45336 5686 45392
rect 5742 45336 13794 45392
rect 5681 45334 13794 45336
rect 29190 45742 51882 45802
rect 52006 45742 58230 45802
rect 5681 45331 5747 45334
rect 3000 45258 3800 45288
rect 4301 45258 4367 45261
rect 3000 45256 4367 45258
rect 3000 45200 4306 45256
rect 4362 45200 4367 45256
rect 3000 45198 4367 45200
rect 3000 45168 3800 45198
rect 4301 45195 4367 45198
rect 11702 45196 11708 45260
rect 11772 45258 11778 45260
rect 29190 45258 29250 45742
rect 47081 45666 47147 45669
rect 47955 45666 48021 45669
rect 47081 45664 48570 45666
rect 47081 45608 47086 45664
rect 47142 45608 47960 45664
rect 48016 45608 48570 45664
rect 47081 45606 48570 45608
rect 47081 45603 47147 45606
rect 47955 45603 48021 45606
rect 11772 45198 29250 45258
rect 11772 45196 11778 45198
rect 6614 45184 6930 45185
rect 6614 45120 6620 45184
rect 6684 45120 6700 45184
rect 6764 45120 6780 45184
rect 6844 45120 6860 45184
rect 6924 45120 6930 45184
rect 6614 45119 6930 45120
rect 48510 45122 48570 45606
rect 51822 45258 51882 45742
rect 58170 45394 58230 45742
rect 86470 45728 86786 45729
rect 86470 45664 86476 45728
rect 86540 45664 86556 45728
rect 86620 45664 86636 45728
rect 86700 45664 86716 45728
rect 86780 45664 86786 45728
rect 86470 45663 86786 45664
rect 85997 45394 86063 45397
rect 58170 45392 86063 45394
rect 58170 45336 86002 45392
rect 86058 45336 86063 45392
rect 58170 45334 86063 45336
rect 85997 45331 86063 45334
rect 86181 45258 86247 45261
rect 51822 45256 86247 45258
rect 51822 45200 86186 45256
rect 86242 45200 86247 45256
rect 51822 45198 86247 45200
rect 86181 45195 86247 45198
rect 88205 45258 88271 45261
rect 89200 45258 90000 45288
rect 88205 45256 90000 45258
rect 88205 45200 88210 45256
rect 88266 45200 90000 45256
rect 88205 45198 90000 45200
rect 88205 45195 88271 45198
rect 87206 45184 87522 45185
rect 85629 45122 85695 45125
rect 48510 45120 85695 45122
rect 48510 45064 85634 45120
rect 85690 45064 85695 45120
rect 87206 45120 87212 45184
rect 87276 45120 87292 45184
rect 87356 45120 87372 45184
rect 87436 45120 87452 45184
rect 87516 45120 87522 45184
rect 89200 45168 90000 45198
rect 87206 45119 87522 45120
rect 48510 45062 85695 45064
rect 85629 45059 85695 45062
rect 8533 44714 8599 44717
rect 8533 44712 10114 44714
rect 8533 44656 8538 44712
rect 8594 44656 10114 44712
rect 8533 44654 10114 44656
rect 8533 44651 8599 44654
rect 5878 44640 6194 44641
rect 3000 44578 3800 44608
rect 4209 44578 4275 44581
rect 3000 44576 4275 44578
rect 3000 44520 4214 44576
rect 4270 44520 4275 44576
rect 5878 44576 5884 44640
rect 5948 44576 5964 44640
rect 6028 44576 6044 44640
rect 6108 44576 6124 44640
rect 6188 44576 6194 44640
rect 10054 44616 10114 44654
rect 46118 44654 47466 44714
rect 46118 44646 46178 44654
rect 45596 44586 46178 44646
rect 47406 44616 47466 44654
rect 83605 44646 83671 44649
rect 83132 44644 83671 44646
rect 83132 44588 83610 44644
rect 83666 44588 83671 44644
rect 83132 44586 83671 44588
rect 83605 44583 83671 44586
rect 86470 44640 86786 44641
rect 5878 44575 6194 44576
rect 86470 44576 86476 44640
rect 86540 44576 86556 44640
rect 86620 44576 86636 44640
rect 86700 44576 86716 44640
rect 86780 44576 86786 44640
rect 86470 44575 86786 44576
rect 88205 44578 88271 44581
rect 89200 44578 90000 44608
rect 88205 44576 90000 44578
rect 3000 44518 4275 44520
rect 3000 44488 3800 44518
rect 4209 44515 4275 44518
rect 88205 44520 88210 44576
rect 88266 44520 90000 44576
rect 88205 44518 90000 44520
rect 88205 44515 88271 44518
rect 89200 44488 90000 44518
rect 6614 44096 6930 44097
rect 6614 44032 6620 44096
rect 6684 44032 6700 44096
rect 6764 44032 6780 44096
rect 6844 44032 6860 44096
rect 6924 44032 6930 44096
rect 6614 44031 6930 44032
rect 87206 44096 87522 44097
rect 87206 44032 87212 44096
rect 87276 44032 87292 44096
rect 87356 44032 87372 44096
rect 87436 44032 87452 44096
rect 87516 44032 87522 44096
rect 87206 44031 87522 44032
rect 88205 43898 88271 43901
rect 89200 43898 90000 43928
rect 88205 43896 90000 43898
rect 88205 43840 88210 43896
rect 88266 43840 90000 43896
rect 88205 43838 90000 43840
rect 88205 43835 88271 43838
rect 89200 43808 90000 43838
rect 46118 43566 47466 43626
rect 46118 43558 46178 43566
rect 5878 43552 6194 43553
rect 5878 43488 5884 43552
rect 5948 43488 5964 43552
rect 6028 43488 6044 43552
rect 6108 43488 6124 43552
rect 6188 43488 6194 43552
rect 5878 43487 6194 43488
rect 8533 43490 8599 43493
rect 10054 43490 10114 43528
rect 45596 43498 46178 43558
rect 47406 43528 47466 43566
rect 83132 43498 83346 43558
rect 8533 43488 10114 43490
rect 8533 43432 8538 43488
rect 8594 43432 10114 43488
rect 8533 43430 10114 43432
rect 83286 43490 83346 43498
rect 86470 43552 86786 43553
rect 85813 43490 85879 43493
rect 83286 43488 85879 43490
rect 83286 43432 85818 43488
rect 85874 43432 85879 43488
rect 86470 43488 86476 43552
rect 86540 43488 86556 43552
rect 86620 43488 86636 43552
rect 86700 43488 86716 43552
rect 86780 43488 86786 43552
rect 86470 43487 86786 43488
rect 83286 43430 85879 43432
rect 8533 43427 8599 43430
rect 85813 43427 85879 43430
rect 3000 43218 3800 43248
rect 4117 43218 4183 43221
rect 3000 43216 4183 43218
rect 3000 43160 4122 43216
rect 4178 43160 4183 43216
rect 3000 43158 4183 43160
rect 3000 43128 3800 43158
rect 4117 43155 4183 43158
rect 88205 43218 88271 43221
rect 89200 43218 90000 43248
rect 88205 43216 90000 43218
rect 88205 43160 88210 43216
rect 88266 43160 90000 43216
rect 88205 43158 90000 43160
rect 88205 43155 88271 43158
rect 89200 43128 90000 43158
rect 6614 43008 6930 43009
rect 6614 42944 6620 43008
rect 6684 42944 6700 43008
rect 6764 42944 6780 43008
rect 6844 42944 6860 43008
rect 6924 42944 6930 43008
rect 6614 42943 6930 42944
rect 87206 43008 87522 43009
rect 87206 42944 87212 43008
rect 87276 42944 87292 43008
rect 87356 42944 87372 43008
rect 87436 42944 87452 43008
rect 87516 42944 87522 43008
rect 87206 42943 87522 42944
rect 3000 42538 3800 42568
rect 4117 42538 4183 42541
rect 3000 42536 4183 42538
rect 3000 42480 4122 42536
rect 4178 42480 4183 42536
rect 3000 42478 4183 42480
rect 3000 42448 3800 42478
rect 4117 42475 4183 42478
rect 8533 42538 8599 42541
rect 85813 42538 85879 42541
rect 8533 42536 10114 42538
rect 8533 42480 8538 42536
rect 8594 42480 10114 42536
rect 8533 42478 10114 42480
rect 8533 42475 8599 42478
rect 5878 42464 6194 42465
rect 5878 42400 5884 42464
rect 5948 42400 5964 42464
rect 6028 42400 6044 42464
rect 6108 42400 6124 42464
rect 6188 42400 6194 42464
rect 10054 42440 10114 42478
rect 46118 42478 47466 42538
rect 46118 42470 46178 42478
rect 45596 42410 46178 42470
rect 47406 42440 47466 42478
rect 83286 42536 85879 42538
rect 83286 42480 85818 42536
rect 85874 42480 85879 42536
rect 83286 42478 85879 42480
rect 83286 42470 83346 42478
rect 85813 42475 85879 42478
rect 88205 42538 88271 42541
rect 89200 42538 90000 42568
rect 88205 42536 90000 42538
rect 88205 42480 88210 42536
rect 88266 42480 90000 42536
rect 88205 42478 90000 42480
rect 88205 42475 88271 42478
rect 83132 42410 83346 42470
rect 86470 42464 86786 42465
rect 5878 42399 6194 42400
rect 86470 42400 86476 42464
rect 86540 42400 86556 42464
rect 86620 42400 86636 42464
rect 86700 42400 86716 42464
rect 86780 42400 86786 42464
rect 89200 42448 90000 42478
rect 86470 42399 86786 42400
rect 6614 41920 6930 41921
rect 6614 41856 6620 41920
rect 6684 41856 6700 41920
rect 6764 41856 6780 41920
rect 6844 41856 6860 41920
rect 6924 41856 6930 41920
rect 6614 41855 6930 41856
rect 87206 41920 87522 41921
rect 87206 41856 87212 41920
rect 87276 41856 87292 41920
rect 87356 41856 87372 41920
rect 87436 41856 87452 41920
rect 87516 41856 87522 41920
rect 87206 41855 87522 41856
rect 5405 41586 5471 41589
rect 87561 41586 87627 41589
rect 5405 41584 10114 41586
rect 5405 41528 5410 41584
rect 5466 41528 10114 41584
rect 5405 41526 10114 41528
rect 5405 41523 5471 41526
rect 5878 41376 6194 41377
rect 5878 41312 5884 41376
rect 5948 41312 5964 41376
rect 6028 41312 6044 41376
rect 6108 41312 6124 41376
rect 6188 41312 6194 41376
rect 10054 41352 10114 41526
rect 83654 41584 87627 41586
rect 83654 41528 87566 41584
rect 87622 41528 87627 41584
rect 83654 41526 87627 41528
rect 46118 41390 47466 41450
rect 46118 41382 46178 41390
rect 45596 41322 46178 41382
rect 47406 41352 47466 41390
rect 83654 41382 83714 41526
rect 87561 41523 87627 41526
rect 83132 41322 83714 41382
rect 86470 41376 86786 41377
rect 5878 41311 6194 41312
rect 86470 41312 86476 41376
rect 86540 41312 86556 41376
rect 86620 41312 86636 41376
rect 86700 41312 86716 41376
rect 86780 41312 86786 41376
rect 86470 41311 86786 41312
rect 3000 41178 3800 41208
rect 4117 41178 4183 41181
rect 3000 41176 4183 41178
rect 3000 41120 4122 41176
rect 4178 41120 4183 41176
rect 3000 41118 4183 41120
rect 3000 41088 3800 41118
rect 4117 41115 4183 41118
rect 88205 41178 88271 41181
rect 89200 41178 90000 41208
rect 88205 41176 90000 41178
rect 88205 41120 88210 41176
rect 88266 41120 90000 41176
rect 88205 41118 90000 41120
rect 88205 41115 88271 41118
rect 89200 41088 90000 41118
rect 6614 40832 6930 40833
rect 6614 40768 6620 40832
rect 6684 40768 6700 40832
rect 6764 40768 6780 40832
rect 6844 40768 6860 40832
rect 6924 40768 6930 40832
rect 6614 40767 6930 40768
rect 87206 40832 87522 40833
rect 87206 40768 87212 40832
rect 87276 40768 87292 40832
rect 87356 40768 87372 40832
rect 87436 40768 87452 40832
rect 87516 40768 87522 40832
rect 87206 40767 87522 40768
rect 3000 40498 3800 40528
rect 3933 40498 3999 40501
rect 87929 40498 87995 40501
rect 3000 40496 3999 40498
rect 3000 40440 3938 40496
rect 3994 40440 3999 40496
rect 3000 40438 3999 40440
rect 3000 40408 3800 40438
rect 3933 40435 3999 40438
rect 83654 40496 87995 40498
rect 83654 40440 87934 40496
rect 87990 40440 87995 40496
rect 83654 40438 87995 40440
rect 8533 40362 8599 40365
rect 8533 40360 10114 40362
rect 8533 40304 8538 40360
rect 8594 40304 10114 40360
rect 8533 40302 10114 40304
rect 8533 40299 8599 40302
rect 5878 40288 6194 40289
rect 5878 40224 5884 40288
rect 5948 40224 5964 40288
rect 6028 40224 6044 40288
rect 6108 40224 6124 40288
rect 6188 40224 6194 40288
rect 10054 40264 10114 40302
rect 45934 40302 47466 40362
rect 45934 40294 45994 40302
rect 45596 40234 45994 40294
rect 47406 40264 47466 40302
rect 83654 40294 83714 40438
rect 87929 40435 87995 40438
rect 88205 40498 88271 40501
rect 89200 40498 90000 40528
rect 88205 40496 90000 40498
rect 88205 40440 88210 40496
rect 88266 40440 90000 40496
rect 88205 40438 90000 40440
rect 88205 40435 88271 40438
rect 89200 40408 90000 40438
rect 83132 40234 83714 40294
rect 86470 40288 86786 40289
rect 5878 40223 6194 40224
rect 86470 40224 86476 40288
rect 86540 40224 86556 40288
rect 86620 40224 86636 40288
rect 86700 40224 86716 40288
rect 86780 40224 86786 40288
rect 86470 40223 86786 40224
rect 6614 39744 6930 39745
rect 6614 39680 6620 39744
rect 6684 39680 6700 39744
rect 6764 39680 6780 39744
rect 6844 39680 6860 39744
rect 6924 39680 6930 39744
rect 6614 39679 6930 39680
rect 87206 39744 87522 39745
rect 87206 39680 87212 39744
rect 87276 39680 87292 39744
rect 87356 39680 87372 39744
rect 87436 39680 87452 39744
rect 87516 39680 87522 39744
rect 87206 39679 87522 39680
rect 87561 39410 87627 39413
rect 83654 39408 87627 39410
rect 83654 39352 87566 39408
rect 87622 39352 87627 39408
rect 83654 39350 87627 39352
rect 8533 39274 8599 39277
rect 8533 39272 10114 39274
rect 8533 39216 8538 39272
rect 8594 39216 10114 39272
rect 8533 39214 10114 39216
rect 8533 39211 8599 39214
rect 5878 39200 6194 39201
rect 3000 39138 3800 39168
rect 4209 39138 4275 39141
rect 3000 39136 4275 39138
rect 3000 39080 4214 39136
rect 4270 39080 4275 39136
rect 5878 39136 5884 39200
rect 5948 39136 5964 39200
rect 6028 39136 6044 39200
rect 6108 39136 6124 39200
rect 6188 39136 6194 39200
rect 10054 39176 10114 39214
rect 46118 39214 47466 39274
rect 46118 39206 46178 39214
rect 45596 39146 46178 39206
rect 47406 39176 47466 39214
rect 83654 39206 83714 39350
rect 87561 39347 87627 39350
rect 83132 39146 83714 39206
rect 86470 39200 86786 39201
rect 5878 39135 6194 39136
rect 86470 39136 86476 39200
rect 86540 39136 86556 39200
rect 86620 39136 86636 39200
rect 86700 39136 86716 39200
rect 86780 39136 86786 39200
rect 86470 39135 86786 39136
rect 88205 39138 88271 39141
rect 89200 39138 90000 39168
rect 88205 39136 90000 39138
rect 3000 39078 4275 39080
rect 3000 39048 3800 39078
rect 4209 39075 4275 39078
rect 88205 39080 88210 39136
rect 88266 39080 90000 39136
rect 88205 39078 90000 39080
rect 88205 39075 88271 39078
rect 89200 39048 90000 39078
rect 6614 38656 6930 38657
rect 6614 38592 6620 38656
rect 6684 38592 6700 38656
rect 6764 38592 6780 38656
rect 6844 38592 6860 38656
rect 6924 38592 6930 38656
rect 6614 38591 6930 38592
rect 87206 38656 87522 38657
rect 87206 38592 87212 38656
rect 87276 38592 87292 38656
rect 87356 38592 87372 38656
rect 87436 38592 87452 38656
rect 87516 38592 87522 38656
rect 87206 38591 87522 38592
rect 46118 38126 47466 38186
rect 46118 38118 46178 38126
rect 5878 38112 6194 38113
rect 5878 38048 5884 38112
rect 5948 38048 5964 38112
rect 6028 38048 6044 38112
rect 6108 38048 6124 38112
rect 6188 38048 6194 38112
rect 5878 38047 6194 38048
rect 8533 38050 8599 38053
rect 10054 38050 10114 38088
rect 45596 38058 46178 38118
rect 47406 38088 47466 38126
rect 83132 38058 83346 38118
rect 8533 38048 10114 38050
rect 8533 37992 8538 38048
rect 8594 37992 10114 38048
rect 8533 37990 10114 37992
rect 83286 38050 83346 38058
rect 86470 38112 86786 38113
rect 85813 38050 85879 38053
rect 83286 38048 85879 38050
rect 83286 37992 85818 38048
rect 85874 37992 85879 38048
rect 86470 38048 86476 38112
rect 86540 38048 86556 38112
rect 86620 38048 86636 38112
rect 86700 38048 86716 38112
rect 86780 38048 86786 38112
rect 86470 38047 86786 38048
rect 83286 37990 85879 37992
rect 8533 37987 8599 37990
rect 85813 37987 85879 37990
rect 3000 37778 3800 37808
rect 4209 37778 4275 37781
rect 3000 37776 4275 37778
rect 3000 37720 4214 37776
rect 4270 37720 4275 37776
rect 3000 37718 4275 37720
rect 3000 37688 3800 37718
rect 4209 37715 4275 37718
rect 88205 37778 88271 37781
rect 89200 37778 90000 37808
rect 88205 37776 90000 37778
rect 88205 37720 88210 37776
rect 88266 37720 90000 37776
rect 88205 37718 90000 37720
rect 88205 37715 88271 37718
rect 89200 37688 90000 37718
rect 6614 37568 6930 37569
rect 6614 37504 6620 37568
rect 6684 37504 6700 37568
rect 6764 37504 6780 37568
rect 6844 37504 6860 37568
rect 6924 37504 6930 37568
rect 6614 37503 6930 37504
rect 87206 37568 87522 37569
rect 87206 37504 87212 37568
rect 87276 37504 87292 37568
rect 87356 37504 87372 37568
rect 87436 37504 87452 37568
rect 87516 37504 87522 37568
rect 87206 37503 87522 37504
rect 3000 37098 3800 37128
rect 4117 37098 4183 37101
rect 3000 37096 4183 37098
rect 3000 37040 4122 37096
rect 4178 37040 4183 37096
rect 3000 37038 4183 37040
rect 3000 37008 3800 37038
rect 4117 37035 4183 37038
rect 8533 37098 8599 37101
rect 85813 37098 85879 37101
rect 8533 37096 10114 37098
rect 8533 37040 8538 37096
rect 8594 37040 10114 37096
rect 8533 37038 10114 37040
rect 8533 37035 8599 37038
rect 5878 37024 6194 37025
rect 5878 36960 5884 37024
rect 5948 36960 5964 37024
rect 6028 36960 6044 37024
rect 6108 36960 6124 37024
rect 6188 36960 6194 37024
rect 10054 37000 10114 37038
rect 46118 37038 47466 37098
rect 46118 37030 46178 37038
rect 45596 36970 46178 37030
rect 47406 37000 47466 37038
rect 83286 37096 85879 37098
rect 83286 37040 85818 37096
rect 85874 37040 85879 37096
rect 83286 37038 85879 37040
rect 83286 37030 83346 37038
rect 85813 37035 85879 37038
rect 88205 37098 88271 37101
rect 89200 37098 90000 37128
rect 88205 37096 90000 37098
rect 88205 37040 88210 37096
rect 88266 37040 90000 37096
rect 88205 37038 90000 37040
rect 88205 37035 88271 37038
rect 83132 36970 83346 37030
rect 86470 37024 86786 37025
rect 5878 36959 6194 36960
rect 86470 36960 86476 37024
rect 86540 36960 86556 37024
rect 86620 36960 86636 37024
rect 86700 36960 86716 37024
rect 86780 36960 86786 37024
rect 89200 37008 90000 37038
rect 86470 36959 86786 36960
rect 6614 36480 6930 36481
rect 6614 36416 6620 36480
rect 6684 36416 6700 36480
rect 6764 36416 6780 36480
rect 6844 36416 6860 36480
rect 6924 36416 6930 36480
rect 6614 36415 6930 36416
rect 87206 36480 87522 36481
rect 87206 36416 87212 36480
rect 87276 36416 87292 36480
rect 87356 36416 87372 36480
rect 87436 36416 87452 36480
rect 87516 36416 87522 36480
rect 87206 36415 87522 36416
rect 5405 36146 5471 36149
rect 5405 36144 10114 36146
rect 5405 36088 5410 36144
rect 5466 36088 10114 36144
rect 5405 36086 10114 36088
rect 5405 36083 5471 36086
rect 5878 35936 6194 35937
rect 5878 35872 5884 35936
rect 5948 35872 5964 35936
rect 6028 35872 6044 35936
rect 6108 35872 6124 35936
rect 6188 35872 6194 35936
rect 10054 35912 10114 36086
rect 84801 36010 84867 36013
rect 46118 35950 47466 36010
rect 46118 35942 46178 35950
rect 45596 35882 46178 35942
rect 47406 35912 47466 35950
rect 83286 36008 84867 36010
rect 83286 35952 84806 36008
rect 84862 35952 84867 36008
rect 83286 35950 84867 35952
rect 83286 35942 83346 35950
rect 84801 35947 84867 35950
rect 83132 35882 83346 35942
rect 86470 35936 86786 35937
rect 5878 35871 6194 35872
rect 86470 35872 86476 35936
rect 86540 35872 86556 35936
rect 86620 35872 86636 35936
rect 86700 35872 86716 35936
rect 86780 35872 86786 35936
rect 86470 35871 86786 35872
rect 3000 35738 3800 35768
rect 4117 35738 4183 35741
rect 3000 35736 4183 35738
rect 3000 35680 4122 35736
rect 4178 35680 4183 35736
rect 3000 35678 4183 35680
rect 3000 35648 3800 35678
rect 4117 35675 4183 35678
rect 88573 35738 88639 35741
rect 89200 35738 90000 35768
rect 88573 35736 90000 35738
rect 88573 35680 88578 35736
rect 88634 35680 90000 35736
rect 88573 35678 90000 35680
rect 88573 35675 88639 35678
rect 89200 35648 90000 35678
rect 6614 35392 6930 35393
rect 6614 35328 6620 35392
rect 6684 35328 6700 35392
rect 6764 35328 6780 35392
rect 6844 35328 6860 35392
rect 6924 35328 6930 35392
rect 6614 35327 6930 35328
rect 87206 35392 87522 35393
rect 87206 35328 87212 35392
rect 87276 35328 87292 35392
rect 87356 35328 87372 35392
rect 87436 35328 87452 35392
rect 87516 35328 87522 35392
rect 87206 35327 87522 35328
rect 3000 35058 3800 35088
rect 4209 35058 4275 35061
rect 3000 35056 4275 35058
rect 3000 35000 4214 35056
rect 4270 35000 4275 35056
rect 3000 34998 4275 35000
rect 3000 34968 3800 34998
rect 4209 34995 4275 34998
rect 88205 35058 88271 35061
rect 89200 35058 90000 35088
rect 88205 35056 90000 35058
rect 88205 35000 88210 35056
rect 88266 35000 90000 35056
rect 88205 34998 90000 35000
rect 88205 34995 88271 34998
rect 89200 34968 90000 34998
rect 8533 34922 8599 34925
rect 85813 34922 85879 34925
rect 8533 34920 10114 34922
rect 8533 34864 8538 34920
rect 8594 34864 10114 34920
rect 8533 34862 10114 34864
rect 8533 34859 8599 34862
rect 5878 34848 6194 34849
rect 5878 34784 5884 34848
rect 5948 34784 5964 34848
rect 6028 34784 6044 34848
rect 6108 34784 6124 34848
rect 6188 34784 6194 34848
rect 10054 34824 10114 34862
rect 46118 34862 47466 34922
rect 46118 34854 46178 34862
rect 45596 34794 46178 34854
rect 47406 34824 47466 34862
rect 83286 34920 85879 34922
rect 83286 34864 85818 34920
rect 85874 34864 85879 34920
rect 83286 34862 85879 34864
rect 83286 34854 83346 34862
rect 85813 34859 85879 34862
rect 83132 34794 83346 34854
rect 86470 34848 86786 34849
rect 5878 34783 6194 34784
rect 86470 34784 86476 34848
rect 86540 34784 86556 34848
rect 86620 34784 86636 34848
rect 86700 34784 86716 34848
rect 86780 34784 86786 34848
rect 86470 34783 86786 34784
rect 6614 34304 6930 34305
rect 6614 34240 6620 34304
rect 6684 34240 6700 34304
rect 6764 34240 6780 34304
rect 6844 34240 6860 34304
rect 6924 34240 6930 34304
rect 6614 34239 6930 34240
rect 87206 34304 87522 34305
rect 87206 34240 87212 34304
rect 87276 34240 87292 34304
rect 87356 34240 87372 34304
rect 87436 34240 87452 34304
rect 87516 34240 87522 34304
rect 87206 34239 87522 34240
rect 8533 33834 8599 33837
rect 85813 33834 85879 33837
rect 8533 33832 10114 33834
rect 8533 33776 8538 33832
rect 8594 33776 10114 33832
rect 8533 33774 10114 33776
rect 8533 33771 8599 33774
rect 5878 33760 6194 33761
rect 3000 33698 3800 33728
rect 4209 33698 4275 33701
rect 3000 33696 4275 33698
rect 3000 33640 4214 33696
rect 4270 33640 4275 33696
rect 5878 33696 5884 33760
rect 5948 33696 5964 33760
rect 6028 33696 6044 33760
rect 6108 33696 6124 33760
rect 6188 33696 6194 33760
rect 10054 33736 10114 33774
rect 46118 33774 47466 33834
rect 46118 33766 46178 33774
rect 45596 33706 46178 33766
rect 47406 33736 47466 33774
rect 83286 33832 85879 33834
rect 83286 33776 85818 33832
rect 85874 33776 85879 33832
rect 83286 33774 85879 33776
rect 83286 33766 83346 33774
rect 85813 33771 85879 33774
rect 83132 33706 83346 33766
rect 86470 33760 86786 33761
rect 5878 33695 6194 33696
rect 86470 33696 86476 33760
rect 86540 33696 86556 33760
rect 86620 33696 86636 33760
rect 86700 33696 86716 33760
rect 86780 33696 86786 33760
rect 86470 33695 86786 33696
rect 88205 33698 88271 33701
rect 89200 33698 90000 33728
rect 88205 33696 90000 33698
rect 3000 33638 4275 33640
rect 3000 33608 3800 33638
rect 4209 33635 4275 33638
rect 88205 33640 88210 33696
rect 88266 33640 90000 33696
rect 88205 33638 90000 33640
rect 88205 33635 88271 33638
rect 89200 33608 90000 33638
rect 6614 33216 6930 33217
rect 6614 33152 6620 33216
rect 6684 33152 6700 33216
rect 6764 33152 6780 33216
rect 6844 33152 6860 33216
rect 6924 33152 6930 33216
rect 6614 33151 6930 33152
rect 87206 33216 87522 33217
rect 87206 33152 87212 33216
rect 87276 33152 87292 33216
rect 87356 33152 87372 33216
rect 87436 33152 87452 33216
rect 87516 33152 87522 33216
rect 87206 33151 87522 33152
rect 46118 32686 47466 32746
rect 46118 32678 46178 32686
rect 5878 32672 6194 32673
rect 5878 32608 5884 32672
rect 5948 32608 5964 32672
rect 6028 32608 6044 32672
rect 6108 32608 6124 32672
rect 6188 32608 6194 32672
rect 5878 32607 6194 32608
rect 8533 32610 8599 32613
rect 10054 32610 10114 32648
rect 45596 32618 46178 32678
rect 47406 32648 47466 32686
rect 83132 32618 83346 32678
rect 8533 32608 10114 32610
rect 8533 32552 8538 32608
rect 8594 32552 10114 32608
rect 8533 32550 10114 32552
rect 83286 32610 83346 32618
rect 86470 32672 86786 32673
rect 85813 32610 85879 32613
rect 83286 32608 85879 32610
rect 83286 32552 85818 32608
rect 85874 32552 85879 32608
rect 86470 32608 86476 32672
rect 86540 32608 86556 32672
rect 86620 32608 86636 32672
rect 86700 32608 86716 32672
rect 86780 32608 86786 32672
rect 86470 32607 86786 32608
rect 83286 32550 85879 32552
rect 8533 32547 8599 32550
rect 85813 32547 85879 32550
rect 3000 32338 3800 32368
rect 4209 32338 4275 32341
rect 3000 32336 4275 32338
rect 3000 32280 4214 32336
rect 4270 32280 4275 32336
rect 3000 32278 4275 32280
rect 3000 32248 3800 32278
rect 4209 32275 4275 32278
rect 88205 32338 88271 32341
rect 89200 32338 90000 32368
rect 88205 32336 90000 32338
rect 88205 32280 88210 32336
rect 88266 32280 90000 32336
rect 88205 32278 90000 32280
rect 88205 32275 88271 32278
rect 89200 32248 90000 32278
rect 6614 32128 6930 32129
rect 6614 32064 6620 32128
rect 6684 32064 6700 32128
rect 6764 32064 6780 32128
rect 6844 32064 6860 32128
rect 6924 32064 6930 32128
rect 6614 32063 6930 32064
rect 87206 32128 87522 32129
rect 87206 32064 87212 32128
rect 87276 32064 87292 32128
rect 87356 32064 87372 32128
rect 87436 32064 87452 32128
rect 87516 32064 87522 32128
rect 87206 32063 87522 32064
rect 3000 31658 3800 31688
rect 4117 31658 4183 31661
rect 3000 31656 4183 31658
rect 3000 31600 4122 31656
rect 4178 31600 4183 31656
rect 3000 31598 4183 31600
rect 3000 31568 3800 31598
rect 4117 31595 4183 31598
rect 8533 31658 8599 31661
rect 85813 31658 85879 31661
rect 8533 31656 10114 31658
rect 8533 31600 8538 31656
rect 8594 31600 10114 31656
rect 8533 31598 10114 31600
rect 8533 31595 8599 31598
rect 5878 31584 6194 31585
rect 5878 31520 5884 31584
rect 5948 31520 5964 31584
rect 6028 31520 6044 31584
rect 6108 31520 6124 31584
rect 6188 31520 6194 31584
rect 10054 31560 10114 31598
rect 46118 31598 47466 31658
rect 46118 31590 46178 31598
rect 45596 31530 46178 31590
rect 47406 31560 47466 31598
rect 83286 31656 85879 31658
rect 83286 31600 85818 31656
rect 85874 31600 85879 31656
rect 83286 31598 85879 31600
rect 83286 31590 83346 31598
rect 85813 31595 85879 31598
rect 88205 31658 88271 31661
rect 89200 31658 90000 31688
rect 88205 31656 90000 31658
rect 88205 31600 88210 31656
rect 88266 31600 90000 31656
rect 88205 31598 90000 31600
rect 88205 31595 88271 31598
rect 83132 31530 83346 31590
rect 86470 31584 86786 31585
rect 5878 31519 6194 31520
rect 86470 31520 86476 31584
rect 86540 31520 86556 31584
rect 86620 31520 86636 31584
rect 86700 31520 86716 31584
rect 86780 31520 86786 31584
rect 89200 31568 90000 31598
rect 86470 31519 86786 31520
rect 6614 31040 6930 31041
rect 6614 30976 6620 31040
rect 6684 30976 6700 31040
rect 6764 30976 6780 31040
rect 6844 30976 6860 31040
rect 6924 30976 6930 31040
rect 6614 30975 6930 30976
rect 87206 31040 87522 31041
rect 87206 30976 87212 31040
rect 87276 30976 87292 31040
rect 87356 30976 87372 31040
rect 87436 30976 87452 31040
rect 87516 30976 87522 31040
rect 87206 30975 87522 30976
rect 84801 30570 84867 30573
rect 46118 30510 47466 30570
rect 46118 30502 46178 30510
rect 5878 30496 6194 30497
rect 5878 30432 5884 30496
rect 5948 30432 5964 30496
rect 6028 30432 6044 30496
rect 6108 30432 6124 30496
rect 6188 30432 6194 30496
rect 5878 30431 6194 30432
rect 3000 30298 3800 30328
rect 4117 30298 4183 30301
rect 3000 30296 4183 30298
rect 3000 30240 4122 30296
rect 4178 30240 4183 30296
rect 3000 30238 4183 30240
rect 3000 30208 3800 30238
rect 4117 30235 4183 30238
rect 5405 30298 5471 30301
rect 10054 30298 10114 30472
rect 45596 30442 46178 30502
rect 47406 30472 47466 30510
rect 83286 30568 84867 30570
rect 83286 30512 84806 30568
rect 84862 30512 84867 30568
rect 83286 30510 84867 30512
rect 83286 30502 83346 30510
rect 84801 30507 84867 30510
rect 83132 30442 83346 30502
rect 86470 30496 86786 30497
rect 86470 30432 86476 30496
rect 86540 30432 86556 30496
rect 86620 30432 86636 30496
rect 86700 30432 86716 30496
rect 86780 30432 86786 30496
rect 86470 30431 86786 30432
rect 5405 30296 10114 30298
rect 5405 30240 5410 30296
rect 5466 30240 10114 30296
rect 5405 30238 10114 30240
rect 88573 30298 88639 30301
rect 89200 30298 90000 30328
rect 88573 30296 90000 30298
rect 88573 30240 88578 30296
rect 88634 30240 90000 30296
rect 88573 30238 90000 30240
rect 5405 30235 5471 30238
rect 88573 30235 88639 30238
rect 89200 30208 90000 30238
rect 6614 29952 6930 29953
rect 6614 29888 6620 29952
rect 6684 29888 6700 29952
rect 6764 29888 6780 29952
rect 6844 29888 6860 29952
rect 6924 29888 6930 29952
rect 6614 29887 6930 29888
rect 87206 29952 87522 29953
rect 87206 29888 87212 29952
rect 87276 29888 87292 29952
rect 87356 29888 87372 29952
rect 87436 29888 87452 29952
rect 87516 29888 87522 29952
rect 87206 29887 87522 29888
rect 3000 29618 3800 29648
rect 4301 29618 4367 29621
rect 3000 29616 4367 29618
rect 3000 29560 4306 29616
rect 4362 29560 4367 29616
rect 3000 29558 4367 29560
rect 3000 29528 3800 29558
rect 4301 29555 4367 29558
rect 88389 29618 88455 29621
rect 89200 29618 90000 29648
rect 88389 29616 90000 29618
rect 88389 29560 88394 29616
rect 88450 29560 90000 29616
rect 88389 29558 90000 29560
rect 88389 29555 88455 29558
rect 89200 29528 90000 29558
rect 8533 29482 8599 29485
rect 85813 29482 85879 29485
rect 8533 29480 10114 29482
rect 8533 29424 8538 29480
rect 8594 29424 10114 29480
rect 8533 29422 10114 29424
rect 8533 29419 8599 29422
rect 5878 29408 6194 29409
rect 5878 29344 5884 29408
rect 5948 29344 5964 29408
rect 6028 29344 6044 29408
rect 6108 29344 6124 29408
rect 6188 29344 6194 29408
rect 10054 29384 10114 29422
rect 46118 29422 47466 29482
rect 46118 29414 46178 29422
rect 45596 29354 46178 29414
rect 47406 29384 47466 29422
rect 83286 29480 85879 29482
rect 83286 29424 85818 29480
rect 85874 29424 85879 29480
rect 83286 29422 85879 29424
rect 83286 29414 83346 29422
rect 85813 29419 85879 29422
rect 83132 29354 83346 29414
rect 86470 29408 86786 29409
rect 5878 29343 6194 29344
rect 86470 29344 86476 29408
rect 86540 29344 86556 29408
rect 86620 29344 86636 29408
rect 86700 29344 86716 29408
rect 86780 29344 86786 29408
rect 86470 29343 86786 29344
rect 6614 28864 6930 28865
rect 6614 28800 6620 28864
rect 6684 28800 6700 28864
rect 6764 28800 6780 28864
rect 6844 28800 6860 28864
rect 6924 28800 6930 28864
rect 6614 28799 6930 28800
rect 87206 28864 87522 28865
rect 87206 28800 87212 28864
rect 87276 28800 87292 28864
rect 87356 28800 87372 28864
rect 87436 28800 87452 28864
rect 87516 28800 87522 28864
rect 87206 28799 87522 28800
rect 8533 28394 8599 28397
rect 85813 28394 85879 28397
rect 8533 28392 10114 28394
rect 8533 28336 8538 28392
rect 8594 28336 10114 28392
rect 8533 28334 10114 28336
rect 8533 28331 8599 28334
rect 5878 28320 6194 28321
rect 3000 28258 3800 28288
rect 4301 28258 4367 28261
rect 3000 28256 4367 28258
rect 3000 28200 4306 28256
rect 4362 28200 4367 28256
rect 5878 28256 5884 28320
rect 5948 28256 5964 28320
rect 6028 28256 6044 28320
rect 6108 28256 6124 28320
rect 6188 28256 6194 28320
rect 10054 28296 10114 28334
rect 46118 28334 47466 28394
rect 46118 28326 46178 28334
rect 45596 28266 46178 28326
rect 47406 28296 47466 28334
rect 83286 28392 85879 28394
rect 83286 28336 85818 28392
rect 85874 28336 85879 28392
rect 83286 28334 85879 28336
rect 83286 28326 83346 28334
rect 85813 28331 85879 28334
rect 83132 28266 83346 28326
rect 86470 28320 86786 28321
rect 5878 28255 6194 28256
rect 86470 28256 86476 28320
rect 86540 28256 86556 28320
rect 86620 28256 86636 28320
rect 86700 28256 86716 28320
rect 86780 28256 86786 28320
rect 86470 28255 86786 28256
rect 88205 28258 88271 28261
rect 89200 28258 90000 28288
rect 88205 28256 90000 28258
rect 3000 28198 4367 28200
rect 3000 28168 3800 28198
rect 4301 28195 4367 28198
rect 88205 28200 88210 28256
rect 88266 28200 90000 28256
rect 88205 28198 90000 28200
rect 88205 28195 88271 28198
rect 89200 28168 90000 28198
rect 6614 27776 6930 27777
rect 6614 27712 6620 27776
rect 6684 27712 6700 27776
rect 6764 27712 6780 27776
rect 6844 27712 6860 27776
rect 6924 27712 6930 27776
rect 6614 27711 6930 27712
rect 87206 27776 87522 27777
rect 87206 27712 87212 27776
rect 87276 27712 87292 27776
rect 87356 27712 87372 27776
rect 87436 27712 87452 27776
rect 87516 27712 87522 27776
rect 87206 27711 87522 27712
rect 46118 27246 47466 27306
rect 46118 27238 46178 27246
rect 5878 27232 6194 27233
rect 5878 27168 5884 27232
rect 5948 27168 5964 27232
rect 6028 27168 6044 27232
rect 6108 27168 6124 27232
rect 6188 27168 6194 27232
rect 5878 27167 6194 27168
rect 8533 27170 8599 27173
rect 10054 27170 10114 27208
rect 45596 27178 46178 27238
rect 47406 27208 47466 27246
rect 83132 27178 83346 27238
rect 8533 27168 10114 27170
rect 8533 27112 8538 27168
rect 8594 27112 10114 27168
rect 8533 27110 10114 27112
rect 83286 27170 83346 27178
rect 86470 27232 86786 27233
rect 85813 27170 85879 27173
rect 83286 27168 85879 27170
rect 83286 27112 85818 27168
rect 85874 27112 85879 27168
rect 86470 27168 86476 27232
rect 86540 27168 86556 27232
rect 86620 27168 86636 27232
rect 86700 27168 86716 27232
rect 86780 27168 86786 27232
rect 86470 27167 86786 27168
rect 83286 27110 85879 27112
rect 8533 27107 8599 27110
rect 85813 27107 85879 27110
rect 3000 26898 3800 26928
rect 4301 26898 4367 26901
rect 3000 26896 4367 26898
rect 3000 26840 4306 26896
rect 4362 26840 4367 26896
rect 3000 26838 4367 26840
rect 3000 26808 3800 26838
rect 4301 26835 4367 26838
rect 88389 26898 88455 26901
rect 89200 26898 90000 26928
rect 88389 26896 90000 26898
rect 88389 26840 88394 26896
rect 88450 26840 90000 26896
rect 88389 26838 90000 26840
rect 88389 26835 88455 26838
rect 89200 26808 90000 26838
rect 6614 26688 6930 26689
rect 6614 26624 6620 26688
rect 6684 26624 6700 26688
rect 6764 26624 6780 26688
rect 6844 26624 6860 26688
rect 6924 26624 6930 26688
rect 6614 26623 6930 26624
rect 87206 26688 87522 26689
rect 87206 26624 87212 26688
rect 87276 26624 87292 26688
rect 87356 26624 87372 26688
rect 87436 26624 87452 26688
rect 87516 26624 87522 26688
rect 87206 26623 87522 26624
rect 87561 26354 87627 26357
rect 83654 26352 87627 26354
rect 83654 26296 87566 26352
rect 87622 26296 87627 26352
rect 83654 26294 87627 26296
rect 3000 26218 3800 26248
rect 4301 26218 4367 26221
rect 3000 26216 4367 26218
rect 3000 26160 4306 26216
rect 4362 26160 4367 26216
rect 3000 26158 4367 26160
rect 3000 26128 3800 26158
rect 4301 26155 4367 26158
rect 8533 26218 8599 26221
rect 8533 26216 10114 26218
rect 8533 26160 8538 26216
rect 8594 26160 10114 26216
rect 8533 26158 10114 26160
rect 8533 26155 8599 26158
rect 5878 26144 6194 26145
rect 5878 26080 5884 26144
rect 5948 26080 5964 26144
rect 6028 26080 6044 26144
rect 6108 26080 6124 26144
rect 6188 26080 6194 26144
rect 10054 26120 10114 26158
rect 46118 26158 47466 26218
rect 46118 26150 46178 26158
rect 45596 26090 46178 26150
rect 47406 26120 47466 26158
rect 83654 26150 83714 26294
rect 87561 26291 87627 26294
rect 88205 26218 88271 26221
rect 89200 26218 90000 26248
rect 88205 26216 90000 26218
rect 88205 26160 88210 26216
rect 88266 26160 90000 26216
rect 88205 26158 90000 26160
rect 88205 26155 88271 26158
rect 83132 26090 83714 26150
rect 86470 26144 86786 26145
rect 5878 26079 6194 26080
rect 86470 26080 86476 26144
rect 86540 26080 86556 26144
rect 86620 26080 86636 26144
rect 86700 26080 86716 26144
rect 86780 26080 86786 26144
rect 89200 26128 90000 26158
rect 86470 26079 86786 26080
rect 6614 25600 6930 25601
rect 6614 25536 6620 25600
rect 6684 25536 6700 25600
rect 6764 25536 6780 25600
rect 6844 25536 6860 25600
rect 6924 25536 6930 25600
rect 6614 25535 6930 25536
rect 87206 25600 87522 25601
rect 87206 25536 87212 25600
rect 87276 25536 87292 25600
rect 87356 25536 87372 25600
rect 87436 25536 87452 25600
rect 87516 25536 87522 25600
rect 87206 25535 87522 25536
rect 5878 25056 6194 25057
rect 5878 24992 5884 25056
rect 5948 24992 5964 25056
rect 6028 24992 6044 25056
rect 6108 24992 6124 25056
rect 6188 24992 6194 25056
rect 5878 24991 6194 24992
rect 3000 24858 3800 24888
rect 4301 24858 4367 24861
rect 3000 24856 4367 24858
rect 3000 24800 4306 24856
rect 4362 24800 4367 24856
rect 3000 24798 4367 24800
rect 3000 24768 3800 24798
rect 4301 24795 4367 24798
rect 5405 24858 5471 24861
rect 10054 24858 10114 25032
rect 45596 25002 46178 25062
rect 46118 24994 46178 25002
rect 47406 24994 47466 25032
rect 83132 25002 83346 25062
rect 46118 24934 47466 24994
rect 83286 24994 83346 25002
rect 86470 25056 86786 25057
rect 84801 24994 84867 24997
rect 83286 24992 84867 24994
rect 83286 24936 84806 24992
rect 84862 24936 84867 24992
rect 86470 24992 86476 25056
rect 86540 24992 86556 25056
rect 86620 24992 86636 25056
rect 86700 24992 86716 25056
rect 86780 24992 86786 25056
rect 86470 24991 86786 24992
rect 83286 24934 84867 24936
rect 84801 24931 84867 24934
rect 5405 24856 10114 24858
rect 5405 24800 5410 24856
rect 5466 24800 10114 24856
rect 5405 24798 10114 24800
rect 88573 24858 88639 24861
rect 89200 24858 90000 24888
rect 88573 24856 90000 24858
rect 88573 24800 88578 24856
rect 88634 24800 90000 24856
rect 88573 24798 90000 24800
rect 5405 24795 5471 24798
rect 88573 24795 88639 24798
rect 89200 24768 90000 24798
rect 6614 24512 6930 24513
rect 6614 24448 6620 24512
rect 6684 24448 6700 24512
rect 6764 24448 6780 24512
rect 6844 24448 6860 24512
rect 6924 24448 6930 24512
rect 6614 24447 6930 24448
rect 87206 24512 87522 24513
rect 87206 24448 87212 24512
rect 87276 24448 87292 24512
rect 87356 24448 87372 24512
rect 87436 24448 87452 24512
rect 87516 24448 87522 24512
rect 87206 24447 87522 24448
rect 3000 24178 3800 24208
rect 4301 24178 4367 24181
rect 87561 24178 87627 24181
rect 3000 24176 4367 24178
rect 3000 24120 4306 24176
rect 4362 24120 4367 24176
rect 3000 24118 4367 24120
rect 3000 24088 3800 24118
rect 4301 24115 4367 24118
rect 83654 24176 87627 24178
rect 83654 24120 87566 24176
rect 87622 24120 87627 24176
rect 83654 24118 87627 24120
rect 8533 24042 8599 24045
rect 8533 24040 10114 24042
rect 8533 23984 8538 24040
rect 8594 23984 10114 24040
rect 8533 23982 10114 23984
rect 8533 23979 8599 23982
rect 5878 23968 6194 23969
rect 5878 23904 5884 23968
rect 5948 23904 5964 23968
rect 6028 23904 6044 23968
rect 6108 23904 6124 23968
rect 6188 23904 6194 23968
rect 10054 23944 10114 23982
rect 46118 23982 47466 24042
rect 46118 23974 46178 23982
rect 45596 23914 46178 23974
rect 47406 23944 47466 23982
rect 83654 23974 83714 24118
rect 87561 24115 87627 24118
rect 88481 24178 88547 24181
rect 89200 24178 90000 24208
rect 88481 24176 90000 24178
rect 88481 24120 88486 24176
rect 88542 24120 90000 24176
rect 88481 24118 90000 24120
rect 88481 24115 88547 24118
rect 89200 24088 90000 24118
rect 83132 23914 83714 23974
rect 86470 23968 86786 23969
rect 5878 23903 6194 23904
rect 86470 23904 86476 23968
rect 86540 23904 86556 23968
rect 86620 23904 86636 23968
rect 86700 23904 86716 23968
rect 86780 23904 86786 23968
rect 86470 23903 86786 23904
rect 6614 23424 6930 23425
rect 6614 23360 6620 23424
rect 6684 23360 6700 23424
rect 6764 23360 6780 23424
rect 6844 23360 6860 23424
rect 6924 23360 6930 23424
rect 6614 23359 6930 23360
rect 87206 23424 87522 23425
rect 87206 23360 87212 23424
rect 87276 23360 87292 23424
rect 87356 23360 87372 23424
rect 87436 23360 87452 23424
rect 87516 23360 87522 23424
rect 87206 23359 87522 23360
rect 8533 22954 8599 22957
rect 85813 22954 85879 22957
rect 8533 22952 10114 22954
rect 8533 22896 8538 22952
rect 8594 22896 10114 22952
rect 8533 22894 10114 22896
rect 8533 22891 8599 22894
rect 5878 22880 6194 22881
rect 3000 22818 3800 22848
rect 4301 22818 4367 22821
rect 3000 22816 4367 22818
rect 3000 22760 4306 22816
rect 4362 22760 4367 22816
rect 5878 22816 5884 22880
rect 5948 22816 5964 22880
rect 6028 22816 6044 22880
rect 6108 22816 6124 22880
rect 6188 22816 6194 22880
rect 10054 22856 10114 22894
rect 46118 22894 47466 22954
rect 46118 22886 46178 22894
rect 45596 22826 46178 22886
rect 47406 22856 47466 22894
rect 83286 22952 85879 22954
rect 83286 22896 85818 22952
rect 85874 22896 85879 22952
rect 83286 22894 85879 22896
rect 83286 22886 83346 22894
rect 85813 22891 85879 22894
rect 83132 22826 83346 22886
rect 86470 22880 86786 22881
rect 5878 22815 6194 22816
rect 86470 22816 86476 22880
rect 86540 22816 86556 22880
rect 86620 22816 86636 22880
rect 86700 22816 86716 22880
rect 86780 22816 86786 22880
rect 86470 22815 86786 22816
rect 88205 22818 88271 22821
rect 89200 22818 90000 22848
rect 88205 22816 90000 22818
rect 3000 22758 4367 22760
rect 3000 22728 3800 22758
rect 4301 22755 4367 22758
rect 88205 22760 88210 22816
rect 88266 22760 90000 22816
rect 88205 22758 90000 22760
rect 88205 22755 88271 22758
rect 89200 22728 90000 22758
rect 6614 22336 6930 22337
rect 6614 22272 6620 22336
rect 6684 22272 6700 22336
rect 6764 22272 6780 22336
rect 6844 22272 6860 22336
rect 6924 22272 6930 22336
rect 6614 22271 6930 22272
rect 87206 22336 87522 22337
rect 87206 22272 87212 22336
rect 87276 22272 87292 22336
rect 87356 22272 87372 22336
rect 87436 22272 87452 22336
rect 87516 22272 87522 22336
rect 87206 22271 87522 22272
rect 46118 21806 47466 21866
rect 46118 21798 46178 21806
rect 5878 21792 6194 21793
rect 5878 21728 5884 21792
rect 5948 21728 5964 21792
rect 6028 21728 6044 21792
rect 6108 21728 6124 21792
rect 6188 21728 6194 21792
rect 5878 21727 6194 21728
rect 8533 21730 8599 21733
rect 10054 21730 10114 21768
rect 45596 21738 46178 21798
rect 47406 21768 47466 21806
rect 83132 21738 83346 21798
rect 8533 21728 10114 21730
rect 8533 21672 8538 21728
rect 8594 21672 10114 21728
rect 8533 21670 10114 21672
rect 83286 21730 83346 21738
rect 86470 21792 86786 21793
rect 85813 21730 85879 21733
rect 83286 21728 85879 21730
rect 83286 21672 85818 21728
rect 85874 21672 85879 21728
rect 86470 21728 86476 21792
rect 86540 21728 86556 21792
rect 86620 21728 86636 21792
rect 86700 21728 86716 21792
rect 86780 21728 86786 21792
rect 86470 21727 86786 21728
rect 83286 21670 85879 21672
rect 8533 21667 8599 21670
rect 85813 21667 85879 21670
rect 3000 21458 3800 21488
rect 4301 21458 4367 21461
rect 3000 21456 4367 21458
rect 3000 21400 4306 21456
rect 4362 21400 4367 21456
rect 3000 21398 4367 21400
rect 3000 21368 3800 21398
rect 4301 21395 4367 21398
rect 88389 21458 88455 21461
rect 89200 21458 90000 21488
rect 88389 21456 90000 21458
rect 88389 21400 88394 21456
rect 88450 21400 90000 21456
rect 88389 21398 90000 21400
rect 88389 21395 88455 21398
rect 89200 21368 90000 21398
rect 6614 21248 6930 21249
rect 6614 21184 6620 21248
rect 6684 21184 6700 21248
rect 6764 21184 6780 21248
rect 6844 21184 6860 21248
rect 6924 21184 6930 21248
rect 6614 21183 6930 21184
rect 87206 21248 87522 21249
rect 87206 21184 87212 21248
rect 87276 21184 87292 21248
rect 87356 21184 87372 21248
rect 87436 21184 87452 21248
rect 87516 21184 87522 21248
rect 87206 21183 87522 21184
rect 5681 20914 5747 20917
rect 5681 20912 10114 20914
rect 5681 20856 5686 20912
rect 5742 20856 10114 20912
rect 5681 20854 10114 20856
rect 5681 20851 5747 20854
rect 3000 20778 3800 20808
rect 4301 20778 4367 20781
rect 3000 20776 4367 20778
rect 3000 20720 4306 20776
rect 4362 20720 4367 20776
rect 3000 20718 4367 20720
rect 3000 20688 3800 20718
rect 4301 20715 4367 20718
rect 5878 20704 6194 20705
rect 5878 20640 5884 20704
rect 5948 20640 5964 20704
rect 6028 20640 6044 20704
rect 6108 20640 6124 20704
rect 6188 20640 6194 20704
rect 10054 20680 10114 20854
rect 84801 20778 84867 20781
rect 46118 20718 47466 20778
rect 46118 20710 46178 20718
rect 45596 20650 46178 20710
rect 47406 20680 47466 20718
rect 83286 20776 84867 20778
rect 83286 20720 84806 20776
rect 84862 20720 84867 20776
rect 83286 20718 84867 20720
rect 83286 20710 83346 20718
rect 84801 20715 84867 20718
rect 88573 20778 88639 20781
rect 89200 20778 90000 20808
rect 88573 20776 90000 20778
rect 88573 20720 88578 20776
rect 88634 20720 90000 20776
rect 88573 20718 90000 20720
rect 88573 20715 88639 20718
rect 83132 20650 83346 20710
rect 86470 20704 86786 20705
rect 5878 20639 6194 20640
rect 86470 20640 86476 20704
rect 86540 20640 86556 20704
rect 86620 20640 86636 20704
rect 86700 20640 86716 20704
rect 86780 20640 86786 20704
rect 89200 20688 90000 20718
rect 86470 20639 86786 20640
rect 6614 20160 6930 20161
rect 6614 20096 6620 20160
rect 6684 20096 6700 20160
rect 6764 20096 6780 20160
rect 6844 20096 6860 20160
rect 6924 20096 6930 20160
rect 6614 20095 6930 20096
rect 87206 20160 87522 20161
rect 87206 20096 87212 20160
rect 87276 20096 87292 20160
rect 87356 20096 87372 20160
rect 87436 20096 87452 20160
rect 87516 20096 87522 20160
rect 87206 20095 87522 20096
rect 87561 19826 87627 19829
rect 83654 19824 87627 19826
rect 83654 19768 87566 19824
rect 87622 19768 87627 19824
rect 83654 19766 87627 19768
rect 8533 19690 8599 19693
rect 8533 19688 10114 19690
rect 8533 19632 8538 19688
rect 8594 19632 10114 19688
rect 8533 19630 10114 19632
rect 8533 19627 8599 19630
rect 5878 19616 6194 19617
rect 5878 19552 5884 19616
rect 5948 19552 5964 19616
rect 6028 19552 6044 19616
rect 6108 19552 6124 19616
rect 6188 19552 6194 19616
rect 10054 19592 10114 19630
rect 46118 19630 47466 19690
rect 46118 19622 46178 19630
rect 45596 19562 46178 19622
rect 47406 19592 47466 19630
rect 83654 19622 83714 19766
rect 87561 19763 87627 19766
rect 83132 19562 83714 19622
rect 86470 19616 86786 19617
rect 5878 19551 6194 19552
rect 86470 19552 86476 19616
rect 86540 19552 86556 19616
rect 86620 19552 86636 19616
rect 86700 19552 86716 19616
rect 86780 19552 86786 19616
rect 86470 19551 86786 19552
rect 3000 19418 3800 19448
rect 4301 19418 4367 19421
rect 3000 19416 4367 19418
rect 3000 19360 4306 19416
rect 4362 19360 4367 19416
rect 3000 19358 4367 19360
rect 3000 19328 3800 19358
rect 4301 19355 4367 19358
rect 88665 19418 88731 19421
rect 89200 19418 90000 19448
rect 88665 19416 90000 19418
rect 88665 19360 88670 19416
rect 88726 19360 90000 19416
rect 88665 19358 90000 19360
rect 88665 19355 88731 19358
rect 89200 19328 90000 19358
rect 6614 19072 6930 19073
rect 6614 19008 6620 19072
rect 6684 19008 6700 19072
rect 6764 19008 6780 19072
rect 6844 19008 6860 19072
rect 6924 19008 6930 19072
rect 6614 19007 6930 19008
rect 87206 19072 87522 19073
rect 87206 19008 87212 19072
rect 87276 19008 87292 19072
rect 87356 19008 87372 19072
rect 87436 19008 87452 19072
rect 87516 19008 87522 19072
rect 87206 19007 87522 19008
rect 3000 18738 3800 18768
rect 4301 18738 4367 18741
rect 87285 18738 87351 18741
rect 3000 18736 4367 18738
rect 3000 18680 4306 18736
rect 4362 18680 4367 18736
rect 3000 18678 4367 18680
rect 3000 18648 3800 18678
rect 4301 18675 4367 18678
rect 83654 18736 87351 18738
rect 83654 18680 87290 18736
rect 87346 18680 87351 18736
rect 83654 18678 87351 18680
rect 8533 18602 8599 18605
rect 8533 18600 10114 18602
rect 8533 18544 8538 18600
rect 8594 18544 10114 18600
rect 8533 18542 10114 18544
rect 8533 18539 8599 18542
rect 5878 18528 6194 18529
rect 5878 18464 5884 18528
rect 5948 18464 5964 18528
rect 6028 18464 6044 18528
rect 6108 18464 6124 18528
rect 6188 18464 6194 18528
rect 10054 18504 10114 18542
rect 46118 18542 47466 18602
rect 46118 18534 46178 18542
rect 45596 18474 46178 18534
rect 47406 18504 47466 18542
rect 83654 18534 83714 18678
rect 87285 18675 87351 18678
rect 88205 18738 88271 18741
rect 89200 18738 90000 18768
rect 88205 18736 90000 18738
rect 88205 18680 88210 18736
rect 88266 18680 90000 18736
rect 88205 18678 90000 18680
rect 88205 18675 88271 18678
rect 89200 18648 90000 18678
rect 83132 18474 83714 18534
rect 86470 18528 86786 18529
rect 5878 18463 6194 18464
rect 86470 18464 86476 18528
rect 86540 18464 86556 18528
rect 86620 18464 86636 18528
rect 86700 18464 86716 18528
rect 86780 18464 86786 18528
rect 86470 18463 86786 18464
rect 6614 17984 6930 17985
rect 6614 17920 6620 17984
rect 6684 17920 6700 17984
rect 6764 17920 6780 17984
rect 6844 17920 6860 17984
rect 6924 17920 6930 17984
rect 6614 17919 6930 17920
rect 87206 17984 87522 17985
rect 87206 17920 87212 17984
rect 87276 17920 87292 17984
rect 87356 17920 87372 17984
rect 87436 17920 87452 17984
rect 87516 17920 87522 17984
rect 87206 17919 87522 17920
rect 8533 17514 8599 17517
rect 85813 17514 85879 17517
rect 8533 17512 10114 17514
rect 8533 17456 8538 17512
rect 8594 17456 10114 17512
rect 8533 17454 10114 17456
rect 8533 17451 8599 17454
rect 5878 17440 6194 17441
rect 3000 17378 3800 17408
rect 4301 17378 4367 17381
rect 3000 17376 4367 17378
rect 3000 17320 4306 17376
rect 4362 17320 4367 17376
rect 5878 17376 5884 17440
rect 5948 17376 5964 17440
rect 6028 17376 6044 17440
rect 6108 17376 6124 17440
rect 6188 17376 6194 17440
rect 10054 17416 10114 17454
rect 46118 17454 47466 17514
rect 46118 17446 46178 17454
rect 45596 17386 46178 17446
rect 47406 17416 47466 17454
rect 83286 17512 85879 17514
rect 83286 17456 85818 17512
rect 85874 17456 85879 17512
rect 83286 17454 85879 17456
rect 83286 17446 83346 17454
rect 85813 17451 85879 17454
rect 83132 17386 83346 17446
rect 86470 17440 86786 17441
rect 5878 17375 6194 17376
rect 86470 17376 86476 17440
rect 86540 17376 86556 17440
rect 86620 17376 86636 17440
rect 86700 17376 86716 17440
rect 86780 17376 86786 17440
rect 86470 17375 86786 17376
rect 88205 17378 88271 17381
rect 89200 17378 90000 17408
rect 88205 17376 90000 17378
rect 3000 17318 4367 17320
rect 3000 17288 3800 17318
rect 4301 17315 4367 17318
rect 88205 17320 88210 17376
rect 88266 17320 90000 17376
rect 88205 17318 90000 17320
rect 88205 17315 88271 17318
rect 89200 17288 90000 17318
rect 6614 16896 6930 16897
rect 6614 16832 6620 16896
rect 6684 16832 6700 16896
rect 6764 16832 6780 16896
rect 6844 16832 6860 16896
rect 6924 16832 6930 16896
rect 6614 16831 6930 16832
rect 87206 16896 87522 16897
rect 87206 16832 87212 16896
rect 87276 16832 87292 16896
rect 87356 16832 87372 16896
rect 87436 16832 87452 16896
rect 87516 16832 87522 16896
rect 87206 16831 87522 16832
rect 46118 16366 47466 16426
rect 46118 16358 46178 16366
rect 5878 16352 6194 16353
rect 5878 16288 5884 16352
rect 5948 16288 5964 16352
rect 6028 16288 6044 16352
rect 6108 16288 6124 16352
rect 6188 16288 6194 16352
rect 5878 16287 6194 16288
rect 8533 16290 8599 16293
rect 10054 16290 10114 16328
rect 45596 16298 46178 16358
rect 47406 16328 47466 16366
rect 83132 16298 83346 16358
rect 8533 16288 10114 16290
rect 8533 16232 8538 16288
rect 8594 16232 10114 16288
rect 8533 16230 10114 16232
rect 83286 16290 83346 16298
rect 86470 16352 86786 16353
rect 85813 16290 85879 16293
rect 83286 16288 85879 16290
rect 83286 16232 85818 16288
rect 85874 16232 85879 16288
rect 86470 16288 86476 16352
rect 86540 16288 86556 16352
rect 86620 16288 86636 16352
rect 86700 16288 86716 16352
rect 86780 16288 86786 16352
rect 86470 16287 86786 16288
rect 83286 16230 85879 16232
rect 8533 16227 8599 16230
rect 85813 16227 85879 16230
rect 3000 16018 3800 16048
rect 4301 16018 4367 16021
rect 3000 16016 4367 16018
rect 3000 15960 4306 16016
rect 4362 15960 4367 16016
rect 3000 15958 4367 15960
rect 3000 15928 3800 15958
rect 4301 15955 4367 15958
rect 88205 16018 88271 16021
rect 89200 16018 90000 16048
rect 88205 16016 90000 16018
rect 88205 15960 88210 16016
rect 88266 15960 90000 16016
rect 88205 15958 90000 15960
rect 88205 15955 88271 15958
rect 89200 15928 90000 15958
rect 6614 15808 6930 15809
rect 6614 15744 6620 15808
rect 6684 15744 6700 15808
rect 6764 15744 6780 15808
rect 6844 15744 6860 15808
rect 6924 15744 6930 15808
rect 6614 15743 6930 15744
rect 87206 15808 87522 15809
rect 87206 15744 87212 15808
rect 87276 15744 87292 15808
rect 87356 15744 87372 15808
rect 87436 15744 87452 15808
rect 87516 15744 87522 15808
rect 87206 15743 87522 15744
rect 3000 15338 3800 15368
rect 4301 15338 4367 15341
rect 84801 15338 84867 15341
rect 3000 15336 4367 15338
rect 3000 15280 4306 15336
rect 4362 15280 4367 15336
rect 3000 15278 4367 15280
rect 3000 15248 3800 15278
rect 4301 15275 4367 15278
rect 46118 15278 47466 15338
rect 46118 15270 46178 15278
rect 5878 15264 6194 15265
rect 5878 15200 5884 15264
rect 5948 15200 5964 15264
rect 6028 15200 6044 15264
rect 6108 15200 6124 15264
rect 6188 15200 6194 15264
rect 5878 15199 6194 15200
rect 5681 15066 5747 15069
rect 10054 15066 10114 15240
rect 45596 15210 46178 15270
rect 47406 15240 47466 15278
rect 83286 15336 84867 15338
rect 83286 15280 84806 15336
rect 84862 15280 84867 15336
rect 83286 15278 84867 15280
rect 83286 15270 83346 15278
rect 84801 15275 84867 15278
rect 88573 15338 88639 15341
rect 89200 15338 90000 15368
rect 88573 15336 90000 15338
rect 88573 15280 88578 15336
rect 88634 15280 90000 15336
rect 88573 15278 90000 15280
rect 88573 15275 88639 15278
rect 83132 15210 83346 15270
rect 86470 15264 86786 15265
rect 86470 15200 86476 15264
rect 86540 15200 86556 15264
rect 86620 15200 86636 15264
rect 86700 15200 86716 15264
rect 86780 15200 86786 15264
rect 89200 15248 90000 15278
rect 86470 15199 86786 15200
rect 5681 15064 10114 15066
rect 5681 15008 5686 15064
rect 5742 15008 10114 15064
rect 5681 15006 10114 15008
rect 5681 15003 5747 15006
rect 6614 14720 6930 14721
rect 6614 14656 6620 14720
rect 6684 14656 6700 14720
rect 6764 14656 6780 14720
rect 6844 14656 6860 14720
rect 6924 14656 6930 14720
rect 6614 14655 6930 14656
rect 87206 14720 87522 14721
rect 87206 14656 87212 14720
rect 87276 14656 87292 14720
rect 87356 14656 87372 14720
rect 87436 14656 87452 14720
rect 87516 14656 87522 14720
rect 87206 14655 87522 14656
rect 88021 14658 88087 14661
rect 89200 14658 90000 14688
rect 88021 14656 90000 14658
rect 88021 14600 88026 14656
rect 88082 14600 90000 14656
rect 88021 14598 90000 14600
rect 88021 14595 88087 14598
rect 89200 14568 90000 14598
rect 45977 14182 46043 14185
rect 83421 14182 83487 14185
rect 45596 14180 46043 14182
rect 5878 14176 6194 14177
rect 5878 14112 5884 14176
rect 5948 14112 5964 14176
rect 6028 14112 6044 14176
rect 6108 14112 6124 14176
rect 6188 14112 6194 14176
rect 45596 14124 45982 14180
rect 46038 14124 46043 14180
rect 45596 14122 46043 14124
rect 83132 14180 83487 14182
rect 83132 14124 83426 14180
rect 83482 14124 83487 14180
rect 83132 14122 83487 14124
rect 45977 14119 46043 14122
rect 83421 14119 83487 14122
rect 86470 14176 86786 14177
rect 5878 14111 6194 14112
rect 86470 14112 86476 14176
rect 86540 14112 86556 14176
rect 86620 14112 86636 14176
rect 86700 14112 86716 14176
rect 86780 14112 86786 14176
rect 86470 14111 86786 14112
rect 6614 13632 6930 13633
rect 6614 13568 6620 13632
rect 6684 13568 6700 13632
rect 6764 13568 6780 13632
rect 6844 13568 6860 13632
rect 6924 13568 6930 13632
rect 6614 13567 6930 13568
rect 87206 13632 87522 13633
rect 87206 13568 87212 13632
rect 87276 13568 87292 13632
rect 87356 13568 87372 13632
rect 87436 13568 87452 13632
rect 87516 13568 87522 13632
rect 87206 13567 87522 13568
rect 88205 13298 88271 13301
rect 89200 13298 90000 13328
rect 88205 13296 90000 13298
rect 88205 13240 88210 13296
rect 88266 13240 90000 13296
rect 88205 13238 90000 13240
rect 88205 13235 88271 13238
rect 89200 13208 90000 13238
rect 45885 13094 45951 13097
rect 83605 13094 83671 13097
rect 45596 13092 45951 13094
rect 5878 13088 6194 13089
rect 5878 13024 5884 13088
rect 5948 13024 5964 13088
rect 6028 13024 6044 13088
rect 6108 13024 6124 13088
rect 6188 13024 6194 13088
rect 45596 13036 45890 13092
rect 45946 13036 45951 13092
rect 45596 13034 45951 13036
rect 83132 13092 83671 13094
rect 83132 13036 83610 13092
rect 83666 13036 83671 13092
rect 83132 13034 83671 13036
rect 45885 13031 45951 13034
rect 83605 13031 83671 13034
rect 86470 13088 86786 13089
rect 5878 13023 6194 13024
rect 86470 13024 86476 13088
rect 86540 13024 86556 13088
rect 86620 13024 86636 13088
rect 86700 13024 86716 13088
rect 86780 13024 86786 13088
rect 86470 13023 86786 13024
rect 88573 12618 88639 12621
rect 89200 12618 90000 12648
rect 88573 12616 90000 12618
rect 88573 12560 88578 12616
rect 88634 12560 90000 12616
rect 88573 12558 90000 12560
rect 88573 12555 88639 12558
rect 6614 12544 6930 12545
rect 6614 12480 6620 12544
rect 6684 12480 6700 12544
rect 6764 12480 6780 12544
rect 6844 12480 6860 12544
rect 6924 12480 6930 12544
rect 6614 12479 6930 12480
rect 87206 12544 87522 12545
rect 87206 12480 87212 12544
rect 87276 12480 87292 12544
rect 87356 12480 87372 12544
rect 87436 12480 87452 12544
rect 87516 12480 87522 12544
rect 89200 12528 90000 12558
rect 87206 12479 87522 12480
rect 46069 12006 46135 12009
rect 83605 12006 83671 12009
rect 45596 12004 46135 12006
rect 5878 12000 6194 12001
rect 5878 11936 5884 12000
rect 5948 11936 5964 12000
rect 6028 11936 6044 12000
rect 6108 11936 6124 12000
rect 6188 11936 6194 12000
rect 45596 11948 46074 12004
rect 46130 11948 46135 12004
rect 45596 11946 46135 11948
rect 83132 12004 83671 12006
rect 83132 11948 83610 12004
rect 83666 11948 83671 12004
rect 83132 11946 83671 11948
rect 46069 11943 46135 11946
rect 83605 11943 83671 11946
rect 86470 12000 86786 12001
rect 5878 11935 6194 11936
rect 86470 11936 86476 12000
rect 86540 11936 86556 12000
rect 86620 11936 86636 12000
rect 86700 11936 86716 12000
rect 86780 11936 86786 12000
rect 86470 11935 86786 11936
rect 6614 11456 6930 11457
rect 6614 11392 6620 11456
rect 6684 11392 6700 11456
rect 6764 11392 6780 11456
rect 6844 11392 6860 11456
rect 6924 11392 6930 11456
rect 6614 11391 6930 11392
rect 87206 11456 87522 11457
rect 87206 11392 87212 11456
rect 87276 11392 87292 11456
rect 87356 11392 87372 11456
rect 87436 11392 87452 11456
rect 87516 11392 87522 11456
rect 87206 11391 87522 11392
rect 46437 10986 46503 10989
rect 45934 10984 46503 10986
rect 45934 10928 46442 10984
rect 46498 10928 46503 10984
rect 45934 10926 46503 10928
rect 45934 10918 45994 10926
rect 46437 10923 46503 10926
rect 83329 10918 83395 10921
rect 5878 10912 6194 10913
rect 5878 10848 5884 10912
rect 5948 10848 5964 10912
rect 6028 10848 6044 10912
rect 6108 10848 6124 10912
rect 6188 10848 6194 10912
rect 45596 10858 45994 10918
rect 83132 10916 83395 10918
rect 83132 10860 83334 10916
rect 83390 10860 83395 10916
rect 83132 10858 83395 10860
rect 83329 10855 83395 10858
rect 86470 10912 86786 10913
rect 5878 10847 6194 10848
rect 86470 10848 86476 10912
rect 86540 10848 86556 10912
rect 86620 10848 86636 10912
rect 86700 10848 86716 10912
rect 86780 10848 86786 10912
rect 86470 10847 86786 10848
rect 88205 10578 88271 10581
rect 89200 10578 90000 10608
rect 88205 10576 90000 10578
rect 88205 10520 88210 10576
rect 88266 10520 90000 10576
rect 88205 10518 90000 10520
rect 88205 10515 88271 10518
rect 89200 10488 90000 10518
rect 6614 10368 6930 10369
rect 6614 10304 6620 10368
rect 6684 10304 6700 10368
rect 6764 10304 6780 10368
rect 6844 10304 6860 10368
rect 6924 10304 6930 10368
rect 6614 10303 6930 10304
rect 87206 10368 87522 10369
rect 87206 10304 87212 10368
rect 87276 10304 87292 10368
rect 87356 10304 87372 10368
rect 87436 10304 87452 10368
rect 87516 10304 87522 10368
rect 87206 10303 87522 10304
rect 45425 10170 45491 10173
rect 46437 10170 46503 10173
rect 45425 10168 46503 10170
rect 45425 10112 45430 10168
rect 45486 10112 46442 10168
rect 46498 10112 46503 10168
rect 45425 10110 46503 10112
rect 45425 10107 45491 10110
rect 46437 10107 46503 10110
rect 5878 9824 6194 9825
rect 5878 9760 5884 9824
rect 5948 9760 5964 9824
rect 6028 9760 6044 9824
rect 6108 9760 6124 9824
rect 6188 9760 6194 9824
rect 5878 9759 6194 9760
rect 86470 9824 86786 9825
rect 86470 9760 86476 9824
rect 86540 9760 86556 9824
rect 86620 9760 86636 9824
rect 86700 9760 86716 9824
rect 86780 9760 86786 9824
rect 86470 9759 86786 9760
rect 6614 9280 6930 9281
rect 6614 9216 6620 9280
rect 6684 9216 6700 9280
rect 6764 9216 6780 9280
rect 6844 9216 6860 9280
rect 6924 9216 6930 9280
rect 6614 9215 6930 9216
rect 87206 9280 87522 9281
rect 87206 9216 87212 9280
rect 87276 9216 87292 9280
rect 87356 9216 87372 9280
rect 87436 9216 87452 9280
rect 87516 9216 87522 9280
rect 87206 9215 87522 9216
rect 5878 8736 6194 8737
rect 5878 8672 5884 8736
rect 5948 8672 5964 8736
rect 6028 8672 6044 8736
rect 6108 8672 6124 8736
rect 6188 8672 6194 8736
rect 5878 8671 6194 8672
rect 86470 8736 86786 8737
rect 86470 8672 86476 8736
rect 86540 8672 86556 8736
rect 86620 8672 86636 8736
rect 86700 8672 86716 8736
rect 86780 8672 86786 8736
rect 86470 8671 86786 8672
rect 6614 8192 6930 8193
rect 6614 8128 6620 8192
rect 6684 8128 6700 8192
rect 6764 8128 6780 8192
rect 6844 8128 6860 8192
rect 6924 8128 6930 8192
rect 6614 8127 6930 8128
rect 87206 8192 87522 8193
rect 87206 8128 87212 8192
rect 87276 8128 87292 8192
rect 87356 8128 87372 8192
rect 87436 8128 87452 8192
rect 87516 8128 87522 8192
rect 87206 8127 87522 8128
rect 5878 7648 6194 7649
rect 5878 7584 5884 7648
rect 5948 7584 5964 7648
rect 6028 7584 6044 7648
rect 6108 7584 6124 7648
rect 6188 7584 6194 7648
rect 5878 7583 6194 7584
rect 17718 7648 18034 7649
rect 17718 7584 17724 7648
rect 17788 7584 17804 7648
rect 17868 7584 17884 7648
rect 17948 7584 17964 7648
rect 18028 7584 18034 7648
rect 17718 7583 18034 7584
rect 36118 7648 36434 7649
rect 36118 7584 36124 7648
rect 36188 7584 36204 7648
rect 36268 7584 36284 7648
rect 36348 7584 36364 7648
rect 36428 7584 36434 7648
rect 36118 7583 36434 7584
rect 54518 7648 54834 7649
rect 54518 7584 54524 7648
rect 54588 7584 54604 7648
rect 54668 7584 54684 7648
rect 54748 7584 54764 7648
rect 54828 7584 54834 7648
rect 54518 7583 54834 7584
rect 72918 7648 73234 7649
rect 72918 7584 72924 7648
rect 72988 7584 73004 7648
rect 73068 7584 73084 7648
rect 73148 7584 73164 7648
rect 73228 7584 73234 7648
rect 72918 7583 73234 7584
rect 86470 7648 86786 7649
rect 86470 7584 86476 7648
rect 86540 7584 86556 7648
rect 86620 7584 86636 7648
rect 86700 7584 86716 7648
rect 86780 7584 86786 7648
rect 86470 7583 86786 7584
rect 6614 7104 6930 7105
rect 6614 7040 6620 7104
rect 6684 7040 6700 7104
rect 6764 7040 6780 7104
rect 6844 7040 6860 7104
rect 6924 7040 6930 7104
rect 6614 7039 6930 7040
rect 18378 7104 18694 7105
rect 18378 7040 18384 7104
rect 18448 7040 18464 7104
rect 18528 7040 18544 7104
rect 18608 7040 18624 7104
rect 18688 7040 18694 7104
rect 18378 7039 18694 7040
rect 36778 7104 37094 7105
rect 36778 7040 36784 7104
rect 36848 7040 36864 7104
rect 36928 7040 36944 7104
rect 37008 7040 37024 7104
rect 37088 7040 37094 7104
rect 36778 7039 37094 7040
rect 55178 7104 55494 7105
rect 55178 7040 55184 7104
rect 55248 7040 55264 7104
rect 55328 7040 55344 7104
rect 55408 7040 55424 7104
rect 55488 7040 55494 7104
rect 55178 7039 55494 7040
rect 73578 7104 73894 7105
rect 73578 7040 73584 7104
rect 73648 7040 73664 7104
rect 73728 7040 73744 7104
rect 73808 7040 73824 7104
rect 73888 7040 73894 7104
rect 73578 7039 73894 7040
rect 87206 7104 87522 7105
rect 87206 7040 87212 7104
rect 87276 7040 87292 7104
rect 87356 7040 87372 7104
rect 87436 7040 87452 7104
rect 87516 7040 87522 7104
rect 87206 7039 87522 7040
rect 17718 6560 18034 6561
rect 17718 6496 17724 6560
rect 17788 6496 17804 6560
rect 17868 6496 17884 6560
rect 17948 6496 17964 6560
rect 18028 6496 18034 6560
rect 17718 6495 18034 6496
rect 36118 6560 36434 6561
rect 36118 6496 36124 6560
rect 36188 6496 36204 6560
rect 36268 6496 36284 6560
rect 36348 6496 36364 6560
rect 36428 6496 36434 6560
rect 36118 6495 36434 6496
rect 54518 6560 54834 6561
rect 54518 6496 54524 6560
rect 54588 6496 54604 6560
rect 54668 6496 54684 6560
rect 54748 6496 54764 6560
rect 54828 6496 54834 6560
rect 54518 6495 54834 6496
rect 72918 6560 73234 6561
rect 72918 6496 72924 6560
rect 72988 6496 73004 6560
rect 73068 6496 73084 6560
rect 73148 6496 73164 6560
rect 73228 6496 73234 6560
rect 72918 6495 73234 6496
rect 18378 6016 18694 6017
rect 18378 5952 18384 6016
rect 18448 5952 18464 6016
rect 18528 5952 18544 6016
rect 18608 5952 18624 6016
rect 18688 5952 18694 6016
rect 18378 5951 18694 5952
rect 36778 6016 37094 6017
rect 36778 5952 36784 6016
rect 36848 5952 36864 6016
rect 36928 5952 36944 6016
rect 37008 5952 37024 6016
rect 37088 5952 37094 6016
rect 36778 5951 37094 5952
rect 55178 6016 55494 6017
rect 55178 5952 55184 6016
rect 55248 5952 55264 6016
rect 55328 5952 55344 6016
rect 55408 5952 55424 6016
rect 55488 5952 55494 6016
rect 55178 5951 55494 5952
rect 73578 6016 73894 6017
rect 73578 5952 73584 6016
rect 73648 5952 73664 6016
rect 73728 5952 73744 6016
rect 73808 5952 73824 6016
rect 73888 5952 73894 6016
rect 73578 5951 73894 5952
rect 17718 5472 18034 5473
rect 17718 5408 17724 5472
rect 17788 5408 17804 5472
rect 17868 5408 17884 5472
rect 17948 5408 17964 5472
rect 18028 5408 18034 5472
rect 17718 5407 18034 5408
rect 36118 5472 36434 5473
rect 36118 5408 36124 5472
rect 36188 5408 36204 5472
rect 36268 5408 36284 5472
rect 36348 5408 36364 5472
rect 36428 5408 36434 5472
rect 36118 5407 36434 5408
rect 54518 5472 54834 5473
rect 54518 5408 54524 5472
rect 54588 5408 54604 5472
rect 54668 5408 54684 5472
rect 54748 5408 54764 5472
rect 54828 5408 54834 5472
rect 54518 5407 54834 5408
rect 72918 5472 73234 5473
rect 72918 5408 72924 5472
rect 72988 5408 73004 5472
rect 73068 5408 73084 5472
rect 73148 5408 73164 5472
rect 73228 5408 73234 5472
rect 72918 5407 73234 5408
rect 18378 4928 18694 4929
rect 18378 4864 18384 4928
rect 18448 4864 18464 4928
rect 18528 4864 18544 4928
rect 18608 4864 18624 4928
rect 18688 4864 18694 4928
rect 18378 4863 18694 4864
rect 36778 4928 37094 4929
rect 36778 4864 36784 4928
rect 36848 4864 36864 4928
rect 36928 4864 36944 4928
rect 37008 4864 37024 4928
rect 37088 4864 37094 4928
rect 36778 4863 37094 4864
rect 55178 4928 55494 4929
rect 55178 4864 55184 4928
rect 55248 4864 55264 4928
rect 55328 4864 55344 4928
rect 55408 4864 55424 4928
rect 55488 4864 55494 4928
rect 55178 4863 55494 4864
rect 73578 4928 73894 4929
rect 73578 4864 73584 4928
rect 73648 4864 73664 4928
rect 73728 4864 73744 4928
rect 73808 4864 73824 4928
rect 73888 4864 73894 4928
rect 73578 4863 73894 4864
<< via3 >>
rect 18384 87612 18448 87616
rect 18384 87556 18388 87612
rect 18388 87556 18444 87612
rect 18444 87556 18448 87612
rect 18384 87552 18448 87556
rect 18464 87612 18528 87616
rect 18464 87556 18468 87612
rect 18468 87556 18524 87612
rect 18524 87556 18528 87612
rect 18464 87552 18528 87556
rect 18544 87612 18608 87616
rect 18544 87556 18548 87612
rect 18548 87556 18604 87612
rect 18604 87556 18608 87612
rect 18544 87552 18608 87556
rect 18624 87612 18688 87616
rect 18624 87556 18628 87612
rect 18628 87556 18684 87612
rect 18684 87556 18688 87612
rect 18624 87552 18688 87556
rect 36784 87612 36848 87616
rect 36784 87556 36788 87612
rect 36788 87556 36844 87612
rect 36844 87556 36848 87612
rect 36784 87552 36848 87556
rect 36864 87612 36928 87616
rect 36864 87556 36868 87612
rect 36868 87556 36924 87612
rect 36924 87556 36928 87612
rect 36864 87552 36928 87556
rect 36944 87612 37008 87616
rect 36944 87556 36948 87612
rect 36948 87556 37004 87612
rect 37004 87556 37008 87612
rect 36944 87552 37008 87556
rect 37024 87612 37088 87616
rect 37024 87556 37028 87612
rect 37028 87556 37084 87612
rect 37084 87556 37088 87612
rect 37024 87552 37088 87556
rect 55184 87612 55248 87616
rect 55184 87556 55188 87612
rect 55188 87556 55244 87612
rect 55244 87556 55248 87612
rect 55184 87552 55248 87556
rect 55264 87612 55328 87616
rect 55264 87556 55268 87612
rect 55268 87556 55324 87612
rect 55324 87556 55328 87612
rect 55264 87552 55328 87556
rect 55344 87612 55408 87616
rect 55344 87556 55348 87612
rect 55348 87556 55404 87612
rect 55404 87556 55408 87612
rect 55344 87552 55408 87556
rect 55424 87612 55488 87616
rect 55424 87556 55428 87612
rect 55428 87556 55484 87612
rect 55484 87556 55488 87612
rect 55424 87552 55488 87556
rect 73584 87612 73648 87616
rect 73584 87556 73588 87612
rect 73588 87556 73644 87612
rect 73644 87556 73648 87612
rect 73584 87552 73648 87556
rect 73664 87612 73728 87616
rect 73664 87556 73668 87612
rect 73668 87556 73724 87612
rect 73724 87556 73728 87612
rect 73664 87552 73728 87556
rect 73744 87612 73808 87616
rect 73744 87556 73748 87612
rect 73748 87556 73804 87612
rect 73804 87556 73808 87612
rect 73744 87552 73808 87556
rect 73824 87612 73888 87616
rect 73824 87556 73828 87612
rect 73828 87556 73884 87612
rect 73884 87556 73888 87612
rect 73824 87552 73888 87556
rect 17724 87068 17788 87072
rect 17724 87012 17728 87068
rect 17728 87012 17784 87068
rect 17784 87012 17788 87068
rect 17724 87008 17788 87012
rect 17804 87068 17868 87072
rect 17804 87012 17808 87068
rect 17808 87012 17864 87068
rect 17864 87012 17868 87068
rect 17804 87008 17868 87012
rect 17884 87068 17948 87072
rect 17884 87012 17888 87068
rect 17888 87012 17944 87068
rect 17944 87012 17948 87068
rect 17884 87008 17948 87012
rect 17964 87068 18028 87072
rect 17964 87012 17968 87068
rect 17968 87012 18024 87068
rect 18024 87012 18028 87068
rect 17964 87008 18028 87012
rect 36124 87068 36188 87072
rect 36124 87012 36128 87068
rect 36128 87012 36184 87068
rect 36184 87012 36188 87068
rect 36124 87008 36188 87012
rect 36204 87068 36268 87072
rect 36204 87012 36208 87068
rect 36208 87012 36264 87068
rect 36264 87012 36268 87068
rect 36204 87008 36268 87012
rect 36284 87068 36348 87072
rect 36284 87012 36288 87068
rect 36288 87012 36344 87068
rect 36344 87012 36348 87068
rect 36284 87008 36348 87012
rect 36364 87068 36428 87072
rect 36364 87012 36368 87068
rect 36368 87012 36424 87068
rect 36424 87012 36428 87068
rect 36364 87008 36428 87012
rect 54524 87068 54588 87072
rect 54524 87012 54528 87068
rect 54528 87012 54584 87068
rect 54584 87012 54588 87068
rect 54524 87008 54588 87012
rect 54604 87068 54668 87072
rect 54604 87012 54608 87068
rect 54608 87012 54664 87068
rect 54664 87012 54668 87068
rect 54604 87008 54668 87012
rect 54684 87068 54748 87072
rect 54684 87012 54688 87068
rect 54688 87012 54744 87068
rect 54744 87012 54748 87068
rect 54684 87008 54748 87012
rect 54764 87068 54828 87072
rect 54764 87012 54768 87068
rect 54768 87012 54824 87068
rect 54824 87012 54828 87068
rect 54764 87008 54828 87012
rect 72924 87068 72988 87072
rect 72924 87012 72928 87068
rect 72928 87012 72984 87068
rect 72984 87012 72988 87068
rect 72924 87008 72988 87012
rect 73004 87068 73068 87072
rect 73004 87012 73008 87068
rect 73008 87012 73064 87068
rect 73064 87012 73068 87068
rect 73004 87008 73068 87012
rect 73084 87068 73148 87072
rect 73084 87012 73088 87068
rect 73088 87012 73144 87068
rect 73144 87012 73148 87068
rect 73084 87008 73148 87012
rect 73164 87068 73228 87072
rect 73164 87012 73168 87068
rect 73168 87012 73224 87068
rect 73224 87012 73228 87068
rect 73164 87008 73228 87012
rect 18384 86524 18448 86528
rect 18384 86468 18388 86524
rect 18388 86468 18444 86524
rect 18444 86468 18448 86524
rect 18384 86464 18448 86468
rect 18464 86524 18528 86528
rect 18464 86468 18468 86524
rect 18468 86468 18524 86524
rect 18524 86468 18528 86524
rect 18464 86464 18528 86468
rect 18544 86524 18608 86528
rect 18544 86468 18548 86524
rect 18548 86468 18604 86524
rect 18604 86468 18608 86524
rect 18544 86464 18608 86468
rect 18624 86524 18688 86528
rect 18624 86468 18628 86524
rect 18628 86468 18684 86524
rect 18684 86468 18688 86524
rect 18624 86464 18688 86468
rect 36784 86524 36848 86528
rect 36784 86468 36788 86524
rect 36788 86468 36844 86524
rect 36844 86468 36848 86524
rect 36784 86464 36848 86468
rect 36864 86524 36928 86528
rect 36864 86468 36868 86524
rect 36868 86468 36924 86524
rect 36924 86468 36928 86524
rect 36864 86464 36928 86468
rect 36944 86524 37008 86528
rect 36944 86468 36948 86524
rect 36948 86468 37004 86524
rect 37004 86468 37008 86524
rect 36944 86464 37008 86468
rect 37024 86524 37088 86528
rect 37024 86468 37028 86524
rect 37028 86468 37084 86524
rect 37084 86468 37088 86524
rect 37024 86464 37088 86468
rect 55184 86524 55248 86528
rect 55184 86468 55188 86524
rect 55188 86468 55244 86524
rect 55244 86468 55248 86524
rect 55184 86464 55248 86468
rect 55264 86524 55328 86528
rect 55264 86468 55268 86524
rect 55268 86468 55324 86524
rect 55324 86468 55328 86524
rect 55264 86464 55328 86468
rect 55344 86524 55408 86528
rect 55344 86468 55348 86524
rect 55348 86468 55404 86524
rect 55404 86468 55408 86524
rect 55344 86464 55408 86468
rect 55424 86524 55488 86528
rect 55424 86468 55428 86524
rect 55428 86468 55484 86524
rect 55484 86468 55488 86524
rect 55424 86464 55488 86468
rect 73584 86524 73648 86528
rect 73584 86468 73588 86524
rect 73588 86468 73644 86524
rect 73644 86468 73648 86524
rect 73584 86464 73648 86468
rect 73664 86524 73728 86528
rect 73664 86468 73668 86524
rect 73668 86468 73724 86524
rect 73724 86468 73728 86524
rect 73664 86464 73728 86468
rect 73744 86524 73808 86528
rect 73744 86468 73748 86524
rect 73748 86468 73804 86524
rect 73804 86468 73808 86524
rect 73744 86464 73808 86468
rect 73824 86524 73888 86528
rect 73824 86468 73828 86524
rect 73828 86468 73884 86524
rect 73884 86468 73888 86524
rect 73824 86464 73888 86468
rect 17724 85980 17788 85984
rect 17724 85924 17728 85980
rect 17728 85924 17784 85980
rect 17784 85924 17788 85980
rect 17724 85920 17788 85924
rect 17804 85980 17868 85984
rect 17804 85924 17808 85980
rect 17808 85924 17864 85980
rect 17864 85924 17868 85980
rect 17804 85920 17868 85924
rect 17884 85980 17948 85984
rect 17884 85924 17888 85980
rect 17888 85924 17944 85980
rect 17944 85924 17948 85980
rect 17884 85920 17948 85924
rect 17964 85980 18028 85984
rect 17964 85924 17968 85980
rect 17968 85924 18024 85980
rect 18024 85924 18028 85980
rect 17964 85920 18028 85924
rect 36124 85980 36188 85984
rect 36124 85924 36128 85980
rect 36128 85924 36184 85980
rect 36184 85924 36188 85980
rect 36124 85920 36188 85924
rect 36204 85980 36268 85984
rect 36204 85924 36208 85980
rect 36208 85924 36264 85980
rect 36264 85924 36268 85980
rect 36204 85920 36268 85924
rect 36284 85980 36348 85984
rect 36284 85924 36288 85980
rect 36288 85924 36344 85980
rect 36344 85924 36348 85980
rect 36284 85920 36348 85924
rect 36364 85980 36428 85984
rect 36364 85924 36368 85980
rect 36368 85924 36424 85980
rect 36424 85924 36428 85980
rect 36364 85920 36428 85924
rect 54524 85980 54588 85984
rect 54524 85924 54528 85980
rect 54528 85924 54584 85980
rect 54584 85924 54588 85980
rect 54524 85920 54588 85924
rect 54604 85980 54668 85984
rect 54604 85924 54608 85980
rect 54608 85924 54664 85980
rect 54664 85924 54668 85980
rect 54604 85920 54668 85924
rect 54684 85980 54748 85984
rect 54684 85924 54688 85980
rect 54688 85924 54744 85980
rect 54744 85924 54748 85980
rect 54684 85920 54748 85924
rect 54764 85980 54828 85984
rect 54764 85924 54768 85980
rect 54768 85924 54824 85980
rect 54824 85924 54828 85980
rect 54764 85920 54828 85924
rect 72924 85980 72988 85984
rect 72924 85924 72928 85980
rect 72928 85924 72984 85980
rect 72984 85924 72988 85980
rect 72924 85920 72988 85924
rect 73004 85980 73068 85984
rect 73004 85924 73008 85980
rect 73008 85924 73064 85980
rect 73064 85924 73068 85980
rect 73004 85920 73068 85924
rect 73084 85980 73148 85984
rect 73084 85924 73088 85980
rect 73088 85924 73144 85980
rect 73144 85924 73148 85980
rect 73084 85920 73148 85924
rect 73164 85980 73228 85984
rect 73164 85924 73168 85980
rect 73168 85924 73224 85980
rect 73224 85924 73228 85980
rect 73164 85920 73228 85924
rect 18384 85436 18448 85440
rect 18384 85380 18388 85436
rect 18388 85380 18444 85436
rect 18444 85380 18448 85436
rect 18384 85376 18448 85380
rect 18464 85436 18528 85440
rect 18464 85380 18468 85436
rect 18468 85380 18524 85436
rect 18524 85380 18528 85436
rect 18464 85376 18528 85380
rect 18544 85436 18608 85440
rect 18544 85380 18548 85436
rect 18548 85380 18604 85436
rect 18604 85380 18608 85436
rect 18544 85376 18608 85380
rect 18624 85436 18688 85440
rect 18624 85380 18628 85436
rect 18628 85380 18684 85436
rect 18684 85380 18688 85436
rect 18624 85376 18688 85380
rect 36784 85436 36848 85440
rect 36784 85380 36788 85436
rect 36788 85380 36844 85436
rect 36844 85380 36848 85436
rect 36784 85376 36848 85380
rect 36864 85436 36928 85440
rect 36864 85380 36868 85436
rect 36868 85380 36924 85436
rect 36924 85380 36928 85436
rect 36864 85376 36928 85380
rect 36944 85436 37008 85440
rect 36944 85380 36948 85436
rect 36948 85380 37004 85436
rect 37004 85380 37008 85436
rect 36944 85376 37008 85380
rect 37024 85436 37088 85440
rect 37024 85380 37028 85436
rect 37028 85380 37084 85436
rect 37084 85380 37088 85436
rect 37024 85376 37088 85380
rect 55184 85436 55248 85440
rect 55184 85380 55188 85436
rect 55188 85380 55244 85436
rect 55244 85380 55248 85436
rect 55184 85376 55248 85380
rect 55264 85436 55328 85440
rect 55264 85380 55268 85436
rect 55268 85380 55324 85436
rect 55324 85380 55328 85436
rect 55264 85376 55328 85380
rect 55344 85436 55408 85440
rect 55344 85380 55348 85436
rect 55348 85380 55404 85436
rect 55404 85380 55408 85436
rect 55344 85376 55408 85380
rect 55424 85436 55488 85440
rect 55424 85380 55428 85436
rect 55428 85380 55484 85436
rect 55484 85380 55488 85436
rect 55424 85376 55488 85380
rect 73584 85436 73648 85440
rect 73584 85380 73588 85436
rect 73588 85380 73644 85436
rect 73644 85380 73648 85436
rect 73584 85376 73648 85380
rect 73664 85436 73728 85440
rect 73664 85380 73668 85436
rect 73668 85380 73724 85436
rect 73724 85380 73728 85436
rect 73664 85376 73728 85380
rect 73744 85436 73808 85440
rect 73744 85380 73748 85436
rect 73748 85380 73804 85436
rect 73804 85380 73808 85436
rect 73744 85376 73808 85380
rect 73824 85436 73888 85440
rect 73824 85380 73828 85436
rect 73828 85380 73884 85436
rect 73884 85380 73888 85436
rect 73824 85376 73888 85380
rect 5884 84892 5948 84896
rect 5884 84836 5888 84892
rect 5888 84836 5944 84892
rect 5944 84836 5948 84892
rect 5884 84832 5948 84836
rect 5964 84892 6028 84896
rect 5964 84836 5968 84892
rect 5968 84836 6024 84892
rect 6024 84836 6028 84892
rect 5964 84832 6028 84836
rect 6044 84892 6108 84896
rect 6044 84836 6048 84892
rect 6048 84836 6104 84892
rect 6104 84836 6108 84892
rect 6044 84832 6108 84836
rect 6124 84892 6188 84896
rect 6124 84836 6128 84892
rect 6128 84836 6184 84892
rect 6184 84836 6188 84892
rect 6124 84832 6188 84836
rect 17724 84892 17788 84896
rect 17724 84836 17728 84892
rect 17728 84836 17784 84892
rect 17784 84836 17788 84892
rect 17724 84832 17788 84836
rect 17804 84892 17868 84896
rect 17804 84836 17808 84892
rect 17808 84836 17864 84892
rect 17864 84836 17868 84892
rect 17804 84832 17868 84836
rect 17884 84892 17948 84896
rect 17884 84836 17888 84892
rect 17888 84836 17944 84892
rect 17944 84836 17948 84892
rect 17884 84832 17948 84836
rect 17964 84892 18028 84896
rect 17964 84836 17968 84892
rect 17968 84836 18024 84892
rect 18024 84836 18028 84892
rect 17964 84832 18028 84836
rect 36124 84892 36188 84896
rect 36124 84836 36128 84892
rect 36128 84836 36184 84892
rect 36184 84836 36188 84892
rect 36124 84832 36188 84836
rect 36204 84892 36268 84896
rect 36204 84836 36208 84892
rect 36208 84836 36264 84892
rect 36264 84836 36268 84892
rect 36204 84832 36268 84836
rect 36284 84892 36348 84896
rect 36284 84836 36288 84892
rect 36288 84836 36344 84892
rect 36344 84836 36348 84892
rect 36284 84832 36348 84836
rect 36364 84892 36428 84896
rect 36364 84836 36368 84892
rect 36368 84836 36424 84892
rect 36424 84836 36428 84892
rect 36364 84832 36428 84836
rect 54524 84892 54588 84896
rect 54524 84836 54528 84892
rect 54528 84836 54584 84892
rect 54584 84836 54588 84892
rect 54524 84832 54588 84836
rect 54604 84892 54668 84896
rect 54604 84836 54608 84892
rect 54608 84836 54664 84892
rect 54664 84836 54668 84892
rect 54604 84832 54668 84836
rect 54684 84892 54748 84896
rect 54684 84836 54688 84892
rect 54688 84836 54744 84892
rect 54744 84836 54748 84892
rect 54684 84832 54748 84836
rect 54764 84892 54828 84896
rect 54764 84836 54768 84892
rect 54768 84836 54824 84892
rect 54824 84836 54828 84892
rect 54764 84832 54828 84836
rect 72924 84892 72988 84896
rect 72924 84836 72928 84892
rect 72928 84836 72984 84892
rect 72984 84836 72988 84892
rect 72924 84832 72988 84836
rect 73004 84892 73068 84896
rect 73004 84836 73008 84892
rect 73008 84836 73064 84892
rect 73064 84836 73068 84892
rect 73004 84832 73068 84836
rect 73084 84892 73148 84896
rect 73084 84836 73088 84892
rect 73088 84836 73144 84892
rect 73144 84836 73148 84892
rect 73084 84832 73148 84836
rect 73164 84892 73228 84896
rect 73164 84836 73168 84892
rect 73168 84836 73224 84892
rect 73224 84836 73228 84892
rect 73164 84832 73228 84836
rect 86476 84892 86540 84896
rect 86476 84836 86480 84892
rect 86480 84836 86536 84892
rect 86536 84836 86540 84892
rect 86476 84832 86540 84836
rect 86556 84892 86620 84896
rect 86556 84836 86560 84892
rect 86560 84836 86616 84892
rect 86616 84836 86620 84892
rect 86556 84832 86620 84836
rect 86636 84892 86700 84896
rect 86636 84836 86640 84892
rect 86640 84836 86696 84892
rect 86696 84836 86700 84892
rect 86636 84832 86700 84836
rect 86716 84892 86780 84896
rect 86716 84836 86720 84892
rect 86720 84836 86776 84892
rect 86776 84836 86780 84892
rect 86716 84832 86780 84836
rect 6620 84348 6684 84352
rect 6620 84292 6624 84348
rect 6624 84292 6680 84348
rect 6680 84292 6684 84348
rect 6620 84288 6684 84292
rect 6700 84348 6764 84352
rect 6700 84292 6704 84348
rect 6704 84292 6760 84348
rect 6760 84292 6764 84348
rect 6700 84288 6764 84292
rect 6780 84348 6844 84352
rect 6780 84292 6784 84348
rect 6784 84292 6840 84348
rect 6840 84292 6844 84348
rect 6780 84288 6844 84292
rect 6860 84348 6924 84352
rect 6860 84292 6864 84348
rect 6864 84292 6920 84348
rect 6920 84292 6924 84348
rect 6860 84288 6924 84292
rect 18384 84348 18448 84352
rect 18384 84292 18388 84348
rect 18388 84292 18444 84348
rect 18444 84292 18448 84348
rect 18384 84288 18448 84292
rect 18464 84348 18528 84352
rect 18464 84292 18468 84348
rect 18468 84292 18524 84348
rect 18524 84292 18528 84348
rect 18464 84288 18528 84292
rect 18544 84348 18608 84352
rect 18544 84292 18548 84348
rect 18548 84292 18604 84348
rect 18604 84292 18608 84348
rect 18544 84288 18608 84292
rect 18624 84348 18688 84352
rect 18624 84292 18628 84348
rect 18628 84292 18684 84348
rect 18684 84292 18688 84348
rect 18624 84288 18688 84292
rect 36784 84348 36848 84352
rect 36784 84292 36788 84348
rect 36788 84292 36844 84348
rect 36844 84292 36848 84348
rect 36784 84288 36848 84292
rect 36864 84348 36928 84352
rect 36864 84292 36868 84348
rect 36868 84292 36924 84348
rect 36924 84292 36928 84348
rect 36864 84288 36928 84292
rect 36944 84348 37008 84352
rect 36944 84292 36948 84348
rect 36948 84292 37004 84348
rect 37004 84292 37008 84348
rect 36944 84288 37008 84292
rect 37024 84348 37088 84352
rect 37024 84292 37028 84348
rect 37028 84292 37084 84348
rect 37084 84292 37088 84348
rect 37024 84288 37088 84292
rect 55184 84348 55248 84352
rect 55184 84292 55188 84348
rect 55188 84292 55244 84348
rect 55244 84292 55248 84348
rect 55184 84288 55248 84292
rect 55264 84348 55328 84352
rect 55264 84292 55268 84348
rect 55268 84292 55324 84348
rect 55324 84292 55328 84348
rect 55264 84288 55328 84292
rect 55344 84348 55408 84352
rect 55344 84292 55348 84348
rect 55348 84292 55404 84348
rect 55404 84292 55408 84348
rect 55344 84288 55408 84292
rect 55424 84348 55488 84352
rect 55424 84292 55428 84348
rect 55428 84292 55484 84348
rect 55484 84292 55488 84348
rect 55424 84288 55488 84292
rect 73584 84348 73648 84352
rect 73584 84292 73588 84348
rect 73588 84292 73644 84348
rect 73644 84292 73648 84348
rect 73584 84288 73648 84292
rect 73664 84348 73728 84352
rect 73664 84292 73668 84348
rect 73668 84292 73724 84348
rect 73724 84292 73728 84348
rect 73664 84288 73728 84292
rect 73744 84348 73808 84352
rect 73744 84292 73748 84348
rect 73748 84292 73804 84348
rect 73804 84292 73808 84348
rect 73744 84288 73808 84292
rect 73824 84348 73888 84352
rect 73824 84292 73828 84348
rect 73828 84292 73884 84348
rect 73884 84292 73888 84348
rect 73824 84288 73888 84292
rect 87212 84348 87276 84352
rect 87212 84292 87216 84348
rect 87216 84292 87272 84348
rect 87272 84292 87276 84348
rect 87212 84288 87276 84292
rect 87292 84348 87356 84352
rect 87292 84292 87296 84348
rect 87296 84292 87352 84348
rect 87352 84292 87356 84348
rect 87292 84288 87356 84292
rect 87372 84348 87436 84352
rect 87372 84292 87376 84348
rect 87376 84292 87432 84348
rect 87432 84292 87436 84348
rect 87372 84288 87436 84292
rect 87452 84348 87516 84352
rect 87452 84292 87456 84348
rect 87456 84292 87512 84348
rect 87512 84292 87516 84348
rect 87452 84288 87516 84292
rect 5884 83804 5948 83808
rect 5884 83748 5888 83804
rect 5888 83748 5944 83804
rect 5944 83748 5948 83804
rect 5884 83744 5948 83748
rect 5964 83804 6028 83808
rect 5964 83748 5968 83804
rect 5968 83748 6024 83804
rect 6024 83748 6028 83804
rect 5964 83744 6028 83748
rect 6044 83804 6108 83808
rect 6044 83748 6048 83804
rect 6048 83748 6104 83804
rect 6104 83748 6108 83804
rect 6044 83744 6108 83748
rect 6124 83804 6188 83808
rect 6124 83748 6128 83804
rect 6128 83748 6184 83804
rect 6184 83748 6188 83804
rect 6124 83744 6188 83748
rect 86476 83804 86540 83808
rect 86476 83748 86480 83804
rect 86480 83748 86536 83804
rect 86536 83748 86540 83804
rect 86476 83744 86540 83748
rect 86556 83804 86620 83808
rect 86556 83748 86560 83804
rect 86560 83748 86616 83804
rect 86616 83748 86620 83804
rect 86556 83744 86620 83748
rect 86636 83804 86700 83808
rect 86636 83748 86640 83804
rect 86640 83748 86696 83804
rect 86696 83748 86700 83804
rect 86636 83744 86700 83748
rect 86716 83804 86780 83808
rect 86716 83748 86720 83804
rect 86720 83748 86776 83804
rect 86776 83748 86780 83804
rect 86716 83744 86780 83748
rect 6620 83260 6684 83264
rect 6620 83204 6624 83260
rect 6624 83204 6680 83260
rect 6680 83204 6684 83260
rect 6620 83200 6684 83204
rect 6700 83260 6764 83264
rect 6700 83204 6704 83260
rect 6704 83204 6760 83260
rect 6760 83204 6764 83260
rect 6700 83200 6764 83204
rect 6780 83260 6844 83264
rect 6780 83204 6784 83260
rect 6784 83204 6840 83260
rect 6840 83204 6844 83260
rect 6780 83200 6844 83204
rect 6860 83260 6924 83264
rect 6860 83204 6864 83260
rect 6864 83204 6920 83260
rect 6920 83204 6924 83260
rect 6860 83200 6924 83204
rect 87212 83260 87276 83264
rect 87212 83204 87216 83260
rect 87216 83204 87272 83260
rect 87272 83204 87276 83260
rect 87212 83200 87276 83204
rect 87292 83260 87356 83264
rect 87292 83204 87296 83260
rect 87296 83204 87352 83260
rect 87352 83204 87356 83260
rect 87292 83200 87356 83204
rect 87372 83260 87436 83264
rect 87372 83204 87376 83260
rect 87376 83204 87432 83260
rect 87432 83204 87436 83260
rect 87372 83200 87436 83204
rect 87452 83260 87516 83264
rect 87452 83204 87456 83260
rect 87456 83204 87512 83260
rect 87512 83204 87516 83260
rect 87452 83200 87516 83204
rect 5884 82716 5948 82720
rect 5884 82660 5888 82716
rect 5888 82660 5944 82716
rect 5944 82660 5948 82716
rect 5884 82656 5948 82660
rect 5964 82716 6028 82720
rect 5964 82660 5968 82716
rect 5968 82660 6024 82716
rect 6024 82660 6028 82716
rect 5964 82656 6028 82660
rect 6044 82716 6108 82720
rect 6044 82660 6048 82716
rect 6048 82660 6104 82716
rect 6104 82660 6108 82716
rect 6044 82656 6108 82660
rect 6124 82716 6188 82720
rect 6124 82660 6128 82716
rect 6128 82660 6184 82716
rect 6184 82660 6188 82716
rect 6124 82656 6188 82660
rect 86476 82716 86540 82720
rect 86476 82660 86480 82716
rect 86480 82660 86536 82716
rect 86536 82660 86540 82716
rect 86476 82656 86540 82660
rect 86556 82716 86620 82720
rect 86556 82660 86560 82716
rect 86560 82660 86616 82716
rect 86616 82660 86620 82716
rect 86556 82656 86620 82660
rect 86636 82716 86700 82720
rect 86636 82660 86640 82716
rect 86640 82660 86696 82716
rect 86696 82660 86700 82716
rect 86636 82656 86700 82660
rect 86716 82716 86780 82720
rect 86716 82660 86720 82716
rect 86720 82660 86776 82716
rect 86776 82660 86780 82716
rect 86716 82656 86780 82660
rect 6620 82172 6684 82176
rect 6620 82116 6624 82172
rect 6624 82116 6680 82172
rect 6680 82116 6684 82172
rect 6620 82112 6684 82116
rect 6700 82172 6764 82176
rect 6700 82116 6704 82172
rect 6704 82116 6760 82172
rect 6760 82116 6764 82172
rect 6700 82112 6764 82116
rect 6780 82172 6844 82176
rect 6780 82116 6784 82172
rect 6784 82116 6840 82172
rect 6840 82116 6844 82172
rect 6780 82112 6844 82116
rect 6860 82172 6924 82176
rect 6860 82116 6864 82172
rect 6864 82116 6920 82172
rect 6920 82116 6924 82172
rect 6860 82112 6924 82116
rect 87212 82172 87276 82176
rect 87212 82116 87216 82172
rect 87216 82116 87272 82172
rect 87272 82116 87276 82172
rect 87212 82112 87276 82116
rect 87292 82172 87356 82176
rect 87292 82116 87296 82172
rect 87296 82116 87352 82172
rect 87352 82116 87356 82172
rect 87292 82112 87356 82116
rect 87372 82172 87436 82176
rect 87372 82116 87376 82172
rect 87376 82116 87432 82172
rect 87432 82116 87436 82172
rect 87372 82112 87436 82116
rect 87452 82172 87516 82176
rect 87452 82116 87456 82172
rect 87456 82116 87512 82172
rect 87512 82116 87516 82172
rect 87452 82112 87516 82116
rect 5884 81628 5948 81632
rect 5884 81572 5888 81628
rect 5888 81572 5944 81628
rect 5944 81572 5948 81628
rect 5884 81568 5948 81572
rect 5964 81628 6028 81632
rect 5964 81572 5968 81628
rect 5968 81572 6024 81628
rect 6024 81572 6028 81628
rect 5964 81568 6028 81572
rect 6044 81628 6108 81632
rect 6044 81572 6048 81628
rect 6048 81572 6104 81628
rect 6104 81572 6108 81628
rect 6044 81568 6108 81572
rect 6124 81628 6188 81632
rect 6124 81572 6128 81628
rect 6128 81572 6184 81628
rect 6184 81572 6188 81628
rect 6124 81568 6188 81572
rect 86476 81628 86540 81632
rect 86476 81572 86480 81628
rect 86480 81572 86536 81628
rect 86536 81572 86540 81628
rect 86476 81568 86540 81572
rect 86556 81628 86620 81632
rect 86556 81572 86560 81628
rect 86560 81572 86616 81628
rect 86616 81572 86620 81628
rect 86556 81568 86620 81572
rect 86636 81628 86700 81632
rect 86636 81572 86640 81628
rect 86640 81572 86696 81628
rect 86696 81572 86700 81628
rect 86636 81568 86700 81572
rect 86716 81628 86780 81632
rect 86716 81572 86720 81628
rect 86720 81572 86776 81628
rect 86776 81572 86780 81628
rect 86716 81568 86780 81572
rect 6620 81084 6684 81088
rect 6620 81028 6624 81084
rect 6624 81028 6680 81084
rect 6680 81028 6684 81084
rect 6620 81024 6684 81028
rect 6700 81084 6764 81088
rect 6700 81028 6704 81084
rect 6704 81028 6760 81084
rect 6760 81028 6764 81084
rect 6700 81024 6764 81028
rect 6780 81084 6844 81088
rect 6780 81028 6784 81084
rect 6784 81028 6840 81084
rect 6840 81028 6844 81084
rect 6780 81024 6844 81028
rect 6860 81084 6924 81088
rect 6860 81028 6864 81084
rect 6864 81028 6920 81084
rect 6920 81028 6924 81084
rect 6860 81024 6924 81028
rect 87212 81084 87276 81088
rect 87212 81028 87216 81084
rect 87216 81028 87272 81084
rect 87272 81028 87276 81084
rect 87212 81024 87276 81028
rect 87292 81084 87356 81088
rect 87292 81028 87296 81084
rect 87296 81028 87352 81084
rect 87352 81028 87356 81084
rect 87292 81024 87356 81028
rect 87372 81084 87436 81088
rect 87372 81028 87376 81084
rect 87376 81028 87432 81084
rect 87432 81028 87436 81084
rect 87372 81024 87436 81028
rect 87452 81084 87516 81088
rect 87452 81028 87456 81084
rect 87456 81028 87512 81084
rect 87512 81028 87516 81084
rect 87452 81024 87516 81028
rect 5884 80540 5948 80544
rect 5884 80484 5888 80540
rect 5888 80484 5944 80540
rect 5944 80484 5948 80540
rect 5884 80480 5948 80484
rect 5964 80540 6028 80544
rect 5964 80484 5968 80540
rect 5968 80484 6024 80540
rect 6024 80484 6028 80540
rect 5964 80480 6028 80484
rect 6044 80540 6108 80544
rect 6044 80484 6048 80540
rect 6048 80484 6104 80540
rect 6104 80484 6108 80540
rect 6044 80480 6108 80484
rect 6124 80540 6188 80544
rect 6124 80484 6128 80540
rect 6128 80484 6184 80540
rect 6184 80484 6188 80540
rect 6124 80480 6188 80484
rect 86476 80540 86540 80544
rect 86476 80484 86480 80540
rect 86480 80484 86536 80540
rect 86536 80484 86540 80540
rect 86476 80480 86540 80484
rect 86556 80540 86620 80544
rect 86556 80484 86560 80540
rect 86560 80484 86616 80540
rect 86616 80484 86620 80540
rect 86556 80480 86620 80484
rect 86636 80540 86700 80544
rect 86636 80484 86640 80540
rect 86640 80484 86696 80540
rect 86696 80484 86700 80540
rect 86636 80480 86700 80484
rect 86716 80540 86780 80544
rect 86716 80484 86720 80540
rect 86720 80484 86776 80540
rect 86776 80484 86780 80540
rect 86716 80480 86780 80484
rect 6620 79996 6684 80000
rect 6620 79940 6624 79996
rect 6624 79940 6680 79996
rect 6680 79940 6684 79996
rect 6620 79936 6684 79940
rect 6700 79996 6764 80000
rect 6700 79940 6704 79996
rect 6704 79940 6760 79996
rect 6760 79940 6764 79996
rect 6700 79936 6764 79940
rect 6780 79996 6844 80000
rect 6780 79940 6784 79996
rect 6784 79940 6840 79996
rect 6840 79940 6844 79996
rect 6780 79936 6844 79940
rect 6860 79996 6924 80000
rect 6860 79940 6864 79996
rect 6864 79940 6920 79996
rect 6920 79940 6924 79996
rect 6860 79936 6924 79940
rect 87212 79996 87276 80000
rect 87212 79940 87216 79996
rect 87216 79940 87272 79996
rect 87272 79940 87276 79996
rect 87212 79936 87276 79940
rect 87292 79996 87356 80000
rect 87292 79940 87296 79996
rect 87296 79940 87352 79996
rect 87352 79940 87356 79996
rect 87292 79936 87356 79940
rect 87372 79996 87436 80000
rect 87372 79940 87376 79996
rect 87376 79940 87432 79996
rect 87432 79940 87436 79996
rect 87372 79936 87436 79940
rect 87452 79996 87516 80000
rect 87452 79940 87456 79996
rect 87456 79940 87512 79996
rect 87512 79940 87516 79996
rect 87452 79936 87516 79940
rect 5884 79452 5948 79456
rect 5884 79396 5888 79452
rect 5888 79396 5944 79452
rect 5944 79396 5948 79452
rect 5884 79392 5948 79396
rect 5964 79452 6028 79456
rect 5964 79396 5968 79452
rect 5968 79396 6024 79452
rect 6024 79396 6028 79452
rect 5964 79392 6028 79396
rect 6044 79452 6108 79456
rect 6044 79396 6048 79452
rect 6048 79396 6104 79452
rect 6104 79396 6108 79452
rect 6044 79392 6108 79396
rect 6124 79452 6188 79456
rect 6124 79396 6128 79452
rect 6128 79396 6184 79452
rect 6184 79396 6188 79452
rect 6124 79392 6188 79396
rect 86476 79452 86540 79456
rect 86476 79396 86480 79452
rect 86480 79396 86536 79452
rect 86536 79396 86540 79452
rect 86476 79392 86540 79396
rect 86556 79452 86620 79456
rect 86556 79396 86560 79452
rect 86560 79396 86616 79452
rect 86616 79396 86620 79452
rect 86556 79392 86620 79396
rect 86636 79452 86700 79456
rect 86636 79396 86640 79452
rect 86640 79396 86696 79452
rect 86696 79396 86700 79452
rect 86636 79392 86700 79396
rect 86716 79452 86780 79456
rect 86716 79396 86720 79452
rect 86720 79396 86776 79452
rect 86776 79396 86780 79452
rect 86716 79392 86780 79396
rect 6620 78908 6684 78912
rect 6620 78852 6624 78908
rect 6624 78852 6680 78908
rect 6680 78852 6684 78908
rect 6620 78848 6684 78852
rect 6700 78908 6764 78912
rect 6700 78852 6704 78908
rect 6704 78852 6760 78908
rect 6760 78852 6764 78908
rect 6700 78848 6764 78852
rect 6780 78908 6844 78912
rect 6780 78852 6784 78908
rect 6784 78852 6840 78908
rect 6840 78852 6844 78908
rect 6780 78848 6844 78852
rect 6860 78908 6924 78912
rect 6860 78852 6864 78908
rect 6864 78852 6920 78908
rect 6920 78852 6924 78908
rect 6860 78848 6924 78852
rect 87212 78908 87276 78912
rect 87212 78852 87216 78908
rect 87216 78852 87272 78908
rect 87272 78852 87276 78908
rect 87212 78848 87276 78852
rect 87292 78908 87356 78912
rect 87292 78852 87296 78908
rect 87296 78852 87352 78908
rect 87352 78852 87356 78908
rect 87292 78848 87356 78852
rect 87372 78908 87436 78912
rect 87372 78852 87376 78908
rect 87376 78852 87432 78908
rect 87432 78852 87436 78908
rect 87372 78848 87436 78852
rect 87452 78908 87516 78912
rect 87452 78852 87456 78908
rect 87456 78852 87512 78908
rect 87512 78852 87516 78908
rect 87452 78848 87516 78852
rect 5884 78364 5948 78368
rect 5884 78308 5888 78364
rect 5888 78308 5944 78364
rect 5944 78308 5948 78364
rect 5884 78304 5948 78308
rect 5964 78364 6028 78368
rect 5964 78308 5968 78364
rect 5968 78308 6024 78364
rect 6024 78308 6028 78364
rect 5964 78304 6028 78308
rect 6044 78364 6108 78368
rect 6044 78308 6048 78364
rect 6048 78308 6104 78364
rect 6104 78308 6108 78364
rect 6044 78304 6108 78308
rect 6124 78364 6188 78368
rect 6124 78308 6128 78364
rect 6128 78308 6184 78364
rect 6184 78308 6188 78364
rect 6124 78304 6188 78308
rect 86476 78364 86540 78368
rect 86476 78308 86480 78364
rect 86480 78308 86536 78364
rect 86536 78308 86540 78364
rect 86476 78304 86540 78308
rect 86556 78364 86620 78368
rect 86556 78308 86560 78364
rect 86560 78308 86616 78364
rect 86616 78308 86620 78364
rect 86556 78304 86620 78308
rect 86636 78364 86700 78368
rect 86636 78308 86640 78364
rect 86640 78308 86696 78364
rect 86696 78308 86700 78364
rect 86636 78304 86700 78308
rect 86716 78364 86780 78368
rect 86716 78308 86720 78364
rect 86720 78308 86776 78364
rect 86776 78308 86780 78364
rect 86716 78304 86780 78308
rect 6620 77820 6684 77824
rect 6620 77764 6624 77820
rect 6624 77764 6680 77820
rect 6680 77764 6684 77820
rect 6620 77760 6684 77764
rect 6700 77820 6764 77824
rect 6700 77764 6704 77820
rect 6704 77764 6760 77820
rect 6760 77764 6764 77820
rect 6700 77760 6764 77764
rect 6780 77820 6844 77824
rect 6780 77764 6784 77820
rect 6784 77764 6840 77820
rect 6840 77764 6844 77820
rect 6780 77760 6844 77764
rect 6860 77820 6924 77824
rect 6860 77764 6864 77820
rect 6864 77764 6920 77820
rect 6920 77764 6924 77820
rect 6860 77760 6924 77764
rect 87212 77820 87276 77824
rect 87212 77764 87216 77820
rect 87216 77764 87272 77820
rect 87272 77764 87276 77820
rect 87212 77760 87276 77764
rect 87292 77820 87356 77824
rect 87292 77764 87296 77820
rect 87296 77764 87352 77820
rect 87352 77764 87356 77820
rect 87292 77760 87356 77764
rect 87372 77820 87436 77824
rect 87372 77764 87376 77820
rect 87376 77764 87432 77820
rect 87432 77764 87436 77820
rect 87372 77760 87436 77764
rect 87452 77820 87516 77824
rect 87452 77764 87456 77820
rect 87456 77764 87512 77820
rect 87512 77764 87516 77820
rect 87452 77760 87516 77764
rect 5884 77276 5948 77280
rect 5884 77220 5888 77276
rect 5888 77220 5944 77276
rect 5944 77220 5948 77276
rect 5884 77216 5948 77220
rect 5964 77276 6028 77280
rect 5964 77220 5968 77276
rect 5968 77220 6024 77276
rect 6024 77220 6028 77276
rect 5964 77216 6028 77220
rect 6044 77276 6108 77280
rect 6044 77220 6048 77276
rect 6048 77220 6104 77276
rect 6104 77220 6108 77276
rect 6044 77216 6108 77220
rect 6124 77276 6188 77280
rect 6124 77220 6128 77276
rect 6128 77220 6184 77276
rect 6184 77220 6188 77276
rect 6124 77216 6188 77220
rect 86476 77276 86540 77280
rect 86476 77220 86480 77276
rect 86480 77220 86536 77276
rect 86536 77220 86540 77276
rect 86476 77216 86540 77220
rect 86556 77276 86620 77280
rect 86556 77220 86560 77276
rect 86560 77220 86616 77276
rect 86616 77220 86620 77276
rect 86556 77216 86620 77220
rect 86636 77276 86700 77280
rect 86636 77220 86640 77276
rect 86640 77220 86696 77276
rect 86696 77220 86700 77276
rect 86636 77216 86700 77220
rect 86716 77276 86780 77280
rect 86716 77220 86720 77276
rect 86720 77220 86776 77276
rect 86776 77220 86780 77276
rect 86716 77216 86780 77220
rect 6620 76732 6684 76736
rect 6620 76676 6624 76732
rect 6624 76676 6680 76732
rect 6680 76676 6684 76732
rect 6620 76672 6684 76676
rect 6700 76732 6764 76736
rect 6700 76676 6704 76732
rect 6704 76676 6760 76732
rect 6760 76676 6764 76732
rect 6700 76672 6764 76676
rect 6780 76732 6844 76736
rect 6780 76676 6784 76732
rect 6784 76676 6840 76732
rect 6840 76676 6844 76732
rect 6780 76672 6844 76676
rect 6860 76732 6924 76736
rect 6860 76676 6864 76732
rect 6864 76676 6920 76732
rect 6920 76676 6924 76732
rect 6860 76672 6924 76676
rect 87212 76732 87276 76736
rect 87212 76676 87216 76732
rect 87216 76676 87272 76732
rect 87272 76676 87276 76732
rect 87212 76672 87276 76676
rect 87292 76732 87356 76736
rect 87292 76676 87296 76732
rect 87296 76676 87352 76732
rect 87352 76676 87356 76732
rect 87292 76672 87356 76676
rect 87372 76732 87436 76736
rect 87372 76676 87376 76732
rect 87376 76676 87432 76732
rect 87432 76676 87436 76732
rect 87372 76672 87436 76676
rect 87452 76732 87516 76736
rect 87452 76676 87456 76732
rect 87456 76676 87512 76732
rect 87512 76676 87516 76732
rect 87452 76672 87516 76676
rect 5884 76188 5948 76192
rect 5884 76132 5888 76188
rect 5888 76132 5944 76188
rect 5944 76132 5948 76188
rect 5884 76128 5948 76132
rect 5964 76188 6028 76192
rect 5964 76132 5968 76188
rect 5968 76132 6024 76188
rect 6024 76132 6028 76188
rect 5964 76128 6028 76132
rect 6044 76188 6108 76192
rect 6044 76132 6048 76188
rect 6048 76132 6104 76188
rect 6104 76132 6108 76188
rect 6044 76128 6108 76132
rect 6124 76188 6188 76192
rect 6124 76132 6128 76188
rect 6128 76132 6184 76188
rect 6184 76132 6188 76188
rect 6124 76128 6188 76132
rect 86476 76188 86540 76192
rect 86476 76132 86480 76188
rect 86480 76132 86536 76188
rect 86536 76132 86540 76188
rect 86476 76128 86540 76132
rect 86556 76188 86620 76192
rect 86556 76132 86560 76188
rect 86560 76132 86616 76188
rect 86616 76132 86620 76188
rect 86556 76128 86620 76132
rect 86636 76188 86700 76192
rect 86636 76132 86640 76188
rect 86640 76132 86696 76188
rect 86696 76132 86700 76188
rect 86636 76128 86700 76132
rect 86716 76188 86780 76192
rect 86716 76132 86720 76188
rect 86720 76132 86776 76188
rect 86776 76132 86780 76188
rect 86716 76128 86780 76132
rect 6620 75644 6684 75648
rect 6620 75588 6624 75644
rect 6624 75588 6680 75644
rect 6680 75588 6684 75644
rect 6620 75584 6684 75588
rect 6700 75644 6764 75648
rect 6700 75588 6704 75644
rect 6704 75588 6760 75644
rect 6760 75588 6764 75644
rect 6700 75584 6764 75588
rect 6780 75644 6844 75648
rect 6780 75588 6784 75644
rect 6784 75588 6840 75644
rect 6840 75588 6844 75644
rect 6780 75584 6844 75588
rect 6860 75644 6924 75648
rect 6860 75588 6864 75644
rect 6864 75588 6920 75644
rect 6920 75588 6924 75644
rect 6860 75584 6924 75588
rect 87212 75644 87276 75648
rect 87212 75588 87216 75644
rect 87216 75588 87272 75644
rect 87272 75588 87276 75644
rect 87212 75584 87276 75588
rect 87292 75644 87356 75648
rect 87292 75588 87296 75644
rect 87296 75588 87352 75644
rect 87352 75588 87356 75644
rect 87292 75584 87356 75588
rect 87372 75644 87436 75648
rect 87372 75588 87376 75644
rect 87376 75588 87432 75644
rect 87432 75588 87436 75644
rect 87372 75584 87436 75588
rect 87452 75644 87516 75648
rect 87452 75588 87456 75644
rect 87456 75588 87512 75644
rect 87512 75588 87516 75644
rect 87452 75584 87516 75588
rect 5884 75100 5948 75104
rect 5884 75044 5888 75100
rect 5888 75044 5944 75100
rect 5944 75044 5948 75100
rect 5884 75040 5948 75044
rect 5964 75100 6028 75104
rect 5964 75044 5968 75100
rect 5968 75044 6024 75100
rect 6024 75044 6028 75100
rect 5964 75040 6028 75044
rect 6044 75100 6108 75104
rect 6044 75044 6048 75100
rect 6048 75044 6104 75100
rect 6104 75044 6108 75100
rect 6044 75040 6108 75044
rect 6124 75100 6188 75104
rect 6124 75044 6128 75100
rect 6128 75044 6184 75100
rect 6184 75044 6188 75100
rect 6124 75040 6188 75044
rect 86476 75100 86540 75104
rect 86476 75044 86480 75100
rect 86480 75044 86536 75100
rect 86536 75044 86540 75100
rect 86476 75040 86540 75044
rect 86556 75100 86620 75104
rect 86556 75044 86560 75100
rect 86560 75044 86616 75100
rect 86616 75044 86620 75100
rect 86556 75040 86620 75044
rect 86636 75100 86700 75104
rect 86636 75044 86640 75100
rect 86640 75044 86696 75100
rect 86696 75044 86700 75100
rect 86636 75040 86700 75044
rect 86716 75100 86780 75104
rect 86716 75044 86720 75100
rect 86720 75044 86776 75100
rect 86776 75044 86780 75100
rect 86716 75040 86780 75044
rect 6620 74556 6684 74560
rect 6620 74500 6624 74556
rect 6624 74500 6680 74556
rect 6680 74500 6684 74556
rect 6620 74496 6684 74500
rect 6700 74556 6764 74560
rect 6700 74500 6704 74556
rect 6704 74500 6760 74556
rect 6760 74500 6764 74556
rect 6700 74496 6764 74500
rect 6780 74556 6844 74560
rect 6780 74500 6784 74556
rect 6784 74500 6840 74556
rect 6840 74500 6844 74556
rect 6780 74496 6844 74500
rect 6860 74556 6924 74560
rect 6860 74500 6864 74556
rect 6864 74500 6920 74556
rect 6920 74500 6924 74556
rect 6860 74496 6924 74500
rect 87212 74556 87276 74560
rect 87212 74500 87216 74556
rect 87216 74500 87272 74556
rect 87272 74500 87276 74556
rect 87212 74496 87276 74500
rect 87292 74556 87356 74560
rect 87292 74500 87296 74556
rect 87296 74500 87352 74556
rect 87352 74500 87356 74556
rect 87292 74496 87356 74500
rect 87372 74556 87436 74560
rect 87372 74500 87376 74556
rect 87376 74500 87432 74556
rect 87432 74500 87436 74556
rect 87372 74496 87436 74500
rect 87452 74556 87516 74560
rect 87452 74500 87456 74556
rect 87456 74500 87512 74556
rect 87512 74500 87516 74556
rect 87452 74496 87516 74500
rect 5884 74012 5948 74016
rect 5884 73956 5888 74012
rect 5888 73956 5944 74012
rect 5944 73956 5948 74012
rect 5884 73952 5948 73956
rect 5964 74012 6028 74016
rect 5964 73956 5968 74012
rect 5968 73956 6024 74012
rect 6024 73956 6028 74012
rect 5964 73952 6028 73956
rect 6044 74012 6108 74016
rect 6044 73956 6048 74012
rect 6048 73956 6104 74012
rect 6104 73956 6108 74012
rect 6044 73952 6108 73956
rect 6124 74012 6188 74016
rect 6124 73956 6128 74012
rect 6128 73956 6184 74012
rect 6184 73956 6188 74012
rect 6124 73952 6188 73956
rect 86476 74012 86540 74016
rect 86476 73956 86480 74012
rect 86480 73956 86536 74012
rect 86536 73956 86540 74012
rect 86476 73952 86540 73956
rect 86556 74012 86620 74016
rect 86556 73956 86560 74012
rect 86560 73956 86616 74012
rect 86616 73956 86620 74012
rect 86556 73952 86620 73956
rect 86636 74012 86700 74016
rect 86636 73956 86640 74012
rect 86640 73956 86696 74012
rect 86696 73956 86700 74012
rect 86636 73952 86700 73956
rect 86716 74012 86780 74016
rect 86716 73956 86720 74012
rect 86720 73956 86776 74012
rect 86776 73956 86780 74012
rect 86716 73952 86780 73956
rect 6620 73468 6684 73472
rect 6620 73412 6624 73468
rect 6624 73412 6680 73468
rect 6680 73412 6684 73468
rect 6620 73408 6684 73412
rect 6700 73468 6764 73472
rect 6700 73412 6704 73468
rect 6704 73412 6760 73468
rect 6760 73412 6764 73468
rect 6700 73408 6764 73412
rect 6780 73468 6844 73472
rect 6780 73412 6784 73468
rect 6784 73412 6840 73468
rect 6840 73412 6844 73468
rect 6780 73408 6844 73412
rect 6860 73468 6924 73472
rect 6860 73412 6864 73468
rect 6864 73412 6920 73468
rect 6920 73412 6924 73468
rect 6860 73408 6924 73412
rect 87212 73468 87276 73472
rect 87212 73412 87216 73468
rect 87216 73412 87272 73468
rect 87272 73412 87276 73468
rect 87212 73408 87276 73412
rect 87292 73468 87356 73472
rect 87292 73412 87296 73468
rect 87296 73412 87352 73468
rect 87352 73412 87356 73468
rect 87292 73408 87356 73412
rect 87372 73468 87436 73472
rect 87372 73412 87376 73468
rect 87376 73412 87432 73468
rect 87432 73412 87436 73468
rect 87372 73408 87436 73412
rect 87452 73468 87516 73472
rect 87452 73412 87456 73468
rect 87456 73412 87512 73468
rect 87512 73412 87516 73468
rect 87452 73408 87516 73412
rect 5884 72924 5948 72928
rect 5884 72868 5888 72924
rect 5888 72868 5944 72924
rect 5944 72868 5948 72924
rect 5884 72864 5948 72868
rect 5964 72924 6028 72928
rect 5964 72868 5968 72924
rect 5968 72868 6024 72924
rect 6024 72868 6028 72924
rect 5964 72864 6028 72868
rect 6044 72924 6108 72928
rect 6044 72868 6048 72924
rect 6048 72868 6104 72924
rect 6104 72868 6108 72924
rect 6044 72864 6108 72868
rect 6124 72924 6188 72928
rect 6124 72868 6128 72924
rect 6128 72868 6184 72924
rect 6184 72868 6188 72924
rect 6124 72864 6188 72868
rect 86476 72924 86540 72928
rect 86476 72868 86480 72924
rect 86480 72868 86536 72924
rect 86536 72868 86540 72924
rect 86476 72864 86540 72868
rect 86556 72924 86620 72928
rect 86556 72868 86560 72924
rect 86560 72868 86616 72924
rect 86616 72868 86620 72924
rect 86556 72864 86620 72868
rect 86636 72924 86700 72928
rect 86636 72868 86640 72924
rect 86640 72868 86696 72924
rect 86696 72868 86700 72924
rect 86636 72864 86700 72868
rect 86716 72924 86780 72928
rect 86716 72868 86720 72924
rect 86720 72868 86776 72924
rect 86776 72868 86780 72924
rect 86716 72864 86780 72868
rect 6620 72380 6684 72384
rect 6620 72324 6624 72380
rect 6624 72324 6680 72380
rect 6680 72324 6684 72380
rect 6620 72320 6684 72324
rect 6700 72380 6764 72384
rect 6700 72324 6704 72380
rect 6704 72324 6760 72380
rect 6760 72324 6764 72380
rect 6700 72320 6764 72324
rect 6780 72380 6844 72384
rect 6780 72324 6784 72380
rect 6784 72324 6840 72380
rect 6840 72324 6844 72380
rect 6780 72320 6844 72324
rect 6860 72380 6924 72384
rect 6860 72324 6864 72380
rect 6864 72324 6920 72380
rect 6920 72324 6924 72380
rect 6860 72320 6924 72324
rect 87212 72380 87276 72384
rect 87212 72324 87216 72380
rect 87216 72324 87272 72380
rect 87272 72324 87276 72380
rect 87212 72320 87276 72324
rect 87292 72380 87356 72384
rect 87292 72324 87296 72380
rect 87296 72324 87352 72380
rect 87352 72324 87356 72380
rect 87292 72320 87356 72324
rect 87372 72380 87436 72384
rect 87372 72324 87376 72380
rect 87376 72324 87432 72380
rect 87432 72324 87436 72380
rect 87372 72320 87436 72324
rect 87452 72380 87516 72384
rect 87452 72324 87456 72380
rect 87456 72324 87512 72380
rect 87512 72324 87516 72380
rect 87452 72320 87516 72324
rect 5884 71836 5948 71840
rect 5884 71780 5888 71836
rect 5888 71780 5944 71836
rect 5944 71780 5948 71836
rect 5884 71776 5948 71780
rect 5964 71836 6028 71840
rect 5964 71780 5968 71836
rect 5968 71780 6024 71836
rect 6024 71780 6028 71836
rect 5964 71776 6028 71780
rect 6044 71836 6108 71840
rect 6044 71780 6048 71836
rect 6048 71780 6104 71836
rect 6104 71780 6108 71836
rect 6044 71776 6108 71780
rect 6124 71836 6188 71840
rect 6124 71780 6128 71836
rect 6128 71780 6184 71836
rect 6184 71780 6188 71836
rect 6124 71776 6188 71780
rect 86476 71836 86540 71840
rect 86476 71780 86480 71836
rect 86480 71780 86536 71836
rect 86536 71780 86540 71836
rect 86476 71776 86540 71780
rect 86556 71836 86620 71840
rect 86556 71780 86560 71836
rect 86560 71780 86616 71836
rect 86616 71780 86620 71836
rect 86556 71776 86620 71780
rect 86636 71836 86700 71840
rect 86636 71780 86640 71836
rect 86640 71780 86696 71836
rect 86696 71780 86700 71836
rect 86636 71776 86700 71780
rect 86716 71836 86780 71840
rect 86716 71780 86720 71836
rect 86720 71780 86776 71836
rect 86776 71780 86780 71836
rect 86716 71776 86780 71780
rect 6620 71292 6684 71296
rect 6620 71236 6624 71292
rect 6624 71236 6680 71292
rect 6680 71236 6684 71292
rect 6620 71232 6684 71236
rect 6700 71292 6764 71296
rect 6700 71236 6704 71292
rect 6704 71236 6760 71292
rect 6760 71236 6764 71292
rect 6700 71232 6764 71236
rect 6780 71292 6844 71296
rect 6780 71236 6784 71292
rect 6784 71236 6840 71292
rect 6840 71236 6844 71292
rect 6780 71232 6844 71236
rect 6860 71292 6924 71296
rect 6860 71236 6864 71292
rect 6864 71236 6920 71292
rect 6920 71236 6924 71292
rect 6860 71232 6924 71236
rect 87212 71292 87276 71296
rect 87212 71236 87216 71292
rect 87216 71236 87272 71292
rect 87272 71236 87276 71292
rect 87212 71232 87276 71236
rect 87292 71292 87356 71296
rect 87292 71236 87296 71292
rect 87296 71236 87352 71292
rect 87352 71236 87356 71292
rect 87292 71232 87356 71236
rect 87372 71292 87436 71296
rect 87372 71236 87376 71292
rect 87376 71236 87432 71292
rect 87432 71236 87436 71292
rect 87372 71232 87436 71236
rect 87452 71292 87516 71296
rect 87452 71236 87456 71292
rect 87456 71236 87512 71292
rect 87512 71236 87516 71292
rect 87452 71232 87516 71236
rect 5884 70748 5948 70752
rect 5884 70692 5888 70748
rect 5888 70692 5944 70748
rect 5944 70692 5948 70748
rect 5884 70688 5948 70692
rect 5964 70748 6028 70752
rect 5964 70692 5968 70748
rect 5968 70692 6024 70748
rect 6024 70692 6028 70748
rect 5964 70688 6028 70692
rect 6044 70748 6108 70752
rect 6044 70692 6048 70748
rect 6048 70692 6104 70748
rect 6104 70692 6108 70748
rect 6044 70688 6108 70692
rect 6124 70748 6188 70752
rect 6124 70692 6128 70748
rect 6128 70692 6184 70748
rect 6184 70692 6188 70748
rect 6124 70688 6188 70692
rect 86476 70748 86540 70752
rect 86476 70692 86480 70748
rect 86480 70692 86536 70748
rect 86536 70692 86540 70748
rect 86476 70688 86540 70692
rect 86556 70748 86620 70752
rect 86556 70692 86560 70748
rect 86560 70692 86616 70748
rect 86616 70692 86620 70748
rect 86556 70688 86620 70692
rect 86636 70748 86700 70752
rect 86636 70692 86640 70748
rect 86640 70692 86696 70748
rect 86696 70692 86700 70748
rect 86636 70688 86700 70692
rect 86716 70748 86780 70752
rect 86716 70692 86720 70748
rect 86720 70692 86776 70748
rect 86776 70692 86780 70748
rect 86716 70688 86780 70692
rect 6620 70204 6684 70208
rect 6620 70148 6624 70204
rect 6624 70148 6680 70204
rect 6680 70148 6684 70204
rect 6620 70144 6684 70148
rect 6700 70204 6764 70208
rect 6700 70148 6704 70204
rect 6704 70148 6760 70204
rect 6760 70148 6764 70204
rect 6700 70144 6764 70148
rect 6780 70204 6844 70208
rect 6780 70148 6784 70204
rect 6784 70148 6840 70204
rect 6840 70148 6844 70204
rect 6780 70144 6844 70148
rect 6860 70204 6924 70208
rect 6860 70148 6864 70204
rect 6864 70148 6920 70204
rect 6920 70148 6924 70204
rect 6860 70144 6924 70148
rect 87212 70204 87276 70208
rect 87212 70148 87216 70204
rect 87216 70148 87272 70204
rect 87272 70148 87276 70204
rect 87212 70144 87276 70148
rect 87292 70204 87356 70208
rect 87292 70148 87296 70204
rect 87296 70148 87352 70204
rect 87352 70148 87356 70204
rect 87292 70144 87356 70148
rect 87372 70204 87436 70208
rect 87372 70148 87376 70204
rect 87376 70148 87432 70204
rect 87432 70148 87436 70204
rect 87372 70144 87436 70148
rect 87452 70204 87516 70208
rect 87452 70148 87456 70204
rect 87456 70148 87512 70204
rect 87512 70148 87516 70204
rect 87452 70144 87516 70148
rect 5884 69660 5948 69664
rect 5884 69604 5888 69660
rect 5888 69604 5944 69660
rect 5944 69604 5948 69660
rect 5884 69600 5948 69604
rect 5964 69660 6028 69664
rect 5964 69604 5968 69660
rect 5968 69604 6024 69660
rect 6024 69604 6028 69660
rect 5964 69600 6028 69604
rect 6044 69660 6108 69664
rect 6044 69604 6048 69660
rect 6048 69604 6104 69660
rect 6104 69604 6108 69660
rect 6044 69600 6108 69604
rect 6124 69660 6188 69664
rect 6124 69604 6128 69660
rect 6128 69604 6184 69660
rect 6184 69604 6188 69660
rect 6124 69600 6188 69604
rect 86476 69660 86540 69664
rect 86476 69604 86480 69660
rect 86480 69604 86536 69660
rect 86536 69604 86540 69660
rect 86476 69600 86540 69604
rect 86556 69660 86620 69664
rect 86556 69604 86560 69660
rect 86560 69604 86616 69660
rect 86616 69604 86620 69660
rect 86556 69600 86620 69604
rect 86636 69660 86700 69664
rect 86636 69604 86640 69660
rect 86640 69604 86696 69660
rect 86696 69604 86700 69660
rect 86636 69600 86700 69604
rect 86716 69660 86780 69664
rect 86716 69604 86720 69660
rect 86720 69604 86776 69660
rect 86776 69604 86780 69660
rect 86716 69600 86780 69604
rect 6620 69116 6684 69120
rect 6620 69060 6624 69116
rect 6624 69060 6680 69116
rect 6680 69060 6684 69116
rect 6620 69056 6684 69060
rect 6700 69116 6764 69120
rect 6700 69060 6704 69116
rect 6704 69060 6760 69116
rect 6760 69060 6764 69116
rect 6700 69056 6764 69060
rect 6780 69116 6844 69120
rect 6780 69060 6784 69116
rect 6784 69060 6840 69116
rect 6840 69060 6844 69116
rect 6780 69056 6844 69060
rect 6860 69116 6924 69120
rect 6860 69060 6864 69116
rect 6864 69060 6920 69116
rect 6920 69060 6924 69116
rect 6860 69056 6924 69060
rect 87212 69116 87276 69120
rect 87212 69060 87216 69116
rect 87216 69060 87272 69116
rect 87272 69060 87276 69116
rect 87212 69056 87276 69060
rect 87292 69116 87356 69120
rect 87292 69060 87296 69116
rect 87296 69060 87352 69116
rect 87352 69060 87356 69116
rect 87292 69056 87356 69060
rect 87372 69116 87436 69120
rect 87372 69060 87376 69116
rect 87376 69060 87432 69116
rect 87432 69060 87436 69116
rect 87372 69056 87436 69060
rect 87452 69116 87516 69120
rect 87452 69060 87456 69116
rect 87456 69060 87512 69116
rect 87512 69060 87516 69116
rect 87452 69056 87516 69060
rect 5884 68572 5948 68576
rect 5884 68516 5888 68572
rect 5888 68516 5944 68572
rect 5944 68516 5948 68572
rect 5884 68512 5948 68516
rect 5964 68572 6028 68576
rect 5964 68516 5968 68572
rect 5968 68516 6024 68572
rect 6024 68516 6028 68572
rect 5964 68512 6028 68516
rect 6044 68572 6108 68576
rect 6044 68516 6048 68572
rect 6048 68516 6104 68572
rect 6104 68516 6108 68572
rect 6044 68512 6108 68516
rect 6124 68572 6188 68576
rect 6124 68516 6128 68572
rect 6128 68516 6184 68572
rect 6184 68516 6188 68572
rect 6124 68512 6188 68516
rect 86476 68572 86540 68576
rect 86476 68516 86480 68572
rect 86480 68516 86536 68572
rect 86536 68516 86540 68572
rect 86476 68512 86540 68516
rect 86556 68572 86620 68576
rect 86556 68516 86560 68572
rect 86560 68516 86616 68572
rect 86616 68516 86620 68572
rect 86556 68512 86620 68516
rect 86636 68572 86700 68576
rect 86636 68516 86640 68572
rect 86640 68516 86696 68572
rect 86696 68516 86700 68572
rect 86636 68512 86700 68516
rect 86716 68572 86780 68576
rect 86716 68516 86720 68572
rect 86720 68516 86776 68572
rect 86776 68516 86780 68572
rect 86716 68512 86780 68516
rect 6620 68028 6684 68032
rect 6620 67972 6624 68028
rect 6624 67972 6680 68028
rect 6680 67972 6684 68028
rect 6620 67968 6684 67972
rect 6700 68028 6764 68032
rect 6700 67972 6704 68028
rect 6704 67972 6760 68028
rect 6760 67972 6764 68028
rect 6700 67968 6764 67972
rect 6780 68028 6844 68032
rect 6780 67972 6784 68028
rect 6784 67972 6840 68028
rect 6840 67972 6844 68028
rect 6780 67968 6844 67972
rect 6860 68028 6924 68032
rect 6860 67972 6864 68028
rect 6864 67972 6920 68028
rect 6920 67972 6924 68028
rect 6860 67968 6924 67972
rect 87212 68028 87276 68032
rect 87212 67972 87216 68028
rect 87216 67972 87272 68028
rect 87272 67972 87276 68028
rect 87212 67968 87276 67972
rect 87292 68028 87356 68032
rect 87292 67972 87296 68028
rect 87296 67972 87352 68028
rect 87352 67972 87356 68028
rect 87292 67968 87356 67972
rect 87372 68028 87436 68032
rect 87372 67972 87376 68028
rect 87376 67972 87432 68028
rect 87432 67972 87436 68028
rect 87372 67968 87436 67972
rect 87452 68028 87516 68032
rect 87452 67972 87456 68028
rect 87456 67972 87512 68028
rect 87512 67972 87516 68028
rect 87452 67968 87516 67972
rect 5884 67484 5948 67488
rect 5884 67428 5888 67484
rect 5888 67428 5944 67484
rect 5944 67428 5948 67484
rect 5884 67424 5948 67428
rect 5964 67484 6028 67488
rect 5964 67428 5968 67484
rect 5968 67428 6024 67484
rect 6024 67428 6028 67484
rect 5964 67424 6028 67428
rect 6044 67484 6108 67488
rect 6044 67428 6048 67484
rect 6048 67428 6104 67484
rect 6104 67428 6108 67484
rect 6044 67424 6108 67428
rect 6124 67484 6188 67488
rect 6124 67428 6128 67484
rect 6128 67428 6184 67484
rect 6184 67428 6188 67484
rect 6124 67424 6188 67428
rect 86476 67484 86540 67488
rect 86476 67428 86480 67484
rect 86480 67428 86536 67484
rect 86536 67428 86540 67484
rect 86476 67424 86540 67428
rect 86556 67484 86620 67488
rect 86556 67428 86560 67484
rect 86560 67428 86616 67484
rect 86616 67428 86620 67484
rect 86556 67424 86620 67428
rect 86636 67484 86700 67488
rect 86636 67428 86640 67484
rect 86640 67428 86696 67484
rect 86696 67428 86700 67484
rect 86636 67424 86700 67428
rect 86716 67484 86780 67488
rect 86716 67428 86720 67484
rect 86720 67428 86776 67484
rect 86776 67428 86780 67484
rect 86716 67424 86780 67428
rect 6620 66940 6684 66944
rect 6620 66884 6624 66940
rect 6624 66884 6680 66940
rect 6680 66884 6684 66940
rect 6620 66880 6684 66884
rect 6700 66940 6764 66944
rect 6700 66884 6704 66940
rect 6704 66884 6760 66940
rect 6760 66884 6764 66940
rect 6700 66880 6764 66884
rect 6780 66940 6844 66944
rect 6780 66884 6784 66940
rect 6784 66884 6840 66940
rect 6840 66884 6844 66940
rect 6780 66880 6844 66884
rect 6860 66940 6924 66944
rect 6860 66884 6864 66940
rect 6864 66884 6920 66940
rect 6920 66884 6924 66940
rect 6860 66880 6924 66884
rect 87212 66940 87276 66944
rect 87212 66884 87216 66940
rect 87216 66884 87272 66940
rect 87272 66884 87276 66940
rect 87212 66880 87276 66884
rect 87292 66940 87356 66944
rect 87292 66884 87296 66940
rect 87296 66884 87352 66940
rect 87352 66884 87356 66940
rect 87292 66880 87356 66884
rect 87372 66940 87436 66944
rect 87372 66884 87376 66940
rect 87376 66884 87432 66940
rect 87432 66884 87436 66940
rect 87372 66880 87436 66884
rect 87452 66940 87516 66944
rect 87452 66884 87456 66940
rect 87456 66884 87512 66940
rect 87512 66884 87516 66940
rect 87452 66880 87516 66884
rect 5884 66396 5948 66400
rect 5884 66340 5888 66396
rect 5888 66340 5944 66396
rect 5944 66340 5948 66396
rect 5884 66336 5948 66340
rect 5964 66396 6028 66400
rect 5964 66340 5968 66396
rect 5968 66340 6024 66396
rect 6024 66340 6028 66396
rect 5964 66336 6028 66340
rect 6044 66396 6108 66400
rect 6044 66340 6048 66396
rect 6048 66340 6104 66396
rect 6104 66340 6108 66396
rect 6044 66336 6108 66340
rect 6124 66396 6188 66400
rect 6124 66340 6128 66396
rect 6128 66340 6184 66396
rect 6184 66340 6188 66396
rect 6124 66336 6188 66340
rect 86476 66396 86540 66400
rect 86476 66340 86480 66396
rect 86480 66340 86536 66396
rect 86536 66340 86540 66396
rect 86476 66336 86540 66340
rect 86556 66396 86620 66400
rect 86556 66340 86560 66396
rect 86560 66340 86616 66396
rect 86616 66340 86620 66396
rect 86556 66336 86620 66340
rect 86636 66396 86700 66400
rect 86636 66340 86640 66396
rect 86640 66340 86696 66396
rect 86696 66340 86700 66396
rect 86636 66336 86700 66340
rect 86716 66396 86780 66400
rect 86716 66340 86720 66396
rect 86720 66340 86776 66396
rect 86776 66340 86780 66396
rect 86716 66336 86780 66340
rect 6620 65852 6684 65856
rect 6620 65796 6624 65852
rect 6624 65796 6680 65852
rect 6680 65796 6684 65852
rect 6620 65792 6684 65796
rect 6700 65852 6764 65856
rect 6700 65796 6704 65852
rect 6704 65796 6760 65852
rect 6760 65796 6764 65852
rect 6700 65792 6764 65796
rect 6780 65852 6844 65856
rect 6780 65796 6784 65852
rect 6784 65796 6840 65852
rect 6840 65796 6844 65852
rect 6780 65792 6844 65796
rect 6860 65852 6924 65856
rect 6860 65796 6864 65852
rect 6864 65796 6920 65852
rect 6920 65796 6924 65852
rect 6860 65792 6924 65796
rect 87212 65852 87276 65856
rect 87212 65796 87216 65852
rect 87216 65796 87272 65852
rect 87272 65796 87276 65852
rect 87212 65792 87276 65796
rect 87292 65852 87356 65856
rect 87292 65796 87296 65852
rect 87296 65796 87352 65852
rect 87352 65796 87356 65852
rect 87292 65792 87356 65796
rect 87372 65852 87436 65856
rect 87372 65796 87376 65852
rect 87376 65796 87432 65852
rect 87432 65796 87436 65852
rect 87372 65792 87436 65796
rect 87452 65852 87516 65856
rect 87452 65796 87456 65852
rect 87456 65796 87512 65852
rect 87512 65796 87516 65852
rect 87452 65792 87516 65796
rect 5884 65308 5948 65312
rect 5884 65252 5888 65308
rect 5888 65252 5944 65308
rect 5944 65252 5948 65308
rect 5884 65248 5948 65252
rect 5964 65308 6028 65312
rect 5964 65252 5968 65308
rect 5968 65252 6024 65308
rect 6024 65252 6028 65308
rect 5964 65248 6028 65252
rect 6044 65308 6108 65312
rect 6044 65252 6048 65308
rect 6048 65252 6104 65308
rect 6104 65252 6108 65308
rect 6044 65248 6108 65252
rect 6124 65308 6188 65312
rect 6124 65252 6128 65308
rect 6128 65252 6184 65308
rect 6184 65252 6188 65308
rect 6124 65248 6188 65252
rect 86476 65308 86540 65312
rect 86476 65252 86480 65308
rect 86480 65252 86536 65308
rect 86536 65252 86540 65308
rect 86476 65248 86540 65252
rect 86556 65308 86620 65312
rect 86556 65252 86560 65308
rect 86560 65252 86616 65308
rect 86616 65252 86620 65308
rect 86556 65248 86620 65252
rect 86636 65308 86700 65312
rect 86636 65252 86640 65308
rect 86640 65252 86696 65308
rect 86696 65252 86700 65308
rect 86636 65248 86700 65252
rect 86716 65308 86780 65312
rect 86716 65252 86720 65308
rect 86720 65252 86776 65308
rect 86776 65252 86780 65308
rect 86716 65248 86780 65252
rect 6620 64764 6684 64768
rect 6620 64708 6624 64764
rect 6624 64708 6680 64764
rect 6680 64708 6684 64764
rect 6620 64704 6684 64708
rect 6700 64764 6764 64768
rect 6700 64708 6704 64764
rect 6704 64708 6760 64764
rect 6760 64708 6764 64764
rect 6700 64704 6764 64708
rect 6780 64764 6844 64768
rect 6780 64708 6784 64764
rect 6784 64708 6840 64764
rect 6840 64708 6844 64764
rect 6780 64704 6844 64708
rect 6860 64764 6924 64768
rect 6860 64708 6864 64764
rect 6864 64708 6920 64764
rect 6920 64708 6924 64764
rect 6860 64704 6924 64708
rect 87212 64764 87276 64768
rect 87212 64708 87216 64764
rect 87216 64708 87272 64764
rect 87272 64708 87276 64764
rect 87212 64704 87276 64708
rect 87292 64764 87356 64768
rect 87292 64708 87296 64764
rect 87296 64708 87352 64764
rect 87352 64708 87356 64764
rect 87292 64704 87356 64708
rect 87372 64764 87436 64768
rect 87372 64708 87376 64764
rect 87376 64708 87432 64764
rect 87432 64708 87436 64764
rect 87372 64704 87436 64708
rect 87452 64764 87516 64768
rect 87452 64708 87456 64764
rect 87456 64708 87512 64764
rect 87512 64708 87516 64764
rect 87452 64704 87516 64708
rect 5884 64220 5948 64224
rect 5884 64164 5888 64220
rect 5888 64164 5944 64220
rect 5944 64164 5948 64220
rect 5884 64160 5948 64164
rect 5964 64220 6028 64224
rect 5964 64164 5968 64220
rect 5968 64164 6024 64220
rect 6024 64164 6028 64220
rect 5964 64160 6028 64164
rect 6044 64220 6108 64224
rect 6044 64164 6048 64220
rect 6048 64164 6104 64220
rect 6104 64164 6108 64220
rect 6044 64160 6108 64164
rect 6124 64220 6188 64224
rect 6124 64164 6128 64220
rect 6128 64164 6184 64220
rect 6184 64164 6188 64220
rect 6124 64160 6188 64164
rect 86476 64220 86540 64224
rect 86476 64164 86480 64220
rect 86480 64164 86536 64220
rect 86536 64164 86540 64220
rect 86476 64160 86540 64164
rect 86556 64220 86620 64224
rect 86556 64164 86560 64220
rect 86560 64164 86616 64220
rect 86616 64164 86620 64220
rect 86556 64160 86620 64164
rect 86636 64220 86700 64224
rect 86636 64164 86640 64220
rect 86640 64164 86696 64220
rect 86696 64164 86700 64220
rect 86636 64160 86700 64164
rect 86716 64220 86780 64224
rect 86716 64164 86720 64220
rect 86720 64164 86776 64220
rect 86776 64164 86780 64220
rect 86716 64160 86780 64164
rect 6620 63676 6684 63680
rect 6620 63620 6624 63676
rect 6624 63620 6680 63676
rect 6680 63620 6684 63676
rect 6620 63616 6684 63620
rect 6700 63676 6764 63680
rect 6700 63620 6704 63676
rect 6704 63620 6760 63676
rect 6760 63620 6764 63676
rect 6700 63616 6764 63620
rect 6780 63676 6844 63680
rect 6780 63620 6784 63676
rect 6784 63620 6840 63676
rect 6840 63620 6844 63676
rect 6780 63616 6844 63620
rect 6860 63676 6924 63680
rect 6860 63620 6864 63676
rect 6864 63620 6920 63676
rect 6920 63620 6924 63676
rect 6860 63616 6924 63620
rect 87212 63676 87276 63680
rect 87212 63620 87216 63676
rect 87216 63620 87272 63676
rect 87272 63620 87276 63676
rect 87212 63616 87276 63620
rect 87292 63676 87356 63680
rect 87292 63620 87296 63676
rect 87296 63620 87352 63676
rect 87352 63620 87356 63676
rect 87292 63616 87356 63620
rect 87372 63676 87436 63680
rect 87372 63620 87376 63676
rect 87376 63620 87432 63676
rect 87432 63620 87436 63676
rect 87372 63616 87436 63620
rect 87452 63676 87516 63680
rect 87452 63620 87456 63676
rect 87456 63620 87512 63676
rect 87512 63620 87516 63676
rect 87452 63616 87516 63620
rect 5884 63132 5948 63136
rect 5884 63076 5888 63132
rect 5888 63076 5944 63132
rect 5944 63076 5948 63132
rect 5884 63072 5948 63076
rect 5964 63132 6028 63136
rect 5964 63076 5968 63132
rect 5968 63076 6024 63132
rect 6024 63076 6028 63132
rect 5964 63072 6028 63076
rect 6044 63132 6108 63136
rect 6044 63076 6048 63132
rect 6048 63076 6104 63132
rect 6104 63076 6108 63132
rect 6044 63072 6108 63076
rect 6124 63132 6188 63136
rect 6124 63076 6128 63132
rect 6128 63076 6184 63132
rect 6184 63076 6188 63132
rect 6124 63072 6188 63076
rect 86476 63132 86540 63136
rect 86476 63076 86480 63132
rect 86480 63076 86536 63132
rect 86536 63076 86540 63132
rect 86476 63072 86540 63076
rect 86556 63132 86620 63136
rect 86556 63076 86560 63132
rect 86560 63076 86616 63132
rect 86616 63076 86620 63132
rect 86556 63072 86620 63076
rect 86636 63132 86700 63136
rect 86636 63076 86640 63132
rect 86640 63076 86696 63132
rect 86696 63076 86700 63132
rect 86636 63072 86700 63076
rect 86716 63132 86780 63136
rect 86716 63076 86720 63132
rect 86720 63076 86776 63132
rect 86776 63076 86780 63132
rect 86716 63072 86780 63076
rect 6620 62588 6684 62592
rect 6620 62532 6624 62588
rect 6624 62532 6680 62588
rect 6680 62532 6684 62588
rect 6620 62528 6684 62532
rect 6700 62588 6764 62592
rect 6700 62532 6704 62588
rect 6704 62532 6760 62588
rect 6760 62532 6764 62588
rect 6700 62528 6764 62532
rect 6780 62588 6844 62592
rect 6780 62532 6784 62588
rect 6784 62532 6840 62588
rect 6840 62532 6844 62588
rect 6780 62528 6844 62532
rect 6860 62588 6924 62592
rect 6860 62532 6864 62588
rect 6864 62532 6920 62588
rect 6920 62532 6924 62588
rect 6860 62528 6924 62532
rect 87212 62588 87276 62592
rect 87212 62532 87216 62588
rect 87216 62532 87272 62588
rect 87272 62532 87276 62588
rect 87212 62528 87276 62532
rect 87292 62588 87356 62592
rect 87292 62532 87296 62588
rect 87296 62532 87352 62588
rect 87352 62532 87356 62588
rect 87292 62528 87356 62532
rect 87372 62588 87436 62592
rect 87372 62532 87376 62588
rect 87376 62532 87432 62588
rect 87432 62532 87436 62588
rect 87372 62528 87436 62532
rect 87452 62588 87516 62592
rect 87452 62532 87456 62588
rect 87456 62532 87512 62588
rect 87512 62532 87516 62588
rect 87452 62528 87516 62532
rect 5884 62044 5948 62048
rect 5884 61988 5888 62044
rect 5888 61988 5944 62044
rect 5944 61988 5948 62044
rect 5884 61984 5948 61988
rect 5964 62044 6028 62048
rect 5964 61988 5968 62044
rect 5968 61988 6024 62044
rect 6024 61988 6028 62044
rect 5964 61984 6028 61988
rect 6044 62044 6108 62048
rect 6044 61988 6048 62044
rect 6048 61988 6104 62044
rect 6104 61988 6108 62044
rect 6044 61984 6108 61988
rect 6124 62044 6188 62048
rect 6124 61988 6128 62044
rect 6128 61988 6184 62044
rect 6184 61988 6188 62044
rect 6124 61984 6188 61988
rect 86476 62044 86540 62048
rect 86476 61988 86480 62044
rect 86480 61988 86536 62044
rect 86536 61988 86540 62044
rect 86476 61984 86540 61988
rect 86556 62044 86620 62048
rect 86556 61988 86560 62044
rect 86560 61988 86616 62044
rect 86616 61988 86620 62044
rect 86556 61984 86620 61988
rect 86636 62044 86700 62048
rect 86636 61988 86640 62044
rect 86640 61988 86696 62044
rect 86696 61988 86700 62044
rect 86636 61984 86700 61988
rect 86716 62044 86780 62048
rect 86716 61988 86720 62044
rect 86720 61988 86776 62044
rect 86776 61988 86780 62044
rect 86716 61984 86780 61988
rect 6620 61500 6684 61504
rect 6620 61444 6624 61500
rect 6624 61444 6680 61500
rect 6680 61444 6684 61500
rect 6620 61440 6684 61444
rect 6700 61500 6764 61504
rect 6700 61444 6704 61500
rect 6704 61444 6760 61500
rect 6760 61444 6764 61500
rect 6700 61440 6764 61444
rect 6780 61500 6844 61504
rect 6780 61444 6784 61500
rect 6784 61444 6840 61500
rect 6840 61444 6844 61500
rect 6780 61440 6844 61444
rect 6860 61500 6924 61504
rect 6860 61444 6864 61500
rect 6864 61444 6920 61500
rect 6920 61444 6924 61500
rect 6860 61440 6924 61444
rect 87212 61500 87276 61504
rect 87212 61444 87216 61500
rect 87216 61444 87272 61500
rect 87272 61444 87276 61500
rect 87212 61440 87276 61444
rect 87292 61500 87356 61504
rect 87292 61444 87296 61500
rect 87296 61444 87352 61500
rect 87352 61444 87356 61500
rect 87292 61440 87356 61444
rect 87372 61500 87436 61504
rect 87372 61444 87376 61500
rect 87376 61444 87432 61500
rect 87432 61444 87436 61500
rect 87372 61440 87436 61444
rect 87452 61500 87516 61504
rect 87452 61444 87456 61500
rect 87456 61444 87512 61500
rect 87512 61444 87516 61500
rect 87452 61440 87516 61444
rect 5884 60956 5948 60960
rect 5884 60900 5888 60956
rect 5888 60900 5944 60956
rect 5944 60900 5948 60956
rect 5884 60896 5948 60900
rect 5964 60956 6028 60960
rect 5964 60900 5968 60956
rect 5968 60900 6024 60956
rect 6024 60900 6028 60956
rect 5964 60896 6028 60900
rect 6044 60956 6108 60960
rect 6044 60900 6048 60956
rect 6048 60900 6104 60956
rect 6104 60900 6108 60956
rect 6044 60896 6108 60900
rect 6124 60956 6188 60960
rect 6124 60900 6128 60956
rect 6128 60900 6184 60956
rect 6184 60900 6188 60956
rect 6124 60896 6188 60900
rect 86476 60956 86540 60960
rect 86476 60900 86480 60956
rect 86480 60900 86536 60956
rect 86536 60900 86540 60956
rect 86476 60896 86540 60900
rect 86556 60956 86620 60960
rect 86556 60900 86560 60956
rect 86560 60900 86616 60956
rect 86616 60900 86620 60956
rect 86556 60896 86620 60900
rect 86636 60956 86700 60960
rect 86636 60900 86640 60956
rect 86640 60900 86696 60956
rect 86696 60900 86700 60956
rect 86636 60896 86700 60900
rect 86716 60956 86780 60960
rect 86716 60900 86720 60956
rect 86720 60900 86776 60956
rect 86776 60900 86780 60956
rect 86716 60896 86780 60900
rect 6620 60412 6684 60416
rect 6620 60356 6624 60412
rect 6624 60356 6680 60412
rect 6680 60356 6684 60412
rect 6620 60352 6684 60356
rect 6700 60412 6764 60416
rect 6700 60356 6704 60412
rect 6704 60356 6760 60412
rect 6760 60356 6764 60412
rect 6700 60352 6764 60356
rect 6780 60412 6844 60416
rect 6780 60356 6784 60412
rect 6784 60356 6840 60412
rect 6840 60356 6844 60412
rect 6780 60352 6844 60356
rect 6860 60412 6924 60416
rect 6860 60356 6864 60412
rect 6864 60356 6920 60412
rect 6920 60356 6924 60412
rect 6860 60352 6924 60356
rect 87212 60412 87276 60416
rect 87212 60356 87216 60412
rect 87216 60356 87272 60412
rect 87272 60356 87276 60412
rect 87212 60352 87276 60356
rect 87292 60412 87356 60416
rect 87292 60356 87296 60412
rect 87296 60356 87352 60412
rect 87352 60356 87356 60412
rect 87292 60352 87356 60356
rect 87372 60412 87436 60416
rect 87372 60356 87376 60412
rect 87376 60356 87432 60412
rect 87432 60356 87436 60412
rect 87372 60352 87436 60356
rect 87452 60412 87516 60416
rect 87452 60356 87456 60412
rect 87456 60356 87512 60412
rect 87512 60356 87516 60412
rect 87452 60352 87516 60356
rect 5884 59868 5948 59872
rect 5884 59812 5888 59868
rect 5888 59812 5944 59868
rect 5944 59812 5948 59868
rect 5884 59808 5948 59812
rect 5964 59868 6028 59872
rect 5964 59812 5968 59868
rect 5968 59812 6024 59868
rect 6024 59812 6028 59868
rect 5964 59808 6028 59812
rect 6044 59868 6108 59872
rect 6044 59812 6048 59868
rect 6048 59812 6104 59868
rect 6104 59812 6108 59868
rect 6044 59808 6108 59812
rect 6124 59868 6188 59872
rect 6124 59812 6128 59868
rect 6128 59812 6184 59868
rect 6184 59812 6188 59868
rect 6124 59808 6188 59812
rect 86476 59868 86540 59872
rect 86476 59812 86480 59868
rect 86480 59812 86536 59868
rect 86536 59812 86540 59868
rect 86476 59808 86540 59812
rect 86556 59868 86620 59872
rect 86556 59812 86560 59868
rect 86560 59812 86616 59868
rect 86616 59812 86620 59868
rect 86556 59808 86620 59812
rect 86636 59868 86700 59872
rect 86636 59812 86640 59868
rect 86640 59812 86696 59868
rect 86696 59812 86700 59868
rect 86636 59808 86700 59812
rect 86716 59868 86780 59872
rect 86716 59812 86720 59868
rect 86720 59812 86776 59868
rect 86776 59812 86780 59868
rect 86716 59808 86780 59812
rect 6620 59324 6684 59328
rect 6620 59268 6624 59324
rect 6624 59268 6680 59324
rect 6680 59268 6684 59324
rect 6620 59264 6684 59268
rect 6700 59324 6764 59328
rect 6700 59268 6704 59324
rect 6704 59268 6760 59324
rect 6760 59268 6764 59324
rect 6700 59264 6764 59268
rect 6780 59324 6844 59328
rect 6780 59268 6784 59324
rect 6784 59268 6840 59324
rect 6840 59268 6844 59324
rect 6780 59264 6844 59268
rect 6860 59324 6924 59328
rect 6860 59268 6864 59324
rect 6864 59268 6920 59324
rect 6920 59268 6924 59324
rect 6860 59264 6924 59268
rect 87212 59324 87276 59328
rect 87212 59268 87216 59324
rect 87216 59268 87272 59324
rect 87272 59268 87276 59324
rect 87212 59264 87276 59268
rect 87292 59324 87356 59328
rect 87292 59268 87296 59324
rect 87296 59268 87352 59324
rect 87352 59268 87356 59324
rect 87292 59264 87356 59268
rect 87372 59324 87436 59328
rect 87372 59268 87376 59324
rect 87376 59268 87432 59324
rect 87432 59268 87436 59324
rect 87372 59264 87436 59268
rect 87452 59324 87516 59328
rect 87452 59268 87456 59324
rect 87456 59268 87512 59324
rect 87512 59268 87516 59324
rect 87452 59264 87516 59268
rect 5884 58780 5948 58784
rect 5884 58724 5888 58780
rect 5888 58724 5944 58780
rect 5944 58724 5948 58780
rect 5884 58720 5948 58724
rect 5964 58780 6028 58784
rect 5964 58724 5968 58780
rect 5968 58724 6024 58780
rect 6024 58724 6028 58780
rect 5964 58720 6028 58724
rect 6044 58780 6108 58784
rect 6044 58724 6048 58780
rect 6048 58724 6104 58780
rect 6104 58724 6108 58780
rect 6044 58720 6108 58724
rect 6124 58780 6188 58784
rect 6124 58724 6128 58780
rect 6128 58724 6184 58780
rect 6184 58724 6188 58780
rect 6124 58720 6188 58724
rect 86476 58780 86540 58784
rect 86476 58724 86480 58780
rect 86480 58724 86536 58780
rect 86536 58724 86540 58780
rect 86476 58720 86540 58724
rect 86556 58780 86620 58784
rect 86556 58724 86560 58780
rect 86560 58724 86616 58780
rect 86616 58724 86620 58780
rect 86556 58720 86620 58724
rect 86636 58780 86700 58784
rect 86636 58724 86640 58780
rect 86640 58724 86696 58780
rect 86696 58724 86700 58780
rect 86636 58720 86700 58724
rect 86716 58780 86780 58784
rect 86716 58724 86720 58780
rect 86720 58724 86776 58780
rect 86776 58724 86780 58780
rect 86716 58720 86780 58724
rect 6620 58236 6684 58240
rect 6620 58180 6624 58236
rect 6624 58180 6680 58236
rect 6680 58180 6684 58236
rect 6620 58176 6684 58180
rect 6700 58236 6764 58240
rect 6700 58180 6704 58236
rect 6704 58180 6760 58236
rect 6760 58180 6764 58236
rect 6700 58176 6764 58180
rect 6780 58236 6844 58240
rect 6780 58180 6784 58236
rect 6784 58180 6840 58236
rect 6840 58180 6844 58236
rect 6780 58176 6844 58180
rect 6860 58236 6924 58240
rect 6860 58180 6864 58236
rect 6864 58180 6920 58236
rect 6920 58180 6924 58236
rect 6860 58176 6924 58180
rect 87212 58236 87276 58240
rect 87212 58180 87216 58236
rect 87216 58180 87272 58236
rect 87272 58180 87276 58236
rect 87212 58176 87276 58180
rect 87292 58236 87356 58240
rect 87292 58180 87296 58236
rect 87296 58180 87352 58236
rect 87352 58180 87356 58236
rect 87292 58176 87356 58180
rect 87372 58236 87436 58240
rect 87372 58180 87376 58236
rect 87376 58180 87432 58236
rect 87432 58180 87436 58236
rect 87372 58176 87436 58180
rect 87452 58236 87516 58240
rect 87452 58180 87456 58236
rect 87456 58180 87512 58236
rect 87512 58180 87516 58236
rect 87452 58176 87516 58180
rect 5884 57692 5948 57696
rect 5884 57636 5888 57692
rect 5888 57636 5944 57692
rect 5944 57636 5948 57692
rect 5884 57632 5948 57636
rect 5964 57692 6028 57696
rect 5964 57636 5968 57692
rect 5968 57636 6024 57692
rect 6024 57636 6028 57692
rect 5964 57632 6028 57636
rect 6044 57692 6108 57696
rect 6044 57636 6048 57692
rect 6048 57636 6104 57692
rect 6104 57636 6108 57692
rect 6044 57632 6108 57636
rect 6124 57692 6188 57696
rect 6124 57636 6128 57692
rect 6128 57636 6184 57692
rect 6184 57636 6188 57692
rect 6124 57632 6188 57636
rect 86476 57692 86540 57696
rect 86476 57636 86480 57692
rect 86480 57636 86536 57692
rect 86536 57636 86540 57692
rect 86476 57632 86540 57636
rect 86556 57692 86620 57696
rect 86556 57636 86560 57692
rect 86560 57636 86616 57692
rect 86616 57636 86620 57692
rect 86556 57632 86620 57636
rect 86636 57692 86700 57696
rect 86636 57636 86640 57692
rect 86640 57636 86696 57692
rect 86696 57636 86700 57692
rect 86636 57632 86700 57636
rect 86716 57692 86780 57696
rect 86716 57636 86720 57692
rect 86720 57636 86776 57692
rect 86776 57636 86780 57692
rect 86716 57632 86780 57636
rect 6620 57148 6684 57152
rect 6620 57092 6624 57148
rect 6624 57092 6680 57148
rect 6680 57092 6684 57148
rect 6620 57088 6684 57092
rect 6700 57148 6764 57152
rect 6700 57092 6704 57148
rect 6704 57092 6760 57148
rect 6760 57092 6764 57148
rect 6700 57088 6764 57092
rect 6780 57148 6844 57152
rect 6780 57092 6784 57148
rect 6784 57092 6840 57148
rect 6840 57092 6844 57148
rect 6780 57088 6844 57092
rect 6860 57148 6924 57152
rect 6860 57092 6864 57148
rect 6864 57092 6920 57148
rect 6920 57092 6924 57148
rect 6860 57088 6924 57092
rect 87212 57148 87276 57152
rect 87212 57092 87216 57148
rect 87216 57092 87272 57148
rect 87272 57092 87276 57148
rect 87212 57088 87276 57092
rect 87292 57148 87356 57152
rect 87292 57092 87296 57148
rect 87296 57092 87352 57148
rect 87352 57092 87356 57148
rect 87292 57088 87356 57092
rect 87372 57148 87436 57152
rect 87372 57092 87376 57148
rect 87376 57092 87432 57148
rect 87432 57092 87436 57148
rect 87372 57088 87436 57092
rect 87452 57148 87516 57152
rect 87452 57092 87456 57148
rect 87456 57092 87512 57148
rect 87512 57092 87516 57148
rect 87452 57088 87516 57092
rect 5884 56604 5948 56608
rect 5884 56548 5888 56604
rect 5888 56548 5944 56604
rect 5944 56548 5948 56604
rect 5884 56544 5948 56548
rect 5964 56604 6028 56608
rect 5964 56548 5968 56604
rect 5968 56548 6024 56604
rect 6024 56548 6028 56604
rect 5964 56544 6028 56548
rect 6044 56604 6108 56608
rect 6044 56548 6048 56604
rect 6048 56548 6104 56604
rect 6104 56548 6108 56604
rect 6044 56544 6108 56548
rect 6124 56604 6188 56608
rect 6124 56548 6128 56604
rect 6128 56548 6184 56604
rect 6184 56548 6188 56604
rect 6124 56544 6188 56548
rect 86476 56604 86540 56608
rect 86476 56548 86480 56604
rect 86480 56548 86536 56604
rect 86536 56548 86540 56604
rect 86476 56544 86540 56548
rect 86556 56604 86620 56608
rect 86556 56548 86560 56604
rect 86560 56548 86616 56604
rect 86616 56548 86620 56604
rect 86556 56544 86620 56548
rect 86636 56604 86700 56608
rect 86636 56548 86640 56604
rect 86640 56548 86696 56604
rect 86696 56548 86700 56604
rect 86636 56544 86700 56548
rect 86716 56604 86780 56608
rect 86716 56548 86720 56604
rect 86720 56548 86776 56604
rect 86776 56548 86780 56604
rect 86716 56544 86780 56548
rect 6620 56060 6684 56064
rect 6620 56004 6624 56060
rect 6624 56004 6680 56060
rect 6680 56004 6684 56060
rect 6620 56000 6684 56004
rect 6700 56060 6764 56064
rect 6700 56004 6704 56060
rect 6704 56004 6760 56060
rect 6760 56004 6764 56060
rect 6700 56000 6764 56004
rect 6780 56060 6844 56064
rect 6780 56004 6784 56060
rect 6784 56004 6840 56060
rect 6840 56004 6844 56060
rect 6780 56000 6844 56004
rect 6860 56060 6924 56064
rect 6860 56004 6864 56060
rect 6864 56004 6920 56060
rect 6920 56004 6924 56060
rect 6860 56000 6924 56004
rect 87212 56060 87276 56064
rect 87212 56004 87216 56060
rect 87216 56004 87272 56060
rect 87272 56004 87276 56060
rect 87212 56000 87276 56004
rect 87292 56060 87356 56064
rect 87292 56004 87296 56060
rect 87296 56004 87352 56060
rect 87352 56004 87356 56060
rect 87292 56000 87356 56004
rect 87372 56060 87436 56064
rect 87372 56004 87376 56060
rect 87376 56004 87432 56060
rect 87432 56004 87436 56060
rect 87372 56000 87436 56004
rect 87452 56060 87516 56064
rect 87452 56004 87456 56060
rect 87456 56004 87512 56060
rect 87512 56004 87516 56060
rect 87452 56000 87516 56004
rect 5884 55516 5948 55520
rect 5884 55460 5888 55516
rect 5888 55460 5944 55516
rect 5944 55460 5948 55516
rect 5884 55456 5948 55460
rect 5964 55516 6028 55520
rect 5964 55460 5968 55516
rect 5968 55460 6024 55516
rect 6024 55460 6028 55516
rect 5964 55456 6028 55460
rect 6044 55516 6108 55520
rect 6044 55460 6048 55516
rect 6048 55460 6104 55516
rect 6104 55460 6108 55516
rect 6044 55456 6108 55460
rect 6124 55516 6188 55520
rect 6124 55460 6128 55516
rect 6128 55460 6184 55516
rect 6184 55460 6188 55516
rect 6124 55456 6188 55460
rect 86476 55516 86540 55520
rect 86476 55460 86480 55516
rect 86480 55460 86536 55516
rect 86536 55460 86540 55516
rect 86476 55456 86540 55460
rect 86556 55516 86620 55520
rect 86556 55460 86560 55516
rect 86560 55460 86616 55516
rect 86616 55460 86620 55516
rect 86556 55456 86620 55460
rect 86636 55516 86700 55520
rect 86636 55460 86640 55516
rect 86640 55460 86696 55516
rect 86696 55460 86700 55516
rect 86636 55456 86700 55460
rect 86716 55516 86780 55520
rect 86716 55460 86720 55516
rect 86720 55460 86776 55516
rect 86776 55460 86780 55516
rect 86716 55456 86780 55460
rect 6620 54972 6684 54976
rect 6620 54916 6624 54972
rect 6624 54916 6680 54972
rect 6680 54916 6684 54972
rect 6620 54912 6684 54916
rect 6700 54972 6764 54976
rect 6700 54916 6704 54972
rect 6704 54916 6760 54972
rect 6760 54916 6764 54972
rect 6700 54912 6764 54916
rect 6780 54972 6844 54976
rect 6780 54916 6784 54972
rect 6784 54916 6840 54972
rect 6840 54916 6844 54972
rect 6780 54912 6844 54916
rect 6860 54972 6924 54976
rect 6860 54916 6864 54972
rect 6864 54916 6920 54972
rect 6920 54916 6924 54972
rect 6860 54912 6924 54916
rect 87212 54972 87276 54976
rect 87212 54916 87216 54972
rect 87216 54916 87272 54972
rect 87272 54916 87276 54972
rect 87212 54912 87276 54916
rect 87292 54972 87356 54976
rect 87292 54916 87296 54972
rect 87296 54916 87352 54972
rect 87352 54916 87356 54972
rect 87292 54912 87356 54916
rect 87372 54972 87436 54976
rect 87372 54916 87376 54972
rect 87376 54916 87432 54972
rect 87432 54916 87436 54972
rect 87372 54912 87436 54916
rect 87452 54972 87516 54976
rect 87452 54916 87456 54972
rect 87456 54916 87512 54972
rect 87512 54916 87516 54972
rect 87452 54912 87516 54916
rect 5884 54428 5948 54432
rect 5884 54372 5888 54428
rect 5888 54372 5944 54428
rect 5944 54372 5948 54428
rect 5884 54368 5948 54372
rect 5964 54428 6028 54432
rect 5964 54372 5968 54428
rect 5968 54372 6024 54428
rect 6024 54372 6028 54428
rect 5964 54368 6028 54372
rect 6044 54428 6108 54432
rect 6044 54372 6048 54428
rect 6048 54372 6104 54428
rect 6104 54372 6108 54428
rect 6044 54368 6108 54372
rect 6124 54428 6188 54432
rect 6124 54372 6128 54428
rect 6128 54372 6184 54428
rect 6184 54372 6188 54428
rect 6124 54368 6188 54372
rect 86476 54428 86540 54432
rect 86476 54372 86480 54428
rect 86480 54372 86536 54428
rect 86536 54372 86540 54428
rect 86476 54368 86540 54372
rect 86556 54428 86620 54432
rect 86556 54372 86560 54428
rect 86560 54372 86616 54428
rect 86616 54372 86620 54428
rect 86556 54368 86620 54372
rect 86636 54428 86700 54432
rect 86636 54372 86640 54428
rect 86640 54372 86696 54428
rect 86696 54372 86700 54428
rect 86636 54368 86700 54372
rect 86716 54428 86780 54432
rect 86716 54372 86720 54428
rect 86720 54372 86776 54428
rect 86776 54372 86780 54428
rect 86716 54368 86780 54372
rect 6620 53884 6684 53888
rect 6620 53828 6624 53884
rect 6624 53828 6680 53884
rect 6680 53828 6684 53884
rect 6620 53824 6684 53828
rect 6700 53884 6764 53888
rect 6700 53828 6704 53884
rect 6704 53828 6760 53884
rect 6760 53828 6764 53884
rect 6700 53824 6764 53828
rect 6780 53884 6844 53888
rect 6780 53828 6784 53884
rect 6784 53828 6840 53884
rect 6840 53828 6844 53884
rect 6780 53824 6844 53828
rect 6860 53884 6924 53888
rect 6860 53828 6864 53884
rect 6864 53828 6920 53884
rect 6920 53828 6924 53884
rect 6860 53824 6924 53828
rect 87212 53884 87276 53888
rect 87212 53828 87216 53884
rect 87216 53828 87272 53884
rect 87272 53828 87276 53884
rect 87212 53824 87276 53828
rect 87292 53884 87356 53888
rect 87292 53828 87296 53884
rect 87296 53828 87352 53884
rect 87352 53828 87356 53884
rect 87292 53824 87356 53828
rect 87372 53884 87436 53888
rect 87372 53828 87376 53884
rect 87376 53828 87432 53884
rect 87432 53828 87436 53884
rect 87372 53824 87436 53828
rect 87452 53884 87516 53888
rect 87452 53828 87456 53884
rect 87456 53828 87512 53884
rect 87512 53828 87516 53884
rect 87452 53824 87516 53828
rect 5884 53340 5948 53344
rect 5884 53284 5888 53340
rect 5888 53284 5944 53340
rect 5944 53284 5948 53340
rect 5884 53280 5948 53284
rect 5964 53340 6028 53344
rect 5964 53284 5968 53340
rect 5968 53284 6024 53340
rect 6024 53284 6028 53340
rect 5964 53280 6028 53284
rect 6044 53340 6108 53344
rect 6044 53284 6048 53340
rect 6048 53284 6104 53340
rect 6104 53284 6108 53340
rect 6044 53280 6108 53284
rect 6124 53340 6188 53344
rect 6124 53284 6128 53340
rect 6128 53284 6184 53340
rect 6184 53284 6188 53340
rect 6124 53280 6188 53284
rect 86476 53340 86540 53344
rect 86476 53284 86480 53340
rect 86480 53284 86536 53340
rect 86536 53284 86540 53340
rect 86476 53280 86540 53284
rect 86556 53340 86620 53344
rect 86556 53284 86560 53340
rect 86560 53284 86616 53340
rect 86616 53284 86620 53340
rect 86556 53280 86620 53284
rect 86636 53340 86700 53344
rect 86636 53284 86640 53340
rect 86640 53284 86696 53340
rect 86696 53284 86700 53340
rect 86636 53280 86700 53284
rect 86716 53340 86780 53344
rect 86716 53284 86720 53340
rect 86720 53284 86776 53340
rect 86776 53284 86780 53340
rect 86716 53280 86780 53284
rect 6620 52796 6684 52800
rect 6620 52740 6624 52796
rect 6624 52740 6680 52796
rect 6680 52740 6684 52796
rect 6620 52736 6684 52740
rect 6700 52796 6764 52800
rect 6700 52740 6704 52796
rect 6704 52740 6760 52796
rect 6760 52740 6764 52796
rect 6700 52736 6764 52740
rect 6780 52796 6844 52800
rect 6780 52740 6784 52796
rect 6784 52740 6840 52796
rect 6840 52740 6844 52796
rect 6780 52736 6844 52740
rect 6860 52796 6924 52800
rect 6860 52740 6864 52796
rect 6864 52740 6920 52796
rect 6920 52740 6924 52796
rect 6860 52736 6924 52740
rect 87212 52796 87276 52800
rect 87212 52740 87216 52796
rect 87216 52740 87272 52796
rect 87272 52740 87276 52796
rect 87212 52736 87276 52740
rect 87292 52796 87356 52800
rect 87292 52740 87296 52796
rect 87296 52740 87352 52796
rect 87352 52740 87356 52796
rect 87292 52736 87356 52740
rect 87372 52796 87436 52800
rect 87372 52740 87376 52796
rect 87376 52740 87432 52796
rect 87432 52740 87436 52796
rect 87372 52736 87436 52740
rect 87452 52796 87516 52800
rect 87452 52740 87456 52796
rect 87456 52740 87512 52796
rect 87512 52740 87516 52796
rect 87452 52736 87516 52740
rect 5884 52252 5948 52256
rect 5884 52196 5888 52252
rect 5888 52196 5944 52252
rect 5944 52196 5948 52252
rect 5884 52192 5948 52196
rect 5964 52252 6028 52256
rect 5964 52196 5968 52252
rect 5968 52196 6024 52252
rect 6024 52196 6028 52252
rect 5964 52192 6028 52196
rect 6044 52252 6108 52256
rect 6044 52196 6048 52252
rect 6048 52196 6104 52252
rect 6104 52196 6108 52252
rect 6044 52192 6108 52196
rect 6124 52252 6188 52256
rect 6124 52196 6128 52252
rect 6128 52196 6184 52252
rect 6184 52196 6188 52252
rect 6124 52192 6188 52196
rect 86476 52252 86540 52256
rect 86476 52196 86480 52252
rect 86480 52196 86536 52252
rect 86536 52196 86540 52252
rect 86476 52192 86540 52196
rect 86556 52252 86620 52256
rect 86556 52196 86560 52252
rect 86560 52196 86616 52252
rect 86616 52196 86620 52252
rect 86556 52192 86620 52196
rect 86636 52252 86700 52256
rect 86636 52196 86640 52252
rect 86640 52196 86696 52252
rect 86696 52196 86700 52252
rect 86636 52192 86700 52196
rect 86716 52252 86780 52256
rect 86716 52196 86720 52252
rect 86720 52196 86776 52252
rect 86776 52196 86780 52252
rect 86716 52192 86780 52196
rect 6620 51708 6684 51712
rect 6620 51652 6624 51708
rect 6624 51652 6680 51708
rect 6680 51652 6684 51708
rect 6620 51648 6684 51652
rect 6700 51708 6764 51712
rect 6700 51652 6704 51708
rect 6704 51652 6760 51708
rect 6760 51652 6764 51708
rect 6700 51648 6764 51652
rect 6780 51708 6844 51712
rect 6780 51652 6784 51708
rect 6784 51652 6840 51708
rect 6840 51652 6844 51708
rect 6780 51648 6844 51652
rect 6860 51708 6924 51712
rect 6860 51652 6864 51708
rect 6864 51652 6920 51708
rect 6920 51652 6924 51708
rect 6860 51648 6924 51652
rect 87212 51708 87276 51712
rect 87212 51652 87216 51708
rect 87216 51652 87272 51708
rect 87272 51652 87276 51708
rect 87212 51648 87276 51652
rect 87292 51708 87356 51712
rect 87292 51652 87296 51708
rect 87296 51652 87352 51708
rect 87352 51652 87356 51708
rect 87292 51648 87356 51652
rect 87372 51708 87436 51712
rect 87372 51652 87376 51708
rect 87376 51652 87432 51708
rect 87432 51652 87436 51708
rect 87372 51648 87436 51652
rect 87452 51708 87516 51712
rect 87452 51652 87456 51708
rect 87456 51652 87512 51708
rect 87512 51652 87516 51708
rect 87452 51648 87516 51652
rect 5884 51164 5948 51168
rect 5884 51108 5888 51164
rect 5888 51108 5944 51164
rect 5944 51108 5948 51164
rect 5884 51104 5948 51108
rect 5964 51164 6028 51168
rect 5964 51108 5968 51164
rect 5968 51108 6024 51164
rect 6024 51108 6028 51164
rect 5964 51104 6028 51108
rect 6044 51164 6108 51168
rect 6044 51108 6048 51164
rect 6048 51108 6104 51164
rect 6104 51108 6108 51164
rect 6044 51104 6108 51108
rect 6124 51164 6188 51168
rect 6124 51108 6128 51164
rect 6128 51108 6184 51164
rect 6184 51108 6188 51164
rect 6124 51104 6188 51108
rect 86476 51164 86540 51168
rect 86476 51108 86480 51164
rect 86480 51108 86536 51164
rect 86536 51108 86540 51164
rect 86476 51104 86540 51108
rect 86556 51164 86620 51168
rect 86556 51108 86560 51164
rect 86560 51108 86616 51164
rect 86616 51108 86620 51164
rect 86556 51104 86620 51108
rect 86636 51164 86700 51168
rect 86636 51108 86640 51164
rect 86640 51108 86696 51164
rect 86696 51108 86700 51164
rect 86636 51104 86700 51108
rect 86716 51164 86780 51168
rect 86716 51108 86720 51164
rect 86720 51108 86776 51164
rect 86776 51108 86780 51164
rect 86716 51104 86780 51108
rect 6620 50620 6684 50624
rect 6620 50564 6624 50620
rect 6624 50564 6680 50620
rect 6680 50564 6684 50620
rect 6620 50560 6684 50564
rect 6700 50620 6764 50624
rect 6700 50564 6704 50620
rect 6704 50564 6760 50620
rect 6760 50564 6764 50620
rect 6700 50560 6764 50564
rect 6780 50620 6844 50624
rect 6780 50564 6784 50620
rect 6784 50564 6840 50620
rect 6840 50564 6844 50620
rect 6780 50560 6844 50564
rect 6860 50620 6924 50624
rect 6860 50564 6864 50620
rect 6864 50564 6920 50620
rect 6920 50564 6924 50620
rect 6860 50560 6924 50564
rect 87212 50620 87276 50624
rect 87212 50564 87216 50620
rect 87216 50564 87272 50620
rect 87272 50564 87276 50620
rect 87212 50560 87276 50564
rect 87292 50620 87356 50624
rect 87292 50564 87296 50620
rect 87296 50564 87352 50620
rect 87352 50564 87356 50620
rect 87292 50560 87356 50564
rect 87372 50620 87436 50624
rect 87372 50564 87376 50620
rect 87376 50564 87432 50620
rect 87432 50564 87436 50620
rect 87372 50560 87436 50564
rect 87452 50620 87516 50624
rect 87452 50564 87456 50620
rect 87456 50564 87512 50620
rect 87512 50564 87516 50620
rect 87452 50560 87516 50564
rect 5884 50076 5948 50080
rect 5884 50020 5888 50076
rect 5888 50020 5944 50076
rect 5944 50020 5948 50076
rect 5884 50016 5948 50020
rect 5964 50076 6028 50080
rect 5964 50020 5968 50076
rect 5968 50020 6024 50076
rect 6024 50020 6028 50076
rect 5964 50016 6028 50020
rect 6044 50076 6108 50080
rect 6044 50020 6048 50076
rect 6048 50020 6104 50076
rect 6104 50020 6108 50076
rect 6044 50016 6108 50020
rect 6124 50076 6188 50080
rect 6124 50020 6128 50076
rect 6128 50020 6184 50076
rect 6184 50020 6188 50076
rect 6124 50016 6188 50020
rect 86476 50076 86540 50080
rect 86476 50020 86480 50076
rect 86480 50020 86536 50076
rect 86536 50020 86540 50076
rect 86476 50016 86540 50020
rect 86556 50076 86620 50080
rect 86556 50020 86560 50076
rect 86560 50020 86616 50076
rect 86616 50020 86620 50076
rect 86556 50016 86620 50020
rect 86636 50076 86700 50080
rect 86636 50020 86640 50076
rect 86640 50020 86696 50076
rect 86696 50020 86700 50076
rect 86636 50016 86700 50020
rect 86716 50076 86780 50080
rect 86716 50020 86720 50076
rect 86720 50020 86776 50076
rect 86776 50020 86780 50076
rect 86716 50016 86780 50020
rect 6620 49532 6684 49536
rect 6620 49476 6624 49532
rect 6624 49476 6680 49532
rect 6680 49476 6684 49532
rect 6620 49472 6684 49476
rect 6700 49532 6764 49536
rect 6700 49476 6704 49532
rect 6704 49476 6760 49532
rect 6760 49476 6764 49532
rect 6700 49472 6764 49476
rect 6780 49532 6844 49536
rect 6780 49476 6784 49532
rect 6784 49476 6840 49532
rect 6840 49476 6844 49532
rect 6780 49472 6844 49476
rect 6860 49532 6924 49536
rect 6860 49476 6864 49532
rect 6864 49476 6920 49532
rect 6920 49476 6924 49532
rect 6860 49472 6924 49476
rect 87212 49532 87276 49536
rect 87212 49476 87216 49532
rect 87216 49476 87272 49532
rect 87272 49476 87276 49532
rect 87212 49472 87276 49476
rect 87292 49532 87356 49536
rect 87292 49476 87296 49532
rect 87296 49476 87352 49532
rect 87352 49476 87356 49532
rect 87292 49472 87356 49476
rect 87372 49532 87436 49536
rect 87372 49476 87376 49532
rect 87376 49476 87432 49532
rect 87432 49476 87436 49532
rect 87372 49472 87436 49476
rect 87452 49532 87516 49536
rect 87452 49476 87456 49532
rect 87456 49476 87512 49532
rect 87512 49476 87516 49532
rect 87452 49472 87516 49476
rect 5884 48988 5948 48992
rect 5884 48932 5888 48988
rect 5888 48932 5944 48988
rect 5944 48932 5948 48988
rect 5884 48928 5948 48932
rect 5964 48988 6028 48992
rect 5964 48932 5968 48988
rect 5968 48932 6024 48988
rect 6024 48932 6028 48988
rect 5964 48928 6028 48932
rect 6044 48988 6108 48992
rect 6044 48932 6048 48988
rect 6048 48932 6104 48988
rect 6104 48932 6108 48988
rect 6044 48928 6108 48932
rect 6124 48988 6188 48992
rect 6124 48932 6128 48988
rect 6128 48932 6184 48988
rect 6184 48932 6188 48988
rect 6124 48928 6188 48932
rect 86476 48988 86540 48992
rect 86476 48932 86480 48988
rect 86480 48932 86536 48988
rect 86536 48932 86540 48988
rect 86476 48928 86540 48932
rect 86556 48988 86620 48992
rect 86556 48932 86560 48988
rect 86560 48932 86616 48988
rect 86616 48932 86620 48988
rect 86556 48928 86620 48932
rect 86636 48988 86700 48992
rect 86636 48932 86640 48988
rect 86640 48932 86696 48988
rect 86696 48932 86700 48988
rect 86636 48928 86700 48932
rect 86716 48988 86780 48992
rect 86716 48932 86720 48988
rect 86720 48932 86776 48988
rect 86776 48932 86780 48988
rect 86716 48928 86780 48932
rect 6620 48444 6684 48448
rect 6620 48388 6624 48444
rect 6624 48388 6680 48444
rect 6680 48388 6684 48444
rect 6620 48384 6684 48388
rect 6700 48444 6764 48448
rect 6700 48388 6704 48444
rect 6704 48388 6760 48444
rect 6760 48388 6764 48444
rect 6700 48384 6764 48388
rect 6780 48444 6844 48448
rect 6780 48388 6784 48444
rect 6784 48388 6840 48444
rect 6840 48388 6844 48444
rect 6780 48384 6844 48388
rect 6860 48444 6924 48448
rect 6860 48388 6864 48444
rect 6864 48388 6920 48444
rect 6920 48388 6924 48444
rect 6860 48384 6924 48388
rect 87212 48444 87276 48448
rect 87212 48388 87216 48444
rect 87216 48388 87272 48444
rect 87272 48388 87276 48444
rect 87212 48384 87276 48388
rect 87292 48444 87356 48448
rect 87292 48388 87296 48444
rect 87296 48388 87352 48444
rect 87352 48388 87356 48444
rect 87292 48384 87356 48388
rect 87372 48444 87436 48448
rect 87372 48388 87376 48444
rect 87376 48388 87432 48444
rect 87432 48388 87436 48444
rect 87372 48384 87436 48388
rect 87452 48444 87516 48448
rect 87452 48388 87456 48444
rect 87456 48388 87512 48444
rect 87512 48388 87516 48444
rect 87452 48384 87516 48388
rect 5884 47900 5948 47904
rect 5884 47844 5888 47900
rect 5888 47844 5944 47900
rect 5944 47844 5948 47900
rect 5884 47840 5948 47844
rect 5964 47900 6028 47904
rect 5964 47844 5968 47900
rect 5968 47844 6024 47900
rect 6024 47844 6028 47900
rect 5964 47840 6028 47844
rect 6044 47900 6108 47904
rect 6044 47844 6048 47900
rect 6048 47844 6104 47900
rect 6104 47844 6108 47900
rect 6044 47840 6108 47844
rect 6124 47900 6188 47904
rect 6124 47844 6128 47900
rect 6128 47844 6184 47900
rect 6184 47844 6188 47900
rect 6124 47840 6188 47844
rect 86476 47900 86540 47904
rect 86476 47844 86480 47900
rect 86480 47844 86536 47900
rect 86536 47844 86540 47900
rect 86476 47840 86540 47844
rect 86556 47900 86620 47904
rect 86556 47844 86560 47900
rect 86560 47844 86616 47900
rect 86616 47844 86620 47900
rect 86556 47840 86620 47844
rect 86636 47900 86700 47904
rect 86636 47844 86640 47900
rect 86640 47844 86696 47900
rect 86696 47844 86700 47900
rect 86636 47840 86700 47844
rect 86716 47900 86780 47904
rect 86716 47844 86720 47900
rect 86720 47844 86776 47900
rect 86776 47844 86780 47900
rect 86716 47840 86780 47844
rect 6620 47356 6684 47360
rect 6620 47300 6624 47356
rect 6624 47300 6680 47356
rect 6680 47300 6684 47356
rect 6620 47296 6684 47300
rect 6700 47356 6764 47360
rect 6700 47300 6704 47356
rect 6704 47300 6760 47356
rect 6760 47300 6764 47356
rect 6700 47296 6764 47300
rect 6780 47356 6844 47360
rect 6780 47300 6784 47356
rect 6784 47300 6840 47356
rect 6840 47300 6844 47356
rect 6780 47296 6844 47300
rect 6860 47356 6924 47360
rect 6860 47300 6864 47356
rect 6864 47300 6920 47356
rect 6920 47300 6924 47356
rect 6860 47296 6924 47300
rect 87212 47356 87276 47360
rect 87212 47300 87216 47356
rect 87216 47300 87272 47356
rect 87272 47300 87276 47356
rect 87212 47296 87276 47300
rect 87292 47356 87356 47360
rect 87292 47300 87296 47356
rect 87296 47300 87352 47356
rect 87352 47300 87356 47356
rect 87292 47296 87356 47300
rect 87372 47356 87436 47360
rect 87372 47300 87376 47356
rect 87376 47300 87432 47356
rect 87432 47300 87436 47356
rect 87372 47296 87436 47300
rect 87452 47356 87516 47360
rect 87452 47300 87456 47356
rect 87456 47300 87512 47356
rect 87512 47300 87516 47356
rect 87452 47296 87516 47300
rect 5884 46812 5948 46816
rect 5884 46756 5888 46812
rect 5888 46756 5944 46812
rect 5944 46756 5948 46812
rect 5884 46752 5948 46756
rect 5964 46812 6028 46816
rect 5964 46756 5968 46812
rect 5968 46756 6024 46812
rect 6024 46756 6028 46812
rect 5964 46752 6028 46756
rect 6044 46812 6108 46816
rect 6044 46756 6048 46812
rect 6048 46756 6104 46812
rect 6104 46756 6108 46812
rect 6044 46752 6108 46756
rect 6124 46812 6188 46816
rect 6124 46756 6128 46812
rect 6128 46756 6184 46812
rect 6184 46756 6188 46812
rect 6124 46752 6188 46756
rect 86476 46812 86540 46816
rect 86476 46756 86480 46812
rect 86480 46756 86536 46812
rect 86536 46756 86540 46812
rect 86476 46752 86540 46756
rect 86556 46812 86620 46816
rect 86556 46756 86560 46812
rect 86560 46756 86616 46812
rect 86616 46756 86620 46812
rect 86556 46752 86620 46756
rect 86636 46812 86700 46816
rect 86636 46756 86640 46812
rect 86640 46756 86696 46812
rect 86696 46756 86700 46812
rect 86636 46752 86700 46756
rect 86716 46812 86780 46816
rect 86716 46756 86720 46812
rect 86720 46756 86776 46812
rect 86776 46756 86780 46812
rect 86716 46752 86780 46756
rect 6620 46268 6684 46272
rect 6620 46212 6624 46268
rect 6624 46212 6680 46268
rect 6680 46212 6684 46268
rect 6620 46208 6684 46212
rect 6700 46268 6764 46272
rect 6700 46212 6704 46268
rect 6704 46212 6760 46268
rect 6760 46212 6764 46268
rect 6700 46208 6764 46212
rect 6780 46268 6844 46272
rect 6780 46212 6784 46268
rect 6784 46212 6840 46268
rect 6840 46212 6844 46268
rect 6780 46208 6844 46212
rect 6860 46268 6924 46272
rect 6860 46212 6864 46268
rect 6864 46212 6920 46268
rect 6920 46212 6924 46268
rect 6860 46208 6924 46212
rect 87212 46268 87276 46272
rect 87212 46212 87216 46268
rect 87216 46212 87272 46268
rect 87272 46212 87276 46268
rect 87212 46208 87276 46212
rect 87292 46268 87356 46272
rect 87292 46212 87296 46268
rect 87296 46212 87352 46268
rect 87352 46212 87356 46268
rect 87292 46208 87356 46212
rect 87372 46268 87436 46272
rect 87372 46212 87376 46268
rect 87376 46212 87432 46268
rect 87432 46212 87436 46268
rect 87372 46208 87436 46212
rect 87452 46268 87516 46272
rect 87452 46212 87456 46268
rect 87456 46212 87512 46268
rect 87512 46212 87516 46268
rect 87452 46208 87516 46212
rect 11708 45740 11772 45804
rect 5884 45724 5948 45728
rect 5884 45668 5888 45724
rect 5888 45668 5944 45724
rect 5944 45668 5948 45724
rect 5884 45664 5948 45668
rect 5964 45724 6028 45728
rect 5964 45668 5968 45724
rect 5968 45668 6024 45724
rect 6024 45668 6028 45724
rect 5964 45664 6028 45668
rect 6044 45724 6108 45728
rect 6044 45668 6048 45724
rect 6048 45668 6104 45724
rect 6104 45668 6108 45724
rect 6044 45664 6108 45668
rect 6124 45724 6188 45728
rect 6124 45668 6128 45724
rect 6128 45668 6184 45724
rect 6184 45668 6188 45724
rect 6124 45664 6188 45668
rect 11708 45196 11772 45260
rect 6620 45180 6684 45184
rect 6620 45124 6624 45180
rect 6624 45124 6680 45180
rect 6680 45124 6684 45180
rect 6620 45120 6684 45124
rect 6700 45180 6764 45184
rect 6700 45124 6704 45180
rect 6704 45124 6760 45180
rect 6760 45124 6764 45180
rect 6700 45120 6764 45124
rect 6780 45180 6844 45184
rect 6780 45124 6784 45180
rect 6784 45124 6840 45180
rect 6840 45124 6844 45180
rect 6780 45120 6844 45124
rect 6860 45180 6924 45184
rect 6860 45124 6864 45180
rect 6864 45124 6920 45180
rect 6920 45124 6924 45180
rect 6860 45120 6924 45124
rect 86476 45724 86540 45728
rect 86476 45668 86480 45724
rect 86480 45668 86536 45724
rect 86536 45668 86540 45724
rect 86476 45664 86540 45668
rect 86556 45724 86620 45728
rect 86556 45668 86560 45724
rect 86560 45668 86616 45724
rect 86616 45668 86620 45724
rect 86556 45664 86620 45668
rect 86636 45724 86700 45728
rect 86636 45668 86640 45724
rect 86640 45668 86696 45724
rect 86696 45668 86700 45724
rect 86636 45664 86700 45668
rect 86716 45724 86780 45728
rect 86716 45668 86720 45724
rect 86720 45668 86776 45724
rect 86776 45668 86780 45724
rect 86716 45664 86780 45668
rect 87212 45180 87276 45184
rect 87212 45124 87216 45180
rect 87216 45124 87272 45180
rect 87272 45124 87276 45180
rect 87212 45120 87276 45124
rect 87292 45180 87356 45184
rect 87292 45124 87296 45180
rect 87296 45124 87352 45180
rect 87352 45124 87356 45180
rect 87292 45120 87356 45124
rect 87372 45180 87436 45184
rect 87372 45124 87376 45180
rect 87376 45124 87432 45180
rect 87432 45124 87436 45180
rect 87372 45120 87436 45124
rect 87452 45180 87516 45184
rect 87452 45124 87456 45180
rect 87456 45124 87512 45180
rect 87512 45124 87516 45180
rect 87452 45120 87516 45124
rect 5884 44636 5948 44640
rect 5884 44580 5888 44636
rect 5888 44580 5944 44636
rect 5944 44580 5948 44636
rect 5884 44576 5948 44580
rect 5964 44636 6028 44640
rect 5964 44580 5968 44636
rect 5968 44580 6024 44636
rect 6024 44580 6028 44636
rect 5964 44576 6028 44580
rect 6044 44636 6108 44640
rect 6044 44580 6048 44636
rect 6048 44580 6104 44636
rect 6104 44580 6108 44636
rect 6044 44576 6108 44580
rect 6124 44636 6188 44640
rect 6124 44580 6128 44636
rect 6128 44580 6184 44636
rect 6184 44580 6188 44636
rect 6124 44576 6188 44580
rect 86476 44636 86540 44640
rect 86476 44580 86480 44636
rect 86480 44580 86536 44636
rect 86536 44580 86540 44636
rect 86476 44576 86540 44580
rect 86556 44636 86620 44640
rect 86556 44580 86560 44636
rect 86560 44580 86616 44636
rect 86616 44580 86620 44636
rect 86556 44576 86620 44580
rect 86636 44636 86700 44640
rect 86636 44580 86640 44636
rect 86640 44580 86696 44636
rect 86696 44580 86700 44636
rect 86636 44576 86700 44580
rect 86716 44636 86780 44640
rect 86716 44580 86720 44636
rect 86720 44580 86776 44636
rect 86776 44580 86780 44636
rect 86716 44576 86780 44580
rect 6620 44092 6684 44096
rect 6620 44036 6624 44092
rect 6624 44036 6680 44092
rect 6680 44036 6684 44092
rect 6620 44032 6684 44036
rect 6700 44092 6764 44096
rect 6700 44036 6704 44092
rect 6704 44036 6760 44092
rect 6760 44036 6764 44092
rect 6700 44032 6764 44036
rect 6780 44092 6844 44096
rect 6780 44036 6784 44092
rect 6784 44036 6840 44092
rect 6840 44036 6844 44092
rect 6780 44032 6844 44036
rect 6860 44092 6924 44096
rect 6860 44036 6864 44092
rect 6864 44036 6920 44092
rect 6920 44036 6924 44092
rect 6860 44032 6924 44036
rect 87212 44092 87276 44096
rect 87212 44036 87216 44092
rect 87216 44036 87272 44092
rect 87272 44036 87276 44092
rect 87212 44032 87276 44036
rect 87292 44092 87356 44096
rect 87292 44036 87296 44092
rect 87296 44036 87352 44092
rect 87352 44036 87356 44092
rect 87292 44032 87356 44036
rect 87372 44092 87436 44096
rect 87372 44036 87376 44092
rect 87376 44036 87432 44092
rect 87432 44036 87436 44092
rect 87372 44032 87436 44036
rect 87452 44092 87516 44096
rect 87452 44036 87456 44092
rect 87456 44036 87512 44092
rect 87512 44036 87516 44092
rect 87452 44032 87516 44036
rect 5884 43548 5948 43552
rect 5884 43492 5888 43548
rect 5888 43492 5944 43548
rect 5944 43492 5948 43548
rect 5884 43488 5948 43492
rect 5964 43548 6028 43552
rect 5964 43492 5968 43548
rect 5968 43492 6024 43548
rect 6024 43492 6028 43548
rect 5964 43488 6028 43492
rect 6044 43548 6108 43552
rect 6044 43492 6048 43548
rect 6048 43492 6104 43548
rect 6104 43492 6108 43548
rect 6044 43488 6108 43492
rect 6124 43548 6188 43552
rect 6124 43492 6128 43548
rect 6128 43492 6184 43548
rect 6184 43492 6188 43548
rect 6124 43488 6188 43492
rect 86476 43548 86540 43552
rect 86476 43492 86480 43548
rect 86480 43492 86536 43548
rect 86536 43492 86540 43548
rect 86476 43488 86540 43492
rect 86556 43548 86620 43552
rect 86556 43492 86560 43548
rect 86560 43492 86616 43548
rect 86616 43492 86620 43548
rect 86556 43488 86620 43492
rect 86636 43548 86700 43552
rect 86636 43492 86640 43548
rect 86640 43492 86696 43548
rect 86696 43492 86700 43548
rect 86636 43488 86700 43492
rect 86716 43548 86780 43552
rect 86716 43492 86720 43548
rect 86720 43492 86776 43548
rect 86776 43492 86780 43548
rect 86716 43488 86780 43492
rect 6620 43004 6684 43008
rect 6620 42948 6624 43004
rect 6624 42948 6680 43004
rect 6680 42948 6684 43004
rect 6620 42944 6684 42948
rect 6700 43004 6764 43008
rect 6700 42948 6704 43004
rect 6704 42948 6760 43004
rect 6760 42948 6764 43004
rect 6700 42944 6764 42948
rect 6780 43004 6844 43008
rect 6780 42948 6784 43004
rect 6784 42948 6840 43004
rect 6840 42948 6844 43004
rect 6780 42944 6844 42948
rect 6860 43004 6924 43008
rect 6860 42948 6864 43004
rect 6864 42948 6920 43004
rect 6920 42948 6924 43004
rect 6860 42944 6924 42948
rect 87212 43004 87276 43008
rect 87212 42948 87216 43004
rect 87216 42948 87272 43004
rect 87272 42948 87276 43004
rect 87212 42944 87276 42948
rect 87292 43004 87356 43008
rect 87292 42948 87296 43004
rect 87296 42948 87352 43004
rect 87352 42948 87356 43004
rect 87292 42944 87356 42948
rect 87372 43004 87436 43008
rect 87372 42948 87376 43004
rect 87376 42948 87432 43004
rect 87432 42948 87436 43004
rect 87372 42944 87436 42948
rect 87452 43004 87516 43008
rect 87452 42948 87456 43004
rect 87456 42948 87512 43004
rect 87512 42948 87516 43004
rect 87452 42944 87516 42948
rect 5884 42460 5948 42464
rect 5884 42404 5888 42460
rect 5888 42404 5944 42460
rect 5944 42404 5948 42460
rect 5884 42400 5948 42404
rect 5964 42460 6028 42464
rect 5964 42404 5968 42460
rect 5968 42404 6024 42460
rect 6024 42404 6028 42460
rect 5964 42400 6028 42404
rect 6044 42460 6108 42464
rect 6044 42404 6048 42460
rect 6048 42404 6104 42460
rect 6104 42404 6108 42460
rect 6044 42400 6108 42404
rect 6124 42460 6188 42464
rect 6124 42404 6128 42460
rect 6128 42404 6184 42460
rect 6184 42404 6188 42460
rect 6124 42400 6188 42404
rect 86476 42460 86540 42464
rect 86476 42404 86480 42460
rect 86480 42404 86536 42460
rect 86536 42404 86540 42460
rect 86476 42400 86540 42404
rect 86556 42460 86620 42464
rect 86556 42404 86560 42460
rect 86560 42404 86616 42460
rect 86616 42404 86620 42460
rect 86556 42400 86620 42404
rect 86636 42460 86700 42464
rect 86636 42404 86640 42460
rect 86640 42404 86696 42460
rect 86696 42404 86700 42460
rect 86636 42400 86700 42404
rect 86716 42460 86780 42464
rect 86716 42404 86720 42460
rect 86720 42404 86776 42460
rect 86776 42404 86780 42460
rect 86716 42400 86780 42404
rect 6620 41916 6684 41920
rect 6620 41860 6624 41916
rect 6624 41860 6680 41916
rect 6680 41860 6684 41916
rect 6620 41856 6684 41860
rect 6700 41916 6764 41920
rect 6700 41860 6704 41916
rect 6704 41860 6760 41916
rect 6760 41860 6764 41916
rect 6700 41856 6764 41860
rect 6780 41916 6844 41920
rect 6780 41860 6784 41916
rect 6784 41860 6840 41916
rect 6840 41860 6844 41916
rect 6780 41856 6844 41860
rect 6860 41916 6924 41920
rect 6860 41860 6864 41916
rect 6864 41860 6920 41916
rect 6920 41860 6924 41916
rect 6860 41856 6924 41860
rect 87212 41916 87276 41920
rect 87212 41860 87216 41916
rect 87216 41860 87272 41916
rect 87272 41860 87276 41916
rect 87212 41856 87276 41860
rect 87292 41916 87356 41920
rect 87292 41860 87296 41916
rect 87296 41860 87352 41916
rect 87352 41860 87356 41916
rect 87292 41856 87356 41860
rect 87372 41916 87436 41920
rect 87372 41860 87376 41916
rect 87376 41860 87432 41916
rect 87432 41860 87436 41916
rect 87372 41856 87436 41860
rect 87452 41916 87516 41920
rect 87452 41860 87456 41916
rect 87456 41860 87512 41916
rect 87512 41860 87516 41916
rect 87452 41856 87516 41860
rect 5884 41372 5948 41376
rect 5884 41316 5888 41372
rect 5888 41316 5944 41372
rect 5944 41316 5948 41372
rect 5884 41312 5948 41316
rect 5964 41372 6028 41376
rect 5964 41316 5968 41372
rect 5968 41316 6024 41372
rect 6024 41316 6028 41372
rect 5964 41312 6028 41316
rect 6044 41372 6108 41376
rect 6044 41316 6048 41372
rect 6048 41316 6104 41372
rect 6104 41316 6108 41372
rect 6044 41312 6108 41316
rect 6124 41372 6188 41376
rect 6124 41316 6128 41372
rect 6128 41316 6184 41372
rect 6184 41316 6188 41372
rect 6124 41312 6188 41316
rect 86476 41372 86540 41376
rect 86476 41316 86480 41372
rect 86480 41316 86536 41372
rect 86536 41316 86540 41372
rect 86476 41312 86540 41316
rect 86556 41372 86620 41376
rect 86556 41316 86560 41372
rect 86560 41316 86616 41372
rect 86616 41316 86620 41372
rect 86556 41312 86620 41316
rect 86636 41372 86700 41376
rect 86636 41316 86640 41372
rect 86640 41316 86696 41372
rect 86696 41316 86700 41372
rect 86636 41312 86700 41316
rect 86716 41372 86780 41376
rect 86716 41316 86720 41372
rect 86720 41316 86776 41372
rect 86776 41316 86780 41372
rect 86716 41312 86780 41316
rect 6620 40828 6684 40832
rect 6620 40772 6624 40828
rect 6624 40772 6680 40828
rect 6680 40772 6684 40828
rect 6620 40768 6684 40772
rect 6700 40828 6764 40832
rect 6700 40772 6704 40828
rect 6704 40772 6760 40828
rect 6760 40772 6764 40828
rect 6700 40768 6764 40772
rect 6780 40828 6844 40832
rect 6780 40772 6784 40828
rect 6784 40772 6840 40828
rect 6840 40772 6844 40828
rect 6780 40768 6844 40772
rect 6860 40828 6924 40832
rect 6860 40772 6864 40828
rect 6864 40772 6920 40828
rect 6920 40772 6924 40828
rect 6860 40768 6924 40772
rect 87212 40828 87276 40832
rect 87212 40772 87216 40828
rect 87216 40772 87272 40828
rect 87272 40772 87276 40828
rect 87212 40768 87276 40772
rect 87292 40828 87356 40832
rect 87292 40772 87296 40828
rect 87296 40772 87352 40828
rect 87352 40772 87356 40828
rect 87292 40768 87356 40772
rect 87372 40828 87436 40832
rect 87372 40772 87376 40828
rect 87376 40772 87432 40828
rect 87432 40772 87436 40828
rect 87372 40768 87436 40772
rect 87452 40828 87516 40832
rect 87452 40772 87456 40828
rect 87456 40772 87512 40828
rect 87512 40772 87516 40828
rect 87452 40768 87516 40772
rect 5884 40284 5948 40288
rect 5884 40228 5888 40284
rect 5888 40228 5944 40284
rect 5944 40228 5948 40284
rect 5884 40224 5948 40228
rect 5964 40284 6028 40288
rect 5964 40228 5968 40284
rect 5968 40228 6024 40284
rect 6024 40228 6028 40284
rect 5964 40224 6028 40228
rect 6044 40284 6108 40288
rect 6044 40228 6048 40284
rect 6048 40228 6104 40284
rect 6104 40228 6108 40284
rect 6044 40224 6108 40228
rect 6124 40284 6188 40288
rect 6124 40228 6128 40284
rect 6128 40228 6184 40284
rect 6184 40228 6188 40284
rect 6124 40224 6188 40228
rect 86476 40284 86540 40288
rect 86476 40228 86480 40284
rect 86480 40228 86536 40284
rect 86536 40228 86540 40284
rect 86476 40224 86540 40228
rect 86556 40284 86620 40288
rect 86556 40228 86560 40284
rect 86560 40228 86616 40284
rect 86616 40228 86620 40284
rect 86556 40224 86620 40228
rect 86636 40284 86700 40288
rect 86636 40228 86640 40284
rect 86640 40228 86696 40284
rect 86696 40228 86700 40284
rect 86636 40224 86700 40228
rect 86716 40284 86780 40288
rect 86716 40228 86720 40284
rect 86720 40228 86776 40284
rect 86776 40228 86780 40284
rect 86716 40224 86780 40228
rect 6620 39740 6684 39744
rect 6620 39684 6624 39740
rect 6624 39684 6680 39740
rect 6680 39684 6684 39740
rect 6620 39680 6684 39684
rect 6700 39740 6764 39744
rect 6700 39684 6704 39740
rect 6704 39684 6760 39740
rect 6760 39684 6764 39740
rect 6700 39680 6764 39684
rect 6780 39740 6844 39744
rect 6780 39684 6784 39740
rect 6784 39684 6840 39740
rect 6840 39684 6844 39740
rect 6780 39680 6844 39684
rect 6860 39740 6924 39744
rect 6860 39684 6864 39740
rect 6864 39684 6920 39740
rect 6920 39684 6924 39740
rect 6860 39680 6924 39684
rect 87212 39740 87276 39744
rect 87212 39684 87216 39740
rect 87216 39684 87272 39740
rect 87272 39684 87276 39740
rect 87212 39680 87276 39684
rect 87292 39740 87356 39744
rect 87292 39684 87296 39740
rect 87296 39684 87352 39740
rect 87352 39684 87356 39740
rect 87292 39680 87356 39684
rect 87372 39740 87436 39744
rect 87372 39684 87376 39740
rect 87376 39684 87432 39740
rect 87432 39684 87436 39740
rect 87372 39680 87436 39684
rect 87452 39740 87516 39744
rect 87452 39684 87456 39740
rect 87456 39684 87512 39740
rect 87512 39684 87516 39740
rect 87452 39680 87516 39684
rect 5884 39196 5948 39200
rect 5884 39140 5888 39196
rect 5888 39140 5944 39196
rect 5944 39140 5948 39196
rect 5884 39136 5948 39140
rect 5964 39196 6028 39200
rect 5964 39140 5968 39196
rect 5968 39140 6024 39196
rect 6024 39140 6028 39196
rect 5964 39136 6028 39140
rect 6044 39196 6108 39200
rect 6044 39140 6048 39196
rect 6048 39140 6104 39196
rect 6104 39140 6108 39196
rect 6044 39136 6108 39140
rect 6124 39196 6188 39200
rect 6124 39140 6128 39196
rect 6128 39140 6184 39196
rect 6184 39140 6188 39196
rect 6124 39136 6188 39140
rect 86476 39196 86540 39200
rect 86476 39140 86480 39196
rect 86480 39140 86536 39196
rect 86536 39140 86540 39196
rect 86476 39136 86540 39140
rect 86556 39196 86620 39200
rect 86556 39140 86560 39196
rect 86560 39140 86616 39196
rect 86616 39140 86620 39196
rect 86556 39136 86620 39140
rect 86636 39196 86700 39200
rect 86636 39140 86640 39196
rect 86640 39140 86696 39196
rect 86696 39140 86700 39196
rect 86636 39136 86700 39140
rect 86716 39196 86780 39200
rect 86716 39140 86720 39196
rect 86720 39140 86776 39196
rect 86776 39140 86780 39196
rect 86716 39136 86780 39140
rect 6620 38652 6684 38656
rect 6620 38596 6624 38652
rect 6624 38596 6680 38652
rect 6680 38596 6684 38652
rect 6620 38592 6684 38596
rect 6700 38652 6764 38656
rect 6700 38596 6704 38652
rect 6704 38596 6760 38652
rect 6760 38596 6764 38652
rect 6700 38592 6764 38596
rect 6780 38652 6844 38656
rect 6780 38596 6784 38652
rect 6784 38596 6840 38652
rect 6840 38596 6844 38652
rect 6780 38592 6844 38596
rect 6860 38652 6924 38656
rect 6860 38596 6864 38652
rect 6864 38596 6920 38652
rect 6920 38596 6924 38652
rect 6860 38592 6924 38596
rect 87212 38652 87276 38656
rect 87212 38596 87216 38652
rect 87216 38596 87272 38652
rect 87272 38596 87276 38652
rect 87212 38592 87276 38596
rect 87292 38652 87356 38656
rect 87292 38596 87296 38652
rect 87296 38596 87352 38652
rect 87352 38596 87356 38652
rect 87292 38592 87356 38596
rect 87372 38652 87436 38656
rect 87372 38596 87376 38652
rect 87376 38596 87432 38652
rect 87432 38596 87436 38652
rect 87372 38592 87436 38596
rect 87452 38652 87516 38656
rect 87452 38596 87456 38652
rect 87456 38596 87512 38652
rect 87512 38596 87516 38652
rect 87452 38592 87516 38596
rect 5884 38108 5948 38112
rect 5884 38052 5888 38108
rect 5888 38052 5944 38108
rect 5944 38052 5948 38108
rect 5884 38048 5948 38052
rect 5964 38108 6028 38112
rect 5964 38052 5968 38108
rect 5968 38052 6024 38108
rect 6024 38052 6028 38108
rect 5964 38048 6028 38052
rect 6044 38108 6108 38112
rect 6044 38052 6048 38108
rect 6048 38052 6104 38108
rect 6104 38052 6108 38108
rect 6044 38048 6108 38052
rect 6124 38108 6188 38112
rect 6124 38052 6128 38108
rect 6128 38052 6184 38108
rect 6184 38052 6188 38108
rect 6124 38048 6188 38052
rect 86476 38108 86540 38112
rect 86476 38052 86480 38108
rect 86480 38052 86536 38108
rect 86536 38052 86540 38108
rect 86476 38048 86540 38052
rect 86556 38108 86620 38112
rect 86556 38052 86560 38108
rect 86560 38052 86616 38108
rect 86616 38052 86620 38108
rect 86556 38048 86620 38052
rect 86636 38108 86700 38112
rect 86636 38052 86640 38108
rect 86640 38052 86696 38108
rect 86696 38052 86700 38108
rect 86636 38048 86700 38052
rect 86716 38108 86780 38112
rect 86716 38052 86720 38108
rect 86720 38052 86776 38108
rect 86776 38052 86780 38108
rect 86716 38048 86780 38052
rect 6620 37564 6684 37568
rect 6620 37508 6624 37564
rect 6624 37508 6680 37564
rect 6680 37508 6684 37564
rect 6620 37504 6684 37508
rect 6700 37564 6764 37568
rect 6700 37508 6704 37564
rect 6704 37508 6760 37564
rect 6760 37508 6764 37564
rect 6700 37504 6764 37508
rect 6780 37564 6844 37568
rect 6780 37508 6784 37564
rect 6784 37508 6840 37564
rect 6840 37508 6844 37564
rect 6780 37504 6844 37508
rect 6860 37564 6924 37568
rect 6860 37508 6864 37564
rect 6864 37508 6920 37564
rect 6920 37508 6924 37564
rect 6860 37504 6924 37508
rect 87212 37564 87276 37568
rect 87212 37508 87216 37564
rect 87216 37508 87272 37564
rect 87272 37508 87276 37564
rect 87212 37504 87276 37508
rect 87292 37564 87356 37568
rect 87292 37508 87296 37564
rect 87296 37508 87352 37564
rect 87352 37508 87356 37564
rect 87292 37504 87356 37508
rect 87372 37564 87436 37568
rect 87372 37508 87376 37564
rect 87376 37508 87432 37564
rect 87432 37508 87436 37564
rect 87372 37504 87436 37508
rect 87452 37564 87516 37568
rect 87452 37508 87456 37564
rect 87456 37508 87512 37564
rect 87512 37508 87516 37564
rect 87452 37504 87516 37508
rect 5884 37020 5948 37024
rect 5884 36964 5888 37020
rect 5888 36964 5944 37020
rect 5944 36964 5948 37020
rect 5884 36960 5948 36964
rect 5964 37020 6028 37024
rect 5964 36964 5968 37020
rect 5968 36964 6024 37020
rect 6024 36964 6028 37020
rect 5964 36960 6028 36964
rect 6044 37020 6108 37024
rect 6044 36964 6048 37020
rect 6048 36964 6104 37020
rect 6104 36964 6108 37020
rect 6044 36960 6108 36964
rect 6124 37020 6188 37024
rect 6124 36964 6128 37020
rect 6128 36964 6184 37020
rect 6184 36964 6188 37020
rect 6124 36960 6188 36964
rect 86476 37020 86540 37024
rect 86476 36964 86480 37020
rect 86480 36964 86536 37020
rect 86536 36964 86540 37020
rect 86476 36960 86540 36964
rect 86556 37020 86620 37024
rect 86556 36964 86560 37020
rect 86560 36964 86616 37020
rect 86616 36964 86620 37020
rect 86556 36960 86620 36964
rect 86636 37020 86700 37024
rect 86636 36964 86640 37020
rect 86640 36964 86696 37020
rect 86696 36964 86700 37020
rect 86636 36960 86700 36964
rect 86716 37020 86780 37024
rect 86716 36964 86720 37020
rect 86720 36964 86776 37020
rect 86776 36964 86780 37020
rect 86716 36960 86780 36964
rect 6620 36476 6684 36480
rect 6620 36420 6624 36476
rect 6624 36420 6680 36476
rect 6680 36420 6684 36476
rect 6620 36416 6684 36420
rect 6700 36476 6764 36480
rect 6700 36420 6704 36476
rect 6704 36420 6760 36476
rect 6760 36420 6764 36476
rect 6700 36416 6764 36420
rect 6780 36476 6844 36480
rect 6780 36420 6784 36476
rect 6784 36420 6840 36476
rect 6840 36420 6844 36476
rect 6780 36416 6844 36420
rect 6860 36476 6924 36480
rect 6860 36420 6864 36476
rect 6864 36420 6920 36476
rect 6920 36420 6924 36476
rect 6860 36416 6924 36420
rect 87212 36476 87276 36480
rect 87212 36420 87216 36476
rect 87216 36420 87272 36476
rect 87272 36420 87276 36476
rect 87212 36416 87276 36420
rect 87292 36476 87356 36480
rect 87292 36420 87296 36476
rect 87296 36420 87352 36476
rect 87352 36420 87356 36476
rect 87292 36416 87356 36420
rect 87372 36476 87436 36480
rect 87372 36420 87376 36476
rect 87376 36420 87432 36476
rect 87432 36420 87436 36476
rect 87372 36416 87436 36420
rect 87452 36476 87516 36480
rect 87452 36420 87456 36476
rect 87456 36420 87512 36476
rect 87512 36420 87516 36476
rect 87452 36416 87516 36420
rect 5884 35932 5948 35936
rect 5884 35876 5888 35932
rect 5888 35876 5944 35932
rect 5944 35876 5948 35932
rect 5884 35872 5948 35876
rect 5964 35932 6028 35936
rect 5964 35876 5968 35932
rect 5968 35876 6024 35932
rect 6024 35876 6028 35932
rect 5964 35872 6028 35876
rect 6044 35932 6108 35936
rect 6044 35876 6048 35932
rect 6048 35876 6104 35932
rect 6104 35876 6108 35932
rect 6044 35872 6108 35876
rect 6124 35932 6188 35936
rect 6124 35876 6128 35932
rect 6128 35876 6184 35932
rect 6184 35876 6188 35932
rect 6124 35872 6188 35876
rect 86476 35932 86540 35936
rect 86476 35876 86480 35932
rect 86480 35876 86536 35932
rect 86536 35876 86540 35932
rect 86476 35872 86540 35876
rect 86556 35932 86620 35936
rect 86556 35876 86560 35932
rect 86560 35876 86616 35932
rect 86616 35876 86620 35932
rect 86556 35872 86620 35876
rect 86636 35932 86700 35936
rect 86636 35876 86640 35932
rect 86640 35876 86696 35932
rect 86696 35876 86700 35932
rect 86636 35872 86700 35876
rect 86716 35932 86780 35936
rect 86716 35876 86720 35932
rect 86720 35876 86776 35932
rect 86776 35876 86780 35932
rect 86716 35872 86780 35876
rect 6620 35388 6684 35392
rect 6620 35332 6624 35388
rect 6624 35332 6680 35388
rect 6680 35332 6684 35388
rect 6620 35328 6684 35332
rect 6700 35388 6764 35392
rect 6700 35332 6704 35388
rect 6704 35332 6760 35388
rect 6760 35332 6764 35388
rect 6700 35328 6764 35332
rect 6780 35388 6844 35392
rect 6780 35332 6784 35388
rect 6784 35332 6840 35388
rect 6840 35332 6844 35388
rect 6780 35328 6844 35332
rect 6860 35388 6924 35392
rect 6860 35332 6864 35388
rect 6864 35332 6920 35388
rect 6920 35332 6924 35388
rect 6860 35328 6924 35332
rect 87212 35388 87276 35392
rect 87212 35332 87216 35388
rect 87216 35332 87272 35388
rect 87272 35332 87276 35388
rect 87212 35328 87276 35332
rect 87292 35388 87356 35392
rect 87292 35332 87296 35388
rect 87296 35332 87352 35388
rect 87352 35332 87356 35388
rect 87292 35328 87356 35332
rect 87372 35388 87436 35392
rect 87372 35332 87376 35388
rect 87376 35332 87432 35388
rect 87432 35332 87436 35388
rect 87372 35328 87436 35332
rect 87452 35388 87516 35392
rect 87452 35332 87456 35388
rect 87456 35332 87512 35388
rect 87512 35332 87516 35388
rect 87452 35328 87516 35332
rect 5884 34844 5948 34848
rect 5884 34788 5888 34844
rect 5888 34788 5944 34844
rect 5944 34788 5948 34844
rect 5884 34784 5948 34788
rect 5964 34844 6028 34848
rect 5964 34788 5968 34844
rect 5968 34788 6024 34844
rect 6024 34788 6028 34844
rect 5964 34784 6028 34788
rect 6044 34844 6108 34848
rect 6044 34788 6048 34844
rect 6048 34788 6104 34844
rect 6104 34788 6108 34844
rect 6044 34784 6108 34788
rect 6124 34844 6188 34848
rect 6124 34788 6128 34844
rect 6128 34788 6184 34844
rect 6184 34788 6188 34844
rect 6124 34784 6188 34788
rect 86476 34844 86540 34848
rect 86476 34788 86480 34844
rect 86480 34788 86536 34844
rect 86536 34788 86540 34844
rect 86476 34784 86540 34788
rect 86556 34844 86620 34848
rect 86556 34788 86560 34844
rect 86560 34788 86616 34844
rect 86616 34788 86620 34844
rect 86556 34784 86620 34788
rect 86636 34844 86700 34848
rect 86636 34788 86640 34844
rect 86640 34788 86696 34844
rect 86696 34788 86700 34844
rect 86636 34784 86700 34788
rect 86716 34844 86780 34848
rect 86716 34788 86720 34844
rect 86720 34788 86776 34844
rect 86776 34788 86780 34844
rect 86716 34784 86780 34788
rect 6620 34300 6684 34304
rect 6620 34244 6624 34300
rect 6624 34244 6680 34300
rect 6680 34244 6684 34300
rect 6620 34240 6684 34244
rect 6700 34300 6764 34304
rect 6700 34244 6704 34300
rect 6704 34244 6760 34300
rect 6760 34244 6764 34300
rect 6700 34240 6764 34244
rect 6780 34300 6844 34304
rect 6780 34244 6784 34300
rect 6784 34244 6840 34300
rect 6840 34244 6844 34300
rect 6780 34240 6844 34244
rect 6860 34300 6924 34304
rect 6860 34244 6864 34300
rect 6864 34244 6920 34300
rect 6920 34244 6924 34300
rect 6860 34240 6924 34244
rect 87212 34300 87276 34304
rect 87212 34244 87216 34300
rect 87216 34244 87272 34300
rect 87272 34244 87276 34300
rect 87212 34240 87276 34244
rect 87292 34300 87356 34304
rect 87292 34244 87296 34300
rect 87296 34244 87352 34300
rect 87352 34244 87356 34300
rect 87292 34240 87356 34244
rect 87372 34300 87436 34304
rect 87372 34244 87376 34300
rect 87376 34244 87432 34300
rect 87432 34244 87436 34300
rect 87372 34240 87436 34244
rect 87452 34300 87516 34304
rect 87452 34244 87456 34300
rect 87456 34244 87512 34300
rect 87512 34244 87516 34300
rect 87452 34240 87516 34244
rect 5884 33756 5948 33760
rect 5884 33700 5888 33756
rect 5888 33700 5944 33756
rect 5944 33700 5948 33756
rect 5884 33696 5948 33700
rect 5964 33756 6028 33760
rect 5964 33700 5968 33756
rect 5968 33700 6024 33756
rect 6024 33700 6028 33756
rect 5964 33696 6028 33700
rect 6044 33756 6108 33760
rect 6044 33700 6048 33756
rect 6048 33700 6104 33756
rect 6104 33700 6108 33756
rect 6044 33696 6108 33700
rect 6124 33756 6188 33760
rect 6124 33700 6128 33756
rect 6128 33700 6184 33756
rect 6184 33700 6188 33756
rect 6124 33696 6188 33700
rect 86476 33756 86540 33760
rect 86476 33700 86480 33756
rect 86480 33700 86536 33756
rect 86536 33700 86540 33756
rect 86476 33696 86540 33700
rect 86556 33756 86620 33760
rect 86556 33700 86560 33756
rect 86560 33700 86616 33756
rect 86616 33700 86620 33756
rect 86556 33696 86620 33700
rect 86636 33756 86700 33760
rect 86636 33700 86640 33756
rect 86640 33700 86696 33756
rect 86696 33700 86700 33756
rect 86636 33696 86700 33700
rect 86716 33756 86780 33760
rect 86716 33700 86720 33756
rect 86720 33700 86776 33756
rect 86776 33700 86780 33756
rect 86716 33696 86780 33700
rect 6620 33212 6684 33216
rect 6620 33156 6624 33212
rect 6624 33156 6680 33212
rect 6680 33156 6684 33212
rect 6620 33152 6684 33156
rect 6700 33212 6764 33216
rect 6700 33156 6704 33212
rect 6704 33156 6760 33212
rect 6760 33156 6764 33212
rect 6700 33152 6764 33156
rect 6780 33212 6844 33216
rect 6780 33156 6784 33212
rect 6784 33156 6840 33212
rect 6840 33156 6844 33212
rect 6780 33152 6844 33156
rect 6860 33212 6924 33216
rect 6860 33156 6864 33212
rect 6864 33156 6920 33212
rect 6920 33156 6924 33212
rect 6860 33152 6924 33156
rect 87212 33212 87276 33216
rect 87212 33156 87216 33212
rect 87216 33156 87272 33212
rect 87272 33156 87276 33212
rect 87212 33152 87276 33156
rect 87292 33212 87356 33216
rect 87292 33156 87296 33212
rect 87296 33156 87352 33212
rect 87352 33156 87356 33212
rect 87292 33152 87356 33156
rect 87372 33212 87436 33216
rect 87372 33156 87376 33212
rect 87376 33156 87432 33212
rect 87432 33156 87436 33212
rect 87372 33152 87436 33156
rect 87452 33212 87516 33216
rect 87452 33156 87456 33212
rect 87456 33156 87512 33212
rect 87512 33156 87516 33212
rect 87452 33152 87516 33156
rect 5884 32668 5948 32672
rect 5884 32612 5888 32668
rect 5888 32612 5944 32668
rect 5944 32612 5948 32668
rect 5884 32608 5948 32612
rect 5964 32668 6028 32672
rect 5964 32612 5968 32668
rect 5968 32612 6024 32668
rect 6024 32612 6028 32668
rect 5964 32608 6028 32612
rect 6044 32668 6108 32672
rect 6044 32612 6048 32668
rect 6048 32612 6104 32668
rect 6104 32612 6108 32668
rect 6044 32608 6108 32612
rect 6124 32668 6188 32672
rect 6124 32612 6128 32668
rect 6128 32612 6184 32668
rect 6184 32612 6188 32668
rect 6124 32608 6188 32612
rect 86476 32668 86540 32672
rect 86476 32612 86480 32668
rect 86480 32612 86536 32668
rect 86536 32612 86540 32668
rect 86476 32608 86540 32612
rect 86556 32668 86620 32672
rect 86556 32612 86560 32668
rect 86560 32612 86616 32668
rect 86616 32612 86620 32668
rect 86556 32608 86620 32612
rect 86636 32668 86700 32672
rect 86636 32612 86640 32668
rect 86640 32612 86696 32668
rect 86696 32612 86700 32668
rect 86636 32608 86700 32612
rect 86716 32668 86780 32672
rect 86716 32612 86720 32668
rect 86720 32612 86776 32668
rect 86776 32612 86780 32668
rect 86716 32608 86780 32612
rect 6620 32124 6684 32128
rect 6620 32068 6624 32124
rect 6624 32068 6680 32124
rect 6680 32068 6684 32124
rect 6620 32064 6684 32068
rect 6700 32124 6764 32128
rect 6700 32068 6704 32124
rect 6704 32068 6760 32124
rect 6760 32068 6764 32124
rect 6700 32064 6764 32068
rect 6780 32124 6844 32128
rect 6780 32068 6784 32124
rect 6784 32068 6840 32124
rect 6840 32068 6844 32124
rect 6780 32064 6844 32068
rect 6860 32124 6924 32128
rect 6860 32068 6864 32124
rect 6864 32068 6920 32124
rect 6920 32068 6924 32124
rect 6860 32064 6924 32068
rect 87212 32124 87276 32128
rect 87212 32068 87216 32124
rect 87216 32068 87272 32124
rect 87272 32068 87276 32124
rect 87212 32064 87276 32068
rect 87292 32124 87356 32128
rect 87292 32068 87296 32124
rect 87296 32068 87352 32124
rect 87352 32068 87356 32124
rect 87292 32064 87356 32068
rect 87372 32124 87436 32128
rect 87372 32068 87376 32124
rect 87376 32068 87432 32124
rect 87432 32068 87436 32124
rect 87372 32064 87436 32068
rect 87452 32124 87516 32128
rect 87452 32068 87456 32124
rect 87456 32068 87512 32124
rect 87512 32068 87516 32124
rect 87452 32064 87516 32068
rect 5884 31580 5948 31584
rect 5884 31524 5888 31580
rect 5888 31524 5944 31580
rect 5944 31524 5948 31580
rect 5884 31520 5948 31524
rect 5964 31580 6028 31584
rect 5964 31524 5968 31580
rect 5968 31524 6024 31580
rect 6024 31524 6028 31580
rect 5964 31520 6028 31524
rect 6044 31580 6108 31584
rect 6044 31524 6048 31580
rect 6048 31524 6104 31580
rect 6104 31524 6108 31580
rect 6044 31520 6108 31524
rect 6124 31580 6188 31584
rect 6124 31524 6128 31580
rect 6128 31524 6184 31580
rect 6184 31524 6188 31580
rect 6124 31520 6188 31524
rect 86476 31580 86540 31584
rect 86476 31524 86480 31580
rect 86480 31524 86536 31580
rect 86536 31524 86540 31580
rect 86476 31520 86540 31524
rect 86556 31580 86620 31584
rect 86556 31524 86560 31580
rect 86560 31524 86616 31580
rect 86616 31524 86620 31580
rect 86556 31520 86620 31524
rect 86636 31580 86700 31584
rect 86636 31524 86640 31580
rect 86640 31524 86696 31580
rect 86696 31524 86700 31580
rect 86636 31520 86700 31524
rect 86716 31580 86780 31584
rect 86716 31524 86720 31580
rect 86720 31524 86776 31580
rect 86776 31524 86780 31580
rect 86716 31520 86780 31524
rect 6620 31036 6684 31040
rect 6620 30980 6624 31036
rect 6624 30980 6680 31036
rect 6680 30980 6684 31036
rect 6620 30976 6684 30980
rect 6700 31036 6764 31040
rect 6700 30980 6704 31036
rect 6704 30980 6760 31036
rect 6760 30980 6764 31036
rect 6700 30976 6764 30980
rect 6780 31036 6844 31040
rect 6780 30980 6784 31036
rect 6784 30980 6840 31036
rect 6840 30980 6844 31036
rect 6780 30976 6844 30980
rect 6860 31036 6924 31040
rect 6860 30980 6864 31036
rect 6864 30980 6920 31036
rect 6920 30980 6924 31036
rect 6860 30976 6924 30980
rect 87212 31036 87276 31040
rect 87212 30980 87216 31036
rect 87216 30980 87272 31036
rect 87272 30980 87276 31036
rect 87212 30976 87276 30980
rect 87292 31036 87356 31040
rect 87292 30980 87296 31036
rect 87296 30980 87352 31036
rect 87352 30980 87356 31036
rect 87292 30976 87356 30980
rect 87372 31036 87436 31040
rect 87372 30980 87376 31036
rect 87376 30980 87432 31036
rect 87432 30980 87436 31036
rect 87372 30976 87436 30980
rect 87452 31036 87516 31040
rect 87452 30980 87456 31036
rect 87456 30980 87512 31036
rect 87512 30980 87516 31036
rect 87452 30976 87516 30980
rect 5884 30492 5948 30496
rect 5884 30436 5888 30492
rect 5888 30436 5944 30492
rect 5944 30436 5948 30492
rect 5884 30432 5948 30436
rect 5964 30492 6028 30496
rect 5964 30436 5968 30492
rect 5968 30436 6024 30492
rect 6024 30436 6028 30492
rect 5964 30432 6028 30436
rect 6044 30492 6108 30496
rect 6044 30436 6048 30492
rect 6048 30436 6104 30492
rect 6104 30436 6108 30492
rect 6044 30432 6108 30436
rect 6124 30492 6188 30496
rect 6124 30436 6128 30492
rect 6128 30436 6184 30492
rect 6184 30436 6188 30492
rect 6124 30432 6188 30436
rect 86476 30492 86540 30496
rect 86476 30436 86480 30492
rect 86480 30436 86536 30492
rect 86536 30436 86540 30492
rect 86476 30432 86540 30436
rect 86556 30492 86620 30496
rect 86556 30436 86560 30492
rect 86560 30436 86616 30492
rect 86616 30436 86620 30492
rect 86556 30432 86620 30436
rect 86636 30492 86700 30496
rect 86636 30436 86640 30492
rect 86640 30436 86696 30492
rect 86696 30436 86700 30492
rect 86636 30432 86700 30436
rect 86716 30492 86780 30496
rect 86716 30436 86720 30492
rect 86720 30436 86776 30492
rect 86776 30436 86780 30492
rect 86716 30432 86780 30436
rect 6620 29948 6684 29952
rect 6620 29892 6624 29948
rect 6624 29892 6680 29948
rect 6680 29892 6684 29948
rect 6620 29888 6684 29892
rect 6700 29948 6764 29952
rect 6700 29892 6704 29948
rect 6704 29892 6760 29948
rect 6760 29892 6764 29948
rect 6700 29888 6764 29892
rect 6780 29948 6844 29952
rect 6780 29892 6784 29948
rect 6784 29892 6840 29948
rect 6840 29892 6844 29948
rect 6780 29888 6844 29892
rect 6860 29948 6924 29952
rect 6860 29892 6864 29948
rect 6864 29892 6920 29948
rect 6920 29892 6924 29948
rect 6860 29888 6924 29892
rect 87212 29948 87276 29952
rect 87212 29892 87216 29948
rect 87216 29892 87272 29948
rect 87272 29892 87276 29948
rect 87212 29888 87276 29892
rect 87292 29948 87356 29952
rect 87292 29892 87296 29948
rect 87296 29892 87352 29948
rect 87352 29892 87356 29948
rect 87292 29888 87356 29892
rect 87372 29948 87436 29952
rect 87372 29892 87376 29948
rect 87376 29892 87432 29948
rect 87432 29892 87436 29948
rect 87372 29888 87436 29892
rect 87452 29948 87516 29952
rect 87452 29892 87456 29948
rect 87456 29892 87512 29948
rect 87512 29892 87516 29948
rect 87452 29888 87516 29892
rect 5884 29404 5948 29408
rect 5884 29348 5888 29404
rect 5888 29348 5944 29404
rect 5944 29348 5948 29404
rect 5884 29344 5948 29348
rect 5964 29404 6028 29408
rect 5964 29348 5968 29404
rect 5968 29348 6024 29404
rect 6024 29348 6028 29404
rect 5964 29344 6028 29348
rect 6044 29404 6108 29408
rect 6044 29348 6048 29404
rect 6048 29348 6104 29404
rect 6104 29348 6108 29404
rect 6044 29344 6108 29348
rect 6124 29404 6188 29408
rect 6124 29348 6128 29404
rect 6128 29348 6184 29404
rect 6184 29348 6188 29404
rect 6124 29344 6188 29348
rect 86476 29404 86540 29408
rect 86476 29348 86480 29404
rect 86480 29348 86536 29404
rect 86536 29348 86540 29404
rect 86476 29344 86540 29348
rect 86556 29404 86620 29408
rect 86556 29348 86560 29404
rect 86560 29348 86616 29404
rect 86616 29348 86620 29404
rect 86556 29344 86620 29348
rect 86636 29404 86700 29408
rect 86636 29348 86640 29404
rect 86640 29348 86696 29404
rect 86696 29348 86700 29404
rect 86636 29344 86700 29348
rect 86716 29404 86780 29408
rect 86716 29348 86720 29404
rect 86720 29348 86776 29404
rect 86776 29348 86780 29404
rect 86716 29344 86780 29348
rect 6620 28860 6684 28864
rect 6620 28804 6624 28860
rect 6624 28804 6680 28860
rect 6680 28804 6684 28860
rect 6620 28800 6684 28804
rect 6700 28860 6764 28864
rect 6700 28804 6704 28860
rect 6704 28804 6760 28860
rect 6760 28804 6764 28860
rect 6700 28800 6764 28804
rect 6780 28860 6844 28864
rect 6780 28804 6784 28860
rect 6784 28804 6840 28860
rect 6840 28804 6844 28860
rect 6780 28800 6844 28804
rect 6860 28860 6924 28864
rect 6860 28804 6864 28860
rect 6864 28804 6920 28860
rect 6920 28804 6924 28860
rect 6860 28800 6924 28804
rect 87212 28860 87276 28864
rect 87212 28804 87216 28860
rect 87216 28804 87272 28860
rect 87272 28804 87276 28860
rect 87212 28800 87276 28804
rect 87292 28860 87356 28864
rect 87292 28804 87296 28860
rect 87296 28804 87352 28860
rect 87352 28804 87356 28860
rect 87292 28800 87356 28804
rect 87372 28860 87436 28864
rect 87372 28804 87376 28860
rect 87376 28804 87432 28860
rect 87432 28804 87436 28860
rect 87372 28800 87436 28804
rect 87452 28860 87516 28864
rect 87452 28804 87456 28860
rect 87456 28804 87512 28860
rect 87512 28804 87516 28860
rect 87452 28800 87516 28804
rect 5884 28316 5948 28320
rect 5884 28260 5888 28316
rect 5888 28260 5944 28316
rect 5944 28260 5948 28316
rect 5884 28256 5948 28260
rect 5964 28316 6028 28320
rect 5964 28260 5968 28316
rect 5968 28260 6024 28316
rect 6024 28260 6028 28316
rect 5964 28256 6028 28260
rect 6044 28316 6108 28320
rect 6044 28260 6048 28316
rect 6048 28260 6104 28316
rect 6104 28260 6108 28316
rect 6044 28256 6108 28260
rect 6124 28316 6188 28320
rect 6124 28260 6128 28316
rect 6128 28260 6184 28316
rect 6184 28260 6188 28316
rect 6124 28256 6188 28260
rect 86476 28316 86540 28320
rect 86476 28260 86480 28316
rect 86480 28260 86536 28316
rect 86536 28260 86540 28316
rect 86476 28256 86540 28260
rect 86556 28316 86620 28320
rect 86556 28260 86560 28316
rect 86560 28260 86616 28316
rect 86616 28260 86620 28316
rect 86556 28256 86620 28260
rect 86636 28316 86700 28320
rect 86636 28260 86640 28316
rect 86640 28260 86696 28316
rect 86696 28260 86700 28316
rect 86636 28256 86700 28260
rect 86716 28316 86780 28320
rect 86716 28260 86720 28316
rect 86720 28260 86776 28316
rect 86776 28260 86780 28316
rect 86716 28256 86780 28260
rect 6620 27772 6684 27776
rect 6620 27716 6624 27772
rect 6624 27716 6680 27772
rect 6680 27716 6684 27772
rect 6620 27712 6684 27716
rect 6700 27772 6764 27776
rect 6700 27716 6704 27772
rect 6704 27716 6760 27772
rect 6760 27716 6764 27772
rect 6700 27712 6764 27716
rect 6780 27772 6844 27776
rect 6780 27716 6784 27772
rect 6784 27716 6840 27772
rect 6840 27716 6844 27772
rect 6780 27712 6844 27716
rect 6860 27772 6924 27776
rect 6860 27716 6864 27772
rect 6864 27716 6920 27772
rect 6920 27716 6924 27772
rect 6860 27712 6924 27716
rect 87212 27772 87276 27776
rect 87212 27716 87216 27772
rect 87216 27716 87272 27772
rect 87272 27716 87276 27772
rect 87212 27712 87276 27716
rect 87292 27772 87356 27776
rect 87292 27716 87296 27772
rect 87296 27716 87352 27772
rect 87352 27716 87356 27772
rect 87292 27712 87356 27716
rect 87372 27772 87436 27776
rect 87372 27716 87376 27772
rect 87376 27716 87432 27772
rect 87432 27716 87436 27772
rect 87372 27712 87436 27716
rect 87452 27772 87516 27776
rect 87452 27716 87456 27772
rect 87456 27716 87512 27772
rect 87512 27716 87516 27772
rect 87452 27712 87516 27716
rect 5884 27228 5948 27232
rect 5884 27172 5888 27228
rect 5888 27172 5944 27228
rect 5944 27172 5948 27228
rect 5884 27168 5948 27172
rect 5964 27228 6028 27232
rect 5964 27172 5968 27228
rect 5968 27172 6024 27228
rect 6024 27172 6028 27228
rect 5964 27168 6028 27172
rect 6044 27228 6108 27232
rect 6044 27172 6048 27228
rect 6048 27172 6104 27228
rect 6104 27172 6108 27228
rect 6044 27168 6108 27172
rect 6124 27228 6188 27232
rect 6124 27172 6128 27228
rect 6128 27172 6184 27228
rect 6184 27172 6188 27228
rect 6124 27168 6188 27172
rect 86476 27228 86540 27232
rect 86476 27172 86480 27228
rect 86480 27172 86536 27228
rect 86536 27172 86540 27228
rect 86476 27168 86540 27172
rect 86556 27228 86620 27232
rect 86556 27172 86560 27228
rect 86560 27172 86616 27228
rect 86616 27172 86620 27228
rect 86556 27168 86620 27172
rect 86636 27228 86700 27232
rect 86636 27172 86640 27228
rect 86640 27172 86696 27228
rect 86696 27172 86700 27228
rect 86636 27168 86700 27172
rect 86716 27228 86780 27232
rect 86716 27172 86720 27228
rect 86720 27172 86776 27228
rect 86776 27172 86780 27228
rect 86716 27168 86780 27172
rect 6620 26684 6684 26688
rect 6620 26628 6624 26684
rect 6624 26628 6680 26684
rect 6680 26628 6684 26684
rect 6620 26624 6684 26628
rect 6700 26684 6764 26688
rect 6700 26628 6704 26684
rect 6704 26628 6760 26684
rect 6760 26628 6764 26684
rect 6700 26624 6764 26628
rect 6780 26684 6844 26688
rect 6780 26628 6784 26684
rect 6784 26628 6840 26684
rect 6840 26628 6844 26684
rect 6780 26624 6844 26628
rect 6860 26684 6924 26688
rect 6860 26628 6864 26684
rect 6864 26628 6920 26684
rect 6920 26628 6924 26684
rect 6860 26624 6924 26628
rect 87212 26684 87276 26688
rect 87212 26628 87216 26684
rect 87216 26628 87272 26684
rect 87272 26628 87276 26684
rect 87212 26624 87276 26628
rect 87292 26684 87356 26688
rect 87292 26628 87296 26684
rect 87296 26628 87352 26684
rect 87352 26628 87356 26684
rect 87292 26624 87356 26628
rect 87372 26684 87436 26688
rect 87372 26628 87376 26684
rect 87376 26628 87432 26684
rect 87432 26628 87436 26684
rect 87372 26624 87436 26628
rect 87452 26684 87516 26688
rect 87452 26628 87456 26684
rect 87456 26628 87512 26684
rect 87512 26628 87516 26684
rect 87452 26624 87516 26628
rect 5884 26140 5948 26144
rect 5884 26084 5888 26140
rect 5888 26084 5944 26140
rect 5944 26084 5948 26140
rect 5884 26080 5948 26084
rect 5964 26140 6028 26144
rect 5964 26084 5968 26140
rect 5968 26084 6024 26140
rect 6024 26084 6028 26140
rect 5964 26080 6028 26084
rect 6044 26140 6108 26144
rect 6044 26084 6048 26140
rect 6048 26084 6104 26140
rect 6104 26084 6108 26140
rect 6044 26080 6108 26084
rect 6124 26140 6188 26144
rect 6124 26084 6128 26140
rect 6128 26084 6184 26140
rect 6184 26084 6188 26140
rect 6124 26080 6188 26084
rect 86476 26140 86540 26144
rect 86476 26084 86480 26140
rect 86480 26084 86536 26140
rect 86536 26084 86540 26140
rect 86476 26080 86540 26084
rect 86556 26140 86620 26144
rect 86556 26084 86560 26140
rect 86560 26084 86616 26140
rect 86616 26084 86620 26140
rect 86556 26080 86620 26084
rect 86636 26140 86700 26144
rect 86636 26084 86640 26140
rect 86640 26084 86696 26140
rect 86696 26084 86700 26140
rect 86636 26080 86700 26084
rect 86716 26140 86780 26144
rect 86716 26084 86720 26140
rect 86720 26084 86776 26140
rect 86776 26084 86780 26140
rect 86716 26080 86780 26084
rect 6620 25596 6684 25600
rect 6620 25540 6624 25596
rect 6624 25540 6680 25596
rect 6680 25540 6684 25596
rect 6620 25536 6684 25540
rect 6700 25596 6764 25600
rect 6700 25540 6704 25596
rect 6704 25540 6760 25596
rect 6760 25540 6764 25596
rect 6700 25536 6764 25540
rect 6780 25596 6844 25600
rect 6780 25540 6784 25596
rect 6784 25540 6840 25596
rect 6840 25540 6844 25596
rect 6780 25536 6844 25540
rect 6860 25596 6924 25600
rect 6860 25540 6864 25596
rect 6864 25540 6920 25596
rect 6920 25540 6924 25596
rect 6860 25536 6924 25540
rect 87212 25596 87276 25600
rect 87212 25540 87216 25596
rect 87216 25540 87272 25596
rect 87272 25540 87276 25596
rect 87212 25536 87276 25540
rect 87292 25596 87356 25600
rect 87292 25540 87296 25596
rect 87296 25540 87352 25596
rect 87352 25540 87356 25596
rect 87292 25536 87356 25540
rect 87372 25596 87436 25600
rect 87372 25540 87376 25596
rect 87376 25540 87432 25596
rect 87432 25540 87436 25596
rect 87372 25536 87436 25540
rect 87452 25596 87516 25600
rect 87452 25540 87456 25596
rect 87456 25540 87512 25596
rect 87512 25540 87516 25596
rect 87452 25536 87516 25540
rect 5884 25052 5948 25056
rect 5884 24996 5888 25052
rect 5888 24996 5944 25052
rect 5944 24996 5948 25052
rect 5884 24992 5948 24996
rect 5964 25052 6028 25056
rect 5964 24996 5968 25052
rect 5968 24996 6024 25052
rect 6024 24996 6028 25052
rect 5964 24992 6028 24996
rect 6044 25052 6108 25056
rect 6044 24996 6048 25052
rect 6048 24996 6104 25052
rect 6104 24996 6108 25052
rect 6044 24992 6108 24996
rect 6124 25052 6188 25056
rect 6124 24996 6128 25052
rect 6128 24996 6184 25052
rect 6184 24996 6188 25052
rect 6124 24992 6188 24996
rect 86476 25052 86540 25056
rect 86476 24996 86480 25052
rect 86480 24996 86536 25052
rect 86536 24996 86540 25052
rect 86476 24992 86540 24996
rect 86556 25052 86620 25056
rect 86556 24996 86560 25052
rect 86560 24996 86616 25052
rect 86616 24996 86620 25052
rect 86556 24992 86620 24996
rect 86636 25052 86700 25056
rect 86636 24996 86640 25052
rect 86640 24996 86696 25052
rect 86696 24996 86700 25052
rect 86636 24992 86700 24996
rect 86716 25052 86780 25056
rect 86716 24996 86720 25052
rect 86720 24996 86776 25052
rect 86776 24996 86780 25052
rect 86716 24992 86780 24996
rect 6620 24508 6684 24512
rect 6620 24452 6624 24508
rect 6624 24452 6680 24508
rect 6680 24452 6684 24508
rect 6620 24448 6684 24452
rect 6700 24508 6764 24512
rect 6700 24452 6704 24508
rect 6704 24452 6760 24508
rect 6760 24452 6764 24508
rect 6700 24448 6764 24452
rect 6780 24508 6844 24512
rect 6780 24452 6784 24508
rect 6784 24452 6840 24508
rect 6840 24452 6844 24508
rect 6780 24448 6844 24452
rect 6860 24508 6924 24512
rect 6860 24452 6864 24508
rect 6864 24452 6920 24508
rect 6920 24452 6924 24508
rect 6860 24448 6924 24452
rect 87212 24508 87276 24512
rect 87212 24452 87216 24508
rect 87216 24452 87272 24508
rect 87272 24452 87276 24508
rect 87212 24448 87276 24452
rect 87292 24508 87356 24512
rect 87292 24452 87296 24508
rect 87296 24452 87352 24508
rect 87352 24452 87356 24508
rect 87292 24448 87356 24452
rect 87372 24508 87436 24512
rect 87372 24452 87376 24508
rect 87376 24452 87432 24508
rect 87432 24452 87436 24508
rect 87372 24448 87436 24452
rect 87452 24508 87516 24512
rect 87452 24452 87456 24508
rect 87456 24452 87512 24508
rect 87512 24452 87516 24508
rect 87452 24448 87516 24452
rect 5884 23964 5948 23968
rect 5884 23908 5888 23964
rect 5888 23908 5944 23964
rect 5944 23908 5948 23964
rect 5884 23904 5948 23908
rect 5964 23964 6028 23968
rect 5964 23908 5968 23964
rect 5968 23908 6024 23964
rect 6024 23908 6028 23964
rect 5964 23904 6028 23908
rect 6044 23964 6108 23968
rect 6044 23908 6048 23964
rect 6048 23908 6104 23964
rect 6104 23908 6108 23964
rect 6044 23904 6108 23908
rect 6124 23964 6188 23968
rect 6124 23908 6128 23964
rect 6128 23908 6184 23964
rect 6184 23908 6188 23964
rect 6124 23904 6188 23908
rect 86476 23964 86540 23968
rect 86476 23908 86480 23964
rect 86480 23908 86536 23964
rect 86536 23908 86540 23964
rect 86476 23904 86540 23908
rect 86556 23964 86620 23968
rect 86556 23908 86560 23964
rect 86560 23908 86616 23964
rect 86616 23908 86620 23964
rect 86556 23904 86620 23908
rect 86636 23964 86700 23968
rect 86636 23908 86640 23964
rect 86640 23908 86696 23964
rect 86696 23908 86700 23964
rect 86636 23904 86700 23908
rect 86716 23964 86780 23968
rect 86716 23908 86720 23964
rect 86720 23908 86776 23964
rect 86776 23908 86780 23964
rect 86716 23904 86780 23908
rect 6620 23420 6684 23424
rect 6620 23364 6624 23420
rect 6624 23364 6680 23420
rect 6680 23364 6684 23420
rect 6620 23360 6684 23364
rect 6700 23420 6764 23424
rect 6700 23364 6704 23420
rect 6704 23364 6760 23420
rect 6760 23364 6764 23420
rect 6700 23360 6764 23364
rect 6780 23420 6844 23424
rect 6780 23364 6784 23420
rect 6784 23364 6840 23420
rect 6840 23364 6844 23420
rect 6780 23360 6844 23364
rect 6860 23420 6924 23424
rect 6860 23364 6864 23420
rect 6864 23364 6920 23420
rect 6920 23364 6924 23420
rect 6860 23360 6924 23364
rect 87212 23420 87276 23424
rect 87212 23364 87216 23420
rect 87216 23364 87272 23420
rect 87272 23364 87276 23420
rect 87212 23360 87276 23364
rect 87292 23420 87356 23424
rect 87292 23364 87296 23420
rect 87296 23364 87352 23420
rect 87352 23364 87356 23420
rect 87292 23360 87356 23364
rect 87372 23420 87436 23424
rect 87372 23364 87376 23420
rect 87376 23364 87432 23420
rect 87432 23364 87436 23420
rect 87372 23360 87436 23364
rect 87452 23420 87516 23424
rect 87452 23364 87456 23420
rect 87456 23364 87512 23420
rect 87512 23364 87516 23420
rect 87452 23360 87516 23364
rect 5884 22876 5948 22880
rect 5884 22820 5888 22876
rect 5888 22820 5944 22876
rect 5944 22820 5948 22876
rect 5884 22816 5948 22820
rect 5964 22876 6028 22880
rect 5964 22820 5968 22876
rect 5968 22820 6024 22876
rect 6024 22820 6028 22876
rect 5964 22816 6028 22820
rect 6044 22876 6108 22880
rect 6044 22820 6048 22876
rect 6048 22820 6104 22876
rect 6104 22820 6108 22876
rect 6044 22816 6108 22820
rect 6124 22876 6188 22880
rect 6124 22820 6128 22876
rect 6128 22820 6184 22876
rect 6184 22820 6188 22876
rect 6124 22816 6188 22820
rect 86476 22876 86540 22880
rect 86476 22820 86480 22876
rect 86480 22820 86536 22876
rect 86536 22820 86540 22876
rect 86476 22816 86540 22820
rect 86556 22876 86620 22880
rect 86556 22820 86560 22876
rect 86560 22820 86616 22876
rect 86616 22820 86620 22876
rect 86556 22816 86620 22820
rect 86636 22876 86700 22880
rect 86636 22820 86640 22876
rect 86640 22820 86696 22876
rect 86696 22820 86700 22876
rect 86636 22816 86700 22820
rect 86716 22876 86780 22880
rect 86716 22820 86720 22876
rect 86720 22820 86776 22876
rect 86776 22820 86780 22876
rect 86716 22816 86780 22820
rect 6620 22332 6684 22336
rect 6620 22276 6624 22332
rect 6624 22276 6680 22332
rect 6680 22276 6684 22332
rect 6620 22272 6684 22276
rect 6700 22332 6764 22336
rect 6700 22276 6704 22332
rect 6704 22276 6760 22332
rect 6760 22276 6764 22332
rect 6700 22272 6764 22276
rect 6780 22332 6844 22336
rect 6780 22276 6784 22332
rect 6784 22276 6840 22332
rect 6840 22276 6844 22332
rect 6780 22272 6844 22276
rect 6860 22332 6924 22336
rect 6860 22276 6864 22332
rect 6864 22276 6920 22332
rect 6920 22276 6924 22332
rect 6860 22272 6924 22276
rect 87212 22332 87276 22336
rect 87212 22276 87216 22332
rect 87216 22276 87272 22332
rect 87272 22276 87276 22332
rect 87212 22272 87276 22276
rect 87292 22332 87356 22336
rect 87292 22276 87296 22332
rect 87296 22276 87352 22332
rect 87352 22276 87356 22332
rect 87292 22272 87356 22276
rect 87372 22332 87436 22336
rect 87372 22276 87376 22332
rect 87376 22276 87432 22332
rect 87432 22276 87436 22332
rect 87372 22272 87436 22276
rect 87452 22332 87516 22336
rect 87452 22276 87456 22332
rect 87456 22276 87512 22332
rect 87512 22276 87516 22332
rect 87452 22272 87516 22276
rect 5884 21788 5948 21792
rect 5884 21732 5888 21788
rect 5888 21732 5944 21788
rect 5944 21732 5948 21788
rect 5884 21728 5948 21732
rect 5964 21788 6028 21792
rect 5964 21732 5968 21788
rect 5968 21732 6024 21788
rect 6024 21732 6028 21788
rect 5964 21728 6028 21732
rect 6044 21788 6108 21792
rect 6044 21732 6048 21788
rect 6048 21732 6104 21788
rect 6104 21732 6108 21788
rect 6044 21728 6108 21732
rect 6124 21788 6188 21792
rect 6124 21732 6128 21788
rect 6128 21732 6184 21788
rect 6184 21732 6188 21788
rect 6124 21728 6188 21732
rect 86476 21788 86540 21792
rect 86476 21732 86480 21788
rect 86480 21732 86536 21788
rect 86536 21732 86540 21788
rect 86476 21728 86540 21732
rect 86556 21788 86620 21792
rect 86556 21732 86560 21788
rect 86560 21732 86616 21788
rect 86616 21732 86620 21788
rect 86556 21728 86620 21732
rect 86636 21788 86700 21792
rect 86636 21732 86640 21788
rect 86640 21732 86696 21788
rect 86696 21732 86700 21788
rect 86636 21728 86700 21732
rect 86716 21788 86780 21792
rect 86716 21732 86720 21788
rect 86720 21732 86776 21788
rect 86776 21732 86780 21788
rect 86716 21728 86780 21732
rect 6620 21244 6684 21248
rect 6620 21188 6624 21244
rect 6624 21188 6680 21244
rect 6680 21188 6684 21244
rect 6620 21184 6684 21188
rect 6700 21244 6764 21248
rect 6700 21188 6704 21244
rect 6704 21188 6760 21244
rect 6760 21188 6764 21244
rect 6700 21184 6764 21188
rect 6780 21244 6844 21248
rect 6780 21188 6784 21244
rect 6784 21188 6840 21244
rect 6840 21188 6844 21244
rect 6780 21184 6844 21188
rect 6860 21244 6924 21248
rect 6860 21188 6864 21244
rect 6864 21188 6920 21244
rect 6920 21188 6924 21244
rect 6860 21184 6924 21188
rect 87212 21244 87276 21248
rect 87212 21188 87216 21244
rect 87216 21188 87272 21244
rect 87272 21188 87276 21244
rect 87212 21184 87276 21188
rect 87292 21244 87356 21248
rect 87292 21188 87296 21244
rect 87296 21188 87352 21244
rect 87352 21188 87356 21244
rect 87292 21184 87356 21188
rect 87372 21244 87436 21248
rect 87372 21188 87376 21244
rect 87376 21188 87432 21244
rect 87432 21188 87436 21244
rect 87372 21184 87436 21188
rect 87452 21244 87516 21248
rect 87452 21188 87456 21244
rect 87456 21188 87512 21244
rect 87512 21188 87516 21244
rect 87452 21184 87516 21188
rect 5884 20700 5948 20704
rect 5884 20644 5888 20700
rect 5888 20644 5944 20700
rect 5944 20644 5948 20700
rect 5884 20640 5948 20644
rect 5964 20700 6028 20704
rect 5964 20644 5968 20700
rect 5968 20644 6024 20700
rect 6024 20644 6028 20700
rect 5964 20640 6028 20644
rect 6044 20700 6108 20704
rect 6044 20644 6048 20700
rect 6048 20644 6104 20700
rect 6104 20644 6108 20700
rect 6044 20640 6108 20644
rect 6124 20700 6188 20704
rect 6124 20644 6128 20700
rect 6128 20644 6184 20700
rect 6184 20644 6188 20700
rect 6124 20640 6188 20644
rect 86476 20700 86540 20704
rect 86476 20644 86480 20700
rect 86480 20644 86536 20700
rect 86536 20644 86540 20700
rect 86476 20640 86540 20644
rect 86556 20700 86620 20704
rect 86556 20644 86560 20700
rect 86560 20644 86616 20700
rect 86616 20644 86620 20700
rect 86556 20640 86620 20644
rect 86636 20700 86700 20704
rect 86636 20644 86640 20700
rect 86640 20644 86696 20700
rect 86696 20644 86700 20700
rect 86636 20640 86700 20644
rect 86716 20700 86780 20704
rect 86716 20644 86720 20700
rect 86720 20644 86776 20700
rect 86776 20644 86780 20700
rect 86716 20640 86780 20644
rect 6620 20156 6684 20160
rect 6620 20100 6624 20156
rect 6624 20100 6680 20156
rect 6680 20100 6684 20156
rect 6620 20096 6684 20100
rect 6700 20156 6764 20160
rect 6700 20100 6704 20156
rect 6704 20100 6760 20156
rect 6760 20100 6764 20156
rect 6700 20096 6764 20100
rect 6780 20156 6844 20160
rect 6780 20100 6784 20156
rect 6784 20100 6840 20156
rect 6840 20100 6844 20156
rect 6780 20096 6844 20100
rect 6860 20156 6924 20160
rect 6860 20100 6864 20156
rect 6864 20100 6920 20156
rect 6920 20100 6924 20156
rect 6860 20096 6924 20100
rect 87212 20156 87276 20160
rect 87212 20100 87216 20156
rect 87216 20100 87272 20156
rect 87272 20100 87276 20156
rect 87212 20096 87276 20100
rect 87292 20156 87356 20160
rect 87292 20100 87296 20156
rect 87296 20100 87352 20156
rect 87352 20100 87356 20156
rect 87292 20096 87356 20100
rect 87372 20156 87436 20160
rect 87372 20100 87376 20156
rect 87376 20100 87432 20156
rect 87432 20100 87436 20156
rect 87372 20096 87436 20100
rect 87452 20156 87516 20160
rect 87452 20100 87456 20156
rect 87456 20100 87512 20156
rect 87512 20100 87516 20156
rect 87452 20096 87516 20100
rect 5884 19612 5948 19616
rect 5884 19556 5888 19612
rect 5888 19556 5944 19612
rect 5944 19556 5948 19612
rect 5884 19552 5948 19556
rect 5964 19612 6028 19616
rect 5964 19556 5968 19612
rect 5968 19556 6024 19612
rect 6024 19556 6028 19612
rect 5964 19552 6028 19556
rect 6044 19612 6108 19616
rect 6044 19556 6048 19612
rect 6048 19556 6104 19612
rect 6104 19556 6108 19612
rect 6044 19552 6108 19556
rect 6124 19612 6188 19616
rect 6124 19556 6128 19612
rect 6128 19556 6184 19612
rect 6184 19556 6188 19612
rect 6124 19552 6188 19556
rect 86476 19612 86540 19616
rect 86476 19556 86480 19612
rect 86480 19556 86536 19612
rect 86536 19556 86540 19612
rect 86476 19552 86540 19556
rect 86556 19612 86620 19616
rect 86556 19556 86560 19612
rect 86560 19556 86616 19612
rect 86616 19556 86620 19612
rect 86556 19552 86620 19556
rect 86636 19612 86700 19616
rect 86636 19556 86640 19612
rect 86640 19556 86696 19612
rect 86696 19556 86700 19612
rect 86636 19552 86700 19556
rect 86716 19612 86780 19616
rect 86716 19556 86720 19612
rect 86720 19556 86776 19612
rect 86776 19556 86780 19612
rect 86716 19552 86780 19556
rect 6620 19068 6684 19072
rect 6620 19012 6624 19068
rect 6624 19012 6680 19068
rect 6680 19012 6684 19068
rect 6620 19008 6684 19012
rect 6700 19068 6764 19072
rect 6700 19012 6704 19068
rect 6704 19012 6760 19068
rect 6760 19012 6764 19068
rect 6700 19008 6764 19012
rect 6780 19068 6844 19072
rect 6780 19012 6784 19068
rect 6784 19012 6840 19068
rect 6840 19012 6844 19068
rect 6780 19008 6844 19012
rect 6860 19068 6924 19072
rect 6860 19012 6864 19068
rect 6864 19012 6920 19068
rect 6920 19012 6924 19068
rect 6860 19008 6924 19012
rect 87212 19068 87276 19072
rect 87212 19012 87216 19068
rect 87216 19012 87272 19068
rect 87272 19012 87276 19068
rect 87212 19008 87276 19012
rect 87292 19068 87356 19072
rect 87292 19012 87296 19068
rect 87296 19012 87352 19068
rect 87352 19012 87356 19068
rect 87292 19008 87356 19012
rect 87372 19068 87436 19072
rect 87372 19012 87376 19068
rect 87376 19012 87432 19068
rect 87432 19012 87436 19068
rect 87372 19008 87436 19012
rect 87452 19068 87516 19072
rect 87452 19012 87456 19068
rect 87456 19012 87512 19068
rect 87512 19012 87516 19068
rect 87452 19008 87516 19012
rect 5884 18524 5948 18528
rect 5884 18468 5888 18524
rect 5888 18468 5944 18524
rect 5944 18468 5948 18524
rect 5884 18464 5948 18468
rect 5964 18524 6028 18528
rect 5964 18468 5968 18524
rect 5968 18468 6024 18524
rect 6024 18468 6028 18524
rect 5964 18464 6028 18468
rect 6044 18524 6108 18528
rect 6044 18468 6048 18524
rect 6048 18468 6104 18524
rect 6104 18468 6108 18524
rect 6044 18464 6108 18468
rect 6124 18524 6188 18528
rect 6124 18468 6128 18524
rect 6128 18468 6184 18524
rect 6184 18468 6188 18524
rect 6124 18464 6188 18468
rect 86476 18524 86540 18528
rect 86476 18468 86480 18524
rect 86480 18468 86536 18524
rect 86536 18468 86540 18524
rect 86476 18464 86540 18468
rect 86556 18524 86620 18528
rect 86556 18468 86560 18524
rect 86560 18468 86616 18524
rect 86616 18468 86620 18524
rect 86556 18464 86620 18468
rect 86636 18524 86700 18528
rect 86636 18468 86640 18524
rect 86640 18468 86696 18524
rect 86696 18468 86700 18524
rect 86636 18464 86700 18468
rect 86716 18524 86780 18528
rect 86716 18468 86720 18524
rect 86720 18468 86776 18524
rect 86776 18468 86780 18524
rect 86716 18464 86780 18468
rect 6620 17980 6684 17984
rect 6620 17924 6624 17980
rect 6624 17924 6680 17980
rect 6680 17924 6684 17980
rect 6620 17920 6684 17924
rect 6700 17980 6764 17984
rect 6700 17924 6704 17980
rect 6704 17924 6760 17980
rect 6760 17924 6764 17980
rect 6700 17920 6764 17924
rect 6780 17980 6844 17984
rect 6780 17924 6784 17980
rect 6784 17924 6840 17980
rect 6840 17924 6844 17980
rect 6780 17920 6844 17924
rect 6860 17980 6924 17984
rect 6860 17924 6864 17980
rect 6864 17924 6920 17980
rect 6920 17924 6924 17980
rect 6860 17920 6924 17924
rect 87212 17980 87276 17984
rect 87212 17924 87216 17980
rect 87216 17924 87272 17980
rect 87272 17924 87276 17980
rect 87212 17920 87276 17924
rect 87292 17980 87356 17984
rect 87292 17924 87296 17980
rect 87296 17924 87352 17980
rect 87352 17924 87356 17980
rect 87292 17920 87356 17924
rect 87372 17980 87436 17984
rect 87372 17924 87376 17980
rect 87376 17924 87432 17980
rect 87432 17924 87436 17980
rect 87372 17920 87436 17924
rect 87452 17980 87516 17984
rect 87452 17924 87456 17980
rect 87456 17924 87512 17980
rect 87512 17924 87516 17980
rect 87452 17920 87516 17924
rect 5884 17436 5948 17440
rect 5884 17380 5888 17436
rect 5888 17380 5944 17436
rect 5944 17380 5948 17436
rect 5884 17376 5948 17380
rect 5964 17436 6028 17440
rect 5964 17380 5968 17436
rect 5968 17380 6024 17436
rect 6024 17380 6028 17436
rect 5964 17376 6028 17380
rect 6044 17436 6108 17440
rect 6044 17380 6048 17436
rect 6048 17380 6104 17436
rect 6104 17380 6108 17436
rect 6044 17376 6108 17380
rect 6124 17436 6188 17440
rect 6124 17380 6128 17436
rect 6128 17380 6184 17436
rect 6184 17380 6188 17436
rect 6124 17376 6188 17380
rect 86476 17436 86540 17440
rect 86476 17380 86480 17436
rect 86480 17380 86536 17436
rect 86536 17380 86540 17436
rect 86476 17376 86540 17380
rect 86556 17436 86620 17440
rect 86556 17380 86560 17436
rect 86560 17380 86616 17436
rect 86616 17380 86620 17436
rect 86556 17376 86620 17380
rect 86636 17436 86700 17440
rect 86636 17380 86640 17436
rect 86640 17380 86696 17436
rect 86696 17380 86700 17436
rect 86636 17376 86700 17380
rect 86716 17436 86780 17440
rect 86716 17380 86720 17436
rect 86720 17380 86776 17436
rect 86776 17380 86780 17436
rect 86716 17376 86780 17380
rect 6620 16892 6684 16896
rect 6620 16836 6624 16892
rect 6624 16836 6680 16892
rect 6680 16836 6684 16892
rect 6620 16832 6684 16836
rect 6700 16892 6764 16896
rect 6700 16836 6704 16892
rect 6704 16836 6760 16892
rect 6760 16836 6764 16892
rect 6700 16832 6764 16836
rect 6780 16892 6844 16896
rect 6780 16836 6784 16892
rect 6784 16836 6840 16892
rect 6840 16836 6844 16892
rect 6780 16832 6844 16836
rect 6860 16892 6924 16896
rect 6860 16836 6864 16892
rect 6864 16836 6920 16892
rect 6920 16836 6924 16892
rect 6860 16832 6924 16836
rect 87212 16892 87276 16896
rect 87212 16836 87216 16892
rect 87216 16836 87272 16892
rect 87272 16836 87276 16892
rect 87212 16832 87276 16836
rect 87292 16892 87356 16896
rect 87292 16836 87296 16892
rect 87296 16836 87352 16892
rect 87352 16836 87356 16892
rect 87292 16832 87356 16836
rect 87372 16892 87436 16896
rect 87372 16836 87376 16892
rect 87376 16836 87432 16892
rect 87432 16836 87436 16892
rect 87372 16832 87436 16836
rect 87452 16892 87516 16896
rect 87452 16836 87456 16892
rect 87456 16836 87512 16892
rect 87512 16836 87516 16892
rect 87452 16832 87516 16836
rect 5884 16348 5948 16352
rect 5884 16292 5888 16348
rect 5888 16292 5944 16348
rect 5944 16292 5948 16348
rect 5884 16288 5948 16292
rect 5964 16348 6028 16352
rect 5964 16292 5968 16348
rect 5968 16292 6024 16348
rect 6024 16292 6028 16348
rect 5964 16288 6028 16292
rect 6044 16348 6108 16352
rect 6044 16292 6048 16348
rect 6048 16292 6104 16348
rect 6104 16292 6108 16348
rect 6044 16288 6108 16292
rect 6124 16348 6188 16352
rect 6124 16292 6128 16348
rect 6128 16292 6184 16348
rect 6184 16292 6188 16348
rect 6124 16288 6188 16292
rect 86476 16348 86540 16352
rect 86476 16292 86480 16348
rect 86480 16292 86536 16348
rect 86536 16292 86540 16348
rect 86476 16288 86540 16292
rect 86556 16348 86620 16352
rect 86556 16292 86560 16348
rect 86560 16292 86616 16348
rect 86616 16292 86620 16348
rect 86556 16288 86620 16292
rect 86636 16348 86700 16352
rect 86636 16292 86640 16348
rect 86640 16292 86696 16348
rect 86696 16292 86700 16348
rect 86636 16288 86700 16292
rect 86716 16348 86780 16352
rect 86716 16292 86720 16348
rect 86720 16292 86776 16348
rect 86776 16292 86780 16348
rect 86716 16288 86780 16292
rect 6620 15804 6684 15808
rect 6620 15748 6624 15804
rect 6624 15748 6680 15804
rect 6680 15748 6684 15804
rect 6620 15744 6684 15748
rect 6700 15804 6764 15808
rect 6700 15748 6704 15804
rect 6704 15748 6760 15804
rect 6760 15748 6764 15804
rect 6700 15744 6764 15748
rect 6780 15804 6844 15808
rect 6780 15748 6784 15804
rect 6784 15748 6840 15804
rect 6840 15748 6844 15804
rect 6780 15744 6844 15748
rect 6860 15804 6924 15808
rect 6860 15748 6864 15804
rect 6864 15748 6920 15804
rect 6920 15748 6924 15804
rect 6860 15744 6924 15748
rect 87212 15804 87276 15808
rect 87212 15748 87216 15804
rect 87216 15748 87272 15804
rect 87272 15748 87276 15804
rect 87212 15744 87276 15748
rect 87292 15804 87356 15808
rect 87292 15748 87296 15804
rect 87296 15748 87352 15804
rect 87352 15748 87356 15804
rect 87292 15744 87356 15748
rect 87372 15804 87436 15808
rect 87372 15748 87376 15804
rect 87376 15748 87432 15804
rect 87432 15748 87436 15804
rect 87372 15744 87436 15748
rect 87452 15804 87516 15808
rect 87452 15748 87456 15804
rect 87456 15748 87512 15804
rect 87512 15748 87516 15804
rect 87452 15744 87516 15748
rect 5884 15260 5948 15264
rect 5884 15204 5888 15260
rect 5888 15204 5944 15260
rect 5944 15204 5948 15260
rect 5884 15200 5948 15204
rect 5964 15260 6028 15264
rect 5964 15204 5968 15260
rect 5968 15204 6024 15260
rect 6024 15204 6028 15260
rect 5964 15200 6028 15204
rect 6044 15260 6108 15264
rect 6044 15204 6048 15260
rect 6048 15204 6104 15260
rect 6104 15204 6108 15260
rect 6044 15200 6108 15204
rect 6124 15260 6188 15264
rect 6124 15204 6128 15260
rect 6128 15204 6184 15260
rect 6184 15204 6188 15260
rect 6124 15200 6188 15204
rect 86476 15260 86540 15264
rect 86476 15204 86480 15260
rect 86480 15204 86536 15260
rect 86536 15204 86540 15260
rect 86476 15200 86540 15204
rect 86556 15260 86620 15264
rect 86556 15204 86560 15260
rect 86560 15204 86616 15260
rect 86616 15204 86620 15260
rect 86556 15200 86620 15204
rect 86636 15260 86700 15264
rect 86636 15204 86640 15260
rect 86640 15204 86696 15260
rect 86696 15204 86700 15260
rect 86636 15200 86700 15204
rect 86716 15260 86780 15264
rect 86716 15204 86720 15260
rect 86720 15204 86776 15260
rect 86776 15204 86780 15260
rect 86716 15200 86780 15204
rect 6620 14716 6684 14720
rect 6620 14660 6624 14716
rect 6624 14660 6680 14716
rect 6680 14660 6684 14716
rect 6620 14656 6684 14660
rect 6700 14716 6764 14720
rect 6700 14660 6704 14716
rect 6704 14660 6760 14716
rect 6760 14660 6764 14716
rect 6700 14656 6764 14660
rect 6780 14716 6844 14720
rect 6780 14660 6784 14716
rect 6784 14660 6840 14716
rect 6840 14660 6844 14716
rect 6780 14656 6844 14660
rect 6860 14716 6924 14720
rect 6860 14660 6864 14716
rect 6864 14660 6920 14716
rect 6920 14660 6924 14716
rect 6860 14656 6924 14660
rect 87212 14716 87276 14720
rect 87212 14660 87216 14716
rect 87216 14660 87272 14716
rect 87272 14660 87276 14716
rect 87212 14656 87276 14660
rect 87292 14716 87356 14720
rect 87292 14660 87296 14716
rect 87296 14660 87352 14716
rect 87352 14660 87356 14716
rect 87292 14656 87356 14660
rect 87372 14716 87436 14720
rect 87372 14660 87376 14716
rect 87376 14660 87432 14716
rect 87432 14660 87436 14716
rect 87372 14656 87436 14660
rect 87452 14716 87516 14720
rect 87452 14660 87456 14716
rect 87456 14660 87512 14716
rect 87512 14660 87516 14716
rect 87452 14656 87516 14660
rect 5884 14172 5948 14176
rect 5884 14116 5888 14172
rect 5888 14116 5944 14172
rect 5944 14116 5948 14172
rect 5884 14112 5948 14116
rect 5964 14172 6028 14176
rect 5964 14116 5968 14172
rect 5968 14116 6024 14172
rect 6024 14116 6028 14172
rect 5964 14112 6028 14116
rect 6044 14172 6108 14176
rect 6044 14116 6048 14172
rect 6048 14116 6104 14172
rect 6104 14116 6108 14172
rect 6044 14112 6108 14116
rect 6124 14172 6188 14176
rect 6124 14116 6128 14172
rect 6128 14116 6184 14172
rect 6184 14116 6188 14172
rect 6124 14112 6188 14116
rect 86476 14172 86540 14176
rect 86476 14116 86480 14172
rect 86480 14116 86536 14172
rect 86536 14116 86540 14172
rect 86476 14112 86540 14116
rect 86556 14172 86620 14176
rect 86556 14116 86560 14172
rect 86560 14116 86616 14172
rect 86616 14116 86620 14172
rect 86556 14112 86620 14116
rect 86636 14172 86700 14176
rect 86636 14116 86640 14172
rect 86640 14116 86696 14172
rect 86696 14116 86700 14172
rect 86636 14112 86700 14116
rect 86716 14172 86780 14176
rect 86716 14116 86720 14172
rect 86720 14116 86776 14172
rect 86776 14116 86780 14172
rect 86716 14112 86780 14116
rect 6620 13628 6684 13632
rect 6620 13572 6624 13628
rect 6624 13572 6680 13628
rect 6680 13572 6684 13628
rect 6620 13568 6684 13572
rect 6700 13628 6764 13632
rect 6700 13572 6704 13628
rect 6704 13572 6760 13628
rect 6760 13572 6764 13628
rect 6700 13568 6764 13572
rect 6780 13628 6844 13632
rect 6780 13572 6784 13628
rect 6784 13572 6840 13628
rect 6840 13572 6844 13628
rect 6780 13568 6844 13572
rect 6860 13628 6924 13632
rect 6860 13572 6864 13628
rect 6864 13572 6920 13628
rect 6920 13572 6924 13628
rect 6860 13568 6924 13572
rect 87212 13628 87276 13632
rect 87212 13572 87216 13628
rect 87216 13572 87272 13628
rect 87272 13572 87276 13628
rect 87212 13568 87276 13572
rect 87292 13628 87356 13632
rect 87292 13572 87296 13628
rect 87296 13572 87352 13628
rect 87352 13572 87356 13628
rect 87292 13568 87356 13572
rect 87372 13628 87436 13632
rect 87372 13572 87376 13628
rect 87376 13572 87432 13628
rect 87432 13572 87436 13628
rect 87372 13568 87436 13572
rect 87452 13628 87516 13632
rect 87452 13572 87456 13628
rect 87456 13572 87512 13628
rect 87512 13572 87516 13628
rect 87452 13568 87516 13572
rect 5884 13084 5948 13088
rect 5884 13028 5888 13084
rect 5888 13028 5944 13084
rect 5944 13028 5948 13084
rect 5884 13024 5948 13028
rect 5964 13084 6028 13088
rect 5964 13028 5968 13084
rect 5968 13028 6024 13084
rect 6024 13028 6028 13084
rect 5964 13024 6028 13028
rect 6044 13084 6108 13088
rect 6044 13028 6048 13084
rect 6048 13028 6104 13084
rect 6104 13028 6108 13084
rect 6044 13024 6108 13028
rect 6124 13084 6188 13088
rect 6124 13028 6128 13084
rect 6128 13028 6184 13084
rect 6184 13028 6188 13084
rect 6124 13024 6188 13028
rect 86476 13084 86540 13088
rect 86476 13028 86480 13084
rect 86480 13028 86536 13084
rect 86536 13028 86540 13084
rect 86476 13024 86540 13028
rect 86556 13084 86620 13088
rect 86556 13028 86560 13084
rect 86560 13028 86616 13084
rect 86616 13028 86620 13084
rect 86556 13024 86620 13028
rect 86636 13084 86700 13088
rect 86636 13028 86640 13084
rect 86640 13028 86696 13084
rect 86696 13028 86700 13084
rect 86636 13024 86700 13028
rect 86716 13084 86780 13088
rect 86716 13028 86720 13084
rect 86720 13028 86776 13084
rect 86776 13028 86780 13084
rect 86716 13024 86780 13028
rect 6620 12540 6684 12544
rect 6620 12484 6624 12540
rect 6624 12484 6680 12540
rect 6680 12484 6684 12540
rect 6620 12480 6684 12484
rect 6700 12540 6764 12544
rect 6700 12484 6704 12540
rect 6704 12484 6760 12540
rect 6760 12484 6764 12540
rect 6700 12480 6764 12484
rect 6780 12540 6844 12544
rect 6780 12484 6784 12540
rect 6784 12484 6840 12540
rect 6840 12484 6844 12540
rect 6780 12480 6844 12484
rect 6860 12540 6924 12544
rect 6860 12484 6864 12540
rect 6864 12484 6920 12540
rect 6920 12484 6924 12540
rect 6860 12480 6924 12484
rect 87212 12540 87276 12544
rect 87212 12484 87216 12540
rect 87216 12484 87272 12540
rect 87272 12484 87276 12540
rect 87212 12480 87276 12484
rect 87292 12540 87356 12544
rect 87292 12484 87296 12540
rect 87296 12484 87352 12540
rect 87352 12484 87356 12540
rect 87292 12480 87356 12484
rect 87372 12540 87436 12544
rect 87372 12484 87376 12540
rect 87376 12484 87432 12540
rect 87432 12484 87436 12540
rect 87372 12480 87436 12484
rect 87452 12540 87516 12544
rect 87452 12484 87456 12540
rect 87456 12484 87512 12540
rect 87512 12484 87516 12540
rect 87452 12480 87516 12484
rect 5884 11996 5948 12000
rect 5884 11940 5888 11996
rect 5888 11940 5944 11996
rect 5944 11940 5948 11996
rect 5884 11936 5948 11940
rect 5964 11996 6028 12000
rect 5964 11940 5968 11996
rect 5968 11940 6024 11996
rect 6024 11940 6028 11996
rect 5964 11936 6028 11940
rect 6044 11996 6108 12000
rect 6044 11940 6048 11996
rect 6048 11940 6104 11996
rect 6104 11940 6108 11996
rect 6044 11936 6108 11940
rect 6124 11996 6188 12000
rect 6124 11940 6128 11996
rect 6128 11940 6184 11996
rect 6184 11940 6188 11996
rect 6124 11936 6188 11940
rect 86476 11996 86540 12000
rect 86476 11940 86480 11996
rect 86480 11940 86536 11996
rect 86536 11940 86540 11996
rect 86476 11936 86540 11940
rect 86556 11996 86620 12000
rect 86556 11940 86560 11996
rect 86560 11940 86616 11996
rect 86616 11940 86620 11996
rect 86556 11936 86620 11940
rect 86636 11996 86700 12000
rect 86636 11940 86640 11996
rect 86640 11940 86696 11996
rect 86696 11940 86700 11996
rect 86636 11936 86700 11940
rect 86716 11996 86780 12000
rect 86716 11940 86720 11996
rect 86720 11940 86776 11996
rect 86776 11940 86780 11996
rect 86716 11936 86780 11940
rect 6620 11452 6684 11456
rect 6620 11396 6624 11452
rect 6624 11396 6680 11452
rect 6680 11396 6684 11452
rect 6620 11392 6684 11396
rect 6700 11452 6764 11456
rect 6700 11396 6704 11452
rect 6704 11396 6760 11452
rect 6760 11396 6764 11452
rect 6700 11392 6764 11396
rect 6780 11452 6844 11456
rect 6780 11396 6784 11452
rect 6784 11396 6840 11452
rect 6840 11396 6844 11452
rect 6780 11392 6844 11396
rect 6860 11452 6924 11456
rect 6860 11396 6864 11452
rect 6864 11396 6920 11452
rect 6920 11396 6924 11452
rect 6860 11392 6924 11396
rect 87212 11452 87276 11456
rect 87212 11396 87216 11452
rect 87216 11396 87272 11452
rect 87272 11396 87276 11452
rect 87212 11392 87276 11396
rect 87292 11452 87356 11456
rect 87292 11396 87296 11452
rect 87296 11396 87352 11452
rect 87352 11396 87356 11452
rect 87292 11392 87356 11396
rect 87372 11452 87436 11456
rect 87372 11396 87376 11452
rect 87376 11396 87432 11452
rect 87432 11396 87436 11452
rect 87372 11392 87436 11396
rect 87452 11452 87516 11456
rect 87452 11396 87456 11452
rect 87456 11396 87512 11452
rect 87512 11396 87516 11452
rect 87452 11392 87516 11396
rect 5884 10908 5948 10912
rect 5884 10852 5888 10908
rect 5888 10852 5944 10908
rect 5944 10852 5948 10908
rect 5884 10848 5948 10852
rect 5964 10908 6028 10912
rect 5964 10852 5968 10908
rect 5968 10852 6024 10908
rect 6024 10852 6028 10908
rect 5964 10848 6028 10852
rect 6044 10908 6108 10912
rect 6044 10852 6048 10908
rect 6048 10852 6104 10908
rect 6104 10852 6108 10908
rect 6044 10848 6108 10852
rect 6124 10908 6188 10912
rect 6124 10852 6128 10908
rect 6128 10852 6184 10908
rect 6184 10852 6188 10908
rect 6124 10848 6188 10852
rect 86476 10908 86540 10912
rect 86476 10852 86480 10908
rect 86480 10852 86536 10908
rect 86536 10852 86540 10908
rect 86476 10848 86540 10852
rect 86556 10908 86620 10912
rect 86556 10852 86560 10908
rect 86560 10852 86616 10908
rect 86616 10852 86620 10908
rect 86556 10848 86620 10852
rect 86636 10908 86700 10912
rect 86636 10852 86640 10908
rect 86640 10852 86696 10908
rect 86696 10852 86700 10908
rect 86636 10848 86700 10852
rect 86716 10908 86780 10912
rect 86716 10852 86720 10908
rect 86720 10852 86776 10908
rect 86776 10852 86780 10908
rect 86716 10848 86780 10852
rect 6620 10364 6684 10368
rect 6620 10308 6624 10364
rect 6624 10308 6680 10364
rect 6680 10308 6684 10364
rect 6620 10304 6684 10308
rect 6700 10364 6764 10368
rect 6700 10308 6704 10364
rect 6704 10308 6760 10364
rect 6760 10308 6764 10364
rect 6700 10304 6764 10308
rect 6780 10364 6844 10368
rect 6780 10308 6784 10364
rect 6784 10308 6840 10364
rect 6840 10308 6844 10364
rect 6780 10304 6844 10308
rect 6860 10364 6924 10368
rect 6860 10308 6864 10364
rect 6864 10308 6920 10364
rect 6920 10308 6924 10364
rect 6860 10304 6924 10308
rect 87212 10364 87276 10368
rect 87212 10308 87216 10364
rect 87216 10308 87272 10364
rect 87272 10308 87276 10364
rect 87212 10304 87276 10308
rect 87292 10364 87356 10368
rect 87292 10308 87296 10364
rect 87296 10308 87352 10364
rect 87352 10308 87356 10364
rect 87292 10304 87356 10308
rect 87372 10364 87436 10368
rect 87372 10308 87376 10364
rect 87376 10308 87432 10364
rect 87432 10308 87436 10364
rect 87372 10304 87436 10308
rect 87452 10364 87516 10368
rect 87452 10308 87456 10364
rect 87456 10308 87512 10364
rect 87512 10308 87516 10364
rect 87452 10304 87516 10308
rect 5884 9820 5948 9824
rect 5884 9764 5888 9820
rect 5888 9764 5944 9820
rect 5944 9764 5948 9820
rect 5884 9760 5948 9764
rect 5964 9820 6028 9824
rect 5964 9764 5968 9820
rect 5968 9764 6024 9820
rect 6024 9764 6028 9820
rect 5964 9760 6028 9764
rect 6044 9820 6108 9824
rect 6044 9764 6048 9820
rect 6048 9764 6104 9820
rect 6104 9764 6108 9820
rect 6044 9760 6108 9764
rect 6124 9820 6188 9824
rect 6124 9764 6128 9820
rect 6128 9764 6184 9820
rect 6184 9764 6188 9820
rect 6124 9760 6188 9764
rect 86476 9820 86540 9824
rect 86476 9764 86480 9820
rect 86480 9764 86536 9820
rect 86536 9764 86540 9820
rect 86476 9760 86540 9764
rect 86556 9820 86620 9824
rect 86556 9764 86560 9820
rect 86560 9764 86616 9820
rect 86616 9764 86620 9820
rect 86556 9760 86620 9764
rect 86636 9820 86700 9824
rect 86636 9764 86640 9820
rect 86640 9764 86696 9820
rect 86696 9764 86700 9820
rect 86636 9760 86700 9764
rect 86716 9820 86780 9824
rect 86716 9764 86720 9820
rect 86720 9764 86776 9820
rect 86776 9764 86780 9820
rect 86716 9760 86780 9764
rect 6620 9276 6684 9280
rect 6620 9220 6624 9276
rect 6624 9220 6680 9276
rect 6680 9220 6684 9276
rect 6620 9216 6684 9220
rect 6700 9276 6764 9280
rect 6700 9220 6704 9276
rect 6704 9220 6760 9276
rect 6760 9220 6764 9276
rect 6700 9216 6764 9220
rect 6780 9276 6844 9280
rect 6780 9220 6784 9276
rect 6784 9220 6840 9276
rect 6840 9220 6844 9276
rect 6780 9216 6844 9220
rect 6860 9276 6924 9280
rect 6860 9220 6864 9276
rect 6864 9220 6920 9276
rect 6920 9220 6924 9276
rect 6860 9216 6924 9220
rect 87212 9276 87276 9280
rect 87212 9220 87216 9276
rect 87216 9220 87272 9276
rect 87272 9220 87276 9276
rect 87212 9216 87276 9220
rect 87292 9276 87356 9280
rect 87292 9220 87296 9276
rect 87296 9220 87352 9276
rect 87352 9220 87356 9276
rect 87292 9216 87356 9220
rect 87372 9276 87436 9280
rect 87372 9220 87376 9276
rect 87376 9220 87432 9276
rect 87432 9220 87436 9276
rect 87372 9216 87436 9220
rect 87452 9276 87516 9280
rect 87452 9220 87456 9276
rect 87456 9220 87512 9276
rect 87512 9220 87516 9276
rect 87452 9216 87516 9220
rect 5884 8732 5948 8736
rect 5884 8676 5888 8732
rect 5888 8676 5944 8732
rect 5944 8676 5948 8732
rect 5884 8672 5948 8676
rect 5964 8732 6028 8736
rect 5964 8676 5968 8732
rect 5968 8676 6024 8732
rect 6024 8676 6028 8732
rect 5964 8672 6028 8676
rect 6044 8732 6108 8736
rect 6044 8676 6048 8732
rect 6048 8676 6104 8732
rect 6104 8676 6108 8732
rect 6044 8672 6108 8676
rect 6124 8732 6188 8736
rect 6124 8676 6128 8732
rect 6128 8676 6184 8732
rect 6184 8676 6188 8732
rect 6124 8672 6188 8676
rect 86476 8732 86540 8736
rect 86476 8676 86480 8732
rect 86480 8676 86536 8732
rect 86536 8676 86540 8732
rect 86476 8672 86540 8676
rect 86556 8732 86620 8736
rect 86556 8676 86560 8732
rect 86560 8676 86616 8732
rect 86616 8676 86620 8732
rect 86556 8672 86620 8676
rect 86636 8732 86700 8736
rect 86636 8676 86640 8732
rect 86640 8676 86696 8732
rect 86696 8676 86700 8732
rect 86636 8672 86700 8676
rect 86716 8732 86780 8736
rect 86716 8676 86720 8732
rect 86720 8676 86776 8732
rect 86776 8676 86780 8732
rect 86716 8672 86780 8676
rect 6620 8188 6684 8192
rect 6620 8132 6624 8188
rect 6624 8132 6680 8188
rect 6680 8132 6684 8188
rect 6620 8128 6684 8132
rect 6700 8188 6764 8192
rect 6700 8132 6704 8188
rect 6704 8132 6760 8188
rect 6760 8132 6764 8188
rect 6700 8128 6764 8132
rect 6780 8188 6844 8192
rect 6780 8132 6784 8188
rect 6784 8132 6840 8188
rect 6840 8132 6844 8188
rect 6780 8128 6844 8132
rect 6860 8188 6924 8192
rect 6860 8132 6864 8188
rect 6864 8132 6920 8188
rect 6920 8132 6924 8188
rect 6860 8128 6924 8132
rect 87212 8188 87276 8192
rect 87212 8132 87216 8188
rect 87216 8132 87272 8188
rect 87272 8132 87276 8188
rect 87212 8128 87276 8132
rect 87292 8188 87356 8192
rect 87292 8132 87296 8188
rect 87296 8132 87352 8188
rect 87352 8132 87356 8188
rect 87292 8128 87356 8132
rect 87372 8188 87436 8192
rect 87372 8132 87376 8188
rect 87376 8132 87432 8188
rect 87432 8132 87436 8188
rect 87372 8128 87436 8132
rect 87452 8188 87516 8192
rect 87452 8132 87456 8188
rect 87456 8132 87512 8188
rect 87512 8132 87516 8188
rect 87452 8128 87516 8132
rect 5884 7644 5948 7648
rect 5884 7588 5888 7644
rect 5888 7588 5944 7644
rect 5944 7588 5948 7644
rect 5884 7584 5948 7588
rect 5964 7644 6028 7648
rect 5964 7588 5968 7644
rect 5968 7588 6024 7644
rect 6024 7588 6028 7644
rect 5964 7584 6028 7588
rect 6044 7644 6108 7648
rect 6044 7588 6048 7644
rect 6048 7588 6104 7644
rect 6104 7588 6108 7644
rect 6044 7584 6108 7588
rect 6124 7644 6188 7648
rect 6124 7588 6128 7644
rect 6128 7588 6184 7644
rect 6184 7588 6188 7644
rect 6124 7584 6188 7588
rect 17724 7644 17788 7648
rect 17724 7588 17728 7644
rect 17728 7588 17784 7644
rect 17784 7588 17788 7644
rect 17724 7584 17788 7588
rect 17804 7644 17868 7648
rect 17804 7588 17808 7644
rect 17808 7588 17864 7644
rect 17864 7588 17868 7644
rect 17804 7584 17868 7588
rect 17884 7644 17948 7648
rect 17884 7588 17888 7644
rect 17888 7588 17944 7644
rect 17944 7588 17948 7644
rect 17884 7584 17948 7588
rect 17964 7644 18028 7648
rect 17964 7588 17968 7644
rect 17968 7588 18024 7644
rect 18024 7588 18028 7644
rect 17964 7584 18028 7588
rect 36124 7644 36188 7648
rect 36124 7588 36128 7644
rect 36128 7588 36184 7644
rect 36184 7588 36188 7644
rect 36124 7584 36188 7588
rect 36204 7644 36268 7648
rect 36204 7588 36208 7644
rect 36208 7588 36264 7644
rect 36264 7588 36268 7644
rect 36204 7584 36268 7588
rect 36284 7644 36348 7648
rect 36284 7588 36288 7644
rect 36288 7588 36344 7644
rect 36344 7588 36348 7644
rect 36284 7584 36348 7588
rect 36364 7644 36428 7648
rect 36364 7588 36368 7644
rect 36368 7588 36424 7644
rect 36424 7588 36428 7644
rect 36364 7584 36428 7588
rect 54524 7644 54588 7648
rect 54524 7588 54528 7644
rect 54528 7588 54584 7644
rect 54584 7588 54588 7644
rect 54524 7584 54588 7588
rect 54604 7644 54668 7648
rect 54604 7588 54608 7644
rect 54608 7588 54664 7644
rect 54664 7588 54668 7644
rect 54604 7584 54668 7588
rect 54684 7644 54748 7648
rect 54684 7588 54688 7644
rect 54688 7588 54744 7644
rect 54744 7588 54748 7644
rect 54684 7584 54748 7588
rect 54764 7644 54828 7648
rect 54764 7588 54768 7644
rect 54768 7588 54824 7644
rect 54824 7588 54828 7644
rect 54764 7584 54828 7588
rect 72924 7644 72988 7648
rect 72924 7588 72928 7644
rect 72928 7588 72984 7644
rect 72984 7588 72988 7644
rect 72924 7584 72988 7588
rect 73004 7644 73068 7648
rect 73004 7588 73008 7644
rect 73008 7588 73064 7644
rect 73064 7588 73068 7644
rect 73004 7584 73068 7588
rect 73084 7644 73148 7648
rect 73084 7588 73088 7644
rect 73088 7588 73144 7644
rect 73144 7588 73148 7644
rect 73084 7584 73148 7588
rect 73164 7644 73228 7648
rect 73164 7588 73168 7644
rect 73168 7588 73224 7644
rect 73224 7588 73228 7644
rect 73164 7584 73228 7588
rect 86476 7644 86540 7648
rect 86476 7588 86480 7644
rect 86480 7588 86536 7644
rect 86536 7588 86540 7644
rect 86476 7584 86540 7588
rect 86556 7644 86620 7648
rect 86556 7588 86560 7644
rect 86560 7588 86616 7644
rect 86616 7588 86620 7644
rect 86556 7584 86620 7588
rect 86636 7644 86700 7648
rect 86636 7588 86640 7644
rect 86640 7588 86696 7644
rect 86696 7588 86700 7644
rect 86636 7584 86700 7588
rect 86716 7644 86780 7648
rect 86716 7588 86720 7644
rect 86720 7588 86776 7644
rect 86776 7588 86780 7644
rect 86716 7584 86780 7588
rect 6620 7100 6684 7104
rect 6620 7044 6624 7100
rect 6624 7044 6680 7100
rect 6680 7044 6684 7100
rect 6620 7040 6684 7044
rect 6700 7100 6764 7104
rect 6700 7044 6704 7100
rect 6704 7044 6760 7100
rect 6760 7044 6764 7100
rect 6700 7040 6764 7044
rect 6780 7100 6844 7104
rect 6780 7044 6784 7100
rect 6784 7044 6840 7100
rect 6840 7044 6844 7100
rect 6780 7040 6844 7044
rect 6860 7100 6924 7104
rect 6860 7044 6864 7100
rect 6864 7044 6920 7100
rect 6920 7044 6924 7100
rect 6860 7040 6924 7044
rect 18384 7100 18448 7104
rect 18384 7044 18388 7100
rect 18388 7044 18444 7100
rect 18444 7044 18448 7100
rect 18384 7040 18448 7044
rect 18464 7100 18528 7104
rect 18464 7044 18468 7100
rect 18468 7044 18524 7100
rect 18524 7044 18528 7100
rect 18464 7040 18528 7044
rect 18544 7100 18608 7104
rect 18544 7044 18548 7100
rect 18548 7044 18604 7100
rect 18604 7044 18608 7100
rect 18544 7040 18608 7044
rect 18624 7100 18688 7104
rect 18624 7044 18628 7100
rect 18628 7044 18684 7100
rect 18684 7044 18688 7100
rect 18624 7040 18688 7044
rect 36784 7100 36848 7104
rect 36784 7044 36788 7100
rect 36788 7044 36844 7100
rect 36844 7044 36848 7100
rect 36784 7040 36848 7044
rect 36864 7100 36928 7104
rect 36864 7044 36868 7100
rect 36868 7044 36924 7100
rect 36924 7044 36928 7100
rect 36864 7040 36928 7044
rect 36944 7100 37008 7104
rect 36944 7044 36948 7100
rect 36948 7044 37004 7100
rect 37004 7044 37008 7100
rect 36944 7040 37008 7044
rect 37024 7100 37088 7104
rect 37024 7044 37028 7100
rect 37028 7044 37084 7100
rect 37084 7044 37088 7100
rect 37024 7040 37088 7044
rect 55184 7100 55248 7104
rect 55184 7044 55188 7100
rect 55188 7044 55244 7100
rect 55244 7044 55248 7100
rect 55184 7040 55248 7044
rect 55264 7100 55328 7104
rect 55264 7044 55268 7100
rect 55268 7044 55324 7100
rect 55324 7044 55328 7100
rect 55264 7040 55328 7044
rect 55344 7100 55408 7104
rect 55344 7044 55348 7100
rect 55348 7044 55404 7100
rect 55404 7044 55408 7100
rect 55344 7040 55408 7044
rect 55424 7100 55488 7104
rect 55424 7044 55428 7100
rect 55428 7044 55484 7100
rect 55484 7044 55488 7100
rect 55424 7040 55488 7044
rect 73584 7100 73648 7104
rect 73584 7044 73588 7100
rect 73588 7044 73644 7100
rect 73644 7044 73648 7100
rect 73584 7040 73648 7044
rect 73664 7100 73728 7104
rect 73664 7044 73668 7100
rect 73668 7044 73724 7100
rect 73724 7044 73728 7100
rect 73664 7040 73728 7044
rect 73744 7100 73808 7104
rect 73744 7044 73748 7100
rect 73748 7044 73804 7100
rect 73804 7044 73808 7100
rect 73744 7040 73808 7044
rect 73824 7100 73888 7104
rect 73824 7044 73828 7100
rect 73828 7044 73884 7100
rect 73884 7044 73888 7100
rect 73824 7040 73888 7044
rect 87212 7100 87276 7104
rect 87212 7044 87216 7100
rect 87216 7044 87272 7100
rect 87272 7044 87276 7100
rect 87212 7040 87276 7044
rect 87292 7100 87356 7104
rect 87292 7044 87296 7100
rect 87296 7044 87352 7100
rect 87352 7044 87356 7100
rect 87292 7040 87356 7044
rect 87372 7100 87436 7104
rect 87372 7044 87376 7100
rect 87376 7044 87432 7100
rect 87432 7044 87436 7100
rect 87372 7040 87436 7044
rect 87452 7100 87516 7104
rect 87452 7044 87456 7100
rect 87456 7044 87512 7100
rect 87512 7044 87516 7100
rect 87452 7040 87516 7044
rect 17724 6556 17788 6560
rect 17724 6500 17728 6556
rect 17728 6500 17784 6556
rect 17784 6500 17788 6556
rect 17724 6496 17788 6500
rect 17804 6556 17868 6560
rect 17804 6500 17808 6556
rect 17808 6500 17864 6556
rect 17864 6500 17868 6556
rect 17804 6496 17868 6500
rect 17884 6556 17948 6560
rect 17884 6500 17888 6556
rect 17888 6500 17944 6556
rect 17944 6500 17948 6556
rect 17884 6496 17948 6500
rect 17964 6556 18028 6560
rect 17964 6500 17968 6556
rect 17968 6500 18024 6556
rect 18024 6500 18028 6556
rect 17964 6496 18028 6500
rect 36124 6556 36188 6560
rect 36124 6500 36128 6556
rect 36128 6500 36184 6556
rect 36184 6500 36188 6556
rect 36124 6496 36188 6500
rect 36204 6556 36268 6560
rect 36204 6500 36208 6556
rect 36208 6500 36264 6556
rect 36264 6500 36268 6556
rect 36204 6496 36268 6500
rect 36284 6556 36348 6560
rect 36284 6500 36288 6556
rect 36288 6500 36344 6556
rect 36344 6500 36348 6556
rect 36284 6496 36348 6500
rect 36364 6556 36428 6560
rect 36364 6500 36368 6556
rect 36368 6500 36424 6556
rect 36424 6500 36428 6556
rect 36364 6496 36428 6500
rect 54524 6556 54588 6560
rect 54524 6500 54528 6556
rect 54528 6500 54584 6556
rect 54584 6500 54588 6556
rect 54524 6496 54588 6500
rect 54604 6556 54668 6560
rect 54604 6500 54608 6556
rect 54608 6500 54664 6556
rect 54664 6500 54668 6556
rect 54604 6496 54668 6500
rect 54684 6556 54748 6560
rect 54684 6500 54688 6556
rect 54688 6500 54744 6556
rect 54744 6500 54748 6556
rect 54684 6496 54748 6500
rect 54764 6556 54828 6560
rect 54764 6500 54768 6556
rect 54768 6500 54824 6556
rect 54824 6500 54828 6556
rect 54764 6496 54828 6500
rect 72924 6556 72988 6560
rect 72924 6500 72928 6556
rect 72928 6500 72984 6556
rect 72984 6500 72988 6556
rect 72924 6496 72988 6500
rect 73004 6556 73068 6560
rect 73004 6500 73008 6556
rect 73008 6500 73064 6556
rect 73064 6500 73068 6556
rect 73004 6496 73068 6500
rect 73084 6556 73148 6560
rect 73084 6500 73088 6556
rect 73088 6500 73144 6556
rect 73144 6500 73148 6556
rect 73084 6496 73148 6500
rect 73164 6556 73228 6560
rect 73164 6500 73168 6556
rect 73168 6500 73224 6556
rect 73224 6500 73228 6556
rect 73164 6496 73228 6500
rect 18384 6012 18448 6016
rect 18384 5956 18388 6012
rect 18388 5956 18444 6012
rect 18444 5956 18448 6012
rect 18384 5952 18448 5956
rect 18464 6012 18528 6016
rect 18464 5956 18468 6012
rect 18468 5956 18524 6012
rect 18524 5956 18528 6012
rect 18464 5952 18528 5956
rect 18544 6012 18608 6016
rect 18544 5956 18548 6012
rect 18548 5956 18604 6012
rect 18604 5956 18608 6012
rect 18544 5952 18608 5956
rect 18624 6012 18688 6016
rect 18624 5956 18628 6012
rect 18628 5956 18684 6012
rect 18684 5956 18688 6012
rect 18624 5952 18688 5956
rect 36784 6012 36848 6016
rect 36784 5956 36788 6012
rect 36788 5956 36844 6012
rect 36844 5956 36848 6012
rect 36784 5952 36848 5956
rect 36864 6012 36928 6016
rect 36864 5956 36868 6012
rect 36868 5956 36924 6012
rect 36924 5956 36928 6012
rect 36864 5952 36928 5956
rect 36944 6012 37008 6016
rect 36944 5956 36948 6012
rect 36948 5956 37004 6012
rect 37004 5956 37008 6012
rect 36944 5952 37008 5956
rect 37024 6012 37088 6016
rect 37024 5956 37028 6012
rect 37028 5956 37084 6012
rect 37084 5956 37088 6012
rect 37024 5952 37088 5956
rect 55184 6012 55248 6016
rect 55184 5956 55188 6012
rect 55188 5956 55244 6012
rect 55244 5956 55248 6012
rect 55184 5952 55248 5956
rect 55264 6012 55328 6016
rect 55264 5956 55268 6012
rect 55268 5956 55324 6012
rect 55324 5956 55328 6012
rect 55264 5952 55328 5956
rect 55344 6012 55408 6016
rect 55344 5956 55348 6012
rect 55348 5956 55404 6012
rect 55404 5956 55408 6012
rect 55344 5952 55408 5956
rect 55424 6012 55488 6016
rect 55424 5956 55428 6012
rect 55428 5956 55484 6012
rect 55484 5956 55488 6012
rect 55424 5952 55488 5956
rect 73584 6012 73648 6016
rect 73584 5956 73588 6012
rect 73588 5956 73644 6012
rect 73644 5956 73648 6012
rect 73584 5952 73648 5956
rect 73664 6012 73728 6016
rect 73664 5956 73668 6012
rect 73668 5956 73724 6012
rect 73724 5956 73728 6012
rect 73664 5952 73728 5956
rect 73744 6012 73808 6016
rect 73744 5956 73748 6012
rect 73748 5956 73804 6012
rect 73804 5956 73808 6012
rect 73744 5952 73808 5956
rect 73824 6012 73888 6016
rect 73824 5956 73828 6012
rect 73828 5956 73884 6012
rect 73884 5956 73888 6012
rect 73824 5952 73888 5956
rect 17724 5468 17788 5472
rect 17724 5412 17728 5468
rect 17728 5412 17784 5468
rect 17784 5412 17788 5468
rect 17724 5408 17788 5412
rect 17804 5468 17868 5472
rect 17804 5412 17808 5468
rect 17808 5412 17864 5468
rect 17864 5412 17868 5468
rect 17804 5408 17868 5412
rect 17884 5468 17948 5472
rect 17884 5412 17888 5468
rect 17888 5412 17944 5468
rect 17944 5412 17948 5468
rect 17884 5408 17948 5412
rect 17964 5468 18028 5472
rect 17964 5412 17968 5468
rect 17968 5412 18024 5468
rect 18024 5412 18028 5468
rect 17964 5408 18028 5412
rect 36124 5468 36188 5472
rect 36124 5412 36128 5468
rect 36128 5412 36184 5468
rect 36184 5412 36188 5468
rect 36124 5408 36188 5412
rect 36204 5468 36268 5472
rect 36204 5412 36208 5468
rect 36208 5412 36264 5468
rect 36264 5412 36268 5468
rect 36204 5408 36268 5412
rect 36284 5468 36348 5472
rect 36284 5412 36288 5468
rect 36288 5412 36344 5468
rect 36344 5412 36348 5468
rect 36284 5408 36348 5412
rect 36364 5468 36428 5472
rect 36364 5412 36368 5468
rect 36368 5412 36424 5468
rect 36424 5412 36428 5468
rect 36364 5408 36428 5412
rect 54524 5468 54588 5472
rect 54524 5412 54528 5468
rect 54528 5412 54584 5468
rect 54584 5412 54588 5468
rect 54524 5408 54588 5412
rect 54604 5468 54668 5472
rect 54604 5412 54608 5468
rect 54608 5412 54664 5468
rect 54664 5412 54668 5468
rect 54604 5408 54668 5412
rect 54684 5468 54748 5472
rect 54684 5412 54688 5468
rect 54688 5412 54744 5468
rect 54744 5412 54748 5468
rect 54684 5408 54748 5412
rect 54764 5468 54828 5472
rect 54764 5412 54768 5468
rect 54768 5412 54824 5468
rect 54824 5412 54828 5468
rect 54764 5408 54828 5412
rect 72924 5468 72988 5472
rect 72924 5412 72928 5468
rect 72928 5412 72984 5468
rect 72984 5412 72988 5468
rect 72924 5408 72988 5412
rect 73004 5468 73068 5472
rect 73004 5412 73008 5468
rect 73008 5412 73064 5468
rect 73064 5412 73068 5468
rect 73004 5408 73068 5412
rect 73084 5468 73148 5472
rect 73084 5412 73088 5468
rect 73088 5412 73144 5468
rect 73144 5412 73148 5468
rect 73084 5408 73148 5412
rect 73164 5468 73228 5472
rect 73164 5412 73168 5468
rect 73168 5412 73224 5468
rect 73224 5412 73228 5468
rect 73164 5408 73228 5412
rect 18384 4924 18448 4928
rect 18384 4868 18388 4924
rect 18388 4868 18444 4924
rect 18444 4868 18448 4924
rect 18384 4864 18448 4868
rect 18464 4924 18528 4928
rect 18464 4868 18468 4924
rect 18468 4868 18524 4924
rect 18524 4868 18528 4924
rect 18464 4864 18528 4868
rect 18544 4924 18608 4928
rect 18544 4868 18548 4924
rect 18548 4868 18604 4924
rect 18604 4868 18608 4924
rect 18544 4864 18608 4868
rect 18624 4924 18688 4928
rect 18624 4868 18628 4924
rect 18628 4868 18684 4924
rect 18684 4868 18688 4924
rect 18624 4864 18688 4868
rect 36784 4924 36848 4928
rect 36784 4868 36788 4924
rect 36788 4868 36844 4924
rect 36844 4868 36848 4924
rect 36784 4864 36848 4868
rect 36864 4924 36928 4928
rect 36864 4868 36868 4924
rect 36868 4868 36924 4924
rect 36924 4868 36928 4924
rect 36864 4864 36928 4868
rect 36944 4924 37008 4928
rect 36944 4868 36948 4924
rect 36948 4868 37004 4924
rect 37004 4868 37008 4924
rect 36944 4864 37008 4868
rect 37024 4924 37088 4928
rect 37024 4868 37028 4924
rect 37028 4868 37084 4924
rect 37084 4868 37088 4924
rect 37024 4864 37088 4868
rect 55184 4924 55248 4928
rect 55184 4868 55188 4924
rect 55188 4868 55244 4924
rect 55244 4868 55248 4924
rect 55184 4864 55248 4868
rect 55264 4924 55328 4928
rect 55264 4868 55268 4924
rect 55268 4868 55324 4924
rect 55324 4868 55328 4924
rect 55264 4864 55328 4868
rect 55344 4924 55408 4928
rect 55344 4868 55348 4924
rect 55348 4868 55404 4924
rect 55404 4868 55408 4924
rect 55344 4864 55408 4868
rect 55424 4924 55488 4928
rect 55424 4868 55428 4924
rect 55428 4868 55484 4924
rect 55484 4868 55488 4924
rect 55424 4864 55488 4868
rect 73584 4924 73648 4928
rect 73584 4868 73588 4924
rect 73588 4868 73644 4924
rect 73644 4868 73648 4924
rect 73584 4864 73648 4868
rect 73664 4924 73728 4928
rect 73664 4868 73668 4924
rect 73668 4868 73724 4924
rect 73724 4868 73728 4924
rect 73664 4864 73728 4868
rect 73744 4924 73808 4928
rect 73744 4868 73748 4924
rect 73748 4868 73804 4924
rect 73804 4868 73808 4924
rect 73744 4864 73808 4868
rect 73824 4924 73888 4928
rect 73824 4868 73828 4924
rect 73828 4868 73884 4924
rect 73884 4868 73888 4924
rect 73824 4864 73888 4868
<< metal4 >>
rect 2696 89722 3016 89764
rect 2696 89486 2738 89722
rect 2974 89486 3016 89722
rect 2696 73874 3016 89486
rect 2696 73638 2738 73874
rect 2974 73638 3016 73874
rect 2696 55474 3016 73638
rect 2696 55238 2738 55474
rect 2974 55238 3016 55474
rect 2696 37074 3016 55238
rect 2696 36838 2738 37074
rect 2974 36838 3016 37074
rect 2696 18674 3016 36838
rect 2696 18438 2738 18674
rect 2974 18438 3016 18674
rect 2696 2994 3016 18438
rect 3356 89062 3676 89104
rect 3356 88826 3398 89062
rect 3634 88826 3676 89062
rect 3356 73214 3676 88826
rect 17716 89062 18036 89764
rect 17716 88826 17758 89062
rect 17994 88826 18036 89062
rect 17716 87072 18036 88826
rect 17716 87008 17724 87072
rect 17788 87008 17804 87072
rect 17868 87008 17884 87072
rect 17948 87008 17964 87072
rect 18028 87008 18036 87072
rect 17716 85984 18036 87008
rect 17716 85920 17724 85984
rect 17788 85920 17804 85984
rect 17868 85920 17884 85984
rect 17948 85920 17964 85984
rect 18028 85920 18036 85984
rect 3356 72978 3398 73214
rect 3634 72978 3676 73214
rect 3356 54814 3676 72978
rect 3356 54578 3398 54814
rect 3634 54578 3676 54814
rect 3356 36414 3676 54578
rect 3356 36178 3398 36414
rect 3634 36178 3676 36414
rect 3356 18014 3676 36178
rect 3356 17778 3398 18014
rect 3634 17778 3676 18014
rect 3356 3654 3676 17778
rect 5876 84896 6196 84912
rect 5876 84832 5884 84896
rect 5948 84832 5964 84896
rect 6028 84832 6044 84896
rect 6108 84832 6124 84896
rect 6188 84832 6196 84896
rect 5876 83808 6196 84832
rect 5876 83744 5884 83808
rect 5948 83744 5964 83808
rect 6028 83744 6044 83808
rect 6108 83744 6124 83808
rect 6188 83744 6196 83808
rect 5876 82720 6196 83744
rect 5876 82656 5884 82720
rect 5948 82656 5964 82720
rect 6028 82656 6044 82720
rect 6108 82656 6124 82720
rect 6188 82656 6196 82720
rect 5876 81632 6196 82656
rect 5876 81568 5884 81632
rect 5948 81568 5964 81632
rect 6028 81568 6044 81632
rect 6108 81568 6124 81632
rect 6188 81568 6196 81632
rect 5876 80544 6196 81568
rect 5876 80480 5884 80544
rect 5948 80480 5964 80544
rect 6028 80480 6044 80544
rect 6108 80480 6124 80544
rect 6188 80480 6196 80544
rect 5876 79456 6196 80480
rect 5876 79392 5884 79456
rect 5948 79392 5964 79456
rect 6028 79392 6044 79456
rect 6108 79392 6124 79456
rect 6188 79392 6196 79456
rect 5876 78368 6196 79392
rect 5876 78304 5884 78368
rect 5948 78304 5964 78368
rect 6028 78304 6044 78368
rect 6108 78304 6124 78368
rect 6188 78304 6196 78368
rect 5876 77280 6196 78304
rect 5876 77216 5884 77280
rect 5948 77216 5964 77280
rect 6028 77216 6044 77280
rect 6108 77216 6124 77280
rect 6188 77216 6196 77280
rect 5876 76192 6196 77216
rect 5876 76128 5884 76192
rect 5948 76128 5964 76192
rect 6028 76128 6044 76192
rect 6108 76128 6124 76192
rect 6188 76128 6196 76192
rect 5876 75104 6196 76128
rect 5876 75040 5884 75104
rect 5948 75040 5964 75104
rect 6028 75040 6044 75104
rect 6108 75040 6124 75104
rect 6188 75040 6196 75104
rect 5876 74016 6196 75040
rect 5876 73952 5884 74016
rect 5948 73952 5964 74016
rect 6028 73952 6044 74016
rect 6108 73952 6124 74016
rect 6188 73952 6196 74016
rect 5876 73214 6196 73952
rect 5876 72978 5918 73214
rect 6154 72978 6196 73214
rect 5876 72928 6196 72978
rect 5876 72864 5884 72928
rect 5948 72864 5964 72928
rect 6028 72864 6044 72928
rect 6108 72864 6124 72928
rect 6188 72864 6196 72928
rect 5876 71840 6196 72864
rect 5876 71776 5884 71840
rect 5948 71776 5964 71840
rect 6028 71776 6044 71840
rect 6108 71776 6124 71840
rect 6188 71776 6196 71840
rect 5876 70752 6196 71776
rect 5876 70688 5884 70752
rect 5948 70688 5964 70752
rect 6028 70688 6044 70752
rect 6108 70688 6124 70752
rect 6188 70688 6196 70752
rect 5876 69664 6196 70688
rect 5876 69600 5884 69664
rect 5948 69600 5964 69664
rect 6028 69600 6044 69664
rect 6108 69600 6124 69664
rect 6188 69600 6196 69664
rect 5876 68576 6196 69600
rect 5876 68512 5884 68576
rect 5948 68512 5964 68576
rect 6028 68512 6044 68576
rect 6108 68512 6124 68576
rect 6188 68512 6196 68576
rect 5876 67488 6196 68512
rect 5876 67424 5884 67488
rect 5948 67424 5964 67488
rect 6028 67424 6044 67488
rect 6108 67424 6124 67488
rect 6188 67424 6196 67488
rect 5876 66400 6196 67424
rect 5876 66336 5884 66400
rect 5948 66336 5964 66400
rect 6028 66336 6044 66400
rect 6108 66336 6124 66400
rect 6188 66336 6196 66400
rect 5876 65312 6196 66336
rect 5876 65248 5884 65312
rect 5948 65248 5964 65312
rect 6028 65248 6044 65312
rect 6108 65248 6124 65312
rect 6188 65248 6196 65312
rect 5876 64224 6196 65248
rect 5876 64160 5884 64224
rect 5948 64160 5964 64224
rect 6028 64160 6044 64224
rect 6108 64160 6124 64224
rect 6188 64160 6196 64224
rect 5876 63136 6196 64160
rect 5876 63072 5884 63136
rect 5948 63072 5964 63136
rect 6028 63072 6044 63136
rect 6108 63072 6124 63136
rect 6188 63072 6196 63136
rect 5876 62048 6196 63072
rect 5876 61984 5884 62048
rect 5948 61984 5964 62048
rect 6028 61984 6044 62048
rect 6108 61984 6124 62048
rect 6188 61984 6196 62048
rect 5876 60960 6196 61984
rect 5876 60896 5884 60960
rect 5948 60896 5964 60960
rect 6028 60896 6044 60960
rect 6108 60896 6124 60960
rect 6188 60896 6196 60960
rect 5876 59872 6196 60896
rect 5876 59808 5884 59872
rect 5948 59808 5964 59872
rect 6028 59808 6044 59872
rect 6108 59808 6124 59872
rect 6188 59808 6196 59872
rect 5876 58784 6196 59808
rect 5876 58720 5884 58784
rect 5948 58720 5964 58784
rect 6028 58720 6044 58784
rect 6108 58720 6124 58784
rect 6188 58720 6196 58784
rect 5876 57696 6196 58720
rect 5876 57632 5884 57696
rect 5948 57632 5964 57696
rect 6028 57632 6044 57696
rect 6108 57632 6124 57696
rect 6188 57632 6196 57696
rect 5876 56608 6196 57632
rect 5876 56544 5884 56608
rect 5948 56544 5964 56608
rect 6028 56544 6044 56608
rect 6108 56544 6124 56608
rect 6188 56544 6196 56608
rect 5876 55520 6196 56544
rect 5876 55456 5884 55520
rect 5948 55456 5964 55520
rect 6028 55456 6044 55520
rect 6108 55456 6124 55520
rect 6188 55456 6196 55520
rect 5876 54814 6196 55456
rect 5876 54578 5918 54814
rect 6154 54578 6196 54814
rect 5876 54432 6196 54578
rect 5876 54368 5884 54432
rect 5948 54368 5964 54432
rect 6028 54368 6044 54432
rect 6108 54368 6124 54432
rect 6188 54368 6196 54432
rect 5876 53344 6196 54368
rect 5876 53280 5884 53344
rect 5948 53280 5964 53344
rect 6028 53280 6044 53344
rect 6108 53280 6124 53344
rect 6188 53280 6196 53344
rect 5876 52256 6196 53280
rect 5876 52192 5884 52256
rect 5948 52192 5964 52256
rect 6028 52192 6044 52256
rect 6108 52192 6124 52256
rect 6188 52192 6196 52256
rect 5876 51168 6196 52192
rect 5876 51104 5884 51168
rect 5948 51104 5964 51168
rect 6028 51104 6044 51168
rect 6108 51104 6124 51168
rect 6188 51104 6196 51168
rect 5876 50080 6196 51104
rect 5876 50016 5884 50080
rect 5948 50016 5964 50080
rect 6028 50016 6044 50080
rect 6108 50016 6124 50080
rect 6188 50016 6196 50080
rect 5876 48992 6196 50016
rect 5876 48928 5884 48992
rect 5948 48928 5964 48992
rect 6028 48928 6044 48992
rect 6108 48928 6124 48992
rect 6188 48928 6196 48992
rect 5876 47904 6196 48928
rect 5876 47840 5884 47904
rect 5948 47840 5964 47904
rect 6028 47840 6044 47904
rect 6108 47840 6124 47904
rect 6188 47840 6196 47904
rect 5876 46816 6196 47840
rect 5876 46752 5884 46816
rect 5948 46752 5964 46816
rect 6028 46752 6044 46816
rect 6108 46752 6124 46816
rect 6188 46752 6196 46816
rect 5876 45728 6196 46752
rect 5876 45664 5884 45728
rect 5948 45664 5964 45728
rect 6028 45664 6044 45728
rect 6108 45664 6124 45728
rect 6188 45664 6196 45728
rect 5876 44640 6196 45664
rect 5876 44576 5884 44640
rect 5948 44576 5964 44640
rect 6028 44576 6044 44640
rect 6108 44576 6124 44640
rect 6188 44576 6196 44640
rect 5876 43552 6196 44576
rect 5876 43488 5884 43552
rect 5948 43488 5964 43552
rect 6028 43488 6044 43552
rect 6108 43488 6124 43552
rect 6188 43488 6196 43552
rect 5876 42464 6196 43488
rect 5876 42400 5884 42464
rect 5948 42400 5964 42464
rect 6028 42400 6044 42464
rect 6108 42400 6124 42464
rect 6188 42400 6196 42464
rect 5876 41376 6196 42400
rect 5876 41312 5884 41376
rect 5948 41312 5964 41376
rect 6028 41312 6044 41376
rect 6108 41312 6124 41376
rect 6188 41312 6196 41376
rect 5876 40288 6196 41312
rect 5876 40224 5884 40288
rect 5948 40224 5964 40288
rect 6028 40224 6044 40288
rect 6108 40224 6124 40288
rect 6188 40224 6196 40288
rect 5876 39200 6196 40224
rect 5876 39136 5884 39200
rect 5948 39136 5964 39200
rect 6028 39136 6044 39200
rect 6108 39136 6124 39200
rect 6188 39136 6196 39200
rect 5876 38112 6196 39136
rect 5876 38048 5884 38112
rect 5948 38048 5964 38112
rect 6028 38048 6044 38112
rect 6108 38048 6124 38112
rect 6188 38048 6196 38112
rect 5876 37024 6196 38048
rect 5876 36960 5884 37024
rect 5948 36960 5964 37024
rect 6028 36960 6044 37024
rect 6108 36960 6124 37024
rect 6188 36960 6196 37024
rect 5876 36414 6196 36960
rect 5876 36178 5918 36414
rect 6154 36178 6196 36414
rect 5876 35936 6196 36178
rect 5876 35872 5884 35936
rect 5948 35872 5964 35936
rect 6028 35872 6044 35936
rect 6108 35872 6124 35936
rect 6188 35872 6196 35936
rect 5876 34848 6196 35872
rect 5876 34784 5884 34848
rect 5948 34784 5964 34848
rect 6028 34784 6044 34848
rect 6108 34784 6124 34848
rect 6188 34784 6196 34848
rect 5876 33760 6196 34784
rect 5876 33696 5884 33760
rect 5948 33696 5964 33760
rect 6028 33696 6044 33760
rect 6108 33696 6124 33760
rect 6188 33696 6196 33760
rect 5876 32672 6196 33696
rect 5876 32608 5884 32672
rect 5948 32608 5964 32672
rect 6028 32608 6044 32672
rect 6108 32608 6124 32672
rect 6188 32608 6196 32672
rect 5876 31584 6196 32608
rect 5876 31520 5884 31584
rect 5948 31520 5964 31584
rect 6028 31520 6044 31584
rect 6108 31520 6124 31584
rect 6188 31520 6196 31584
rect 5876 30496 6196 31520
rect 5876 30432 5884 30496
rect 5948 30432 5964 30496
rect 6028 30432 6044 30496
rect 6108 30432 6124 30496
rect 6188 30432 6196 30496
rect 5876 29408 6196 30432
rect 5876 29344 5884 29408
rect 5948 29344 5964 29408
rect 6028 29344 6044 29408
rect 6108 29344 6124 29408
rect 6188 29344 6196 29408
rect 5876 28320 6196 29344
rect 5876 28256 5884 28320
rect 5948 28256 5964 28320
rect 6028 28256 6044 28320
rect 6108 28256 6124 28320
rect 6188 28256 6196 28320
rect 5876 27232 6196 28256
rect 5876 27168 5884 27232
rect 5948 27168 5964 27232
rect 6028 27168 6044 27232
rect 6108 27168 6124 27232
rect 6188 27168 6196 27232
rect 5876 26144 6196 27168
rect 5876 26080 5884 26144
rect 5948 26080 5964 26144
rect 6028 26080 6044 26144
rect 6108 26080 6124 26144
rect 6188 26080 6196 26144
rect 5876 25056 6196 26080
rect 5876 24992 5884 25056
rect 5948 24992 5964 25056
rect 6028 24992 6044 25056
rect 6108 24992 6124 25056
rect 6188 24992 6196 25056
rect 5876 23968 6196 24992
rect 5876 23904 5884 23968
rect 5948 23904 5964 23968
rect 6028 23904 6044 23968
rect 6108 23904 6124 23968
rect 6188 23904 6196 23968
rect 5876 22880 6196 23904
rect 5876 22816 5884 22880
rect 5948 22816 5964 22880
rect 6028 22816 6044 22880
rect 6108 22816 6124 22880
rect 6188 22816 6196 22880
rect 5876 21792 6196 22816
rect 5876 21728 5884 21792
rect 5948 21728 5964 21792
rect 6028 21728 6044 21792
rect 6108 21728 6124 21792
rect 6188 21728 6196 21792
rect 5876 20704 6196 21728
rect 5876 20640 5884 20704
rect 5948 20640 5964 20704
rect 6028 20640 6044 20704
rect 6108 20640 6124 20704
rect 6188 20640 6196 20704
rect 5876 19616 6196 20640
rect 5876 19552 5884 19616
rect 5948 19552 5964 19616
rect 6028 19552 6044 19616
rect 6108 19552 6124 19616
rect 6188 19552 6196 19616
rect 5876 18528 6196 19552
rect 5876 18464 5884 18528
rect 5948 18464 5964 18528
rect 6028 18464 6044 18528
rect 6108 18464 6124 18528
rect 6188 18464 6196 18528
rect 5876 18014 6196 18464
rect 5876 17778 5918 18014
rect 6154 17778 6196 18014
rect 5876 17440 6196 17778
rect 5876 17376 5884 17440
rect 5948 17376 5964 17440
rect 6028 17376 6044 17440
rect 6108 17376 6124 17440
rect 6188 17376 6196 17440
rect 5876 16352 6196 17376
rect 5876 16288 5884 16352
rect 5948 16288 5964 16352
rect 6028 16288 6044 16352
rect 6108 16288 6124 16352
rect 6188 16288 6196 16352
rect 5876 15264 6196 16288
rect 5876 15200 5884 15264
rect 5948 15200 5964 15264
rect 6028 15200 6044 15264
rect 6108 15200 6124 15264
rect 6188 15200 6196 15264
rect 5876 14176 6196 15200
rect 5876 14112 5884 14176
rect 5948 14112 5964 14176
rect 6028 14112 6044 14176
rect 6108 14112 6124 14176
rect 6188 14112 6196 14176
rect 5876 13088 6196 14112
rect 5876 13024 5884 13088
rect 5948 13024 5964 13088
rect 6028 13024 6044 13088
rect 6108 13024 6124 13088
rect 6188 13024 6196 13088
rect 5876 12000 6196 13024
rect 5876 11936 5884 12000
rect 5948 11936 5964 12000
rect 6028 11936 6044 12000
rect 6108 11936 6124 12000
rect 6188 11936 6196 12000
rect 5876 10912 6196 11936
rect 5876 10848 5884 10912
rect 5948 10848 5964 10912
rect 6028 10848 6044 10912
rect 6108 10848 6124 10912
rect 6188 10848 6196 10912
rect 5876 9824 6196 10848
rect 5876 9760 5884 9824
rect 5948 9760 5964 9824
rect 6028 9760 6044 9824
rect 6108 9760 6124 9824
rect 6188 9760 6196 9824
rect 5876 8736 6196 9760
rect 5876 8672 5884 8736
rect 5948 8672 5964 8736
rect 6028 8672 6044 8736
rect 6108 8672 6124 8736
rect 6188 8672 6196 8736
rect 5876 7648 6196 8672
rect 5876 7584 5884 7648
rect 5948 7584 5964 7648
rect 6028 7584 6044 7648
rect 6108 7584 6124 7648
rect 6188 7584 6196 7648
rect 5876 7024 6196 7584
rect 6612 84352 6932 84912
rect 6612 84288 6620 84352
rect 6684 84288 6700 84352
rect 6764 84288 6780 84352
rect 6844 84288 6860 84352
rect 6924 84288 6932 84352
rect 6612 83264 6932 84288
rect 6612 83200 6620 83264
rect 6684 83200 6700 83264
rect 6764 83200 6780 83264
rect 6844 83200 6860 83264
rect 6924 83200 6932 83264
rect 6612 82176 6932 83200
rect 6612 82112 6620 82176
rect 6684 82112 6700 82176
rect 6764 82112 6780 82176
rect 6844 82112 6860 82176
rect 6924 82112 6932 82176
rect 6612 81088 6932 82112
rect 6612 81024 6620 81088
rect 6684 81024 6700 81088
rect 6764 81024 6780 81088
rect 6844 81024 6860 81088
rect 6924 81024 6932 81088
rect 17716 84896 18036 85920
rect 17716 84832 17724 84896
rect 17788 84832 17804 84896
rect 17868 84832 17884 84896
rect 17948 84832 17964 84896
rect 18028 84832 18036 84896
rect 17716 81029 18036 84832
rect 18376 89722 18696 89764
rect 18376 89486 18418 89722
rect 18654 89486 18696 89722
rect 18376 87616 18696 89486
rect 18376 87552 18384 87616
rect 18448 87552 18464 87616
rect 18528 87552 18544 87616
rect 18608 87552 18624 87616
rect 18688 87552 18696 87616
rect 18376 86528 18696 87552
rect 18376 86464 18384 86528
rect 18448 86464 18464 86528
rect 18528 86464 18544 86528
rect 18608 86464 18624 86528
rect 18688 86464 18696 86528
rect 18376 85440 18696 86464
rect 18376 85376 18384 85440
rect 18448 85376 18464 85440
rect 18528 85376 18544 85440
rect 18608 85376 18624 85440
rect 18688 85376 18696 85440
rect 18376 84352 18696 85376
rect 18376 84288 18384 84352
rect 18448 84288 18464 84352
rect 18528 84288 18544 84352
rect 18608 84288 18624 84352
rect 18688 84288 18696 84352
rect 18376 81029 18696 84288
rect 36116 89062 36436 89764
rect 36116 88826 36158 89062
rect 36394 88826 36436 89062
rect 36116 87072 36436 88826
rect 36116 87008 36124 87072
rect 36188 87008 36204 87072
rect 36268 87008 36284 87072
rect 36348 87008 36364 87072
rect 36428 87008 36436 87072
rect 36116 85984 36436 87008
rect 36116 85920 36124 85984
rect 36188 85920 36204 85984
rect 36268 85920 36284 85984
rect 36348 85920 36364 85984
rect 36428 85920 36436 85984
rect 36116 84896 36436 85920
rect 36116 84832 36124 84896
rect 36188 84832 36204 84896
rect 36268 84832 36284 84896
rect 36348 84832 36364 84896
rect 36428 84832 36436 84896
rect 36116 81029 36436 84832
rect 36776 89722 37096 89764
rect 36776 89486 36818 89722
rect 37054 89486 37096 89722
rect 36776 87616 37096 89486
rect 36776 87552 36784 87616
rect 36848 87552 36864 87616
rect 36928 87552 36944 87616
rect 37008 87552 37024 87616
rect 37088 87552 37096 87616
rect 36776 86528 37096 87552
rect 36776 86464 36784 86528
rect 36848 86464 36864 86528
rect 36928 86464 36944 86528
rect 37008 86464 37024 86528
rect 37088 86464 37096 86528
rect 36776 85440 37096 86464
rect 36776 85376 36784 85440
rect 36848 85376 36864 85440
rect 36928 85376 36944 85440
rect 37008 85376 37024 85440
rect 37088 85376 37096 85440
rect 36776 84352 37096 85376
rect 36776 84288 36784 84352
rect 36848 84288 36864 84352
rect 36928 84288 36944 84352
rect 37008 84288 37024 84352
rect 37088 84288 37096 84352
rect 36776 81029 37096 84288
rect 54516 89062 54836 89764
rect 54516 88826 54558 89062
rect 54794 88826 54836 89062
rect 54516 87072 54836 88826
rect 54516 87008 54524 87072
rect 54588 87008 54604 87072
rect 54668 87008 54684 87072
rect 54748 87008 54764 87072
rect 54828 87008 54836 87072
rect 54516 85984 54836 87008
rect 54516 85920 54524 85984
rect 54588 85920 54604 85984
rect 54668 85920 54684 85984
rect 54748 85920 54764 85984
rect 54828 85920 54836 85984
rect 54516 84896 54836 85920
rect 54516 84832 54524 84896
rect 54588 84832 54604 84896
rect 54668 84832 54684 84896
rect 54748 84832 54764 84896
rect 54828 84832 54836 84896
rect 54516 81029 54836 84832
rect 55176 89722 55496 89764
rect 55176 89486 55218 89722
rect 55454 89486 55496 89722
rect 55176 87616 55496 89486
rect 55176 87552 55184 87616
rect 55248 87552 55264 87616
rect 55328 87552 55344 87616
rect 55408 87552 55424 87616
rect 55488 87552 55496 87616
rect 55176 86528 55496 87552
rect 55176 86464 55184 86528
rect 55248 86464 55264 86528
rect 55328 86464 55344 86528
rect 55408 86464 55424 86528
rect 55488 86464 55496 86528
rect 55176 85440 55496 86464
rect 55176 85376 55184 85440
rect 55248 85376 55264 85440
rect 55328 85376 55344 85440
rect 55408 85376 55424 85440
rect 55488 85376 55496 85440
rect 55176 84352 55496 85376
rect 55176 84288 55184 84352
rect 55248 84288 55264 84352
rect 55328 84288 55344 84352
rect 55408 84288 55424 84352
rect 55488 84288 55496 84352
rect 55176 81029 55496 84288
rect 72916 89062 73236 89764
rect 72916 88826 72958 89062
rect 73194 88826 73236 89062
rect 72916 87072 73236 88826
rect 72916 87008 72924 87072
rect 72988 87008 73004 87072
rect 73068 87008 73084 87072
rect 73148 87008 73164 87072
rect 73228 87008 73236 87072
rect 72916 85984 73236 87008
rect 72916 85920 72924 85984
rect 72988 85920 73004 85984
rect 73068 85920 73084 85984
rect 73148 85920 73164 85984
rect 73228 85920 73236 85984
rect 72916 84896 73236 85920
rect 72916 84832 72924 84896
rect 72988 84832 73004 84896
rect 73068 84832 73084 84896
rect 73148 84832 73164 84896
rect 73228 84832 73236 84896
rect 72916 81029 73236 84832
rect 73576 89722 73896 89764
rect 73576 89486 73618 89722
rect 73854 89486 73896 89722
rect 73576 87616 73896 89486
rect 90456 89722 90776 89764
rect 90456 89486 90498 89722
rect 90734 89486 90776 89722
rect 73576 87552 73584 87616
rect 73648 87552 73664 87616
rect 73728 87552 73744 87616
rect 73808 87552 73824 87616
rect 73888 87552 73896 87616
rect 73576 86528 73896 87552
rect 73576 86464 73584 86528
rect 73648 86464 73664 86528
rect 73728 86464 73744 86528
rect 73808 86464 73824 86528
rect 73888 86464 73896 86528
rect 73576 85440 73896 86464
rect 73576 85376 73584 85440
rect 73648 85376 73664 85440
rect 73728 85376 73744 85440
rect 73808 85376 73824 85440
rect 73888 85376 73896 85440
rect 73576 84352 73896 85376
rect 89796 89062 90116 89104
rect 89796 88826 89838 89062
rect 90074 88826 90116 89062
rect 73576 84288 73584 84352
rect 73648 84288 73664 84352
rect 73728 84288 73744 84352
rect 73808 84288 73824 84352
rect 73888 84288 73896 84352
rect 73576 81029 73896 84288
rect 86468 84896 86788 84912
rect 86468 84832 86476 84896
rect 86540 84832 86556 84896
rect 86620 84832 86636 84896
rect 86700 84832 86716 84896
rect 86780 84832 86788 84896
rect 86468 83808 86788 84832
rect 86468 83744 86476 83808
rect 86540 83744 86556 83808
rect 86620 83744 86636 83808
rect 86700 83744 86716 83808
rect 86780 83744 86788 83808
rect 86468 82720 86788 83744
rect 86468 82656 86476 82720
rect 86540 82656 86556 82720
rect 86620 82656 86636 82720
rect 86700 82656 86716 82720
rect 86780 82656 86788 82720
rect 86468 81632 86788 82656
rect 86468 81568 86476 81632
rect 86540 81568 86556 81632
rect 86620 81568 86636 81632
rect 86700 81568 86716 81632
rect 86780 81568 86788 81632
rect 6612 80000 6932 81024
rect 11144 80630 11186 80866
rect 11422 80630 11464 80866
rect 43744 80630 43786 80866
rect 44022 80630 44064 80866
rect 48544 80630 48586 80866
rect 48822 80630 48864 80866
rect 81144 80630 81186 80866
rect 81422 80630 81464 80866
rect 86468 80544 86788 81568
rect 86468 80480 86476 80544
rect 86540 80480 86556 80544
rect 86620 80480 86636 80544
rect 86700 80480 86716 80544
rect 86780 80480 86788 80544
rect 6612 79936 6620 80000
rect 6684 79936 6700 80000
rect 6764 79936 6780 80000
rect 6844 79936 6860 80000
rect 6924 79936 6932 80000
rect 10484 79970 10526 80206
rect 10762 79970 10804 80206
rect 43084 79970 43126 80206
rect 43362 79970 43404 80206
rect 47884 79970 47926 80206
rect 48162 79970 48204 80206
rect 80484 79970 80526 80206
rect 80762 79970 80804 80206
rect 6612 78912 6932 79936
rect 6612 78848 6620 78912
rect 6684 78848 6700 78912
rect 6764 78848 6780 78912
rect 6844 78848 6860 78912
rect 6924 78848 6932 78912
rect 6612 77824 6932 78848
rect 6612 77760 6620 77824
rect 6684 77760 6700 77824
rect 6764 77760 6780 77824
rect 6844 77760 6860 77824
rect 6924 77760 6932 77824
rect 6612 76736 6932 77760
rect 6612 76672 6620 76736
rect 6684 76672 6700 76736
rect 6764 76672 6780 76736
rect 6844 76672 6860 76736
rect 6924 76672 6932 76736
rect 6612 75648 6932 76672
rect 6612 75584 6620 75648
rect 6684 75584 6700 75648
rect 6764 75584 6780 75648
rect 6844 75584 6860 75648
rect 6924 75584 6932 75648
rect 6612 74560 6932 75584
rect 6612 74496 6620 74560
rect 6684 74496 6700 74560
rect 6764 74496 6780 74560
rect 6844 74496 6860 74560
rect 6924 74496 6932 74560
rect 6612 73874 6932 74496
rect 86468 79456 86788 80480
rect 86468 79392 86476 79456
rect 86540 79392 86556 79456
rect 86620 79392 86636 79456
rect 86700 79392 86716 79456
rect 86780 79392 86788 79456
rect 86468 78368 86788 79392
rect 86468 78304 86476 78368
rect 86540 78304 86556 78368
rect 86620 78304 86636 78368
rect 86700 78304 86716 78368
rect 86780 78304 86788 78368
rect 86468 77280 86788 78304
rect 86468 77216 86476 77280
rect 86540 77216 86556 77280
rect 86620 77216 86636 77280
rect 86700 77216 86716 77280
rect 86780 77216 86788 77280
rect 86468 76192 86788 77216
rect 86468 76128 86476 76192
rect 86540 76128 86556 76192
rect 86620 76128 86636 76192
rect 86700 76128 86716 76192
rect 86780 76128 86788 76192
rect 86468 75104 86788 76128
rect 86468 75040 86476 75104
rect 86540 75040 86556 75104
rect 86620 75040 86636 75104
rect 86700 75040 86716 75104
rect 86780 75040 86788 75104
rect 86468 74016 86788 75040
rect 86468 73952 86476 74016
rect 86540 73952 86556 74016
rect 86620 73952 86636 74016
rect 86700 73952 86716 74016
rect 86780 73952 86788 74016
rect 6612 73638 6654 73874
rect 6890 73638 6932 73874
rect 11144 73638 11186 73874
rect 11422 73638 11464 73874
rect 43744 73638 43786 73874
rect 44022 73638 44064 73874
rect 48544 73638 48586 73874
rect 48822 73638 48864 73874
rect 81144 73638 81186 73874
rect 81422 73638 81464 73874
rect 6612 73472 6932 73638
rect 6612 73408 6620 73472
rect 6684 73408 6700 73472
rect 6764 73408 6780 73472
rect 6844 73408 6860 73472
rect 6924 73408 6932 73472
rect 6612 72384 6932 73408
rect 86468 73214 86788 73952
rect 10484 72978 10526 73214
rect 10762 72978 10804 73214
rect 43084 72978 43126 73214
rect 43362 72978 43404 73214
rect 47884 72978 47926 73214
rect 48162 72978 48204 73214
rect 80484 72978 80526 73214
rect 80762 72978 80804 73214
rect 86468 72978 86510 73214
rect 86746 72978 86788 73214
rect 6612 72320 6620 72384
rect 6684 72320 6700 72384
rect 6764 72320 6780 72384
rect 6844 72320 6860 72384
rect 6924 72320 6932 72384
rect 6612 71296 6932 72320
rect 6612 71232 6620 71296
rect 6684 71232 6700 71296
rect 6764 71232 6780 71296
rect 6844 71232 6860 71296
rect 6924 71232 6932 71296
rect 6612 70208 6932 71232
rect 6612 70144 6620 70208
rect 6684 70144 6700 70208
rect 6764 70144 6780 70208
rect 6844 70144 6860 70208
rect 6924 70144 6932 70208
rect 6612 69120 6932 70144
rect 6612 69056 6620 69120
rect 6684 69056 6700 69120
rect 6764 69056 6780 69120
rect 6844 69056 6860 69120
rect 6924 69056 6932 69120
rect 6612 68032 6932 69056
rect 6612 67968 6620 68032
rect 6684 67968 6700 68032
rect 6764 67968 6780 68032
rect 6844 67968 6860 68032
rect 6924 67968 6932 68032
rect 6612 66944 6932 67968
rect 6612 66880 6620 66944
rect 6684 66880 6700 66944
rect 6764 66880 6780 66944
rect 6844 66880 6860 66944
rect 6924 66880 6932 66944
rect 6612 65856 6932 66880
rect 6612 65792 6620 65856
rect 6684 65792 6700 65856
rect 6764 65792 6780 65856
rect 6844 65792 6860 65856
rect 6924 65792 6932 65856
rect 6612 64768 6932 65792
rect 6612 64704 6620 64768
rect 6684 64704 6700 64768
rect 6764 64704 6780 64768
rect 6844 64704 6860 64768
rect 6924 64704 6932 64768
rect 6612 63680 6932 64704
rect 6612 63616 6620 63680
rect 6684 63616 6700 63680
rect 6764 63616 6780 63680
rect 6844 63616 6860 63680
rect 6924 63616 6932 63680
rect 6612 62592 6932 63616
rect 6612 62528 6620 62592
rect 6684 62528 6700 62592
rect 6764 62528 6780 62592
rect 6844 62528 6860 62592
rect 6924 62528 6932 62592
rect 6612 61504 6932 62528
rect 6612 61440 6620 61504
rect 6684 61440 6700 61504
rect 6764 61440 6780 61504
rect 6844 61440 6860 61504
rect 6924 61440 6932 61504
rect 6612 60416 6932 61440
rect 6612 60352 6620 60416
rect 6684 60352 6700 60416
rect 6764 60352 6780 60416
rect 6844 60352 6860 60416
rect 6924 60352 6932 60416
rect 6612 59328 6932 60352
rect 6612 59264 6620 59328
rect 6684 59264 6700 59328
rect 6764 59264 6780 59328
rect 6844 59264 6860 59328
rect 6924 59264 6932 59328
rect 6612 58240 6932 59264
rect 6612 58176 6620 58240
rect 6684 58176 6700 58240
rect 6764 58176 6780 58240
rect 6844 58176 6860 58240
rect 6924 58176 6932 58240
rect 6612 57152 6932 58176
rect 6612 57088 6620 57152
rect 6684 57088 6700 57152
rect 6764 57088 6780 57152
rect 6844 57088 6860 57152
rect 6924 57088 6932 57152
rect 6612 56064 6932 57088
rect 6612 56000 6620 56064
rect 6684 56000 6700 56064
rect 6764 56000 6780 56064
rect 6844 56000 6860 56064
rect 6924 56000 6932 56064
rect 6612 55474 6932 56000
rect 86468 72928 86788 72978
rect 86468 72864 86476 72928
rect 86540 72864 86556 72928
rect 86620 72864 86636 72928
rect 86700 72864 86716 72928
rect 86780 72864 86788 72928
rect 86468 71840 86788 72864
rect 86468 71776 86476 71840
rect 86540 71776 86556 71840
rect 86620 71776 86636 71840
rect 86700 71776 86716 71840
rect 86780 71776 86788 71840
rect 86468 70752 86788 71776
rect 86468 70688 86476 70752
rect 86540 70688 86556 70752
rect 86620 70688 86636 70752
rect 86700 70688 86716 70752
rect 86780 70688 86788 70752
rect 86468 69664 86788 70688
rect 86468 69600 86476 69664
rect 86540 69600 86556 69664
rect 86620 69600 86636 69664
rect 86700 69600 86716 69664
rect 86780 69600 86788 69664
rect 86468 68576 86788 69600
rect 86468 68512 86476 68576
rect 86540 68512 86556 68576
rect 86620 68512 86636 68576
rect 86700 68512 86716 68576
rect 86780 68512 86788 68576
rect 86468 67488 86788 68512
rect 86468 67424 86476 67488
rect 86540 67424 86556 67488
rect 86620 67424 86636 67488
rect 86700 67424 86716 67488
rect 86780 67424 86788 67488
rect 86468 66400 86788 67424
rect 86468 66336 86476 66400
rect 86540 66336 86556 66400
rect 86620 66336 86636 66400
rect 86700 66336 86716 66400
rect 86780 66336 86788 66400
rect 86468 65312 86788 66336
rect 86468 65248 86476 65312
rect 86540 65248 86556 65312
rect 86620 65248 86636 65312
rect 86700 65248 86716 65312
rect 86780 65248 86788 65312
rect 86468 64224 86788 65248
rect 86468 64160 86476 64224
rect 86540 64160 86556 64224
rect 86620 64160 86636 64224
rect 86700 64160 86716 64224
rect 86780 64160 86788 64224
rect 86468 63136 86788 64160
rect 86468 63072 86476 63136
rect 86540 63072 86556 63136
rect 86620 63072 86636 63136
rect 86700 63072 86716 63136
rect 86780 63072 86788 63136
rect 86468 62048 86788 63072
rect 86468 61984 86476 62048
rect 86540 61984 86556 62048
rect 86620 61984 86636 62048
rect 86700 61984 86716 62048
rect 86780 61984 86788 62048
rect 86468 60960 86788 61984
rect 86468 60896 86476 60960
rect 86540 60896 86556 60960
rect 86620 60896 86636 60960
rect 86700 60896 86716 60960
rect 86780 60896 86788 60960
rect 86468 59872 86788 60896
rect 86468 59808 86476 59872
rect 86540 59808 86556 59872
rect 86620 59808 86636 59872
rect 86700 59808 86716 59872
rect 86780 59808 86788 59872
rect 86468 58784 86788 59808
rect 86468 58720 86476 58784
rect 86540 58720 86556 58784
rect 86620 58720 86636 58784
rect 86700 58720 86716 58784
rect 86780 58720 86788 58784
rect 86468 57696 86788 58720
rect 86468 57632 86476 57696
rect 86540 57632 86556 57696
rect 86620 57632 86636 57696
rect 86700 57632 86716 57696
rect 86780 57632 86788 57696
rect 86468 56608 86788 57632
rect 86468 56544 86476 56608
rect 86540 56544 86556 56608
rect 86620 56544 86636 56608
rect 86700 56544 86716 56608
rect 86780 56544 86788 56608
rect 86468 55520 86788 56544
rect 6612 55238 6654 55474
rect 6890 55238 6932 55474
rect 11144 55238 11186 55474
rect 11422 55238 11464 55474
rect 43744 55238 43786 55474
rect 44022 55238 44064 55474
rect 48544 55238 48586 55474
rect 48822 55238 48864 55474
rect 81144 55238 81186 55474
rect 81422 55238 81464 55474
rect 86468 55456 86476 55520
rect 86540 55456 86556 55520
rect 86620 55456 86636 55520
rect 86700 55456 86716 55520
rect 86780 55456 86788 55520
rect 6612 54976 6932 55238
rect 6612 54912 6620 54976
rect 6684 54912 6700 54976
rect 6764 54912 6780 54976
rect 6844 54912 6860 54976
rect 6924 54912 6932 54976
rect 6612 53888 6932 54912
rect 86468 54814 86788 55456
rect 10484 54578 10526 54814
rect 10762 54578 10804 54814
rect 43084 54578 43126 54814
rect 43362 54578 43404 54814
rect 47884 54578 47926 54814
rect 48162 54578 48204 54814
rect 80484 54578 80526 54814
rect 80762 54578 80804 54814
rect 86468 54578 86510 54814
rect 86746 54578 86788 54814
rect 6612 53824 6620 53888
rect 6684 53824 6700 53888
rect 6764 53824 6780 53888
rect 6844 53824 6860 53888
rect 6924 53824 6932 53888
rect 6612 52800 6932 53824
rect 6612 52736 6620 52800
rect 6684 52736 6700 52800
rect 6764 52736 6780 52800
rect 6844 52736 6860 52800
rect 6924 52736 6932 52800
rect 6612 51712 6932 52736
rect 6612 51648 6620 51712
rect 6684 51648 6700 51712
rect 6764 51648 6780 51712
rect 6844 51648 6860 51712
rect 6924 51648 6932 51712
rect 6612 50624 6932 51648
rect 6612 50560 6620 50624
rect 6684 50560 6700 50624
rect 6764 50560 6780 50624
rect 6844 50560 6860 50624
rect 6924 50560 6932 50624
rect 6612 49536 6932 50560
rect 6612 49472 6620 49536
rect 6684 49472 6700 49536
rect 6764 49472 6780 49536
rect 6844 49472 6860 49536
rect 6924 49472 6932 49536
rect 6612 48448 6932 49472
rect 6612 48384 6620 48448
rect 6684 48384 6700 48448
rect 6764 48384 6780 48448
rect 6844 48384 6860 48448
rect 6924 48384 6932 48448
rect 6612 47360 6932 48384
rect 86468 54432 86788 54578
rect 86468 54368 86476 54432
rect 86540 54368 86556 54432
rect 86620 54368 86636 54432
rect 86700 54368 86716 54432
rect 86780 54368 86788 54432
rect 86468 53344 86788 54368
rect 86468 53280 86476 53344
rect 86540 53280 86556 53344
rect 86620 53280 86636 53344
rect 86700 53280 86716 53344
rect 86780 53280 86788 53344
rect 86468 52256 86788 53280
rect 86468 52192 86476 52256
rect 86540 52192 86556 52256
rect 86620 52192 86636 52256
rect 86700 52192 86716 52256
rect 86780 52192 86788 52256
rect 86468 51168 86788 52192
rect 86468 51104 86476 51168
rect 86540 51104 86556 51168
rect 86620 51104 86636 51168
rect 86700 51104 86716 51168
rect 86780 51104 86788 51168
rect 86468 50080 86788 51104
rect 86468 50016 86476 50080
rect 86540 50016 86556 50080
rect 86620 50016 86636 50080
rect 86700 50016 86716 50080
rect 86780 50016 86788 50080
rect 86468 48992 86788 50016
rect 86468 48928 86476 48992
rect 86540 48928 86556 48992
rect 86620 48928 86636 48992
rect 86700 48928 86716 48992
rect 86780 48928 86788 48992
rect 11144 48030 11186 48266
rect 11422 48030 11464 48266
rect 43744 48030 43786 48266
rect 44022 48030 44064 48266
rect 48544 48030 48586 48266
rect 48822 48030 48864 48266
rect 81144 48030 81186 48266
rect 81422 48030 81464 48266
rect 86468 47904 86788 48928
rect 86468 47840 86476 47904
rect 86540 47840 86556 47904
rect 86620 47840 86636 47904
rect 86700 47840 86716 47904
rect 86780 47840 86788 47904
rect 10484 47370 10526 47606
rect 10762 47370 10804 47606
rect 43084 47370 43126 47606
rect 43362 47370 43404 47606
rect 47884 47370 47926 47606
rect 48162 47370 48204 47606
rect 80484 47370 80526 47606
rect 80762 47370 80804 47606
rect 6612 47296 6620 47360
rect 6684 47296 6700 47360
rect 6764 47296 6780 47360
rect 6844 47296 6860 47360
rect 6924 47296 6932 47360
rect 6612 46272 6932 47296
rect 6612 46208 6620 46272
rect 6684 46208 6700 46272
rect 6764 46208 6780 46272
rect 6844 46208 6860 46272
rect 6924 46208 6932 46272
rect 6612 45184 6932 46208
rect 86468 46816 86788 47840
rect 86468 46752 86476 46816
rect 86540 46752 86556 46816
rect 86620 46752 86636 46816
rect 86700 46752 86716 46816
rect 86780 46752 86788 46816
rect 11707 45804 11773 45805
rect 11707 45740 11708 45804
rect 11772 45740 11773 45804
rect 11707 45739 11773 45740
rect 11710 45261 11770 45739
rect 86468 45728 86788 46752
rect 86468 45664 86476 45728
rect 86540 45664 86556 45728
rect 86620 45664 86636 45728
rect 86700 45664 86716 45728
rect 86780 45664 86788 45728
rect 11707 45260 11773 45261
rect 11707 45196 11708 45260
rect 11772 45196 11773 45260
rect 11707 45195 11773 45196
rect 6612 45120 6620 45184
rect 6684 45120 6700 45184
rect 6764 45120 6780 45184
rect 6844 45120 6860 45184
rect 6924 45120 6932 45184
rect 6612 44096 6932 45120
rect 86468 44640 86788 45664
rect 86468 44576 86476 44640
rect 86540 44576 86556 44640
rect 86620 44576 86636 44640
rect 86700 44576 86716 44640
rect 86780 44576 86788 44640
rect 11144 44230 11186 44466
rect 11422 44230 11464 44466
rect 43744 44230 43786 44466
rect 44022 44230 44064 44466
rect 48544 44230 48586 44466
rect 48822 44230 48864 44466
rect 81144 44230 81186 44466
rect 81422 44230 81464 44466
rect 6612 44032 6620 44096
rect 6684 44032 6700 44096
rect 6764 44032 6780 44096
rect 6844 44032 6860 44096
rect 6924 44032 6932 44096
rect 6612 43008 6932 44032
rect 10484 43570 10526 43806
rect 10762 43570 10804 43806
rect 43084 43570 43126 43806
rect 43362 43570 43404 43806
rect 47884 43570 47926 43806
rect 48162 43570 48204 43806
rect 80484 43570 80526 43806
rect 80762 43570 80804 43806
rect 6612 42944 6620 43008
rect 6684 42944 6700 43008
rect 6764 42944 6780 43008
rect 6844 42944 6860 43008
rect 6924 42944 6932 43008
rect 6612 41920 6932 42944
rect 6612 41856 6620 41920
rect 6684 41856 6700 41920
rect 6764 41856 6780 41920
rect 6844 41856 6860 41920
rect 6924 41856 6932 41920
rect 6612 40832 6932 41856
rect 6612 40768 6620 40832
rect 6684 40768 6700 40832
rect 6764 40768 6780 40832
rect 6844 40768 6860 40832
rect 6924 40768 6932 40832
rect 6612 39744 6932 40768
rect 6612 39680 6620 39744
rect 6684 39680 6700 39744
rect 6764 39680 6780 39744
rect 6844 39680 6860 39744
rect 6924 39680 6932 39744
rect 6612 38656 6932 39680
rect 6612 38592 6620 38656
rect 6684 38592 6700 38656
rect 6764 38592 6780 38656
rect 6844 38592 6860 38656
rect 6924 38592 6932 38656
rect 6612 37568 6932 38592
rect 6612 37504 6620 37568
rect 6684 37504 6700 37568
rect 6764 37504 6780 37568
rect 6844 37504 6860 37568
rect 6924 37504 6932 37568
rect 6612 37074 6932 37504
rect 86468 43552 86788 44576
rect 86468 43488 86476 43552
rect 86540 43488 86556 43552
rect 86620 43488 86636 43552
rect 86700 43488 86716 43552
rect 86780 43488 86788 43552
rect 86468 42464 86788 43488
rect 86468 42400 86476 42464
rect 86540 42400 86556 42464
rect 86620 42400 86636 42464
rect 86700 42400 86716 42464
rect 86780 42400 86788 42464
rect 86468 41376 86788 42400
rect 86468 41312 86476 41376
rect 86540 41312 86556 41376
rect 86620 41312 86636 41376
rect 86700 41312 86716 41376
rect 86780 41312 86788 41376
rect 86468 40288 86788 41312
rect 86468 40224 86476 40288
rect 86540 40224 86556 40288
rect 86620 40224 86636 40288
rect 86700 40224 86716 40288
rect 86780 40224 86788 40288
rect 86468 39200 86788 40224
rect 86468 39136 86476 39200
rect 86540 39136 86556 39200
rect 86620 39136 86636 39200
rect 86700 39136 86716 39200
rect 86780 39136 86788 39200
rect 86468 38112 86788 39136
rect 86468 38048 86476 38112
rect 86540 38048 86556 38112
rect 86620 38048 86636 38112
rect 86700 38048 86716 38112
rect 86780 38048 86788 38112
rect 6612 36838 6654 37074
rect 6890 36838 6932 37074
rect 11144 36838 11186 37074
rect 11422 36838 11464 37074
rect 43744 36838 43786 37074
rect 44022 36838 44064 37074
rect 48544 36838 48586 37074
rect 48822 36838 48864 37074
rect 81144 36838 81186 37074
rect 81422 36838 81464 37074
rect 86468 37024 86788 38048
rect 86468 36960 86476 37024
rect 86540 36960 86556 37024
rect 86620 36960 86636 37024
rect 86700 36960 86716 37024
rect 86780 36960 86788 37024
rect 6612 36480 6932 36838
rect 6612 36416 6620 36480
rect 6684 36416 6700 36480
rect 6764 36416 6780 36480
rect 6844 36416 6860 36480
rect 6924 36416 6932 36480
rect 6612 35392 6932 36416
rect 86468 36414 86788 36960
rect 10484 36178 10526 36414
rect 10762 36178 10804 36414
rect 43084 36178 43126 36414
rect 43362 36178 43404 36414
rect 47884 36178 47926 36414
rect 48162 36178 48204 36414
rect 80484 36178 80526 36414
rect 80762 36178 80804 36414
rect 86468 36178 86510 36414
rect 86746 36178 86788 36414
rect 6612 35328 6620 35392
rect 6684 35328 6700 35392
rect 6764 35328 6780 35392
rect 6844 35328 6860 35392
rect 6924 35328 6932 35392
rect 6612 34304 6932 35328
rect 6612 34240 6620 34304
rect 6684 34240 6700 34304
rect 6764 34240 6780 34304
rect 6844 34240 6860 34304
rect 6924 34240 6932 34304
rect 6612 33216 6932 34240
rect 6612 33152 6620 33216
rect 6684 33152 6700 33216
rect 6764 33152 6780 33216
rect 6844 33152 6860 33216
rect 6924 33152 6932 33216
rect 6612 32128 6932 33152
rect 6612 32064 6620 32128
rect 6684 32064 6700 32128
rect 6764 32064 6780 32128
rect 6844 32064 6860 32128
rect 6924 32064 6932 32128
rect 6612 31040 6932 32064
rect 6612 30976 6620 31040
rect 6684 30976 6700 31040
rect 6764 30976 6780 31040
rect 6844 30976 6860 31040
rect 6924 30976 6932 31040
rect 6612 29952 6932 30976
rect 6612 29888 6620 29952
rect 6684 29888 6700 29952
rect 6764 29888 6780 29952
rect 6844 29888 6860 29952
rect 6924 29888 6932 29952
rect 6612 28864 6932 29888
rect 6612 28800 6620 28864
rect 6684 28800 6700 28864
rect 6764 28800 6780 28864
rect 6844 28800 6860 28864
rect 6924 28800 6932 28864
rect 6612 27776 6932 28800
rect 6612 27712 6620 27776
rect 6684 27712 6700 27776
rect 6764 27712 6780 27776
rect 6844 27712 6860 27776
rect 6924 27712 6932 27776
rect 6612 26688 6932 27712
rect 6612 26624 6620 26688
rect 6684 26624 6700 26688
rect 6764 26624 6780 26688
rect 6844 26624 6860 26688
rect 6924 26624 6932 26688
rect 6612 25600 6932 26624
rect 6612 25536 6620 25600
rect 6684 25536 6700 25600
rect 6764 25536 6780 25600
rect 6844 25536 6860 25600
rect 6924 25536 6932 25600
rect 6612 24512 6932 25536
rect 6612 24448 6620 24512
rect 6684 24448 6700 24512
rect 6764 24448 6780 24512
rect 6844 24448 6860 24512
rect 6924 24448 6932 24512
rect 6612 23424 6932 24448
rect 6612 23360 6620 23424
rect 6684 23360 6700 23424
rect 6764 23360 6780 23424
rect 6844 23360 6860 23424
rect 6924 23360 6932 23424
rect 6612 22336 6932 23360
rect 6612 22272 6620 22336
rect 6684 22272 6700 22336
rect 6764 22272 6780 22336
rect 6844 22272 6860 22336
rect 6924 22272 6932 22336
rect 6612 21248 6932 22272
rect 6612 21184 6620 21248
rect 6684 21184 6700 21248
rect 6764 21184 6780 21248
rect 6844 21184 6860 21248
rect 6924 21184 6932 21248
rect 6612 20160 6932 21184
rect 6612 20096 6620 20160
rect 6684 20096 6700 20160
rect 6764 20096 6780 20160
rect 6844 20096 6860 20160
rect 6924 20096 6932 20160
rect 6612 19072 6932 20096
rect 6612 19008 6620 19072
rect 6684 19008 6700 19072
rect 6764 19008 6780 19072
rect 6844 19008 6860 19072
rect 6924 19008 6932 19072
rect 6612 18674 6932 19008
rect 86468 35936 86788 36178
rect 86468 35872 86476 35936
rect 86540 35872 86556 35936
rect 86620 35872 86636 35936
rect 86700 35872 86716 35936
rect 86780 35872 86788 35936
rect 86468 34848 86788 35872
rect 86468 34784 86476 34848
rect 86540 34784 86556 34848
rect 86620 34784 86636 34848
rect 86700 34784 86716 34848
rect 86780 34784 86788 34848
rect 86468 33760 86788 34784
rect 86468 33696 86476 33760
rect 86540 33696 86556 33760
rect 86620 33696 86636 33760
rect 86700 33696 86716 33760
rect 86780 33696 86788 33760
rect 86468 32672 86788 33696
rect 86468 32608 86476 32672
rect 86540 32608 86556 32672
rect 86620 32608 86636 32672
rect 86700 32608 86716 32672
rect 86780 32608 86788 32672
rect 86468 31584 86788 32608
rect 86468 31520 86476 31584
rect 86540 31520 86556 31584
rect 86620 31520 86636 31584
rect 86700 31520 86716 31584
rect 86780 31520 86788 31584
rect 86468 30496 86788 31520
rect 86468 30432 86476 30496
rect 86540 30432 86556 30496
rect 86620 30432 86636 30496
rect 86700 30432 86716 30496
rect 86780 30432 86788 30496
rect 86468 29408 86788 30432
rect 86468 29344 86476 29408
rect 86540 29344 86556 29408
rect 86620 29344 86636 29408
rect 86700 29344 86716 29408
rect 86780 29344 86788 29408
rect 86468 28320 86788 29344
rect 86468 28256 86476 28320
rect 86540 28256 86556 28320
rect 86620 28256 86636 28320
rect 86700 28256 86716 28320
rect 86780 28256 86788 28320
rect 86468 27232 86788 28256
rect 86468 27168 86476 27232
rect 86540 27168 86556 27232
rect 86620 27168 86636 27232
rect 86700 27168 86716 27232
rect 86780 27168 86788 27232
rect 86468 26144 86788 27168
rect 86468 26080 86476 26144
rect 86540 26080 86556 26144
rect 86620 26080 86636 26144
rect 86700 26080 86716 26144
rect 86780 26080 86788 26144
rect 86468 25056 86788 26080
rect 86468 24992 86476 25056
rect 86540 24992 86556 25056
rect 86620 24992 86636 25056
rect 86700 24992 86716 25056
rect 86780 24992 86788 25056
rect 86468 23968 86788 24992
rect 86468 23904 86476 23968
rect 86540 23904 86556 23968
rect 86620 23904 86636 23968
rect 86700 23904 86716 23968
rect 86780 23904 86788 23968
rect 86468 22880 86788 23904
rect 86468 22816 86476 22880
rect 86540 22816 86556 22880
rect 86620 22816 86636 22880
rect 86700 22816 86716 22880
rect 86780 22816 86788 22880
rect 86468 21792 86788 22816
rect 86468 21728 86476 21792
rect 86540 21728 86556 21792
rect 86620 21728 86636 21792
rect 86700 21728 86716 21792
rect 86780 21728 86788 21792
rect 86468 20704 86788 21728
rect 86468 20640 86476 20704
rect 86540 20640 86556 20704
rect 86620 20640 86636 20704
rect 86700 20640 86716 20704
rect 86780 20640 86788 20704
rect 86468 19616 86788 20640
rect 86468 19552 86476 19616
rect 86540 19552 86556 19616
rect 86620 19552 86636 19616
rect 86700 19552 86716 19616
rect 86780 19552 86788 19616
rect 6612 18438 6654 18674
rect 6890 18438 6932 18674
rect 11144 18438 11186 18674
rect 11422 18438 11464 18674
rect 43744 18438 43786 18674
rect 44022 18438 44064 18674
rect 48544 18438 48586 18674
rect 48822 18438 48864 18674
rect 81144 18438 81186 18674
rect 81422 18438 81464 18674
rect 86468 18528 86788 19552
rect 86468 18464 86476 18528
rect 86540 18464 86556 18528
rect 86620 18464 86636 18528
rect 86700 18464 86716 18528
rect 86780 18464 86788 18528
rect 6612 17984 6932 18438
rect 86468 18014 86788 18464
rect 6612 17920 6620 17984
rect 6684 17920 6700 17984
rect 6764 17920 6780 17984
rect 6844 17920 6860 17984
rect 6924 17920 6932 17984
rect 6612 16896 6932 17920
rect 10484 17778 10526 18014
rect 10762 17778 10804 18014
rect 43084 17778 43126 18014
rect 43362 17778 43404 18014
rect 47884 17778 47926 18014
rect 48162 17778 48204 18014
rect 80484 17778 80526 18014
rect 80762 17778 80804 18014
rect 86468 17778 86510 18014
rect 86746 17778 86788 18014
rect 6612 16832 6620 16896
rect 6684 16832 6700 16896
rect 6764 16832 6780 16896
rect 6844 16832 6860 16896
rect 6924 16832 6932 16896
rect 6612 15808 6932 16832
rect 6612 15744 6620 15808
rect 6684 15744 6700 15808
rect 6764 15744 6780 15808
rect 6844 15744 6860 15808
rect 6924 15744 6932 15808
rect 6612 14720 6932 15744
rect 6612 14656 6620 14720
rect 6684 14656 6700 14720
rect 6764 14656 6780 14720
rect 6844 14656 6860 14720
rect 6924 14656 6932 14720
rect 6612 13632 6932 14656
rect 6612 13568 6620 13632
rect 6684 13568 6700 13632
rect 6764 13568 6780 13632
rect 6844 13568 6860 13632
rect 6924 13568 6932 13632
rect 6612 12544 6932 13568
rect 6612 12480 6620 12544
rect 6684 12480 6700 12544
rect 6764 12480 6780 12544
rect 6844 12480 6860 12544
rect 6924 12480 6932 12544
rect 6612 11456 6932 12480
rect 86468 17440 86788 17778
rect 86468 17376 86476 17440
rect 86540 17376 86556 17440
rect 86620 17376 86636 17440
rect 86700 17376 86716 17440
rect 86780 17376 86788 17440
rect 86468 16352 86788 17376
rect 86468 16288 86476 16352
rect 86540 16288 86556 16352
rect 86620 16288 86636 16352
rect 86700 16288 86716 16352
rect 86780 16288 86788 16352
rect 86468 15264 86788 16288
rect 86468 15200 86476 15264
rect 86540 15200 86556 15264
rect 86620 15200 86636 15264
rect 86700 15200 86716 15264
rect 86780 15200 86788 15264
rect 86468 14176 86788 15200
rect 86468 14112 86476 14176
rect 86540 14112 86556 14176
rect 86620 14112 86636 14176
rect 86700 14112 86716 14176
rect 86780 14112 86788 14176
rect 86468 13088 86788 14112
rect 86468 13024 86476 13088
rect 86540 13024 86556 13088
rect 86620 13024 86636 13088
rect 86700 13024 86716 13088
rect 86780 13024 86788 13088
rect 86468 12000 86788 13024
rect 86468 11936 86476 12000
rect 86540 11936 86556 12000
rect 86620 11936 86636 12000
rect 86700 11936 86716 12000
rect 86780 11936 86788 12000
rect 11144 11630 11186 11866
rect 11422 11630 11464 11866
rect 43744 11630 43786 11866
rect 44022 11630 44064 11866
rect 48544 11630 48586 11866
rect 48822 11630 48864 11866
rect 81144 11630 81186 11866
rect 81422 11630 81464 11866
rect 6612 11392 6620 11456
rect 6684 11392 6700 11456
rect 6764 11392 6780 11456
rect 6844 11392 6860 11456
rect 6924 11392 6932 11456
rect 6612 10368 6932 11392
rect 10484 10970 10526 11206
rect 10762 10970 10804 11206
rect 43084 10970 43126 11206
rect 43362 10970 43404 11206
rect 47884 10970 47926 11206
rect 48162 10970 48204 11206
rect 80484 10970 80526 11206
rect 80762 10970 80804 11206
rect 6612 10304 6620 10368
rect 6684 10304 6700 10368
rect 6764 10304 6780 10368
rect 6844 10304 6860 10368
rect 6924 10304 6932 10368
rect 6612 9280 6932 10304
rect 86468 10912 86788 11936
rect 86468 10848 86476 10912
rect 86540 10848 86556 10912
rect 86620 10848 86636 10912
rect 86700 10848 86716 10912
rect 86780 10848 86788 10912
rect 6612 9216 6620 9280
rect 6684 9216 6700 9280
rect 6764 9216 6780 9280
rect 6844 9216 6860 9280
rect 6924 9216 6932 9280
rect 6612 8192 6932 9216
rect 6612 8128 6620 8192
rect 6684 8128 6700 8192
rect 6764 8128 6780 8192
rect 6844 8128 6860 8192
rect 6924 8128 6932 8192
rect 6612 7104 6932 8128
rect 6612 7040 6620 7104
rect 6684 7040 6700 7104
rect 6764 7040 6780 7104
rect 6844 7040 6860 7104
rect 6924 7040 6932 7104
rect 6612 7024 6932 7040
rect 17716 7648 18036 10187
rect 17716 7584 17724 7648
rect 17788 7584 17804 7648
rect 17868 7584 17884 7648
rect 17948 7584 17964 7648
rect 18028 7584 18036 7648
rect 3356 3418 3398 3654
rect 3634 3418 3676 3654
rect 3356 3376 3676 3418
rect 17716 6560 18036 7584
rect 17716 6496 17724 6560
rect 17788 6496 17804 6560
rect 17868 6496 17884 6560
rect 17948 6496 17964 6560
rect 18028 6496 18036 6560
rect 17716 5472 18036 6496
rect 17716 5408 17724 5472
rect 17788 5408 17804 5472
rect 17868 5408 17884 5472
rect 17948 5408 17964 5472
rect 18028 5408 18036 5472
rect 17716 3654 18036 5408
rect 17716 3418 17758 3654
rect 17994 3418 18036 3654
rect 2696 2758 2738 2994
rect 2974 2758 3016 2994
rect 2696 2716 3016 2758
rect 17716 2716 18036 3418
rect 18376 7104 18696 10187
rect 18376 7040 18384 7104
rect 18448 7040 18464 7104
rect 18528 7040 18544 7104
rect 18608 7040 18624 7104
rect 18688 7040 18696 7104
rect 18376 6016 18696 7040
rect 18376 5952 18384 6016
rect 18448 5952 18464 6016
rect 18528 5952 18544 6016
rect 18608 5952 18624 6016
rect 18688 5952 18696 6016
rect 18376 4928 18696 5952
rect 18376 4864 18384 4928
rect 18448 4864 18464 4928
rect 18528 4864 18544 4928
rect 18608 4864 18624 4928
rect 18688 4864 18696 4928
rect 18376 2994 18696 4864
rect 18376 2758 18418 2994
rect 18654 2758 18696 2994
rect 18376 2716 18696 2758
rect 36116 7648 36436 10187
rect 36116 7584 36124 7648
rect 36188 7584 36204 7648
rect 36268 7584 36284 7648
rect 36348 7584 36364 7648
rect 36428 7584 36436 7648
rect 36116 6560 36436 7584
rect 36116 6496 36124 6560
rect 36188 6496 36204 6560
rect 36268 6496 36284 6560
rect 36348 6496 36364 6560
rect 36428 6496 36436 6560
rect 36116 5472 36436 6496
rect 36116 5408 36124 5472
rect 36188 5408 36204 5472
rect 36268 5408 36284 5472
rect 36348 5408 36364 5472
rect 36428 5408 36436 5472
rect 36116 3654 36436 5408
rect 36116 3418 36158 3654
rect 36394 3418 36436 3654
rect 36116 2716 36436 3418
rect 36776 7104 37096 10187
rect 36776 7040 36784 7104
rect 36848 7040 36864 7104
rect 36928 7040 36944 7104
rect 37008 7040 37024 7104
rect 37088 7040 37096 7104
rect 36776 6016 37096 7040
rect 36776 5952 36784 6016
rect 36848 5952 36864 6016
rect 36928 5952 36944 6016
rect 37008 5952 37024 6016
rect 37088 5952 37096 6016
rect 36776 4928 37096 5952
rect 36776 4864 36784 4928
rect 36848 4864 36864 4928
rect 36928 4864 36944 4928
rect 37008 4864 37024 4928
rect 37088 4864 37096 4928
rect 36776 2994 37096 4864
rect 36776 2758 36818 2994
rect 37054 2758 37096 2994
rect 36776 2716 37096 2758
rect 54516 7648 54836 10187
rect 54516 7584 54524 7648
rect 54588 7584 54604 7648
rect 54668 7584 54684 7648
rect 54748 7584 54764 7648
rect 54828 7584 54836 7648
rect 54516 6560 54836 7584
rect 54516 6496 54524 6560
rect 54588 6496 54604 6560
rect 54668 6496 54684 6560
rect 54748 6496 54764 6560
rect 54828 6496 54836 6560
rect 54516 5472 54836 6496
rect 54516 5408 54524 5472
rect 54588 5408 54604 5472
rect 54668 5408 54684 5472
rect 54748 5408 54764 5472
rect 54828 5408 54836 5472
rect 54516 3654 54836 5408
rect 54516 3418 54558 3654
rect 54794 3418 54836 3654
rect 54516 2716 54836 3418
rect 55176 7104 55496 10187
rect 55176 7040 55184 7104
rect 55248 7040 55264 7104
rect 55328 7040 55344 7104
rect 55408 7040 55424 7104
rect 55488 7040 55496 7104
rect 55176 6016 55496 7040
rect 55176 5952 55184 6016
rect 55248 5952 55264 6016
rect 55328 5952 55344 6016
rect 55408 5952 55424 6016
rect 55488 5952 55496 6016
rect 55176 4928 55496 5952
rect 55176 4864 55184 4928
rect 55248 4864 55264 4928
rect 55328 4864 55344 4928
rect 55408 4864 55424 4928
rect 55488 4864 55496 4928
rect 55176 2994 55496 4864
rect 55176 2758 55218 2994
rect 55454 2758 55496 2994
rect 55176 2716 55496 2758
rect 72916 7648 73236 10187
rect 72916 7584 72924 7648
rect 72988 7584 73004 7648
rect 73068 7584 73084 7648
rect 73148 7584 73164 7648
rect 73228 7584 73236 7648
rect 72916 6560 73236 7584
rect 72916 6496 72924 6560
rect 72988 6496 73004 6560
rect 73068 6496 73084 6560
rect 73148 6496 73164 6560
rect 73228 6496 73236 6560
rect 72916 5472 73236 6496
rect 72916 5408 72924 5472
rect 72988 5408 73004 5472
rect 73068 5408 73084 5472
rect 73148 5408 73164 5472
rect 73228 5408 73236 5472
rect 72916 3654 73236 5408
rect 72916 3418 72958 3654
rect 73194 3418 73236 3654
rect 72916 2716 73236 3418
rect 73576 7104 73896 10187
rect 73576 7040 73584 7104
rect 73648 7040 73664 7104
rect 73728 7040 73744 7104
rect 73808 7040 73824 7104
rect 73888 7040 73896 7104
rect 73576 6016 73896 7040
rect 86468 9824 86788 10848
rect 86468 9760 86476 9824
rect 86540 9760 86556 9824
rect 86620 9760 86636 9824
rect 86700 9760 86716 9824
rect 86780 9760 86788 9824
rect 86468 8736 86788 9760
rect 86468 8672 86476 8736
rect 86540 8672 86556 8736
rect 86620 8672 86636 8736
rect 86700 8672 86716 8736
rect 86780 8672 86788 8736
rect 86468 7648 86788 8672
rect 86468 7584 86476 7648
rect 86540 7584 86556 7648
rect 86620 7584 86636 7648
rect 86700 7584 86716 7648
rect 86780 7584 86788 7648
rect 86468 7024 86788 7584
rect 87204 84352 87524 84912
rect 87204 84288 87212 84352
rect 87276 84288 87292 84352
rect 87356 84288 87372 84352
rect 87436 84288 87452 84352
rect 87516 84288 87524 84352
rect 87204 83264 87524 84288
rect 87204 83200 87212 83264
rect 87276 83200 87292 83264
rect 87356 83200 87372 83264
rect 87436 83200 87452 83264
rect 87516 83200 87524 83264
rect 87204 82176 87524 83200
rect 87204 82112 87212 82176
rect 87276 82112 87292 82176
rect 87356 82112 87372 82176
rect 87436 82112 87452 82176
rect 87516 82112 87524 82176
rect 87204 81088 87524 82112
rect 87204 81024 87212 81088
rect 87276 81024 87292 81088
rect 87356 81024 87372 81088
rect 87436 81024 87452 81088
rect 87516 81024 87524 81088
rect 87204 80000 87524 81024
rect 87204 79936 87212 80000
rect 87276 79936 87292 80000
rect 87356 79936 87372 80000
rect 87436 79936 87452 80000
rect 87516 79936 87524 80000
rect 87204 78912 87524 79936
rect 87204 78848 87212 78912
rect 87276 78848 87292 78912
rect 87356 78848 87372 78912
rect 87436 78848 87452 78912
rect 87516 78848 87524 78912
rect 87204 77824 87524 78848
rect 87204 77760 87212 77824
rect 87276 77760 87292 77824
rect 87356 77760 87372 77824
rect 87436 77760 87452 77824
rect 87516 77760 87524 77824
rect 87204 76736 87524 77760
rect 87204 76672 87212 76736
rect 87276 76672 87292 76736
rect 87356 76672 87372 76736
rect 87436 76672 87452 76736
rect 87516 76672 87524 76736
rect 87204 75648 87524 76672
rect 87204 75584 87212 75648
rect 87276 75584 87292 75648
rect 87356 75584 87372 75648
rect 87436 75584 87452 75648
rect 87516 75584 87524 75648
rect 87204 74560 87524 75584
rect 87204 74496 87212 74560
rect 87276 74496 87292 74560
rect 87356 74496 87372 74560
rect 87436 74496 87452 74560
rect 87516 74496 87524 74560
rect 87204 73874 87524 74496
rect 87204 73638 87246 73874
rect 87482 73638 87524 73874
rect 87204 73472 87524 73638
rect 87204 73408 87212 73472
rect 87276 73408 87292 73472
rect 87356 73408 87372 73472
rect 87436 73408 87452 73472
rect 87516 73408 87524 73472
rect 87204 72384 87524 73408
rect 87204 72320 87212 72384
rect 87276 72320 87292 72384
rect 87356 72320 87372 72384
rect 87436 72320 87452 72384
rect 87516 72320 87524 72384
rect 87204 71296 87524 72320
rect 87204 71232 87212 71296
rect 87276 71232 87292 71296
rect 87356 71232 87372 71296
rect 87436 71232 87452 71296
rect 87516 71232 87524 71296
rect 87204 70208 87524 71232
rect 87204 70144 87212 70208
rect 87276 70144 87292 70208
rect 87356 70144 87372 70208
rect 87436 70144 87452 70208
rect 87516 70144 87524 70208
rect 87204 69120 87524 70144
rect 87204 69056 87212 69120
rect 87276 69056 87292 69120
rect 87356 69056 87372 69120
rect 87436 69056 87452 69120
rect 87516 69056 87524 69120
rect 87204 68032 87524 69056
rect 87204 67968 87212 68032
rect 87276 67968 87292 68032
rect 87356 67968 87372 68032
rect 87436 67968 87452 68032
rect 87516 67968 87524 68032
rect 87204 66944 87524 67968
rect 87204 66880 87212 66944
rect 87276 66880 87292 66944
rect 87356 66880 87372 66944
rect 87436 66880 87452 66944
rect 87516 66880 87524 66944
rect 87204 65856 87524 66880
rect 87204 65792 87212 65856
rect 87276 65792 87292 65856
rect 87356 65792 87372 65856
rect 87436 65792 87452 65856
rect 87516 65792 87524 65856
rect 87204 64768 87524 65792
rect 87204 64704 87212 64768
rect 87276 64704 87292 64768
rect 87356 64704 87372 64768
rect 87436 64704 87452 64768
rect 87516 64704 87524 64768
rect 87204 63680 87524 64704
rect 87204 63616 87212 63680
rect 87276 63616 87292 63680
rect 87356 63616 87372 63680
rect 87436 63616 87452 63680
rect 87516 63616 87524 63680
rect 87204 62592 87524 63616
rect 87204 62528 87212 62592
rect 87276 62528 87292 62592
rect 87356 62528 87372 62592
rect 87436 62528 87452 62592
rect 87516 62528 87524 62592
rect 87204 61504 87524 62528
rect 87204 61440 87212 61504
rect 87276 61440 87292 61504
rect 87356 61440 87372 61504
rect 87436 61440 87452 61504
rect 87516 61440 87524 61504
rect 87204 60416 87524 61440
rect 87204 60352 87212 60416
rect 87276 60352 87292 60416
rect 87356 60352 87372 60416
rect 87436 60352 87452 60416
rect 87516 60352 87524 60416
rect 87204 59328 87524 60352
rect 87204 59264 87212 59328
rect 87276 59264 87292 59328
rect 87356 59264 87372 59328
rect 87436 59264 87452 59328
rect 87516 59264 87524 59328
rect 87204 58240 87524 59264
rect 87204 58176 87212 58240
rect 87276 58176 87292 58240
rect 87356 58176 87372 58240
rect 87436 58176 87452 58240
rect 87516 58176 87524 58240
rect 87204 57152 87524 58176
rect 87204 57088 87212 57152
rect 87276 57088 87292 57152
rect 87356 57088 87372 57152
rect 87436 57088 87452 57152
rect 87516 57088 87524 57152
rect 87204 56064 87524 57088
rect 87204 56000 87212 56064
rect 87276 56000 87292 56064
rect 87356 56000 87372 56064
rect 87436 56000 87452 56064
rect 87516 56000 87524 56064
rect 87204 55474 87524 56000
rect 87204 55238 87246 55474
rect 87482 55238 87524 55474
rect 87204 54976 87524 55238
rect 87204 54912 87212 54976
rect 87276 54912 87292 54976
rect 87356 54912 87372 54976
rect 87436 54912 87452 54976
rect 87516 54912 87524 54976
rect 87204 53888 87524 54912
rect 87204 53824 87212 53888
rect 87276 53824 87292 53888
rect 87356 53824 87372 53888
rect 87436 53824 87452 53888
rect 87516 53824 87524 53888
rect 87204 52800 87524 53824
rect 87204 52736 87212 52800
rect 87276 52736 87292 52800
rect 87356 52736 87372 52800
rect 87436 52736 87452 52800
rect 87516 52736 87524 52800
rect 87204 51712 87524 52736
rect 87204 51648 87212 51712
rect 87276 51648 87292 51712
rect 87356 51648 87372 51712
rect 87436 51648 87452 51712
rect 87516 51648 87524 51712
rect 87204 50624 87524 51648
rect 87204 50560 87212 50624
rect 87276 50560 87292 50624
rect 87356 50560 87372 50624
rect 87436 50560 87452 50624
rect 87516 50560 87524 50624
rect 87204 49536 87524 50560
rect 87204 49472 87212 49536
rect 87276 49472 87292 49536
rect 87356 49472 87372 49536
rect 87436 49472 87452 49536
rect 87516 49472 87524 49536
rect 87204 48448 87524 49472
rect 87204 48384 87212 48448
rect 87276 48384 87292 48448
rect 87356 48384 87372 48448
rect 87436 48384 87452 48448
rect 87516 48384 87524 48448
rect 87204 47360 87524 48384
rect 87204 47296 87212 47360
rect 87276 47296 87292 47360
rect 87356 47296 87372 47360
rect 87436 47296 87452 47360
rect 87516 47296 87524 47360
rect 87204 46272 87524 47296
rect 87204 46208 87212 46272
rect 87276 46208 87292 46272
rect 87356 46208 87372 46272
rect 87436 46208 87452 46272
rect 87516 46208 87524 46272
rect 87204 45184 87524 46208
rect 87204 45120 87212 45184
rect 87276 45120 87292 45184
rect 87356 45120 87372 45184
rect 87436 45120 87452 45184
rect 87516 45120 87524 45184
rect 87204 44096 87524 45120
rect 87204 44032 87212 44096
rect 87276 44032 87292 44096
rect 87356 44032 87372 44096
rect 87436 44032 87452 44096
rect 87516 44032 87524 44096
rect 87204 43008 87524 44032
rect 87204 42944 87212 43008
rect 87276 42944 87292 43008
rect 87356 42944 87372 43008
rect 87436 42944 87452 43008
rect 87516 42944 87524 43008
rect 87204 41920 87524 42944
rect 87204 41856 87212 41920
rect 87276 41856 87292 41920
rect 87356 41856 87372 41920
rect 87436 41856 87452 41920
rect 87516 41856 87524 41920
rect 87204 40832 87524 41856
rect 87204 40768 87212 40832
rect 87276 40768 87292 40832
rect 87356 40768 87372 40832
rect 87436 40768 87452 40832
rect 87516 40768 87524 40832
rect 87204 39744 87524 40768
rect 87204 39680 87212 39744
rect 87276 39680 87292 39744
rect 87356 39680 87372 39744
rect 87436 39680 87452 39744
rect 87516 39680 87524 39744
rect 87204 38656 87524 39680
rect 87204 38592 87212 38656
rect 87276 38592 87292 38656
rect 87356 38592 87372 38656
rect 87436 38592 87452 38656
rect 87516 38592 87524 38656
rect 87204 37568 87524 38592
rect 87204 37504 87212 37568
rect 87276 37504 87292 37568
rect 87356 37504 87372 37568
rect 87436 37504 87452 37568
rect 87516 37504 87524 37568
rect 87204 37074 87524 37504
rect 87204 36838 87246 37074
rect 87482 36838 87524 37074
rect 87204 36480 87524 36838
rect 87204 36416 87212 36480
rect 87276 36416 87292 36480
rect 87356 36416 87372 36480
rect 87436 36416 87452 36480
rect 87516 36416 87524 36480
rect 87204 35392 87524 36416
rect 87204 35328 87212 35392
rect 87276 35328 87292 35392
rect 87356 35328 87372 35392
rect 87436 35328 87452 35392
rect 87516 35328 87524 35392
rect 87204 34304 87524 35328
rect 87204 34240 87212 34304
rect 87276 34240 87292 34304
rect 87356 34240 87372 34304
rect 87436 34240 87452 34304
rect 87516 34240 87524 34304
rect 87204 33216 87524 34240
rect 87204 33152 87212 33216
rect 87276 33152 87292 33216
rect 87356 33152 87372 33216
rect 87436 33152 87452 33216
rect 87516 33152 87524 33216
rect 87204 32128 87524 33152
rect 87204 32064 87212 32128
rect 87276 32064 87292 32128
rect 87356 32064 87372 32128
rect 87436 32064 87452 32128
rect 87516 32064 87524 32128
rect 87204 31040 87524 32064
rect 87204 30976 87212 31040
rect 87276 30976 87292 31040
rect 87356 30976 87372 31040
rect 87436 30976 87452 31040
rect 87516 30976 87524 31040
rect 87204 29952 87524 30976
rect 87204 29888 87212 29952
rect 87276 29888 87292 29952
rect 87356 29888 87372 29952
rect 87436 29888 87452 29952
rect 87516 29888 87524 29952
rect 87204 28864 87524 29888
rect 87204 28800 87212 28864
rect 87276 28800 87292 28864
rect 87356 28800 87372 28864
rect 87436 28800 87452 28864
rect 87516 28800 87524 28864
rect 87204 27776 87524 28800
rect 87204 27712 87212 27776
rect 87276 27712 87292 27776
rect 87356 27712 87372 27776
rect 87436 27712 87452 27776
rect 87516 27712 87524 27776
rect 87204 26688 87524 27712
rect 87204 26624 87212 26688
rect 87276 26624 87292 26688
rect 87356 26624 87372 26688
rect 87436 26624 87452 26688
rect 87516 26624 87524 26688
rect 87204 25600 87524 26624
rect 87204 25536 87212 25600
rect 87276 25536 87292 25600
rect 87356 25536 87372 25600
rect 87436 25536 87452 25600
rect 87516 25536 87524 25600
rect 87204 24512 87524 25536
rect 87204 24448 87212 24512
rect 87276 24448 87292 24512
rect 87356 24448 87372 24512
rect 87436 24448 87452 24512
rect 87516 24448 87524 24512
rect 87204 23424 87524 24448
rect 87204 23360 87212 23424
rect 87276 23360 87292 23424
rect 87356 23360 87372 23424
rect 87436 23360 87452 23424
rect 87516 23360 87524 23424
rect 87204 22336 87524 23360
rect 87204 22272 87212 22336
rect 87276 22272 87292 22336
rect 87356 22272 87372 22336
rect 87436 22272 87452 22336
rect 87516 22272 87524 22336
rect 87204 21248 87524 22272
rect 87204 21184 87212 21248
rect 87276 21184 87292 21248
rect 87356 21184 87372 21248
rect 87436 21184 87452 21248
rect 87516 21184 87524 21248
rect 87204 20160 87524 21184
rect 87204 20096 87212 20160
rect 87276 20096 87292 20160
rect 87356 20096 87372 20160
rect 87436 20096 87452 20160
rect 87516 20096 87524 20160
rect 87204 19072 87524 20096
rect 87204 19008 87212 19072
rect 87276 19008 87292 19072
rect 87356 19008 87372 19072
rect 87436 19008 87452 19072
rect 87516 19008 87524 19072
rect 87204 18674 87524 19008
rect 87204 18438 87246 18674
rect 87482 18438 87524 18674
rect 87204 17984 87524 18438
rect 87204 17920 87212 17984
rect 87276 17920 87292 17984
rect 87356 17920 87372 17984
rect 87436 17920 87452 17984
rect 87516 17920 87524 17984
rect 87204 16896 87524 17920
rect 87204 16832 87212 16896
rect 87276 16832 87292 16896
rect 87356 16832 87372 16896
rect 87436 16832 87452 16896
rect 87516 16832 87524 16896
rect 87204 15808 87524 16832
rect 87204 15744 87212 15808
rect 87276 15744 87292 15808
rect 87356 15744 87372 15808
rect 87436 15744 87452 15808
rect 87516 15744 87524 15808
rect 87204 14720 87524 15744
rect 87204 14656 87212 14720
rect 87276 14656 87292 14720
rect 87356 14656 87372 14720
rect 87436 14656 87452 14720
rect 87516 14656 87524 14720
rect 87204 13632 87524 14656
rect 87204 13568 87212 13632
rect 87276 13568 87292 13632
rect 87356 13568 87372 13632
rect 87436 13568 87452 13632
rect 87516 13568 87524 13632
rect 87204 12544 87524 13568
rect 87204 12480 87212 12544
rect 87276 12480 87292 12544
rect 87356 12480 87372 12544
rect 87436 12480 87452 12544
rect 87516 12480 87524 12544
rect 87204 11456 87524 12480
rect 87204 11392 87212 11456
rect 87276 11392 87292 11456
rect 87356 11392 87372 11456
rect 87436 11392 87452 11456
rect 87516 11392 87524 11456
rect 87204 10368 87524 11392
rect 87204 10304 87212 10368
rect 87276 10304 87292 10368
rect 87356 10304 87372 10368
rect 87436 10304 87452 10368
rect 87516 10304 87524 10368
rect 87204 9280 87524 10304
rect 87204 9216 87212 9280
rect 87276 9216 87292 9280
rect 87356 9216 87372 9280
rect 87436 9216 87452 9280
rect 87516 9216 87524 9280
rect 87204 8192 87524 9216
rect 87204 8128 87212 8192
rect 87276 8128 87292 8192
rect 87356 8128 87372 8192
rect 87436 8128 87452 8192
rect 87516 8128 87524 8192
rect 87204 7104 87524 8128
rect 87204 7040 87212 7104
rect 87276 7040 87292 7104
rect 87356 7040 87372 7104
rect 87436 7040 87452 7104
rect 87516 7040 87524 7104
rect 87204 7024 87524 7040
rect 89796 73214 90116 88826
rect 89796 72978 89838 73214
rect 90074 72978 90116 73214
rect 89796 54814 90116 72978
rect 89796 54578 89838 54814
rect 90074 54578 90116 54814
rect 89796 36414 90116 54578
rect 89796 36178 89838 36414
rect 90074 36178 90116 36414
rect 89796 18014 90116 36178
rect 89796 17778 89838 18014
rect 90074 17778 90116 18014
rect 73576 5952 73584 6016
rect 73648 5952 73664 6016
rect 73728 5952 73744 6016
rect 73808 5952 73824 6016
rect 73888 5952 73896 6016
rect 73576 4928 73896 5952
rect 73576 4864 73584 4928
rect 73648 4864 73664 4928
rect 73728 4864 73744 4928
rect 73808 4864 73824 4928
rect 73888 4864 73896 4928
rect 73576 2994 73896 4864
rect 89796 3654 90116 17778
rect 89796 3418 89838 3654
rect 90074 3418 90116 3654
rect 89796 3376 90116 3418
rect 90456 73874 90776 89486
rect 90456 73638 90498 73874
rect 90734 73638 90776 73874
rect 90456 55474 90776 73638
rect 90456 55238 90498 55474
rect 90734 55238 90776 55474
rect 90456 37074 90776 55238
rect 90456 36838 90498 37074
rect 90734 36838 90776 37074
rect 90456 18674 90776 36838
rect 90456 18438 90498 18674
rect 90734 18438 90776 18674
rect 73576 2758 73618 2994
rect 73854 2758 73896 2994
rect 73576 2716 73896 2758
rect 90456 2994 90776 18438
rect 90456 2758 90498 2994
rect 90734 2758 90776 2994
rect 90456 2716 90776 2758
<< via4 >>
rect 2738 89486 2974 89722
rect 2738 73638 2974 73874
rect 2738 55238 2974 55474
rect 2738 36838 2974 37074
rect 2738 18438 2974 18674
rect 3398 88826 3634 89062
rect 17758 88826 17994 89062
rect 3398 72978 3634 73214
rect 3398 54578 3634 54814
rect 3398 36178 3634 36414
rect 3398 17778 3634 18014
rect 5918 72978 6154 73214
rect 5918 54578 6154 54814
rect 5918 36178 6154 36414
rect 5918 17778 6154 18014
rect 18418 89486 18654 89722
rect 36158 88826 36394 89062
rect 36818 89486 37054 89722
rect 54558 88826 54794 89062
rect 55218 89486 55454 89722
rect 72958 88826 73194 89062
rect 73618 89486 73854 89722
rect 90498 89486 90734 89722
rect 89838 88826 90074 89062
rect 11186 80630 11422 80866
rect 43786 80630 44022 80866
rect 48586 80630 48822 80866
rect 81186 80630 81422 80866
rect 10526 79970 10762 80206
rect 43126 79970 43362 80206
rect 47926 79970 48162 80206
rect 80526 79970 80762 80206
rect 6654 73638 6890 73874
rect 11186 73638 11422 73874
rect 43786 73638 44022 73874
rect 48586 73638 48822 73874
rect 81186 73638 81422 73874
rect 10526 72978 10762 73214
rect 43126 72978 43362 73214
rect 47926 72978 48162 73214
rect 80526 72978 80762 73214
rect 86510 72978 86746 73214
rect 6654 55238 6890 55474
rect 11186 55238 11422 55474
rect 43786 55238 44022 55474
rect 48586 55238 48822 55474
rect 81186 55238 81422 55474
rect 10526 54578 10762 54814
rect 43126 54578 43362 54814
rect 47926 54578 48162 54814
rect 80526 54578 80762 54814
rect 86510 54578 86746 54814
rect 11186 48030 11422 48266
rect 43786 48030 44022 48266
rect 48586 48030 48822 48266
rect 81186 48030 81422 48266
rect 10526 47370 10762 47606
rect 43126 47370 43362 47606
rect 47926 47370 48162 47606
rect 80526 47370 80762 47606
rect 11186 44230 11422 44466
rect 43786 44230 44022 44466
rect 48586 44230 48822 44466
rect 81186 44230 81422 44466
rect 10526 43570 10762 43806
rect 43126 43570 43362 43806
rect 47926 43570 48162 43806
rect 80526 43570 80762 43806
rect 6654 36838 6890 37074
rect 11186 36838 11422 37074
rect 43786 36838 44022 37074
rect 48586 36838 48822 37074
rect 81186 36838 81422 37074
rect 10526 36178 10762 36414
rect 43126 36178 43362 36414
rect 47926 36178 48162 36414
rect 80526 36178 80762 36414
rect 86510 36178 86746 36414
rect 6654 18438 6890 18674
rect 11186 18438 11422 18674
rect 43786 18438 44022 18674
rect 48586 18438 48822 18674
rect 81186 18438 81422 18674
rect 10526 17778 10762 18014
rect 43126 17778 43362 18014
rect 47926 17778 48162 18014
rect 80526 17778 80762 18014
rect 86510 17778 86746 18014
rect 11186 11630 11422 11866
rect 43786 11630 44022 11866
rect 48586 11630 48822 11866
rect 81186 11630 81422 11866
rect 10526 10970 10762 11206
rect 43126 10970 43362 11206
rect 47926 10970 48162 11206
rect 80526 10970 80762 11206
rect 3398 3418 3634 3654
rect 17758 3418 17994 3654
rect 2738 2758 2974 2994
rect 18418 2758 18654 2994
rect 36158 3418 36394 3654
rect 36818 2758 37054 2994
rect 54558 3418 54794 3654
rect 55218 2758 55454 2994
rect 72958 3418 73194 3654
rect 87246 73638 87482 73874
rect 87246 55238 87482 55474
rect 87246 36838 87482 37074
rect 87246 18438 87482 18674
rect 89838 72978 90074 73214
rect 89838 54578 90074 54814
rect 89838 36178 90074 36414
rect 89838 17778 90074 18014
rect 89838 3418 90074 3654
rect 90498 73638 90734 73874
rect 90498 55238 90734 55474
rect 90498 36838 90734 37074
rect 90498 18438 90734 18674
rect 73618 2758 73854 2994
rect 90498 2758 90734 2994
<< metal5 >>
rect 2696 89722 90776 89764
rect 2696 89486 2738 89722
rect 2974 89486 18418 89722
rect 18654 89486 36818 89722
rect 37054 89486 55218 89722
rect 55454 89486 73618 89722
rect 73854 89486 90498 89722
rect 90734 89486 90776 89722
rect 2696 89444 90776 89486
rect 3356 89062 90116 89104
rect 3356 88826 3398 89062
rect 3634 88826 17758 89062
rect 17994 88826 36158 89062
rect 36394 88826 54558 89062
rect 54794 88826 72958 89062
rect 73194 88826 89838 89062
rect 90074 88826 90116 89062
rect 3356 88784 90116 88826
rect 11162 80866 11446 80908
rect 11162 80630 11186 80866
rect 11422 80630 11446 80866
rect 11162 80588 11446 80630
rect 43762 80866 44046 80908
rect 43762 80630 43786 80866
rect 44022 80630 44046 80866
rect 43762 80588 44046 80630
rect 48562 80866 48846 80908
rect 48562 80630 48586 80866
rect 48822 80630 48846 80866
rect 48562 80588 48846 80630
rect 81162 80866 81446 80908
rect 81162 80630 81186 80866
rect 81422 80630 81446 80866
rect 81162 80588 81446 80630
rect 10502 80206 10786 80248
rect 10502 79970 10526 80206
rect 10762 79970 10786 80206
rect 10502 79928 10786 79970
rect 43102 80206 43386 80248
rect 43102 79970 43126 80206
rect 43362 79970 43386 80206
rect 43102 79928 43386 79970
rect 47902 80206 48186 80248
rect 47902 79970 47926 80206
rect 48162 79970 48186 80206
rect 47902 79928 48186 79970
rect 80502 80206 80786 80248
rect 80502 79970 80526 80206
rect 80762 79970 80786 80206
rect 80502 79928 80786 79970
rect 2696 73874 90776 73916
rect 2696 73638 2738 73874
rect 2974 73638 6654 73874
rect 6890 73638 11186 73874
rect 11422 73638 43786 73874
rect 44022 73638 48586 73874
rect 48822 73638 81186 73874
rect 81422 73638 87246 73874
rect 87482 73638 90498 73874
rect 90734 73638 90776 73874
rect 2696 73596 90776 73638
rect 2696 73214 90776 73256
rect 2696 72978 3398 73214
rect 3634 72978 5918 73214
rect 6154 72978 10526 73214
rect 10762 72978 43126 73214
rect 43362 72978 47926 73214
rect 48162 72978 80526 73214
rect 80762 72978 86510 73214
rect 86746 72978 89838 73214
rect 90074 72978 90776 73214
rect 2696 72936 90776 72978
rect 2696 55474 90776 55516
rect 2696 55238 2738 55474
rect 2974 55238 6654 55474
rect 6890 55238 11186 55474
rect 11422 55238 43786 55474
rect 44022 55238 48586 55474
rect 48822 55238 81186 55474
rect 81422 55238 87246 55474
rect 87482 55238 90498 55474
rect 90734 55238 90776 55474
rect 2696 55196 90776 55238
rect 2696 54814 90776 54856
rect 2696 54578 3398 54814
rect 3634 54578 5918 54814
rect 6154 54578 10526 54814
rect 10762 54578 43126 54814
rect 43362 54578 47926 54814
rect 48162 54578 80526 54814
rect 80762 54578 86510 54814
rect 86746 54578 89838 54814
rect 90074 54578 90776 54814
rect 2696 54536 90776 54578
rect 11162 48266 11446 48308
rect 11162 48030 11186 48266
rect 11422 48030 11446 48266
rect 11162 47988 11446 48030
rect 43762 48266 44046 48308
rect 43762 48030 43786 48266
rect 44022 48030 44046 48266
rect 43762 47988 44046 48030
rect 48562 48266 48846 48308
rect 48562 48030 48586 48266
rect 48822 48030 48846 48266
rect 48562 47988 48846 48030
rect 81162 48266 81446 48308
rect 81162 48030 81186 48266
rect 81422 48030 81446 48266
rect 81162 47988 81446 48030
rect 10502 47606 10786 47648
rect 10502 47370 10526 47606
rect 10762 47370 10786 47606
rect 10502 47328 10786 47370
rect 43102 47606 43386 47648
rect 43102 47370 43126 47606
rect 43362 47370 43386 47606
rect 43102 47328 43386 47370
rect 47902 47606 48186 47648
rect 47902 47370 47926 47606
rect 48162 47370 48186 47606
rect 47902 47328 48186 47370
rect 80502 47606 80786 47648
rect 80502 47370 80526 47606
rect 80762 47370 80786 47606
rect 80502 47328 80786 47370
rect 11162 44466 11446 44508
rect 11162 44230 11186 44466
rect 11422 44230 11446 44466
rect 11162 44188 11446 44230
rect 43762 44466 44046 44508
rect 43762 44230 43786 44466
rect 44022 44230 44046 44466
rect 43762 44188 44046 44230
rect 48562 44466 48846 44508
rect 48562 44230 48586 44466
rect 48822 44230 48846 44466
rect 48562 44188 48846 44230
rect 81162 44466 81446 44508
rect 81162 44230 81186 44466
rect 81422 44230 81446 44466
rect 81162 44188 81446 44230
rect 10502 43806 10786 43848
rect 10502 43570 10526 43806
rect 10762 43570 10786 43806
rect 10502 43528 10786 43570
rect 43102 43806 43386 43848
rect 43102 43570 43126 43806
rect 43362 43570 43386 43806
rect 43102 43528 43386 43570
rect 47902 43806 48186 43848
rect 47902 43570 47926 43806
rect 48162 43570 48186 43806
rect 47902 43528 48186 43570
rect 80502 43806 80786 43848
rect 80502 43570 80526 43806
rect 80762 43570 80786 43806
rect 80502 43528 80786 43570
rect 2696 37074 90776 37116
rect 2696 36838 2738 37074
rect 2974 36838 6654 37074
rect 6890 36838 11186 37074
rect 11422 36838 43786 37074
rect 44022 36838 48586 37074
rect 48822 36838 81186 37074
rect 81422 36838 87246 37074
rect 87482 36838 90498 37074
rect 90734 36838 90776 37074
rect 2696 36796 90776 36838
rect 2696 36414 90776 36456
rect 2696 36178 3398 36414
rect 3634 36178 5918 36414
rect 6154 36178 10526 36414
rect 10762 36178 43126 36414
rect 43362 36178 47926 36414
rect 48162 36178 80526 36414
rect 80762 36178 86510 36414
rect 86746 36178 89838 36414
rect 90074 36178 90776 36414
rect 2696 36136 90776 36178
rect 2696 18674 90776 18716
rect 2696 18438 2738 18674
rect 2974 18438 6654 18674
rect 6890 18438 11186 18674
rect 11422 18438 43786 18674
rect 44022 18438 48586 18674
rect 48822 18438 81186 18674
rect 81422 18438 87246 18674
rect 87482 18438 90498 18674
rect 90734 18438 90776 18674
rect 2696 18396 90776 18438
rect 2696 18014 90776 18056
rect 2696 17778 3398 18014
rect 3634 17778 5918 18014
rect 6154 17778 10526 18014
rect 10762 17778 43126 18014
rect 43362 17778 47926 18014
rect 48162 17778 80526 18014
rect 80762 17778 86510 18014
rect 86746 17778 89838 18014
rect 90074 17778 90776 18014
rect 2696 17736 90776 17778
rect 11162 11866 11446 11908
rect 11162 11630 11186 11866
rect 11422 11630 11446 11866
rect 11162 11588 11446 11630
rect 43762 11866 44046 11908
rect 43762 11630 43786 11866
rect 44022 11630 44046 11866
rect 43762 11588 44046 11630
rect 48562 11866 48846 11908
rect 48562 11630 48586 11866
rect 48822 11630 48846 11866
rect 48562 11588 48846 11630
rect 81162 11866 81446 11908
rect 81162 11630 81186 11866
rect 81422 11630 81446 11866
rect 81162 11588 81446 11630
rect 10502 11206 10786 11248
rect 10502 10970 10526 11206
rect 10762 10970 10786 11206
rect 10502 10928 10786 10970
rect 43102 11206 43386 11248
rect 43102 10970 43126 11206
rect 43362 10970 43386 11206
rect 43102 10928 43386 10970
rect 47902 11206 48186 11248
rect 47902 10970 47926 11206
rect 48162 10970 48186 11206
rect 47902 10928 48186 10970
rect 80502 11206 80786 11248
rect 80502 10970 80526 11206
rect 80762 10970 80786 11206
rect 80502 10928 80786 10970
rect 3356 3654 90116 3696
rect 3356 3418 3398 3654
rect 3634 3418 17758 3654
rect 17994 3418 36158 3654
rect 36394 3418 54558 3654
rect 54794 3418 72958 3654
rect 73194 3418 89838 3654
rect 90074 3418 90116 3654
rect 3356 3376 90116 3418
rect 2696 2994 90776 3036
rect 2696 2758 2738 2994
rect 2974 2758 18418 2994
rect 18654 2758 36818 2994
rect 37054 2758 55218 2994
rect 55454 2758 73618 2994
rect 73854 2758 90498 2994
rect 90734 2758 90776 2994
rect 2696 2716 90776 2758
use sky130_fd_sc_hd__diode_2  ANTENNA_cell0_clk
timestamp 18001
transform 1 0 7268 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell0_config_data_out
timestamp 18001
transform -1 0 45540 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell0_config_en
timestamp 18001
transform -1 0 7268 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell0_le_clk
timestamp 18001
transform -1 0 45724 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell0_le_en
timestamp 18001
transform -1 0 45908 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell0_le_nrst
timestamp 18001
transform -1 0 46092 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell0_nrst
timestamp 18001
transform -1 0 7636 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell1_clk
timestamp 18001
transform -1 0 85744 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell1_config_data_in
timestamp 18001
transform -1 0 85928 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell1_config_data_out
timestamp 18001
transform -1 0 85744 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell1_config_en
timestamp 18001
transform -1 0 86112 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell1_le_clk
timestamp 18001
transform 1 0 85560 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell1_le_en
timestamp 18001
transform 1 0 85560 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell1_le_nrst
timestamp 18001
transform 1 0 85560 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell1_nrst
timestamp 18001
transform -1 0 86296 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell2_clk
timestamp 18001
transform -1 0 10764 0 1 84320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell2_config_data_in
timestamp 18001
transform -1 0 14076 0 1 84320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell2_config_data_out
timestamp 18001
transform -1 0 45540 0 1 84320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell2_config_en
timestamp 18001
transform 1 0 12788 0 1 84320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell2_le_clk
timestamp 18001
transform -1 0 45724 0 1 84320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell2_le_en
timestamp 18001
transform -1 0 45908 0 1 84320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell2_le_nrst
timestamp 18001
transform -1 0 46092 0 1 84320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell2_nrst
timestamp 18001
transform 1 0 11684 0 1 84320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell3_clk
timestamp 18001
transform -1 0 48208 0 1 84320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell3_config_data_in
timestamp 18001
transform -1 0 51520 0 1 84320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell3_config_en
timestamp 18001
transform 1 0 50232 0 1 84320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell3_le_clk
timestamp 18001
transform 1 0 85560 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell3_le_en
timestamp 18001
transform 1 0 85560 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell3_le_nrst
timestamp 18001
transform 1 0 85560 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell3_nrst
timestamp 18001
transform 1 0 49128 0 1 84320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 18001
transform 1 0 31004 0 1 84320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_X
timestamp 18001
transform -1 0 31004 0 1 84320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0__f_clk_A
timestamp 18001
transform 1 0 7452 0 -1 64736
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0__f_clk_X
timestamp 18001
transform 1 0 7452 0 -1 63648
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1__f_clk_A
timestamp 18001
transform -1 0 40940 0 1 84320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1__f_clk_X
timestamp 18001
transform -1 0 43056 0 1 84320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 18001
transform -1 0 5612 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 18001
transform -1 0 37720 0 1 86496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_X
timestamp 18001
transform 1 0 37720 0 1 86496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 18001
transform -1 0 88044 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 18001
transform -1 0 88044 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 18001
transform -1 0 88044 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 18001
transform -1 0 87860 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 18001
transform -1 0 87860 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 18001
transform -1 0 87860 0 1 66912
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 18001
transform -1 0 88044 0 -1 68000
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 18001
transform -1 0 87860 0 1 69088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 18001
transform -1 0 87860 0 1 70176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 18001
transform -1 0 88044 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 18001
transform -1 0 87860 0 1 71264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 18001
transform -1 0 87860 0 1 72352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 18001
transform -1 0 88044 0 -1 73440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 18001
transform -1 0 87860 0 1 74528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 18001
transform -1 0 87860 0 1 75616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 18001
transform -1 0 88136 0 1 76704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 18001
transform -1 0 87860 0 1 77792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 18001
transform -1 0 88044 0 -1 78880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 18001
transform -1 0 87860 0 1 79968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 18001
transform -1 0 87860 0 1 81056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 18001
transform -1 0 87860 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 18001
transform -1 0 88044 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 18001
transform -1 0 88044 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 18001
transform -1 0 88044 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 18001
transform -1 0 88044 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 18001
transform -1 0 87860 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 18001
transform -1 0 87952 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 18001
transform -1 0 88320 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 18001
transform -1 0 16652 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 18001
transform -1 0 26680 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 18001
transform -1 0 27324 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 18001
transform -1 0 28612 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 18001
transform -1 0 29900 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 18001
transform -1 0 54280 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 18001
transform -1 0 54096 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 18001
transform -1 0 55016 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 18001
transform -1 0 56304 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 18001
transform -1 0 16836 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 18001
transform -1 0 57592 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 18001
transform -1 0 58236 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 18001
transform -1 0 59524 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 18001
transform -1 0 60812 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 18001
transform -1 0 61456 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 18001
transform -1 0 62744 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 18001
transform -1 0 64032 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 18001
transform -1 0 65320 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 18001
transform -1 0 65964 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 18001
transform -1 0 67252 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 18001
transform -1 0 17664 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 18001
transform -1 0 18952 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 18001
transform -1 0 19596 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 18001
transform -1 0 20884 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 18001
transform -1 0 22172 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 18001
transform -1 0 23460 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 18001
transform -1 0 24104 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 18001
transform -1 0 25392 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 18001
transform -1 0 31188 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 18001
transform -1 0 42136 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 18001
transform -1 0 42780 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 18001
transform -1 0 44068 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 18001
transform -1 0 45356 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 18001
transform -1 0 68540 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 18001
transform -1 0 69184 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 18001
transform -1 0 70472 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 18001
transform -1 0 71760 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 18001
transform -1 0 31832 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 18001
transform -1 0 73048 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 18001
transform -1 0 73692 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 18001
transform -1 0 74980 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 18001
transform -1 0 76268 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 18001
transform -1 0 76912 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 18001
transform -1 0 78200 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 18001
transform -1 0 79488 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 18001
transform -1 0 80776 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input77_A
timestamp 18001
transform -1 0 81420 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input78_A
timestamp 18001
transform -1 0 87860 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 18001
transform -1 0 33120 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 18001
transform -1 0 34408 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input81_A
timestamp 18001
transform -1 0 35052 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input82_A
timestamp 18001
transform -1 0 36340 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input83_A
timestamp 18001
transform -1 0 37628 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input84_A
timestamp 18001
transform -1 0 38916 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input85_A
timestamp 18001
transform -1 0 39560 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input86_A
timestamp 18001
transform -1 0 40848 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input87_A
timestamp 18001
transform -1 0 5612 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input88_A
timestamp 18001
transform -1 0 5612 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input89_A
timestamp 18001
transform -1 0 5612 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input90_A
timestamp 18001
transform -1 0 5612 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input91_A
timestamp 18001
transform -1 0 5612 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input92_A
timestamp 18001
transform -1 0 5612 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input93_A
timestamp 18001
transform -1 0 5612 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input94_A
timestamp 18001
transform -1 0 5612 0 1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input95_A
timestamp 18001
transform -1 0 5612 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input96_A
timestamp 18001
transform -1 0 5612 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input97_A
timestamp 18001
transform -1 0 5612 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input98_A
timestamp 18001
transform -1 0 5612 0 -1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input99_A
timestamp 18001
transform -1 0 5612 0 1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input100_A
timestamp 18001
transform -1 0 5612 0 1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input101_A
timestamp 18001
transform -1 0 5612 0 1 60384
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input102_A
timestamp 18001
transform -1 0 5612 0 1 61472
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input103_A
timestamp 18001
transform -1 0 5612 0 -1 62560
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input104_A
timestamp 18001
transform -1 0 5612 0 1 63648
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input105_A
timestamp 18001
transform -1 0 5612 0 1 64736
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input106_A
timestamp 18001
transform -1 0 5612 0 1 65824
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input107_A
timestamp 18001
transform -1 0 5612 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input108_A
timestamp 18001
transform -1 0 5612 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input109_A
timestamp 18001
transform -1 0 5612 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input110_A
timestamp 18001
transform -1 0 5612 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input111_A
timestamp 18001
transform -1 0 5612 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input112_A
timestamp 18001
transform -1 0 5612 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input113_A
timestamp 18001
transform -1 0 5612 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input114_A
timestamp 18001
transform -1 0 5612 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input115_A
timestamp 18001
transform -1 0 88136 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input115_X
timestamp 18001
transform -1 0 88228 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input116_A
timestamp 18001
transform -1 0 87768 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input116_X
timestamp 18001
transform -1 0 88320 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input117_A
timestamp 18001
transform -1 0 88136 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input117_X
timestamp 18001
transform -1 0 88320 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input118_A
timestamp 18001
transform -1 0 38640 0 1 86496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input118_X
timestamp 18001
transform 1 0 39836 0 -1 87584
box -38 -48 222 592
use fpgacell  cell0
timestamp 0
transform 1 0 10000 0 1 10000
box 0 0 1 1
use fpgacell  cell1
timestamp 0
transform 1 0 47400 0 1 10000
box 0 0 1 1
use fpgacell  cell2
timestamp 0
transform 1 0 10000 0 1 46400
box 0 0 1 1
use fpgacell  cell3
timestamp 0
transform 1 0 47400 0 1 46400
box 0 0 1 1
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 18001
transform -1 0 30636 0 1 84320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 18001
transform -1 0 7452 0 1 63648
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 18001
transform 1 0 41032 0 1 84320
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3
timestamp 1636986456
transform 1 0 5152 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1636986456
transform 1 0 6256 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp 18001
transform 1 0 7360 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1636986456
transform 1 0 7544 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1636986456
transform 1 0 8648 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp 18001
transform 1 0 9752 0 1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1636986456
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1636986456
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 18001
transform 1 0 12328 0 1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1636986456
transform 1 0 12696 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1636986456
transform 1 0 13800 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 18001
transform 1 0 14904 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_117
timestamp 18001
transform 1 0 15640 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_124
timestamp 18001
transform 1 0 16284 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_132
timestamp 18001
transform 1 0 17020 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 18001
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_141
timestamp 18001
transform 1 0 17848 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_147
timestamp 18001
transform 1 0 18400 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_152
timestamp 18001
transform 1 0 18860 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_159
timestamp 18001
transform 1 0 19504 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 18001
transform 1 0 20240 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_173
timestamp 18001
transform 1 0 20792 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_181
timestamp 18001
transform 1 0 21528 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_187
timestamp 18001
transform 1 0 22080 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 18001
transform 1 0 22816 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_201
timestamp 18001
transform 1 0 23368 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_208
timestamp 18001
transform 1 0 24012 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_216
timestamp 18001
transform 1 0 24748 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 18001
transform 1 0 25300 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_225
timestamp 18001
transform 1 0 25576 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_231
timestamp 18001
transform 1 0 26128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_236
timestamp 18001
transform 1 0 26588 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_243
timestamp 18001
transform 1 0 27232 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 18001
transform 1 0 27968 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_257
timestamp 18001
transform 1 0 28520 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_265
timestamp 18001
transform 1 0 29256 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_271
timestamp 18001
transform 1 0 29808 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_279
timestamp 18001
transform 1 0 30544 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_286
timestamp 18001
transform 1 0 31188 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_293
timestamp 18001
transform 1 0 31832 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_301
timestamp 18001
transform 1 0 32568 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 18001
transform 1 0 33120 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_309
timestamp 18001
transform 1 0 33304 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_315
timestamp 18001
transform 1 0 33856 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_321
timestamp 18001
transform 1 0 34408 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_328
timestamp 18001
transform 1 0 35052 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_342
timestamp 18001
transform 1 0 36340 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_350
timestamp 18001
transform 1 0 37076 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_356
timestamp 18001
transform 1 0 37628 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_370
timestamp 18001
transform 1 0 38916 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_377
timestamp 18001
transform 1 0 39560 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_385
timestamp 18001
transform 1 0 40296 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_391
timestamp 18001
transform 1 0 40848 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_393
timestamp 18001
transform 1 0 41032 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_399
timestamp 18001
transform 1 0 41584 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_405
timestamp 18001
transform 1 0 42136 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_412
timestamp 18001
transform 1 0 42780 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_426
timestamp 18001
transform 1 0 44068 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_434
timestamp 18001
transform 1 0 44804 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_440
timestamp 18001
transform 1 0 45356 0 1 4896
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_449
timestamp 1636986456
transform 1 0 46184 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_461
timestamp 1636986456
transform 1 0 47288 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_473
timestamp 18001
transform 1 0 48392 0 1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_477
timestamp 1636986456
transform 1 0 48760 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_489
timestamp 1636986456
transform 1 0 49864 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_501
timestamp 18001
transform 1 0 50968 0 1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_505
timestamp 1636986456
transform 1 0 51336 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_517
timestamp 18001
transform 1 0 52440 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_523
timestamp 18001
transform 1 0 52992 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_530
timestamp 18001
transform 1 0 53636 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_533
timestamp 18001
transform 1 0 53912 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_539
timestamp 18001
transform 1 0 54464 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_544
timestamp 18001
transform 1 0 54924 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_552
timestamp 18001
transform 1 0 55660 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_558
timestamp 18001
transform 1 0 56212 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_561
timestamp 18001
transform 1 0 56488 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_567
timestamp 18001
transform 1 0 57040 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_572
timestamp 18001
transform 1 0 57500 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_579
timestamp 18001
transform 1 0 58144 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_587
timestamp 18001
transform 1 0 58880 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_593
timestamp 18001
transform 1 0 59432 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_601
timestamp 18001
transform 1 0 60168 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_607
timestamp 18001
transform 1 0 60720 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_614
timestamp 18001
transform 1 0 61364 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_617
timestamp 18001
transform 1 0 61640 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_623
timestamp 18001
transform 1 0 62192 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_628
timestamp 18001
transform 1 0 62652 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_636
timestamp 18001
transform 1 0 63388 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_642
timestamp 18001
transform 1 0 63940 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_645
timestamp 18001
transform 1 0 64216 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_651
timestamp 18001
transform 1 0 64768 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_656
timestamp 18001
transform 1 0 65228 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_663
timestamp 18001
transform 1 0 65872 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_671
timestamp 18001
transform 1 0 66608 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_677
timestamp 18001
transform 1 0 67160 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_685
timestamp 18001
transform 1 0 67896 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_692
timestamp 18001
transform 1 0 68540 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_699
timestamp 18001
transform 1 0 69184 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_701
timestamp 18001
transform 1 0 69368 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_707
timestamp 18001
transform 1 0 69920 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_713
timestamp 18001
transform 1 0 70472 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_721
timestamp 18001
transform 1 0 71208 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_727
timestamp 18001
transform 1 0 71760 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_729
timestamp 18001
transform 1 0 71944 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_735
timestamp 18001
transform 1 0 72496 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_741
timestamp 18001
transform 1 0 73048 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_748
timestamp 18001
transform 1 0 73692 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_762
timestamp 18001
transform 1 0 74980 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_770
timestamp 18001
transform 1 0 75716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_776
timestamp 18001
transform 1 0 76268 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_783
timestamp 18001
transform 1 0 76912 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_785
timestamp 18001
transform 1 0 77096 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_791
timestamp 18001
transform 1 0 77648 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_797
timestamp 18001
transform 1 0 78200 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_805
timestamp 18001
transform 1 0 78936 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_811
timestamp 18001
transform 1 0 79488 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_813
timestamp 18001
transform 1 0 79672 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_819
timestamp 18001
transform 1 0 80224 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_825
timestamp 18001
transform 1 0 80776 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_832
timestamp 18001
transform 1 0 81420 0 1 4896
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_841
timestamp 1636986456
transform 1 0 82248 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_853
timestamp 1636986456
transform 1 0 83352 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_865
timestamp 18001
transform 1 0 84456 0 1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_869
timestamp 1636986456
transform 1 0 84824 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_881
timestamp 1636986456
transform 1 0 85928 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_893
timestamp 18001
transform 1 0 87032 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_897
timestamp 18001
transform 1 0 87400 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_905
timestamp 18001
transform 1 0 88136 0 1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1636986456
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1636986456
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1636986456
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1636986456
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 18001
transform 1 0 9568 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 18001
transform 1 0 9936 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1636986456
transform 1 0 10120 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1636986456
transform 1 0 11224 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1636986456
transform 1 0 12328 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1636986456
transform 1 0 13432 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 18001
transform 1 0 14536 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 18001
transform 1 0 15088 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1636986456
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1636986456
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1636986456
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1636986456
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 18001
transform 1 0 19688 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 18001
transform 1 0 20240 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1636986456
transform 1 0 20424 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1636986456
transform 1 0 21528 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1636986456
transform 1 0 22632 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1636986456
transform 1 0 23736 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 18001
transform 1 0 24840 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 18001
transform 1 0 25392 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1636986456
transform 1 0 25576 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1636986456
transform 1 0 26680 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1636986456
transform 1 0 27784 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1636986456
transform 1 0 28888 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 18001
transform 1 0 29992 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 18001
transform 1 0 30544 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1636986456
transform 1 0 30728 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1636986456
transform 1 0 31832 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1636986456
transform 1 0 32936 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1636986456
transform 1 0 34040 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 18001
transform 1 0 35144 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 18001
transform 1 0 35696 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1636986456
transform 1 0 35880 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1636986456
transform 1 0 36984 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1636986456
transform 1 0 38088 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1636986456
transform 1 0 39192 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 18001
transform 1 0 40296 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 18001
transform 1 0 40848 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1636986456
transform 1 0 41032 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_405
timestamp 1636986456
transform 1 0 42136 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_417
timestamp 1636986456
transform 1 0 43240 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_429
timestamp 1636986456
transform 1 0 44344 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 18001
transform 1 0 45448 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 18001
transform 1 0 46000 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_449
timestamp 1636986456
transform 1 0 46184 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_461
timestamp 1636986456
transform 1 0 47288 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_473
timestamp 1636986456
transform 1 0 48392 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_485
timestamp 1636986456
transform 1 0 49496 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_497
timestamp 18001
transform 1 0 50600 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 18001
transform 1 0 51152 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_505
timestamp 1636986456
transform 1 0 51336 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_517
timestamp 1636986456
transform 1 0 52440 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_529
timestamp 1636986456
transform 1 0 53544 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_541
timestamp 1636986456
transform 1 0 54648 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_553
timestamp 18001
transform 1 0 55752 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_559
timestamp 18001
transform 1 0 56304 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_561
timestamp 1636986456
transform 1 0 56488 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_573
timestamp 1636986456
transform 1 0 57592 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_585
timestamp 1636986456
transform 1 0 58696 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_597
timestamp 1636986456
transform 1 0 59800 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_609
timestamp 18001
transform 1 0 60904 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_615
timestamp 18001
transform 1 0 61456 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_617
timestamp 1636986456
transform 1 0 61640 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_629
timestamp 1636986456
transform 1 0 62744 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_641
timestamp 1636986456
transform 1 0 63848 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_653
timestamp 1636986456
transform 1 0 64952 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_665
timestamp 18001
transform 1 0 66056 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_671
timestamp 18001
transform 1 0 66608 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_673
timestamp 1636986456
transform 1 0 66792 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_685
timestamp 1636986456
transform 1 0 67896 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_697
timestamp 1636986456
transform 1 0 69000 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_709
timestamp 1636986456
transform 1 0 70104 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_721
timestamp 18001
transform 1 0 71208 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_727
timestamp 18001
transform 1 0 71760 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_729
timestamp 1636986456
transform 1 0 71944 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_741
timestamp 1636986456
transform 1 0 73048 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_753
timestamp 1636986456
transform 1 0 74152 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_765
timestamp 1636986456
transform 1 0 75256 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_777
timestamp 18001
transform 1 0 76360 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_783
timestamp 18001
transform 1 0 76912 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_785
timestamp 1636986456
transform 1 0 77096 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_797
timestamp 1636986456
transform 1 0 78200 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_809
timestamp 1636986456
transform 1 0 79304 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_821
timestamp 1636986456
transform 1 0 80408 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_833
timestamp 18001
transform 1 0 81512 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_839
timestamp 18001
transform 1 0 82064 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_841
timestamp 1636986456
transform 1 0 82248 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_853
timestamp 1636986456
transform 1 0 83352 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_865
timestamp 1636986456
transform 1 0 84456 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_877
timestamp 1636986456
transform 1 0 85560 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_889
timestamp 18001
transform 1 0 86664 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_895
timestamp 18001
transform 1 0 87216 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_897
timestamp 18001
transform 1 0 87400 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_905
timestamp 18001
transform 1 0 88136 0 -1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1636986456
transform 1 0 5152 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1636986456
transform 1 0 6256 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 18001
transform 1 0 7360 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1636986456
transform 1 0 7544 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1636986456
transform 1 0 8648 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1636986456
transform 1 0 9752 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1636986456
transform 1 0 10856 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 18001
transform 1 0 11960 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 18001
transform 1 0 12512 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1636986456
transform 1 0 12696 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1636986456
transform 1 0 13800 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1636986456
transform 1 0 14904 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1636986456
transform 1 0 16008 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 18001
transform 1 0 17112 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 18001
transform 1 0 17664 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1636986456
transform 1 0 17848 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1636986456
transform 1 0 18952 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1636986456
transform 1 0 20056 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1636986456
transform 1 0 21160 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 18001
transform 1 0 22264 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 18001
transform 1 0 22816 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1636986456
transform 1 0 23000 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1636986456
transform 1 0 24104 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1636986456
transform 1 0 25208 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1636986456
transform 1 0 26312 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 18001
transform 1 0 27416 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 18001
transform 1 0 27968 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1636986456
transform 1 0 28152 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1636986456
transform 1 0 29256 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1636986456
transform 1 0 30360 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1636986456
transform 1 0 31464 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 18001
transform 1 0 32568 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 18001
transform 1 0 33120 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1636986456
transform 1 0 33304 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1636986456
transform 1 0 34408 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1636986456
transform 1 0 35512 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1636986456
transform 1 0 36616 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 18001
transform 1 0 37720 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 18001
transform 1 0 38272 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1636986456
transform 1 0 38456 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1636986456
transform 1 0 39560 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1636986456
transform 1 0 40664 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1636986456
transform 1 0 41768 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 18001
transform 1 0 42872 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 18001
transform 1 0 43424 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1636986456
transform 1 0 43608 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1636986456
transform 1 0 44712 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 1636986456
transform 1 0 45816 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_457
timestamp 1636986456
transform 1 0 46920 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 18001
transform 1 0 48024 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 18001
transform 1 0 48576 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_477
timestamp 1636986456
transform 1 0 48760 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_489
timestamp 1636986456
transform 1 0 49864 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_501
timestamp 1636986456
transform 1 0 50968 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_513
timestamp 1636986456
transform 1 0 52072 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_525
timestamp 18001
transform 1 0 53176 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 18001
transform 1 0 53728 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_533
timestamp 1636986456
transform 1 0 53912 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_545
timestamp 1636986456
transform 1 0 55016 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_557
timestamp 1636986456
transform 1 0 56120 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_569
timestamp 1636986456
transform 1 0 57224 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_581
timestamp 18001
transform 1 0 58328 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 18001
transform 1 0 58880 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_589
timestamp 1636986456
transform 1 0 59064 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_601
timestamp 1636986456
transform 1 0 60168 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_613
timestamp 1636986456
transform 1 0 61272 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_625
timestamp 1636986456
transform 1 0 62376 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_637
timestamp 18001
transform 1 0 63480 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_643
timestamp 18001
transform 1 0 64032 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_645
timestamp 1636986456
transform 1 0 64216 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_657
timestamp 1636986456
transform 1 0 65320 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_669
timestamp 1636986456
transform 1 0 66424 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_681
timestamp 1636986456
transform 1 0 67528 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_693
timestamp 18001
transform 1 0 68632 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_699
timestamp 18001
transform 1 0 69184 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_701
timestamp 1636986456
transform 1 0 69368 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_713
timestamp 1636986456
transform 1 0 70472 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_725
timestamp 1636986456
transform 1 0 71576 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_737
timestamp 1636986456
transform 1 0 72680 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_749
timestamp 18001
transform 1 0 73784 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_755
timestamp 18001
transform 1 0 74336 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_757
timestamp 1636986456
transform 1 0 74520 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_769
timestamp 1636986456
transform 1 0 75624 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_781
timestamp 1636986456
transform 1 0 76728 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_793
timestamp 1636986456
transform 1 0 77832 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_805
timestamp 18001
transform 1 0 78936 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_811
timestamp 18001
transform 1 0 79488 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_813
timestamp 1636986456
transform 1 0 79672 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_825
timestamp 1636986456
transform 1 0 80776 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_837
timestamp 1636986456
transform 1 0 81880 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_849
timestamp 1636986456
transform 1 0 82984 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_861
timestamp 18001
transform 1 0 84088 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_867
timestamp 18001
transform 1 0 84640 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_869
timestamp 1636986456
transform 1 0 84824 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_881
timestamp 1636986456
transform 1 0 85928 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_893
timestamp 1636986456
transform 1 0 87032 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_905
timestamp 18001
transform 1 0 88136 0 1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1636986456
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1636986456
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1636986456
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1636986456
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 18001
transform 1 0 9568 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 18001
transform 1 0 9936 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1636986456
transform 1 0 10120 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1636986456
transform 1 0 11224 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1636986456
transform 1 0 12328 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1636986456
transform 1 0 13432 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 18001
transform 1 0 14536 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 18001
transform 1 0 15088 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1636986456
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1636986456
transform 1 0 16376 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1636986456
transform 1 0 17480 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1636986456
transform 1 0 18584 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 18001
transform 1 0 19688 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 18001
transform 1 0 20240 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1636986456
transform 1 0 20424 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1636986456
transform 1 0 21528 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1636986456
transform 1 0 22632 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1636986456
transform 1 0 23736 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 18001
transform 1 0 24840 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 18001
transform 1 0 25392 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1636986456
transform 1 0 25576 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1636986456
transform 1 0 26680 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1636986456
transform 1 0 27784 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1636986456
transform 1 0 28888 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 18001
transform 1 0 29992 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 18001
transform 1 0 30544 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1636986456
transform 1 0 30728 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1636986456
transform 1 0 31832 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1636986456
transform 1 0 32936 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1636986456
transform 1 0 34040 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 18001
transform 1 0 35144 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 18001
transform 1 0 35696 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1636986456
transform 1 0 35880 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1636986456
transform 1 0 36984 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1636986456
transform 1 0 38088 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1636986456
transform 1 0 39192 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 18001
transform 1 0 40296 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 18001
transform 1 0 40848 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1636986456
transform 1 0 41032 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1636986456
transform 1 0 42136 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1636986456
transform 1 0 43240 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1636986456
transform 1 0 44344 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 18001
transform 1 0 45448 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 18001
transform 1 0 46000 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1636986456
transform 1 0 46184 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1636986456
transform 1 0 47288 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1636986456
transform 1 0 48392 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1636986456
transform 1 0 49496 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 18001
transform 1 0 50600 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 18001
transform 1 0 51152 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_505
timestamp 1636986456
transform 1 0 51336 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_517
timestamp 1636986456
transform 1 0 52440 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_529
timestamp 1636986456
transform 1 0 53544 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_541
timestamp 1636986456
transform 1 0 54648 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_553
timestamp 18001
transform 1 0 55752 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 18001
transform 1 0 56304 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_561
timestamp 1636986456
transform 1 0 56488 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_573
timestamp 1636986456
transform 1 0 57592 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_585
timestamp 1636986456
transform 1 0 58696 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_597
timestamp 1636986456
transform 1 0 59800 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_609
timestamp 18001
transform 1 0 60904 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 18001
transform 1 0 61456 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_617
timestamp 1636986456
transform 1 0 61640 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_629
timestamp 1636986456
transform 1 0 62744 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_641
timestamp 1636986456
transform 1 0 63848 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_653
timestamp 1636986456
transform 1 0 64952 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_665
timestamp 18001
transform 1 0 66056 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_671
timestamp 18001
transform 1 0 66608 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_673
timestamp 1636986456
transform 1 0 66792 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_685
timestamp 1636986456
transform 1 0 67896 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_697
timestamp 1636986456
transform 1 0 69000 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_709
timestamp 1636986456
transform 1 0 70104 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_721
timestamp 18001
transform 1 0 71208 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_727
timestamp 18001
transform 1 0 71760 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_729
timestamp 1636986456
transform 1 0 71944 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_741
timestamp 1636986456
transform 1 0 73048 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_753
timestamp 1636986456
transform 1 0 74152 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_765
timestamp 1636986456
transform 1 0 75256 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_777
timestamp 18001
transform 1 0 76360 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_783
timestamp 18001
transform 1 0 76912 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_785
timestamp 1636986456
transform 1 0 77096 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_797
timestamp 1636986456
transform 1 0 78200 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_809
timestamp 1636986456
transform 1 0 79304 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_821
timestamp 1636986456
transform 1 0 80408 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_833
timestamp 18001
transform 1 0 81512 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_839
timestamp 18001
transform 1 0 82064 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_841
timestamp 1636986456
transform 1 0 82248 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_853
timestamp 1636986456
transform 1 0 83352 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_865
timestamp 1636986456
transform 1 0 84456 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_877
timestamp 1636986456
transform 1 0 85560 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_889
timestamp 18001
transform 1 0 86664 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_895
timestamp 18001
transform 1 0 87216 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_897
timestamp 18001
transform 1 0 87400 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_905
timestamp 18001
transform 1 0 88136 0 -1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1636986456
transform 1 0 5152 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1636986456
transform 1 0 6256 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 18001
transform 1 0 7360 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1636986456
transform 1 0 7544 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1636986456
transform 1 0 8648 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_53
timestamp 18001
transform 1 0 9752 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_57
timestamp 1636986456
transform 1 0 10120 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_69
timestamp 1636986456
transform 1 0 11224 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_81
timestamp 18001
transform 1 0 12328 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1636986456
transform 1 0 12696 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1636986456
transform 1 0 13800 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_109
timestamp 18001
transform 1 0 14904 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_113
timestamp 1636986456
transform 1 0 15272 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_125
timestamp 1636986456
transform 1 0 16376 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_137
timestamp 18001
transform 1 0 17480 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1636986456
transform 1 0 17848 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1636986456
transform 1 0 18952 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_165
timestamp 18001
transform 1 0 20056 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_169
timestamp 1636986456
transform 1 0 20424 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_181
timestamp 1636986456
transform 1 0 21528 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_193
timestamp 18001
transform 1 0 22632 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1636986456
transform 1 0 23000 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1636986456
transform 1 0 24104 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_221
timestamp 18001
transform 1 0 25208 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_225
timestamp 1636986456
transform 1 0 25576 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_237
timestamp 1636986456
transform 1 0 26680 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_249
timestamp 18001
transform 1 0 27784 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1636986456
transform 1 0 28152 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1636986456
transform 1 0 29256 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_277
timestamp 18001
transform 1 0 30360 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_281
timestamp 1636986456
transform 1 0 30728 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_293
timestamp 1636986456
transform 1 0 31832 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_305
timestamp 18001
transform 1 0 32936 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1636986456
transform 1 0 33304 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1636986456
transform 1 0 34408 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_333
timestamp 18001
transform 1 0 35512 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_337
timestamp 1636986456
transform 1 0 35880 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_349
timestamp 1636986456
transform 1 0 36984 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_361
timestamp 18001
transform 1 0 38088 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1636986456
transform 1 0 38456 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1636986456
transform 1 0 39560 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_389
timestamp 18001
transform 1 0 40664 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_393
timestamp 1636986456
transform 1 0 41032 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_405
timestamp 1636986456
transform 1 0 42136 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_417
timestamp 18001
transform 1 0 43240 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1636986456
transform 1 0 43608 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_433
timestamp 18001
transform 1 0 44712 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_439
timestamp 18001
transform 1 0 45264 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_449
timestamp 1636986456
transform 1 0 46184 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_461
timestamp 1636986456
transform 1 0 47288 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_473
timestamp 18001
transform 1 0 48392 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1636986456
transform 1 0 48760 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1636986456
transform 1 0 49864 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_501
timestamp 18001
transform 1 0 50968 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_505
timestamp 1636986456
transform 1 0 51336 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_517
timestamp 1636986456
transform 1 0 52440 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_529
timestamp 18001
transform 1 0 53544 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_533
timestamp 1636986456
transform 1 0 53912 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_545
timestamp 1636986456
transform 1 0 55016 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_557
timestamp 18001
transform 1 0 56120 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_561
timestamp 1636986456
transform 1 0 56488 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_573
timestamp 1636986456
transform 1 0 57592 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_585
timestamp 18001
transform 1 0 58696 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_589
timestamp 1636986456
transform 1 0 59064 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_601
timestamp 1636986456
transform 1 0 60168 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_613
timestamp 18001
transform 1 0 61272 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_617
timestamp 1636986456
transform 1 0 61640 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_629
timestamp 1636986456
transform 1 0 62744 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_641
timestamp 18001
transform 1 0 63848 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_645
timestamp 1636986456
transform 1 0 64216 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_657
timestamp 1636986456
transform 1 0 65320 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_669
timestamp 18001
transform 1 0 66424 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_673
timestamp 1636986456
transform 1 0 66792 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_685
timestamp 1636986456
transform 1 0 67896 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_697
timestamp 18001
transform 1 0 69000 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_701
timestamp 1636986456
transform 1 0 69368 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_713
timestamp 1636986456
transform 1 0 70472 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_725
timestamp 18001
transform 1 0 71576 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_729
timestamp 1636986456
transform 1 0 71944 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_741
timestamp 1636986456
transform 1 0 73048 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_753
timestamp 18001
transform 1 0 74152 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_757
timestamp 1636986456
transform 1 0 74520 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_769
timestamp 1636986456
transform 1 0 75624 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_781
timestamp 18001
transform 1 0 76728 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_785
timestamp 1636986456
transform 1 0 77096 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_797
timestamp 1636986456
transform 1 0 78200 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_809
timestamp 18001
transform 1 0 79304 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_813
timestamp 1636986456
transform 1 0 79672 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_825
timestamp 1636986456
transform 1 0 80776 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_837
timestamp 18001
transform 1 0 81880 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_841
timestamp 1636986456
transform 1 0 82248 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_853
timestamp 1636986456
transform 1 0 83352 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_865
timestamp 18001
transform 1 0 84456 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_869
timestamp 1636986456
transform 1 0 84824 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_881
timestamp 1636986456
transform 1 0 85928 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_893
timestamp 18001
transform 1 0 87032 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_897
timestamp 18001
transform 1 0 87400 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_905
timestamp 18001
transform 1 0 88136 0 1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1636986456
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1636986456
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_27
timestamp 18001
transform 1 0 7360 0 -1 8160
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_877
timestamp 1636986456
transform 1 0 85560 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_889
timestamp 1636986456
transform 1 0 86664 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_901
timestamp 18001
transform 1 0 87768 0 -1 8160
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1636986456
transform 1 0 5152 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1636986456
transform 1 0 6256 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 18001
transform 1 0 7360 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_29
timestamp 18001
transform 1 0 7544 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_877
timestamp 1636986456
transform 1 0 85560 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_889
timestamp 1636986456
transform 1 0 86664 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_901
timestamp 18001
transform 1 0 87768 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_903
timestamp 18001
transform 1 0 87952 0 1 8160
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1636986456
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1636986456
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_27
timestamp 18001
transform 1 0 7360 0 -1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_877
timestamp 1636986456
transform 1 0 85560 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_889
timestamp 1636986456
transform 1 0 86664 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_901
timestamp 18001
transform 1 0 87768 0 -1 9248
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1636986456
transform 1 0 5152 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1636986456
transform 1 0 6256 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 18001
transform 1 0 7360 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_29
timestamp 18001
transform 1 0 7544 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_877
timestamp 1636986456
transform 1 0 85560 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_889
timestamp 1636986456
transform 1 0 86664 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_901
timestamp 18001
transform 1 0 87768 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_903
timestamp 18001
transform 1 0 87952 0 1 9248
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1636986456
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1636986456
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_27
timestamp 18001
transform 1 0 7360 0 -1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_877
timestamp 1636986456
transform 1 0 85560 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_889
timestamp 1636986456
transform 1 0 86664 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_901
timestamp 18001
transform 1 0 87768 0 -1 10336
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1636986456
transform 1 0 5152 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1636986456
transform 1 0 6256 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 18001
transform 1 0 7360 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_29
timestamp 18001
transform 1 0 7544 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_877
timestamp 1636986456
transform 1 0 85560 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_889
timestamp 18001
transform 1 0 86664 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_897
timestamp 18001
transform 1 0 87400 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_903
timestamp 18001
transform 1 0 87952 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1636986456
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1636986456
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_27
timestamp 18001
transform 1 0 7360 0 -1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_879
timestamp 1636986456
transform 1 0 85744 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_891
timestamp 1636986456
transform 1 0 86848 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_903
timestamp 18001
transform 1 0 87952 0 -1 11424
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1636986456
transform 1 0 5152 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1636986456
transform 1 0 6256 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 18001
transform 1 0 7360 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_29
timestamp 18001
transform 1 0 7544 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_877
timestamp 1636986456
transform 1 0 85560 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_889
timestamp 1636986456
transform 1 0 86664 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_901
timestamp 18001
transform 1 0 87768 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_903
timestamp 18001
transform 1 0 87952 0 1 11424
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1636986456
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1636986456
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_27
timestamp 18001
transform 1 0 7360 0 -1 12512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_879
timestamp 1636986456
transform 1 0 85744 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_891
timestamp 1636986456
transform 1 0 86848 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_903
timestamp 18001
transform 1 0 87952 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_906
timestamp 18001
transform 1 0 88228 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1636986456
transform 1 0 5152 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1636986456
transform 1 0 6256 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 18001
transform 1 0 7360 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_29
timestamp 18001
transform 1 0 7544 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_877
timestamp 1636986456
transform 1 0 85560 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_889
timestamp 18001
transform 1 0 86664 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_895
timestamp 18001
transform 1 0 87216 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1636986456
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1636986456
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_27
timestamp 18001
transform 1 0 7360 0 -1 13600
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_879
timestamp 1636986456
transform 1 0 85744 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_891
timestamp 18001
transform 1 0 86848 0 -1 13600
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1636986456
transform 1 0 5152 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1636986456
transform 1 0 6256 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 18001
transform 1 0 7360 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_29
timestamp 18001
transform 1 0 7544 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_877
timestamp 1636986456
transform 1 0 85560 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_889
timestamp 1636986456
transform 1 0 86664 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_901
timestamp 18001
transform 1 0 87768 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_903
timestamp 18001
transform 1 0 87952 0 1 13600
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1636986456
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1636986456
transform 1 0 6256 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_27
timestamp 18001
transform 1 0 7360 0 -1 14688
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_879
timestamp 1636986456
transform 1 0 85744 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_891
timestamp 1636986456
transform 1 0 86848 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_903
timestamp 18001
transform 1 0 87952 0 -1 14688
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1636986456
transform 1 0 5152 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1636986456
transform 1 0 6256 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 18001
transform 1 0 7360 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_29
timestamp 18001
transform 1 0 7544 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_877
timestamp 1636986456
transform 1 0 85560 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_889
timestamp 18001
transform 1 0 86664 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_895
timestamp 18001
transform 1 0 87216 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_8
timestamp 1636986456
transform 1 0 5612 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_20
timestamp 18001
transform 1 0 6716 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_28
timestamp 18001
transform 1 0 7452 0 -1 15776
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_877
timestamp 1636986456
transform 1 0 85560 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_889
timestamp 1636986456
transform 1 0 86664 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_901
timestamp 18001
transform 1 0 87768 0 -1 15776
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_8
timestamp 1636986456
transform 1 0 5612 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_20
timestamp 18001
transform 1 0 6716 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_29
timestamp 18001
transform 1 0 7544 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_877
timestamp 1636986456
transform 1 0 85560 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_889
timestamp 1636986456
transform 1 0 86664 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_901
timestamp 18001
transform 1 0 87768 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1636986456
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1636986456
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_27
timestamp 18001
transform 1 0 7360 0 -1 16864
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_877
timestamp 1636986456
transform 1 0 85560 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_889
timestamp 1636986456
transform 1 0 86664 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_901
timestamp 18001
transform 1 0 87768 0 -1 16864
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1636986456
transform 1 0 5152 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1636986456
transform 1 0 6256 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 18001
transform 1 0 7360 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_29
timestamp 18001
transform 1 0 7544 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_877
timestamp 1636986456
transform 1 0 85560 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_889
timestamp 1636986456
transform 1 0 86664 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_901
timestamp 18001
transform 1 0 87768 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_903
timestamp 18001
transform 1 0 87952 0 1 16864
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_8
timestamp 1636986456
transform 1 0 5612 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_20
timestamp 18001
transform 1 0 6716 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_28
timestamp 18001
transform 1 0 7452 0 -1 17952
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_877
timestamp 1636986456
transform 1 0 85560 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_889
timestamp 1636986456
transform 1 0 86664 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_901
timestamp 18001
transform 1 0 87768 0 -1 17952
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1636986456
transform 1 0 5152 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1636986456
transform 1 0 6256 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 18001
transform 1 0 7360 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_29
timestamp 18001
transform 1 0 7544 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_877
timestamp 1636986456
transform 1 0 85560 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_889
timestamp 1636986456
transform 1 0 86664 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_901
timestamp 18001
transform 1 0 87768 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_903
timestamp 18001
transform 1 0 87952 0 1 17952
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_8
timestamp 1636986456
transform 1 0 5612 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_20
timestamp 18001
transform 1 0 6716 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_28
timestamp 18001
transform 1 0 7452 0 -1 19040
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_877
timestamp 1636986456
transform 1 0 85560 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_889
timestamp 1636986456
transform 1 0 86664 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_901
timestamp 18001
transform 1 0 87768 0 -1 19040
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1636986456
transform 1 0 5152 0 1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1636986456
transform 1 0 6256 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 18001
transform 1 0 7360 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_29
timestamp 18001
transform 1 0 7544 0 1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_877
timestamp 1636986456
transform 1 0 85560 0 1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_889
timestamp 1636986456
transform 1 0 86664 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_901
timestamp 18001
transform 1 0 87768 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_903
timestamp 18001
transform 1 0 87952 0 1 19040
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_8
timestamp 1636986456
transform 1 0 5612 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_20
timestamp 18001
transform 1 0 6716 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_28
timestamp 18001
transform 1 0 7452 0 -1 20128
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_877
timestamp 1636986456
transform 1 0 85560 0 -1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_889
timestamp 1636986456
transform 1 0 86664 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_901
timestamp 18001
transform 1 0 87768 0 -1 20128
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1636986456
transform 1 0 5152 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1636986456
transform 1 0 6256 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 18001
transform 1 0 7360 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_29
timestamp 18001
transform 1 0 7544 0 1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_877
timestamp 1636986456
transform 1 0 85560 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_889
timestamp 1636986456
transform 1 0 86664 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_901
timestamp 18001
transform 1 0 87768 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_903
timestamp 18001
transform 1 0 87952 0 1 20128
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_8
timestamp 1636986456
transform 1 0 5612 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_20
timestamp 18001
transform 1 0 6716 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_28
timestamp 18001
transform 1 0 7452 0 -1 21216
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_877
timestamp 1636986456
transform 1 0 85560 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_889
timestamp 1636986456
transform 1 0 86664 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_901
timestamp 18001
transform 1 0 87768 0 -1 21216
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_8
timestamp 1636986456
transform 1 0 5612 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_20
timestamp 18001
transform 1 0 6716 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_29
timestamp 18001
transform 1 0 7544 0 1 21216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_877
timestamp 1636986456
transform 1 0 85560 0 1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_889
timestamp 1636986456
transform 1 0 86664 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_901
timestamp 18001
transform 1 0 87768 0 1 21216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1636986456
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1636986456
transform 1 0 6256 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_27
timestamp 18001
transform 1 0 7360 0 -1 22304
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_877
timestamp 1636986456
transform 1 0 85560 0 -1 22304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_889
timestamp 1636986456
transform 1 0 86664 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_901
timestamp 18001
transform 1 0 87768 0 -1 22304
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1636986456
transform 1 0 5152 0 1 22304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1636986456
transform 1 0 6256 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 18001
transform 1 0 7360 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_29
timestamp 18001
transform 1 0 7544 0 1 22304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_877
timestamp 1636986456
transform 1 0 85560 0 1 22304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_889
timestamp 1636986456
transform 1 0 86664 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_901
timestamp 18001
transform 1 0 87768 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_903
timestamp 18001
transform 1 0 87952 0 1 22304
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_8
timestamp 1636986456
transform 1 0 5612 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_20
timestamp 18001
transform 1 0 6716 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_28
timestamp 18001
transform 1 0 7452 0 -1 23392
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_877
timestamp 1636986456
transform 1 0 85560 0 -1 23392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_889
timestamp 1636986456
transform 1 0 86664 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_901
timestamp 18001
transform 1 0 87768 0 -1 23392
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1636986456
transform 1 0 5152 0 1 23392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1636986456
transform 1 0 6256 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 18001
transform 1 0 7360 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_29
timestamp 18001
transform 1 0 7544 0 1 23392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_877
timestamp 1636986456
transform 1 0 85560 0 1 23392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_889
timestamp 1636986456
transform 1 0 86664 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_901
timestamp 18001
transform 1 0 87768 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_903
timestamp 18001
transform 1 0 87952 0 1 23392
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_8
timestamp 1636986456
transform 1 0 5612 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_20
timestamp 18001
transform 1 0 6716 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_28
timestamp 18001
transform 1 0 7452 0 -1 24480
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_877
timestamp 1636986456
transform 1 0 85560 0 -1 24480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_889
timestamp 1636986456
transform 1 0 86664 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_901
timestamp 18001
transform 1 0 87768 0 -1 24480
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1636986456
transform 1 0 5152 0 1 24480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1636986456
transform 1 0 6256 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 18001
transform 1 0 7360 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_29
timestamp 18001
transform 1 0 7544 0 1 24480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_877
timestamp 1636986456
transform 1 0 85560 0 1 24480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_889
timestamp 1636986456
transform 1 0 86664 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_901
timestamp 18001
transform 1 0 87768 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_903
timestamp 18001
transform 1 0 87952 0 1 24480
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_8
timestamp 1636986456
transform 1 0 5612 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_20
timestamp 18001
transform 1 0 6716 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_28
timestamp 18001
transform 1 0 7452 0 -1 25568
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_877
timestamp 1636986456
transform 1 0 85560 0 -1 25568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_889
timestamp 1636986456
transform 1 0 86664 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_901
timestamp 18001
transform 1 0 87768 0 -1 25568
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1636986456
transform 1 0 5152 0 1 25568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1636986456
transform 1 0 6256 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 18001
transform 1 0 7360 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_29
timestamp 18001
transform 1 0 7544 0 1 25568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_877
timestamp 1636986456
transform 1 0 85560 0 1 25568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_889
timestamp 1636986456
transform 1 0 86664 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_901
timestamp 18001
transform 1 0 87768 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_903
timestamp 18001
transform 1 0 87952 0 1 25568
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_8
timestamp 1636986456
transform 1 0 5612 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_20
timestamp 18001
transform 1 0 6716 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_28
timestamp 18001
transform 1 0 7452 0 -1 26656
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_877
timestamp 1636986456
transform 1 0 85560 0 -1 26656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_889
timestamp 1636986456
transform 1 0 86664 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_901
timestamp 18001
transform 1 0 87768 0 -1 26656
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_8
timestamp 1636986456
transform 1 0 5612 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_20
timestamp 18001
transform 1 0 6716 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_29
timestamp 18001
transform 1 0 7544 0 1 26656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_877
timestamp 1636986456
transform 1 0 85560 0 1 26656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_889
timestamp 1636986456
transform 1 0 86664 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_901
timestamp 18001
transform 1 0 87768 0 1 26656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1636986456
transform 1 0 5152 0 -1 27744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1636986456
transform 1 0 6256 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_27
timestamp 18001
transform 1 0 7360 0 -1 27744
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_877
timestamp 1636986456
transform 1 0 85560 0 -1 27744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_889
timestamp 1636986456
transform 1 0 86664 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_901
timestamp 18001
transform 1 0 87768 0 -1 27744
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1636986456
transform 1 0 5152 0 1 27744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1636986456
transform 1 0 6256 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 18001
transform 1 0 7360 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_29
timestamp 18001
transform 1 0 7544 0 1 27744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_877
timestamp 1636986456
transform 1 0 85560 0 1 27744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_889
timestamp 1636986456
transform 1 0 86664 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_901
timestamp 18001
transform 1 0 87768 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_903
timestamp 18001
transform 1 0 87952 0 1 27744
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_8
timestamp 1636986456
transform 1 0 5612 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_20
timestamp 18001
transform 1 0 6716 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_28
timestamp 18001
transform 1 0 7452 0 -1 28832
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_877
timestamp 1636986456
transform 1 0 85560 0 -1 28832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_889
timestamp 1636986456
transform 1 0 86664 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_901
timestamp 18001
transform 1 0 87768 0 -1 28832
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1636986456
transform 1 0 5152 0 1 28832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1636986456
transform 1 0 6256 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 18001
transform 1 0 7360 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_44_29
timestamp 18001
transform 1 0 7544 0 1 28832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_877
timestamp 1636986456
transform 1 0 85560 0 1 28832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_889
timestamp 1636986456
transform 1 0 86664 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_901
timestamp 18001
transform 1 0 87768 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_903
timestamp 18001
transform 1 0 87952 0 1 28832
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_8
timestamp 1636986456
transform 1 0 5612 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_20
timestamp 18001
transform 1 0 6716 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_28
timestamp 18001
transform 1 0 7452 0 -1 29920
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_877
timestamp 1636986456
transform 1 0 85560 0 -1 29920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_889
timestamp 1636986456
transform 1 0 86664 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_901
timestamp 18001
transform 1 0 87768 0 -1 29920
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1636986456
transform 1 0 5152 0 1 29920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1636986456
transform 1 0 6256 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 18001
transform 1 0 7360 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_29
timestamp 18001
transform 1 0 7544 0 1 29920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_877
timestamp 1636986456
transform 1 0 85560 0 1 29920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_889
timestamp 1636986456
transform 1 0 86664 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_901
timestamp 18001
transform 1 0 87768 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_903
timestamp 18001
transform 1 0 87952 0 1 29920
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_7
timestamp 1636986456
transform 1 0 5520 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_19
timestamp 18001
transform 1 0 6624 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_27
timestamp 18001
transform 1 0 7360 0 -1 31008
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_877
timestamp 1636986456
transform 1 0 85560 0 -1 31008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_889
timestamp 1636986456
transform 1 0 86664 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_901
timestamp 18001
transform 1 0 87768 0 -1 31008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1636986456
transform 1 0 5152 0 1 31008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1636986456
transform 1 0 6256 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 18001
transform 1 0 7360 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_29
timestamp 18001
transform 1 0 7544 0 1 31008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_877
timestamp 1636986456
transform 1 0 85560 0 1 31008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_889
timestamp 1636986456
transform 1 0 86664 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_901
timestamp 18001
transform 1 0 87768 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_903
timestamp 18001
transform 1 0 87952 0 1 31008
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_7
timestamp 1636986456
transform 1 0 5520 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_19
timestamp 18001
transform 1 0 6624 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_27
timestamp 18001
transform 1 0 7360 0 -1 32096
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_877
timestamp 1636986456
transform 1 0 85560 0 -1 32096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_889
timestamp 1636986456
transform 1 0 86664 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_901
timestamp 18001
transform 1 0 87768 0 -1 32096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_7
timestamp 1636986456
transform 1 0 5520 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_19
timestamp 18001
transform 1 0 6624 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 18001
transform 1 0 7360 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_50_29
timestamp 18001
transform 1 0 7544 0 1 32096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_877
timestamp 1636986456
transform 1 0 85560 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_889
timestamp 18001
transform 1 0 86664 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_897
timestamp 18001
transform 1 0 87400 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_50_903
timestamp 18001
transform 1 0 87952 0 1 32096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1636986456
transform 1 0 5152 0 -1 33184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1636986456
transform 1 0 6256 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_27
timestamp 18001
transform 1 0 7360 0 -1 33184
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_877
timestamp 1636986456
transform 1 0 85560 0 -1 33184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_889
timestamp 1636986456
transform 1 0 86664 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_901
timestamp 18001
transform 1 0 87768 0 -1 33184
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1636986456
transform 1 0 5152 0 1 33184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1636986456
transform 1 0 6256 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 18001
transform 1 0 7360 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_52_29
timestamp 18001
transform 1 0 7544 0 1 33184
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_877
timestamp 1636986456
transform 1 0 85560 0 1 33184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_889
timestamp 1636986456
transform 1 0 86664 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_901
timestamp 18001
transform 1 0 87768 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_903
timestamp 18001
transform 1 0 87952 0 1 33184
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_7
timestamp 1636986456
transform 1 0 5520 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_19
timestamp 18001
transform 1 0 6624 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_27
timestamp 18001
transform 1 0 7360 0 -1 34272
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_877
timestamp 1636986456
transform 1 0 85560 0 -1 34272
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_889
timestamp 1636986456
transform 1 0 86664 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_901
timestamp 18001
transform 1 0 87768 0 -1 34272
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1636986456
transform 1 0 5152 0 1 34272
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1636986456
transform 1 0 6256 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 18001
transform 1 0 7360 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_29
timestamp 18001
transform 1 0 7544 0 1 34272
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_877
timestamp 1636986456
transform 1 0 85560 0 1 34272
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_889
timestamp 1636986456
transform 1 0 86664 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_901
timestamp 18001
transform 1 0 87768 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_903
timestamp 18001
transform 1 0 87952 0 1 34272
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_7
timestamp 1636986456
transform 1 0 5520 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_19
timestamp 18001
transform 1 0 6624 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_27
timestamp 18001
transform 1 0 7360 0 -1 35360
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_877
timestamp 1636986456
transform 1 0 85560 0 -1 35360
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_889
timestamp 1636986456
transform 1 0 86664 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_901
timestamp 18001
transform 1 0 87768 0 -1 35360
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1636986456
transform 1 0 5152 0 1 35360
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1636986456
transform 1 0 6256 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 18001
transform 1 0 7360 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_56_29
timestamp 18001
transform 1 0 7544 0 1 35360
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_877
timestamp 1636986456
transform 1 0 85560 0 1 35360
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_889
timestamp 1636986456
transform 1 0 86664 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_901
timestamp 18001
transform 1 0 87768 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_903
timestamp 18001
transform 1 0 87952 0 1 35360
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_7
timestamp 1636986456
transform 1 0 5520 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_19
timestamp 18001
transform 1 0 6624 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_27
timestamp 18001
transform 1 0 7360 0 -1 36448
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_877
timestamp 1636986456
transform 1 0 85560 0 -1 36448
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_889
timestamp 1636986456
transform 1 0 86664 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_901
timestamp 18001
transform 1 0 87768 0 -1 36448
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1636986456
transform 1 0 5152 0 1 36448
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1636986456
transform 1 0 6256 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 18001
transform 1 0 7360 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_58_29
timestamp 18001
transform 1 0 7544 0 1 36448
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_877
timestamp 1636986456
transform 1 0 85560 0 1 36448
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_889
timestamp 1636986456
transform 1 0 86664 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_901
timestamp 18001
transform 1 0 87768 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_903
timestamp 18001
transform 1 0 87952 0 1 36448
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_7
timestamp 1636986456
transform 1 0 5520 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_19
timestamp 18001
transform 1 0 6624 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_27
timestamp 18001
transform 1 0 7360 0 -1 37536
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_877
timestamp 1636986456
transform 1 0 85560 0 -1 37536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_889
timestamp 1636986456
transform 1 0 86664 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_901
timestamp 18001
transform 1 0 87768 0 -1 37536
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_7
timestamp 1636986456
transform 1 0 5520 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_19
timestamp 18001
transform 1 0 6624 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 18001
transform 1 0 7360 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_60_29
timestamp 18001
transform 1 0 7544 0 1 37536
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_877
timestamp 1636986456
transform 1 0 85560 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_889
timestamp 18001
transform 1 0 86664 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_897
timestamp 18001
transform 1 0 87400 0 1 37536
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1636986456
transform 1 0 5152 0 -1 38624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1636986456
transform 1 0 6256 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_27
timestamp 18001
transform 1 0 7360 0 -1 38624
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_877
timestamp 1636986456
transform 1 0 85560 0 -1 38624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_889
timestamp 1636986456
transform 1 0 86664 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_901
timestamp 18001
transform 1 0 87768 0 -1 38624
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1636986456
transform 1 0 5152 0 1 38624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1636986456
transform 1 0 6256 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 18001
transform 1 0 7360 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_62_29
timestamp 18001
transform 1 0 7544 0 1 38624
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_877
timestamp 1636986456
transform 1 0 85560 0 1 38624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_889
timestamp 1636986456
transform 1 0 86664 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_901
timestamp 18001
transform 1 0 87768 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_903
timestamp 18001
transform 1 0 87952 0 1 38624
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_7
timestamp 1636986456
transform 1 0 5520 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_19
timestamp 18001
transform 1 0 6624 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_27
timestamp 18001
transform 1 0 7360 0 -1 39712
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_877
timestamp 1636986456
transform 1 0 85560 0 -1 39712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_889
timestamp 1636986456
transform 1 0 86664 0 -1 39712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1636986456
transform 1 0 5152 0 1 39712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1636986456
transform 1 0 6256 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 18001
transform 1 0 7360 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_64_29
timestamp 18001
transform 1 0 7544 0 1 39712
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_877
timestamp 1636986456
transform 1 0 85560 0 1 39712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_889
timestamp 1636986456
transform 1 0 86664 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_901
timestamp 18001
transform 1 0 87768 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_903
timestamp 18001
transform 1 0 87952 0 1 39712
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_7
timestamp 1636986456
transform 1 0 5520 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_19
timestamp 18001
transform 1 0 6624 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_27
timestamp 18001
transform 1 0 7360 0 -1 40800
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_65_877
timestamp 1636986456
transform 1 0 85560 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_889
timestamp 18001
transform 1 0 86664 0 -1 40800
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1636986456
transform 1 0 5152 0 1 40800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 1636986456
transform 1 0 6256 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 18001
transform 1 0 7360 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_66_29
timestamp 18001
transform 1 0 7544 0 1 40800
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_877
timestamp 1636986456
transform 1 0 85560 0 1 40800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_889
timestamp 1636986456
transform 1 0 86664 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_901
timestamp 18001
transform 1 0 87768 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_903
timestamp 18001
transform 1 0 87952 0 1 40800
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_7
timestamp 1636986456
transform 1 0 5520 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_19
timestamp 18001
transform 1 0 6624 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_27
timestamp 18001
transform 1 0 7360 0 -1 41888
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_67_877
timestamp 1636986456
transform 1 0 85560 0 -1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_889
timestamp 1636986456
transform 1 0 86664 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_901
timestamp 18001
transform 1 0 87768 0 -1 41888
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1636986456
transform 1 0 5152 0 1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1636986456
transform 1 0 6256 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 18001
transform 1 0 7360 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_68_29
timestamp 18001
transform 1 0 7544 0 1 41888
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_877
timestamp 1636986456
transform 1 0 85560 0 1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_889
timestamp 1636986456
transform 1 0 86664 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_901
timestamp 18001
transform 1 0 87768 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_903
timestamp 18001
transform 1 0 87952 0 1 41888
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_69_7
timestamp 1636986456
transform 1 0 5520 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_19
timestamp 18001
transform 1 0 6624 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_69_27
timestamp 18001
transform 1 0 7360 0 -1 42976
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_69_877
timestamp 1636986456
transform 1 0 85560 0 -1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_889
timestamp 1636986456
transform 1 0 86664 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_901
timestamp 18001
transform 1 0 87768 0 -1 42976
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_7
timestamp 1636986456
transform 1 0 5520 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_19
timestamp 18001
transform 1 0 6624 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 18001
transform 1 0 7360 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_70_29
timestamp 18001
transform 1 0 7544 0 1 42976
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_877
timestamp 1636986456
transform 1 0 85560 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_889
timestamp 18001
transform 1 0 86664 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_70_897
timestamp 18001
transform 1 0 87400 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_70_903
timestamp 18001
transform 1 0 87952 0 1 42976
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1636986456
transform 1 0 5152 0 -1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1636986456
transform 1 0 6256 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_71_27
timestamp 18001
transform 1 0 7360 0 -1 44064
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_71_877
timestamp 1636986456
transform 1 0 85560 0 -1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_889
timestamp 1636986456
transform 1 0 86664 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_901
timestamp 18001
transform 1 0 87768 0 -1 44064
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1636986456
transform 1 0 5152 0 1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1636986456
transform 1 0 6256 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 18001
transform 1 0 7360 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_72_29
timestamp 18001
transform 1 0 7544 0 1 44064
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_877
timestamp 1636986456
transform 1 0 85560 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_889
timestamp 18001
transform 1 0 86664 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_72_897
timestamp 18001
transform 1 0 87400 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_72_903
timestamp 18001
transform 1 0 87952 0 1 44064
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_7
timestamp 1636986456
transform 1 0 5520 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_19
timestamp 18001
transform 1 0 6624 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_27
timestamp 18001
transform 1 0 7360 0 -1 45152
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_877
timestamp 1636986456
transform 1 0 85560 0 -1 45152
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_889
timestamp 1636986456
transform 1 0 86664 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_901
timestamp 18001
transform 1 0 87768 0 -1 45152
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_74_8
timestamp 1636986456
transform 1 0 5612 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_20
timestamp 18001
transform 1 0 6716 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_29
timestamp 18001
transform 1 0 7544 0 1 45152
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_885
timestamp 1636986456
transform 1 0 86296 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_897
timestamp 18001
transform 1 0 87400 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_901
timestamp 18001
transform 1 0 87768 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_74_903
timestamp 18001
transform 1 0 87952 0 1 45152
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_3
timestamp 1636986456
transform 1 0 5152 0 -1 46240
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_15
timestamp 1636986456
transform 1 0 6256 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_27
timestamp 18001
transform 1 0 7360 0 -1 46240
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_75_877
timestamp 1636986456
transform 1 0 85560 0 -1 46240
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_889
timestamp 1636986456
transform 1 0 86664 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_901
timestamp 18001
transform 1 0 87768 0 -1 46240
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1636986456
transform 1 0 5152 0 1 46240
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1636986456
transform 1 0 6256 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 18001
transform 1 0 7360 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_76_29
timestamp 18001
transform 1 0 7544 0 1 46240
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_877
timestamp 1636986456
transform 1 0 85560 0 1 46240
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_889
timestamp 1636986456
transform 1 0 86664 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_901
timestamp 18001
transform 1 0 87768 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_903
timestamp 18001
transform 1 0 87952 0 1 46240
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1636986456
transform 1 0 5152 0 -1 47328
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1636986456
transform 1 0 6256 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_77_27
timestamp 18001
transform 1 0 7360 0 -1 47328
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_77_877
timestamp 1636986456
transform 1 0 85560 0 -1 47328
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_889
timestamp 1636986456
transform 1 0 86664 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_77_901
timestamp 18001
transform 1 0 87768 0 -1 47328
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1636986456
transform 1 0 5152 0 1 47328
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1636986456
transform 1 0 6256 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 18001
transform 1 0 7360 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_78_29
timestamp 18001
transform 1 0 7544 0 1 47328
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_877
timestamp 1636986456
transform 1 0 85560 0 1 47328
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_889
timestamp 1636986456
transform 1 0 86664 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_901
timestamp 18001
transform 1 0 87768 0 1 47328
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1636986456
transform 1 0 5152 0 -1 48416
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1636986456
transform 1 0 6256 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_27
timestamp 18001
transform 1 0 7360 0 -1 48416
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_79_877
timestamp 1636986456
transform 1 0 85560 0 -1 48416
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_889
timestamp 1636986456
transform 1 0 86664 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_901
timestamp 18001
transform 1 0 87768 0 -1 48416
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_3
timestamp 1636986456
transform 1 0 5152 0 1 48416
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 1636986456
transform 1 0 6256 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 18001
transform 1 0 7360 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_80_29
timestamp 18001
transform 1 0 7544 0 1 48416
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_879
timestamp 1636986456
transform 1 0 85744 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_891
timestamp 18001
transform 1 0 86848 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_899
timestamp 18001
transform 1 0 87584 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_80_903
timestamp 18001
transform 1 0 87952 0 1 48416
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1636986456
transform 1 0 5152 0 -1 49504
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1636986456
transform 1 0 6256 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_81_27
timestamp 18001
transform 1 0 7360 0 -1 49504
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_81_877
timestamp 1636986456
transform 1 0 85560 0 -1 49504
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_889
timestamp 1636986456
transform 1 0 86664 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_901
timestamp 18001
transform 1 0 87768 0 -1 49504
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_82_3
timestamp 1636986456
transform 1 0 5152 0 1 49504
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_15
timestamp 1636986456
transform 1 0 6256 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 18001
transform 1 0 7360 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_82_29
timestamp 18001
transform 1 0 7544 0 1 49504
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_879
timestamp 1636986456
transform 1 0 85744 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_891
timestamp 18001
transform 1 0 86848 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_899
timestamp 18001
transform 1 0 87584 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_903
timestamp 18001
transform 1 0 87952 0 1 49504
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_83_3
timestamp 1636986456
transform 1 0 5152 0 -1 50592
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_15
timestamp 1636986456
transform 1 0 6256 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_83_27
timestamp 18001
transform 1 0 7360 0 -1 50592
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_83_877
timestamp 1636986456
transform 1 0 85560 0 -1 50592
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_889
timestamp 1636986456
transform 1 0 86664 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_901
timestamp 18001
transform 1 0 87768 0 -1 50592
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_84_3
timestamp 1636986456
transform 1 0 5152 0 1 50592
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_15
timestamp 1636986456
transform 1 0 6256 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 18001
transform 1 0 7360 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_84_29
timestamp 18001
transform 1 0 7544 0 1 50592
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_879
timestamp 1636986456
transform 1 0 85744 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_891
timestamp 18001
transform 1 0 86848 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_84_899
timestamp 18001
transform 1 0 87584 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_84_903
timestamp 18001
transform 1 0 87952 0 1 50592
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_85_8
timestamp 1636986456
transform 1 0 5612 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_20
timestamp 18001
transform 1 0 6716 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_85_28
timestamp 18001
transform 1 0 7452 0 -1 51680
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_85_877
timestamp 1636986456
transform 1 0 85560 0 -1 51680
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_889
timestamp 1636986456
transform 1 0 86664 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_85_901
timestamp 18001
transform 1 0 87768 0 -1 51680
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_86_3
timestamp 1636986456
transform 1 0 5152 0 1 51680
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_15
timestamp 1636986456
transform 1 0 6256 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 18001
transform 1 0 7360 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_86_29
timestamp 18001
transform 1 0 7544 0 1 51680
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_877
timestamp 1636986456
transform 1 0 85560 0 1 51680
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_889
timestamp 1636986456
transform 1 0 86664 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_901
timestamp 18001
transform 1 0 87768 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_903
timestamp 18001
transform 1 0 87952 0 1 51680
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_87_3
timestamp 1636986456
transform 1 0 5152 0 -1 52768
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_15
timestamp 1636986456
transform 1 0 6256 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_87_27
timestamp 18001
transform 1 0 7360 0 -1 52768
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_87_877
timestamp 1636986456
transform 1 0 85560 0 -1 52768
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_889
timestamp 1636986456
transform 1 0 86664 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_901
timestamp 18001
transform 1 0 87768 0 -1 52768
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_88_8
timestamp 1636986456
transform 1 0 5612 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_20
timestamp 18001
transform 1 0 6716 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_88_29
timestamp 18001
transform 1 0 7544 0 1 52768
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_877
timestamp 1636986456
transform 1 0 85560 0 1 52768
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_889
timestamp 1636986456
transform 1 0 86664 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_901
timestamp 18001
transform 1 0 87768 0 1 52768
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_3
timestamp 1636986456
transform 1 0 5152 0 -1 53856
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_15
timestamp 1636986456
transform 1 0 6256 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_89_27
timestamp 18001
transform 1 0 7360 0 -1 53856
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_89_877
timestamp 1636986456
transform 1 0 85560 0 -1 53856
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_889
timestamp 1636986456
transform 1 0 86664 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_901
timestamp 18001
transform 1 0 87768 0 -1 53856
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_90_8
timestamp 1636986456
transform 1 0 5612 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_90_20
timestamp 18001
transform 1 0 6716 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_90_29
timestamp 18001
transform 1 0 7544 0 1 53856
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_877
timestamp 1636986456
transform 1 0 85560 0 1 53856
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_889
timestamp 1636986456
transform 1 0 86664 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_901
timestamp 18001
transform 1 0 87768 0 1 53856
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_3
timestamp 1636986456
transform 1 0 5152 0 -1 54944
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_15
timestamp 1636986456
transform 1 0 6256 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_91_27
timestamp 18001
transform 1 0 7360 0 -1 54944
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_91_877
timestamp 1636986456
transform 1 0 85560 0 -1 54944
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_889
timestamp 1636986456
transform 1 0 86664 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_901
timestamp 18001
transform 1 0 87768 0 -1 54944
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_92_8
timestamp 1636986456
transform 1 0 5612 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_20
timestamp 18001
transform 1 0 6716 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_92_29
timestamp 18001
transform 1 0 7544 0 1 54944
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_877
timestamp 1636986456
transform 1 0 85560 0 1 54944
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_889
timestamp 1636986456
transform 1 0 86664 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_901
timestamp 18001
transform 1 0 87768 0 1 54944
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_3
timestamp 1636986456
transform 1 0 5152 0 -1 56032
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_15
timestamp 1636986456
transform 1 0 6256 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_93_27
timestamp 18001
transform 1 0 7360 0 -1 56032
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_93_877
timestamp 1636986456
transform 1 0 85560 0 -1 56032
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_889
timestamp 1636986456
transform 1 0 86664 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_901
timestamp 18001
transform 1 0 87768 0 -1 56032
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_94_8
timestamp 1636986456
transform 1 0 5612 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_20
timestamp 18001
transform 1 0 6716 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_94_29
timestamp 18001
transform 1 0 7544 0 1 56032
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_877
timestamp 1636986456
transform 1 0 85560 0 1 56032
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_889
timestamp 1636986456
transform 1 0 86664 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_901
timestamp 18001
transform 1 0 87768 0 1 56032
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_8
timestamp 1636986456
transform 1 0 5612 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_20
timestamp 18001
transform 1 0 6716 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_95_28
timestamp 18001
transform 1 0 7452 0 -1 57120
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_95_877
timestamp 1636986456
transform 1 0 85560 0 -1 57120
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_889
timestamp 1636986456
transform 1 0 86664 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_95_901
timestamp 18001
transform 1 0 87768 0 -1 57120
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_96_3
timestamp 1636986456
transform 1 0 5152 0 1 57120
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_15
timestamp 1636986456
transform 1 0 6256 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_27
timestamp 18001
transform 1 0 7360 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_96_29
timestamp 18001
transform 1 0 7544 0 1 57120
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_877
timestamp 1636986456
transform 1 0 85560 0 1 57120
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_889
timestamp 1636986456
transform 1 0 86664 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_901
timestamp 18001
transform 1 0 87768 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_96_903
timestamp 18001
transform 1 0 87952 0 1 57120
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_97_3
timestamp 1636986456
transform 1 0 5152 0 -1 58208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_15
timestamp 1636986456
transform 1 0 6256 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_97_27
timestamp 18001
transform 1 0 7360 0 -1 58208
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_97_877
timestamp 1636986456
transform 1 0 85560 0 -1 58208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_889
timestamp 1636986456
transform 1 0 86664 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_901
timestamp 18001
transform 1 0 87768 0 -1 58208
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_98_8
timestamp 1636986456
transform 1 0 5612 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_20
timestamp 18001
transform 1 0 6716 0 1 58208
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_98_29
timestamp 18001
transform 1 0 7544 0 1 58208
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_877
timestamp 1636986456
transform 1 0 85560 0 1 58208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_889
timestamp 1636986456
transform 1 0 86664 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_901
timestamp 18001
transform 1 0 87768 0 1 58208
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_3
timestamp 1636986456
transform 1 0 5152 0 -1 59296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_15
timestamp 1636986456
transform 1 0 6256 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_99_27
timestamp 18001
transform 1 0 7360 0 -1 59296
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_99_877
timestamp 1636986456
transform 1 0 85560 0 -1 59296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_889
timestamp 1636986456
transform 1 0 86664 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_901
timestamp 18001
transform 1 0 87768 0 -1 59296
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_100_8
timestamp 1636986456
transform 1 0 5612 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_20
timestamp 18001
transform 1 0 6716 0 1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_100_29
timestamp 18001
transform 1 0 7544 0 1 59296
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_877
timestamp 1636986456
transform 1 0 85560 0 1 59296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_889
timestamp 1636986456
transform 1 0 86664 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_901
timestamp 18001
transform 1 0 87768 0 1 59296
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_3
timestamp 1636986456
transform 1 0 5152 0 -1 60384
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_15
timestamp 1636986456
transform 1 0 6256 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_27
timestamp 18001
transform 1 0 7360 0 -1 60384
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_877
timestamp 1636986456
transform 1 0 85560 0 -1 60384
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_889
timestamp 1636986456
transform 1 0 86664 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_901
timestamp 18001
transform 1 0 87768 0 -1 60384
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_102_8
timestamp 1636986456
transform 1 0 5612 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_102_20
timestamp 18001
transform 1 0 6716 0 1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_102_29
timestamp 18001
transform 1 0 7544 0 1 60384
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_877
timestamp 1636986456
transform 1 0 85560 0 1 60384
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_889
timestamp 1636986456
transform 1 0 86664 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_102_901
timestamp 18001
transform 1 0 87768 0 1 60384
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_3
timestamp 1636986456
transform 1 0 5152 0 -1 61472
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_15
timestamp 1636986456
transform 1 0 6256 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_103_27
timestamp 18001
transform 1 0 7360 0 -1 61472
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_103_877
timestamp 1636986456
transform 1 0 85560 0 -1 61472
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_889
timestamp 1636986456
transform 1 0 86664 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_901
timestamp 18001
transform 1 0 87768 0 -1 61472
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_104_8
timestamp 1636986456
transform 1 0 5612 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_104_20
timestamp 18001
transform 1 0 6716 0 1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_104_29
timestamp 18001
transform 1 0 7544 0 1 61472
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_877
timestamp 1636986456
transform 1 0 85560 0 1 61472
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_889
timestamp 1636986456
transform 1 0 86664 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_104_901
timestamp 18001
transform 1 0 87768 0 1 61472
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_8
timestamp 1636986456
transform 1 0 5612 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_105_20
timestamp 18001
transform 1 0 6716 0 -1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_105_28
timestamp 18001
transform 1 0 7452 0 -1 62560
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_105_877
timestamp 1636986456
transform 1 0 85560 0 -1 62560
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_889
timestamp 1636986456
transform 1 0 86664 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_105_901
timestamp 18001
transform 1 0 87768 0 -1 62560
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_106_3
timestamp 1636986456
transform 1 0 5152 0 1 62560
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_15
timestamp 1636986456
transform 1 0 6256 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_106_27
timestamp 18001
transform 1 0 7360 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_106_29
timestamp 18001
transform 1 0 7544 0 1 62560
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_877
timestamp 1636986456
transform 1 0 85560 0 1 62560
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_889
timestamp 1636986456
transform 1 0 86664 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_106_901
timestamp 18001
transform 1 0 87768 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_106_903
timestamp 18001
transform 1 0 87952 0 1 62560
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_107_3
timestamp 1636986456
transform 1 0 5152 0 -1 63648
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_15
timestamp 1636986456
transform 1 0 6256 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_107_27
timestamp 18001
transform 1 0 7360 0 -1 63648
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_877
timestamp 1636986456
transform 1 0 85560 0 -1 63648
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_889
timestamp 1636986456
transform 1 0 86664 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_901
timestamp 18001
transform 1 0 87768 0 -1 63648
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_29
timestamp 18001
transform 1 0 7544 0 1 63648
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_877
timestamp 1636986456
transform 1 0 85560 0 1 63648
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_889
timestamp 1636986456
transform 1 0 86664 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_108_901
timestamp 18001
transform 1 0 87768 0 1 63648
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_3
timestamp 1636986456
transform 1 0 5152 0 -1 64736
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_15
timestamp 1636986456
transform 1 0 6256 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_109_27
timestamp 18001
transform 1 0 7360 0 -1 64736
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_877
timestamp 1636986456
transform 1 0 85560 0 -1 64736
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_889
timestamp 1636986456
transform 1 0 86664 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_901
timestamp 18001
transform 1 0 87768 0 -1 64736
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_110_8
timestamp 1636986456
transform 1 0 5612 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_110_20
timestamp 18001
transform 1 0 6716 0 1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_110_29
timestamp 18001
transform 1 0 7544 0 1 64736
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_877
timestamp 1636986456
transform 1 0 85560 0 1 64736
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_889
timestamp 1636986456
transform 1 0 86664 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_110_901
timestamp 18001
transform 1 0 87768 0 1 64736
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_3
timestamp 1636986456
transform 1 0 5152 0 -1 65824
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_15
timestamp 1636986456
transform 1 0 6256 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_111_27
timestamp 18001
transform 1 0 7360 0 -1 65824
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_111_877
timestamp 1636986456
transform 1 0 85560 0 -1 65824
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_889
timestamp 1636986456
transform 1 0 86664 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_901
timestamp 18001
transform 1 0 87768 0 -1 65824
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_112_8
timestamp 1636986456
transform 1 0 5612 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_112_20
timestamp 18001
transform 1 0 6716 0 1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_112_29
timestamp 18001
transform 1 0 7544 0 1 65824
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_877
timestamp 1636986456
transform 1 0 85560 0 1 65824
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_889
timestamp 1636986456
transform 1 0 86664 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_112_901
timestamp 18001
transform 1 0 87768 0 1 65824
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_3
timestamp 1636986456
transform 1 0 5152 0 -1 66912
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_15
timestamp 1636986456
transform 1 0 6256 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_113_27
timestamp 18001
transform 1 0 7360 0 -1 66912
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_113_877
timestamp 1636986456
transform 1 0 85560 0 -1 66912
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_889
timestamp 1636986456
transform 1 0 86664 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_901
timestamp 18001
transform 1 0 87768 0 -1 66912
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_114_7
timestamp 1636986456
transform 1 0 5520 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_114_19
timestamp 18001
transform 1 0 6624 0 1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_114_27
timestamp 18001
transform 1 0 7360 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_114_29
timestamp 18001
transform 1 0 7544 0 1 66912
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_877
timestamp 1636986456
transform 1 0 85560 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_114_889
timestamp 18001
transform 1 0 86664 0 1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_114_897
timestamp 18001
transform 1 0 87400 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_114_903
timestamp 18001
transform 1 0 87952 0 1 66912
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_7
timestamp 1636986456
transform 1 0 5520 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_115_19
timestamp 18001
transform 1 0 6624 0 -1 68000
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_115_27
timestamp 18001
transform 1 0 7360 0 -1 68000
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_115_877
timestamp 1636986456
transform 1 0 85560 0 -1 68000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_889
timestamp 1636986456
transform 1 0 86664 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_115_901
timestamp 18001
transform 1 0 87768 0 -1 68000
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_3
timestamp 1636986456
transform 1 0 5152 0 1 68000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_15
timestamp 1636986456
transform 1 0 6256 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_116_27
timestamp 18001
transform 1 0 7360 0 1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_116_29
timestamp 18001
transform 1 0 7544 0 1 68000
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_877
timestamp 1636986456
transform 1 0 85560 0 1 68000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_889
timestamp 1636986456
transform 1 0 86664 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_116_901
timestamp 18001
transform 1 0 87768 0 1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_116_903
timestamp 18001
transform 1 0 87952 0 1 68000
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_117_3
timestamp 1636986456
transform 1 0 5152 0 -1 69088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_15
timestamp 1636986456
transform 1 0 6256 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_27
timestamp 18001
transform 1 0 7360 0 -1 69088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_877
timestamp 1636986456
transform 1 0 85560 0 -1 69088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_889
timestamp 1636986456
transform 1 0 86664 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_901
timestamp 18001
transform 1 0 87768 0 -1 69088
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_118_7
timestamp 1636986456
transform 1 0 5520 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_118_19
timestamp 18001
transform 1 0 6624 0 1 69088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_118_27
timestamp 18001
transform 1 0 7360 0 1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_118_29
timestamp 18001
transform 1 0 7544 0 1 69088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_877
timestamp 1636986456
transform 1 0 85560 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_118_889
timestamp 18001
transform 1 0 86664 0 1 69088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_118_897
timestamp 18001
transform 1 0 87400 0 1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_118_903
timestamp 18001
transform 1 0 87952 0 1 69088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_3
timestamp 1636986456
transform 1 0 5152 0 -1 70176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_15
timestamp 1636986456
transform 1 0 6256 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_119_27
timestamp 18001
transform 1 0 7360 0 -1 70176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_119_877
timestamp 1636986456
transform 1 0 85560 0 -1 70176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_889
timestamp 1636986456
transform 1 0 86664 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_901
timestamp 18001
transform 1 0 87768 0 -1 70176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_120_7
timestamp 1636986456
transform 1 0 5520 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_120_19
timestamp 18001
transform 1 0 6624 0 1 70176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_120_27
timestamp 18001
transform 1 0 7360 0 1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_120_29
timestamp 18001
transform 1 0 7544 0 1 70176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_877
timestamp 1636986456
transform 1 0 85560 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_120_889
timestamp 18001
transform 1 0 86664 0 1 70176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_120_897
timestamp 18001
transform 1 0 87400 0 1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_120_903
timestamp 18001
transform 1 0 87952 0 1 70176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_3
timestamp 1636986456
transform 1 0 5152 0 -1 71264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_15
timestamp 1636986456
transform 1 0 6256 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_121_27
timestamp 18001
transform 1 0 7360 0 -1 71264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_121_877
timestamp 1636986456
transform 1 0 85560 0 -1 71264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_889
timestamp 1636986456
transform 1 0 86664 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_901
timestamp 18001
transform 1 0 87768 0 -1 71264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_122_7
timestamp 1636986456
transform 1 0 5520 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_122_19
timestamp 18001
transform 1 0 6624 0 1 71264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_122_27
timestamp 18001
transform 1 0 7360 0 1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_122_29
timestamp 18001
transform 1 0 7544 0 1 71264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_877
timestamp 1636986456
transform 1 0 85560 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_122_889
timestamp 18001
transform 1 0 86664 0 1 71264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_122_897
timestamp 18001
transform 1 0 87400 0 1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_122_903
timestamp 18001
transform 1 0 87952 0 1 71264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_3
timestamp 1636986456
transform 1 0 5152 0 -1 72352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_15
timestamp 1636986456
transform 1 0 6256 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_27
timestamp 18001
transform 1 0 7360 0 -1 72352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_123_877
timestamp 1636986456
transform 1 0 85560 0 -1 72352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_889
timestamp 1636986456
transform 1 0 86664 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_901
timestamp 18001
transform 1 0 87768 0 -1 72352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_124_7
timestamp 1636986456
transform 1 0 5520 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_124_19
timestamp 18001
transform 1 0 6624 0 1 72352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_124_27
timestamp 18001
transform 1 0 7360 0 1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_124_29
timestamp 18001
transform 1 0 7544 0 1 72352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_877
timestamp 1636986456
transform 1 0 85560 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_124_889
timestamp 18001
transform 1 0 86664 0 1 72352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_124_897
timestamp 18001
transform 1 0 87400 0 1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_124_903
timestamp 18001
transform 1 0 87952 0 1 72352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_7
timestamp 1636986456
transform 1 0 5520 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_125_19
timestamp 18001
transform 1 0 6624 0 -1 73440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_125_27
timestamp 18001
transform 1 0 7360 0 -1 73440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_125_877
timestamp 1636986456
transform 1 0 85560 0 -1 73440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_889
timestamp 1636986456
transform 1 0 86664 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_125_901
timestamp 18001
transform 1 0 87768 0 -1 73440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_3
timestamp 1636986456
transform 1 0 5152 0 1 73440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_15
timestamp 1636986456
transform 1 0 6256 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_126_27
timestamp 18001
transform 1 0 7360 0 1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_126_29
timestamp 18001
transform 1 0 7544 0 1 73440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_877
timestamp 1636986456
transform 1 0 85560 0 1 73440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_889
timestamp 1636986456
transform 1 0 86664 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_126_901
timestamp 18001
transform 1 0 87768 0 1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_126_903
timestamp 18001
transform 1 0 87952 0 1 73440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_127_3
timestamp 1636986456
transform 1 0 5152 0 -1 74528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_15
timestamp 1636986456
transform 1 0 6256 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_127_27
timestamp 18001
transform 1 0 7360 0 -1 74528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_127_877
timestamp 1636986456
transform 1 0 85560 0 -1 74528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_889
timestamp 1636986456
transform 1 0 86664 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_901
timestamp 18001
transform 1 0 87768 0 -1 74528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_128_7
timestamp 1636986456
transform 1 0 5520 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_128_19
timestamp 18001
transform 1 0 6624 0 1 74528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_128_27
timestamp 18001
transform 1 0 7360 0 1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_128_29
timestamp 18001
transform 1 0 7544 0 1 74528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_877
timestamp 1636986456
transform 1 0 85560 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_128_889
timestamp 18001
transform 1 0 86664 0 1 74528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_128_897
timestamp 18001
transform 1 0 87400 0 1 74528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_129_3
timestamp 1636986456
transform 1 0 5152 0 -1 75616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_15
timestamp 1636986456
transform 1 0 6256 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_129_27
timestamp 18001
transform 1 0 7360 0 -1 75616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_129_877
timestamp 1636986456
transform 1 0 85560 0 -1 75616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_889
timestamp 1636986456
transform 1 0 86664 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_901
timestamp 18001
transform 1 0 87768 0 -1 75616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_130_7
timestamp 1636986456
transform 1 0 5520 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_130_19
timestamp 18001
transform 1 0 6624 0 1 75616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_130_27
timestamp 18001
transform 1 0 7360 0 1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_130_29
timestamp 18001
transform 1 0 7544 0 1 75616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_877
timestamp 1636986456
transform 1 0 85560 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_130_889
timestamp 18001
transform 1 0 86664 0 1 75616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_130_897
timestamp 18001
transform 1 0 87400 0 1 75616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_131_3
timestamp 1636986456
transform 1 0 5152 0 -1 76704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_15
timestamp 1636986456
transform 1 0 6256 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_131_27
timestamp 18001
transform 1 0 7360 0 -1 76704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_131_877
timestamp 1636986456
transform 1 0 85560 0 -1 76704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_889
timestamp 1636986456
transform 1 0 86664 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_901
timestamp 18001
transform 1 0 87768 0 -1 76704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_132_7
timestamp 1636986456
transform 1 0 5520 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_132_19
timestamp 18001
transform 1 0 6624 0 1 76704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_132_27
timestamp 18001
transform 1 0 7360 0 1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_132_29
timestamp 18001
transform 1 0 7544 0 1 76704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_877
timestamp 1636986456
transform 1 0 85560 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_132_889
timestamp 18001
transform 1 0 86664 0 1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_132_905
timestamp 18001
transform 1 0 88136 0 1 76704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_133_3
timestamp 1636986456
transform 1 0 5152 0 -1 77792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_15
timestamp 1636986456
transform 1 0 6256 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_133_27
timestamp 18001
transform 1 0 7360 0 -1 77792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_133_877
timestamp 1636986456
transform 1 0 85560 0 -1 77792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_889
timestamp 1636986456
transform 1 0 86664 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_901
timestamp 18001
transform 1 0 87768 0 -1 77792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_134_7
timestamp 1636986456
transform 1 0 5520 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_134_19
timestamp 18001
transform 1 0 6624 0 1 77792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_134_27
timestamp 18001
transform 1 0 7360 0 1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_134_29
timestamp 18001
transform 1 0 7544 0 1 77792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_877
timestamp 1636986456
transform 1 0 85560 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_134_889
timestamp 18001
transform 1 0 86664 0 1 77792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_134_897
timestamp 18001
transform 1 0 87400 0 1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_134_903
timestamp 18001
transform 1 0 87952 0 1 77792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_7
timestamp 1636986456
transform 1 0 5520 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_135_19
timestamp 18001
transform 1 0 6624 0 -1 78880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_135_27
timestamp 18001
transform 1 0 7360 0 -1 78880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_135_877
timestamp 1636986456
transform 1 0 85560 0 -1 78880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_889
timestamp 1636986456
transform 1 0 86664 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_135_901
timestamp 18001
transform 1 0 87768 0 -1 78880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_3
timestamp 1636986456
transform 1 0 5152 0 1 78880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_15
timestamp 1636986456
transform 1 0 6256 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_136_27
timestamp 18001
transform 1 0 7360 0 1 78880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_136_29
timestamp 18001
transform 1 0 7544 0 1 78880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_877
timestamp 1636986456
transform 1 0 85560 0 1 78880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_889
timestamp 1636986456
transform 1 0 86664 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_136_901
timestamp 18001
transform 1 0 87768 0 1 78880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_136_903
timestamp 18001
transform 1 0 87952 0 1 78880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_137_3
timestamp 1636986456
transform 1 0 5152 0 -1 79968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_15
timestamp 1636986456
transform 1 0 6256 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_137_27
timestamp 18001
transform 1 0 7360 0 -1 79968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_137_877
timestamp 1636986456
transform 1 0 85560 0 -1 79968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_889
timestamp 1636986456
transform 1 0 86664 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_901
timestamp 18001
transform 1 0 87768 0 -1 79968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_138_7
timestamp 1636986456
transform 1 0 5520 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_138_19
timestamp 18001
transform 1 0 6624 0 1 79968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_138_27
timestamp 18001
transform 1 0 7360 0 1 79968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_138_29
timestamp 18001
transform 1 0 7544 0 1 79968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_138_877
timestamp 1636986456
transform 1 0 85560 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_138_889
timestamp 18001
transform 1 0 86664 0 1 79968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_138_897
timestamp 18001
transform 1 0 87400 0 1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_138_903
timestamp 18001
transform 1 0 87952 0 1 79968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_139_3
timestamp 1636986456
transform 1 0 5152 0 -1 81056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_15
timestamp 1636986456
transform 1 0 6256 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_139_27
timestamp 18001
transform 1 0 7360 0 -1 81056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_139_877
timestamp 1636986456
transform 1 0 85560 0 -1 81056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_889
timestamp 1636986456
transform 1 0 86664 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_139_901
timestamp 18001
transform 1 0 87768 0 -1 81056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_140_7
timestamp 1636986456
transform 1 0 5520 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_140_19
timestamp 18001
transform 1 0 6624 0 1 81056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_140_27
timestamp 18001
transform 1 0 7360 0 1 81056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_140_29
timestamp 18001
transform 1 0 7544 0 1 81056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_140_877
timestamp 1636986456
transform 1 0 85560 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_140_889
timestamp 18001
transform 1 0 86664 0 1 81056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_140_897
timestamp 18001
transform 1 0 87400 0 1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_140_903
timestamp 18001
transform 1 0 87952 0 1 81056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_141_3
timestamp 1636986456
transform 1 0 5152 0 -1 82144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_15
timestamp 1636986456
transform 1 0 6256 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_141_27
timestamp 18001
transform 1 0 7360 0 -1 82144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_141_877
timestamp 1636986456
transform 1 0 85560 0 -1 82144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_889
timestamp 1636986456
transform 1 0 86664 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_141_901
timestamp 18001
transform 1 0 87768 0 -1 82144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_142_3
timestamp 1636986456
transform 1 0 5152 0 1 82144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_15
timestamp 1636986456
transform 1 0 6256 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_142_27
timestamp 18001
transform 1 0 7360 0 1 82144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_142_29
timestamp 18001
transform 1 0 7544 0 1 82144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_142_877
timestamp 1636986456
transform 1 0 85560 0 1 82144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_889
timestamp 1636986456
transform 1 0 86664 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_142_901
timestamp 18001
transform 1 0 87768 0 1 82144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_142_903
timestamp 18001
transform 1 0 87952 0 1 82144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_143_3
timestamp 1636986456
transform 1 0 5152 0 -1 83232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_15
timestamp 1636986456
transform 1 0 6256 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_143_27
timestamp 18001
transform 1 0 7360 0 -1 83232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_143_877
timestamp 1636986456
transform 1 0 85560 0 -1 83232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_889
timestamp 1636986456
transform 1 0 86664 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_143_901
timestamp 18001
transform 1 0 87768 0 -1 83232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_144_3
timestamp 1636986456
transform 1 0 5152 0 1 83232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_15
timestamp 1636986456
transform 1 0 6256 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_144_27
timestamp 18001
transform 1 0 7360 0 1 83232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_144_29
timestamp 18001
transform 1 0 7544 0 1 83232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_144_877
timestamp 1636986456
transform 1 0 85560 0 1 83232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_889
timestamp 1636986456
transform 1 0 86664 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_144_901
timestamp 18001
transform 1 0 87768 0 1 83232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_144_903
timestamp 18001
transform 1 0 87952 0 1 83232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_145_3
timestamp 1636986456
transform 1 0 5152 0 -1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_15
timestamp 1636986456
transform 1 0 6256 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_145_27
timestamp 18001
transform 1 0 7360 0 -1 84320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_145_877
timestamp 1636986456
transform 1 0 85560 0 -1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_889
timestamp 1636986456
transform 1 0 86664 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_145_901
timestamp 18001
transform 1 0 87768 0 -1 84320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_146_3
timestamp 1636986456
transform 1 0 5152 0 1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_15
timestamp 1636986456
transform 1 0 6256 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_146_27
timestamp 18001
transform 1 0 7360 0 1 84320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_146_29
timestamp 1636986456
transform 1 0 7544 0 1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_41
timestamp 1636986456
transform 1 0 8648 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_146_53
timestamp 18001
transform 1 0 9752 0 1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_146_57
timestamp 18001
transform 1 0 10120 0 1 84320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_146_61
timestamp 18001
transform 1 0 10488 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_146_64
timestamp 18001
transform 1 0 10764 0 1 84320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_146_72
timestamp 18001
transform 1 0 11500 0 1 84320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_146_76
timestamp 18001
transform 1 0 11868 0 1 84320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_146_85
timestamp 18001
transform 1 0 12696 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_146_88
timestamp 18001
transform 1 0 12972 0 1 84320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_146_96
timestamp 18001
transform 1 0 13708 0 1 84320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_146_100
timestamp 1636986456
transform 1 0 14076 0 1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_113
timestamp 1636986456
transform 1 0 15272 0 1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_125
timestamp 1636986456
transform 1 0 16376 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_146_137
timestamp 18001
transform 1 0 17480 0 1 84320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_146_141
timestamp 1636986456
transform 1 0 17848 0 1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_153
timestamp 1636986456
transform 1 0 18952 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_146_165
timestamp 18001
transform 1 0 20056 0 1 84320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_146_169
timestamp 1636986456
transform 1 0 20424 0 1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_181
timestamp 1636986456
transform 1 0 21528 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_146_193
timestamp 18001
transform 1 0 22632 0 1 84320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_146_197
timestamp 1636986456
transform 1 0 23000 0 1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_209
timestamp 1636986456
transform 1 0 24104 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_146_221
timestamp 18001
transform 1 0 25208 0 1 84320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_146_225
timestamp 1636986456
transform 1 0 25576 0 1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_237
timestamp 1636986456
transform 1 0 26680 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_146_249
timestamp 18001
transform 1 0 27784 0 1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_146_253
timestamp 18001
transform 1 0 28152 0 1 84320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_146_259
timestamp 18001
transform 1 0 28704 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_146_281
timestamp 18001
transform 1 0 30728 0 1 84320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_146_286
timestamp 1636986456
transform 1 0 31188 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_146_298
timestamp 18001
transform 1 0 32292 0 1 84320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_146_306
timestamp 18001
transform 1 0 33028 0 1 84320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_146_309
timestamp 1636986456
transform 1 0 33304 0 1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_321
timestamp 1636986456
transform 1 0 34408 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_146_333
timestamp 18001
transform 1 0 35512 0 1 84320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_146_337
timestamp 1636986456
transform 1 0 35880 0 1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_349
timestamp 1636986456
transform 1 0 36984 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_146_361
timestamp 18001
transform 1 0 38088 0 1 84320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_146_365
timestamp 1636986456
transform 1 0 38456 0 1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_377
timestamp 1636986456
transform 1 0 39560 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_146_389
timestamp 18001
transform 1 0 40664 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_146_415
timestamp 18001
transform 1 0 43056 0 1 84320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_146_419
timestamp 18001
transform 1 0 43424 0 1 84320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_146_421
timestamp 1636986456
transform 1 0 43608 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_146_433
timestamp 18001
transform 1 0 44712 0 1 84320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_146_439
timestamp 18001
transform 1 0 45264 0 1 84320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_146_449
timestamp 1636986456
transform 1 0 46184 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_146_461
timestamp 18001
transform 1 0 47288 0 1 84320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_146_471
timestamp 18001
transform 1 0 48208 0 1 84320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_146_475
timestamp 18001
transform 1 0 48576 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_146_477
timestamp 18001
transform 1 0 48760 0 1 84320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_146_483
timestamp 18001
transform 1 0 49312 0 1 84320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_146_491
timestamp 18001
transform 1 0 50048 0 1 84320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_146_495
timestamp 18001
transform 1 0 50416 0 1 84320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_146_503
timestamp 18001
transform 1 0 51152 0 1 84320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_146_507
timestamp 1636986456
transform 1 0 51520 0 1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_519
timestamp 1636986456
transform 1 0 52624 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_146_531
timestamp 18001
transform 1 0 53728 0 1 84320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_146_533
timestamp 1636986456
transform 1 0 53912 0 1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_545
timestamp 1636986456
transform 1 0 55016 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_146_557
timestamp 18001
transform 1 0 56120 0 1 84320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_146_561
timestamp 1636986456
transform 1 0 56488 0 1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_573
timestamp 1636986456
transform 1 0 57592 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_146_585
timestamp 18001
transform 1 0 58696 0 1 84320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_146_589
timestamp 1636986456
transform 1 0 59064 0 1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_601
timestamp 1636986456
transform 1 0 60168 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_146_613
timestamp 18001
transform 1 0 61272 0 1 84320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_146_617
timestamp 1636986456
transform 1 0 61640 0 1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_629
timestamp 1636986456
transform 1 0 62744 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_146_641
timestamp 18001
transform 1 0 63848 0 1 84320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_146_645
timestamp 1636986456
transform 1 0 64216 0 1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_657
timestamp 1636986456
transform 1 0 65320 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_146_669
timestamp 18001
transform 1 0 66424 0 1 84320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_146_673
timestamp 1636986456
transform 1 0 66792 0 1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_685
timestamp 1636986456
transform 1 0 67896 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_146_697
timestamp 18001
transform 1 0 69000 0 1 84320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_146_701
timestamp 1636986456
transform 1 0 69368 0 1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_713
timestamp 1636986456
transform 1 0 70472 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_146_725
timestamp 18001
transform 1 0 71576 0 1 84320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_146_729
timestamp 1636986456
transform 1 0 71944 0 1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_741
timestamp 1636986456
transform 1 0 73048 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_146_753
timestamp 18001
transform 1 0 74152 0 1 84320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_146_757
timestamp 1636986456
transform 1 0 74520 0 1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_769
timestamp 1636986456
transform 1 0 75624 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_146_781
timestamp 18001
transform 1 0 76728 0 1 84320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_146_785
timestamp 1636986456
transform 1 0 77096 0 1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_797
timestamp 1636986456
transform 1 0 78200 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_146_809
timestamp 18001
transform 1 0 79304 0 1 84320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_146_813
timestamp 1636986456
transform 1 0 79672 0 1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_825
timestamp 1636986456
transform 1 0 80776 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_146_837
timestamp 18001
transform 1 0 81880 0 1 84320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_146_841
timestamp 1636986456
transform 1 0 82248 0 1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_853
timestamp 1636986456
transform 1 0 83352 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_146_865
timestamp 18001
transform 1 0 84456 0 1 84320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_146_869
timestamp 1636986456
transform 1 0 84824 0 1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_881
timestamp 1636986456
transform 1 0 85928 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_146_893
timestamp 18001
transform 1 0 87032 0 1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_146_897
timestamp 18001
transform 1 0 87400 0 1 84320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_146_905
timestamp 18001
transform 1 0 88136 0 1 84320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_147_3
timestamp 1636986456
transform 1 0 5152 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_15
timestamp 1636986456
transform 1 0 6256 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_27
timestamp 1636986456
transform 1 0 7360 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_39
timestamp 1636986456
transform 1 0 8464 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_147_51
timestamp 18001
transform 1 0 9568 0 -1 85408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_147_55
timestamp 18001
transform 1 0 9936 0 -1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_57
timestamp 1636986456
transform 1 0 10120 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_69
timestamp 1636986456
transform 1 0 11224 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_81
timestamp 1636986456
transform 1 0 12328 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_93
timestamp 1636986456
transform 1 0 13432 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_105
timestamp 18001
transform 1 0 14536 0 -1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_111
timestamp 18001
transform 1 0 15088 0 -1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_113
timestamp 1636986456
transform 1 0 15272 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_125
timestamp 1636986456
transform 1 0 16376 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_137
timestamp 1636986456
transform 1 0 17480 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_149
timestamp 1636986456
transform 1 0 18584 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_161
timestamp 18001
transform 1 0 19688 0 -1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_167
timestamp 18001
transform 1 0 20240 0 -1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_169
timestamp 1636986456
transform 1 0 20424 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_181
timestamp 1636986456
transform 1 0 21528 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_193
timestamp 1636986456
transform 1 0 22632 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_205
timestamp 1636986456
transform 1 0 23736 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_217
timestamp 18001
transform 1 0 24840 0 -1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_223
timestamp 18001
transform 1 0 25392 0 -1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_225
timestamp 1636986456
transform 1 0 25576 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_237
timestamp 1636986456
transform 1 0 26680 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_249
timestamp 1636986456
transform 1 0 27784 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_261
timestamp 1636986456
transform 1 0 28888 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_273
timestamp 18001
transform 1 0 29992 0 -1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_279
timestamp 18001
transform 1 0 30544 0 -1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_281
timestamp 1636986456
transform 1 0 30728 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_293
timestamp 1636986456
transform 1 0 31832 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_305
timestamp 1636986456
transform 1 0 32936 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_317
timestamp 1636986456
transform 1 0 34040 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_329
timestamp 18001
transform 1 0 35144 0 -1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_335
timestamp 18001
transform 1 0 35696 0 -1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_337
timestamp 1636986456
transform 1 0 35880 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_349
timestamp 1636986456
transform 1 0 36984 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_361
timestamp 1636986456
transform 1 0 38088 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_373
timestamp 1636986456
transform 1 0 39192 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_385
timestamp 18001
transform 1 0 40296 0 -1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_391
timestamp 18001
transform 1 0 40848 0 -1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_393
timestamp 1636986456
transform 1 0 41032 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_405
timestamp 1636986456
transform 1 0 42136 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_417
timestamp 1636986456
transform 1 0 43240 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_429
timestamp 1636986456
transform 1 0 44344 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_441
timestamp 18001
transform 1 0 45448 0 -1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_447
timestamp 18001
transform 1 0 46000 0 -1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_449
timestamp 1636986456
transform 1 0 46184 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_461
timestamp 1636986456
transform 1 0 47288 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_473
timestamp 1636986456
transform 1 0 48392 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_485
timestamp 1636986456
transform 1 0 49496 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_497
timestamp 18001
transform 1 0 50600 0 -1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_503
timestamp 18001
transform 1 0 51152 0 -1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_505
timestamp 1636986456
transform 1 0 51336 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_517
timestamp 1636986456
transform 1 0 52440 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_529
timestamp 1636986456
transform 1 0 53544 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_541
timestamp 1636986456
transform 1 0 54648 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_553
timestamp 18001
transform 1 0 55752 0 -1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_559
timestamp 18001
transform 1 0 56304 0 -1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_561
timestamp 1636986456
transform 1 0 56488 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_573
timestamp 1636986456
transform 1 0 57592 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_585
timestamp 1636986456
transform 1 0 58696 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_597
timestamp 1636986456
transform 1 0 59800 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_609
timestamp 18001
transform 1 0 60904 0 -1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_615
timestamp 18001
transform 1 0 61456 0 -1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_617
timestamp 1636986456
transform 1 0 61640 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_629
timestamp 1636986456
transform 1 0 62744 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_641
timestamp 1636986456
transform 1 0 63848 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_653
timestamp 1636986456
transform 1 0 64952 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_665
timestamp 18001
transform 1 0 66056 0 -1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_671
timestamp 18001
transform 1 0 66608 0 -1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_673
timestamp 1636986456
transform 1 0 66792 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_685
timestamp 1636986456
transform 1 0 67896 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_697
timestamp 1636986456
transform 1 0 69000 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_709
timestamp 1636986456
transform 1 0 70104 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_721
timestamp 18001
transform 1 0 71208 0 -1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_727
timestamp 18001
transform 1 0 71760 0 -1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_729
timestamp 1636986456
transform 1 0 71944 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_741
timestamp 1636986456
transform 1 0 73048 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_753
timestamp 1636986456
transform 1 0 74152 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_765
timestamp 1636986456
transform 1 0 75256 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_777
timestamp 18001
transform 1 0 76360 0 -1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_783
timestamp 18001
transform 1 0 76912 0 -1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_785
timestamp 1636986456
transform 1 0 77096 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_797
timestamp 1636986456
transform 1 0 78200 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_809
timestamp 1636986456
transform 1 0 79304 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_821
timestamp 1636986456
transform 1 0 80408 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_833
timestamp 18001
transform 1 0 81512 0 -1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_839
timestamp 18001
transform 1 0 82064 0 -1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_841
timestamp 1636986456
transform 1 0 82248 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_853
timestamp 1636986456
transform 1 0 83352 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_865
timestamp 1636986456
transform 1 0 84456 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_877
timestamp 1636986456
transform 1 0 85560 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_889
timestamp 18001
transform 1 0 86664 0 -1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_895
timestamp 18001
transform 1 0 87216 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_147_897
timestamp 18001
transform 1 0 87400 0 -1 85408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_147_905
timestamp 18001
transform 1 0 88136 0 -1 85408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_148_3
timestamp 1636986456
transform 1 0 5152 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_15
timestamp 1636986456
transform 1 0 6256 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_148_27
timestamp 18001
transform 1 0 7360 0 1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_29
timestamp 1636986456
transform 1 0 7544 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_41
timestamp 1636986456
transform 1 0 8648 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_53
timestamp 1636986456
transform 1 0 9752 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_65
timestamp 1636986456
transform 1 0 10856 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_77
timestamp 18001
transform 1 0 11960 0 1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_83
timestamp 18001
transform 1 0 12512 0 1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_85
timestamp 1636986456
transform 1 0 12696 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_97
timestamp 1636986456
transform 1 0 13800 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_109
timestamp 1636986456
transform 1 0 14904 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_121
timestamp 1636986456
transform 1 0 16008 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_133
timestamp 18001
transform 1 0 17112 0 1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_139
timestamp 18001
transform 1 0 17664 0 1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_141
timestamp 1636986456
transform 1 0 17848 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_153
timestamp 1636986456
transform 1 0 18952 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_165
timestamp 1636986456
transform 1 0 20056 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_177
timestamp 1636986456
transform 1 0 21160 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_189
timestamp 18001
transform 1 0 22264 0 1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_195
timestamp 18001
transform 1 0 22816 0 1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_197
timestamp 1636986456
transform 1 0 23000 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_209
timestamp 1636986456
transform 1 0 24104 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_221
timestamp 1636986456
transform 1 0 25208 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_233
timestamp 1636986456
transform 1 0 26312 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_245
timestamp 18001
transform 1 0 27416 0 1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_251
timestamp 18001
transform 1 0 27968 0 1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_253
timestamp 1636986456
transform 1 0 28152 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_265
timestamp 1636986456
transform 1 0 29256 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_277
timestamp 1636986456
transform 1 0 30360 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_289
timestamp 1636986456
transform 1 0 31464 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_301
timestamp 18001
transform 1 0 32568 0 1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_307
timestamp 18001
transform 1 0 33120 0 1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_309
timestamp 1636986456
transform 1 0 33304 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_321
timestamp 1636986456
transform 1 0 34408 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_333
timestamp 1636986456
transform 1 0 35512 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_345
timestamp 1636986456
transform 1 0 36616 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_357
timestamp 18001
transform 1 0 37720 0 1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_363
timestamp 18001
transform 1 0 38272 0 1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_365
timestamp 1636986456
transform 1 0 38456 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_377
timestamp 1636986456
transform 1 0 39560 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_389
timestamp 1636986456
transform 1 0 40664 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_401
timestamp 1636986456
transform 1 0 41768 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_413
timestamp 18001
transform 1 0 42872 0 1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_419
timestamp 18001
transform 1 0 43424 0 1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_421
timestamp 1636986456
transform 1 0 43608 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_433
timestamp 1636986456
transform 1 0 44712 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_445
timestamp 1636986456
transform 1 0 45816 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_457
timestamp 1636986456
transform 1 0 46920 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_469
timestamp 18001
transform 1 0 48024 0 1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_475
timestamp 18001
transform 1 0 48576 0 1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_477
timestamp 1636986456
transform 1 0 48760 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_489
timestamp 1636986456
transform 1 0 49864 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_501
timestamp 1636986456
transform 1 0 50968 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_513
timestamp 1636986456
transform 1 0 52072 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_525
timestamp 18001
transform 1 0 53176 0 1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_531
timestamp 18001
transform 1 0 53728 0 1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_533
timestamp 1636986456
transform 1 0 53912 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_545
timestamp 1636986456
transform 1 0 55016 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_557
timestamp 1636986456
transform 1 0 56120 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_569
timestamp 1636986456
transform 1 0 57224 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_581
timestamp 18001
transform 1 0 58328 0 1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_587
timestamp 18001
transform 1 0 58880 0 1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_589
timestamp 1636986456
transform 1 0 59064 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_601
timestamp 1636986456
transform 1 0 60168 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_613
timestamp 1636986456
transform 1 0 61272 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_625
timestamp 1636986456
transform 1 0 62376 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_637
timestamp 18001
transform 1 0 63480 0 1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_643
timestamp 18001
transform 1 0 64032 0 1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_645
timestamp 1636986456
transform 1 0 64216 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_657
timestamp 1636986456
transform 1 0 65320 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_669
timestamp 1636986456
transform 1 0 66424 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_681
timestamp 1636986456
transform 1 0 67528 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_693
timestamp 18001
transform 1 0 68632 0 1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_699
timestamp 18001
transform 1 0 69184 0 1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_701
timestamp 1636986456
transform 1 0 69368 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_713
timestamp 1636986456
transform 1 0 70472 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_725
timestamp 1636986456
transform 1 0 71576 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_737
timestamp 1636986456
transform 1 0 72680 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_749
timestamp 18001
transform 1 0 73784 0 1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_755
timestamp 18001
transform 1 0 74336 0 1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_757
timestamp 1636986456
transform 1 0 74520 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_769
timestamp 1636986456
transform 1 0 75624 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_781
timestamp 1636986456
transform 1 0 76728 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_793
timestamp 1636986456
transform 1 0 77832 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_805
timestamp 18001
transform 1 0 78936 0 1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_811
timestamp 18001
transform 1 0 79488 0 1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_813
timestamp 1636986456
transform 1 0 79672 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_825
timestamp 1636986456
transform 1 0 80776 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_837
timestamp 1636986456
transform 1 0 81880 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_849
timestamp 1636986456
transform 1 0 82984 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_861
timestamp 18001
transform 1 0 84088 0 1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_867
timestamp 18001
transform 1 0 84640 0 1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_869
timestamp 1636986456
transform 1 0 84824 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_881
timestamp 1636986456
transform 1 0 85928 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_893
timestamp 1636986456
transform 1 0 87032 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_148_905
timestamp 18001
transform 1 0 88136 0 1 85408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_149_3
timestamp 1636986456
transform 1 0 5152 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_15
timestamp 1636986456
transform 1 0 6256 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_27
timestamp 1636986456
transform 1 0 7360 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_39
timestamp 1636986456
transform 1 0 8464 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_149_51
timestamp 18001
transform 1 0 9568 0 -1 86496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_149_55
timestamp 18001
transform 1 0 9936 0 -1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_57
timestamp 1636986456
transform 1 0 10120 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_69
timestamp 1636986456
transform 1 0 11224 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_81
timestamp 1636986456
transform 1 0 12328 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_93
timestamp 1636986456
transform 1 0 13432 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_105
timestamp 18001
transform 1 0 14536 0 -1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_111
timestamp 18001
transform 1 0 15088 0 -1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_113
timestamp 1636986456
transform 1 0 15272 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_125
timestamp 1636986456
transform 1 0 16376 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_137
timestamp 1636986456
transform 1 0 17480 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_149
timestamp 1636986456
transform 1 0 18584 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_161
timestamp 18001
transform 1 0 19688 0 -1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_167
timestamp 18001
transform 1 0 20240 0 -1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_169
timestamp 1636986456
transform 1 0 20424 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_181
timestamp 1636986456
transform 1 0 21528 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_193
timestamp 1636986456
transform 1 0 22632 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_205
timestamp 1636986456
transform 1 0 23736 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_217
timestamp 18001
transform 1 0 24840 0 -1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_223
timestamp 18001
transform 1 0 25392 0 -1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_225
timestamp 1636986456
transform 1 0 25576 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_237
timestamp 1636986456
transform 1 0 26680 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_249
timestamp 1636986456
transform 1 0 27784 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_261
timestamp 1636986456
transform 1 0 28888 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_273
timestamp 18001
transform 1 0 29992 0 -1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_279
timestamp 18001
transform 1 0 30544 0 -1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_281
timestamp 1636986456
transform 1 0 30728 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_293
timestamp 1636986456
transform 1 0 31832 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_305
timestamp 1636986456
transform 1 0 32936 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_317
timestamp 1636986456
transform 1 0 34040 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_329
timestamp 18001
transform 1 0 35144 0 -1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_335
timestamp 18001
transform 1 0 35696 0 -1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_337
timestamp 1636986456
transform 1 0 35880 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_349
timestamp 1636986456
transform 1 0 36984 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_361
timestamp 1636986456
transform 1 0 38088 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_373
timestamp 1636986456
transform 1 0 39192 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_385
timestamp 18001
transform 1 0 40296 0 -1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_391
timestamp 18001
transform 1 0 40848 0 -1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_393
timestamp 1636986456
transform 1 0 41032 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_405
timestamp 1636986456
transform 1 0 42136 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_417
timestamp 1636986456
transform 1 0 43240 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_429
timestamp 1636986456
transform 1 0 44344 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_441
timestamp 18001
transform 1 0 45448 0 -1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_447
timestamp 18001
transform 1 0 46000 0 -1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_449
timestamp 1636986456
transform 1 0 46184 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_461
timestamp 1636986456
transform 1 0 47288 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_473
timestamp 1636986456
transform 1 0 48392 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_485
timestamp 1636986456
transform 1 0 49496 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_497
timestamp 18001
transform 1 0 50600 0 -1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_503
timestamp 18001
transform 1 0 51152 0 -1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_505
timestamp 1636986456
transform 1 0 51336 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_517
timestamp 1636986456
transform 1 0 52440 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_529
timestamp 1636986456
transform 1 0 53544 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_541
timestamp 1636986456
transform 1 0 54648 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_553
timestamp 18001
transform 1 0 55752 0 -1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_559
timestamp 18001
transform 1 0 56304 0 -1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_561
timestamp 1636986456
transform 1 0 56488 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_573
timestamp 1636986456
transform 1 0 57592 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_585
timestamp 1636986456
transform 1 0 58696 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_597
timestamp 1636986456
transform 1 0 59800 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_609
timestamp 18001
transform 1 0 60904 0 -1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_615
timestamp 18001
transform 1 0 61456 0 -1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_617
timestamp 1636986456
transform 1 0 61640 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_629
timestamp 1636986456
transform 1 0 62744 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_641
timestamp 1636986456
transform 1 0 63848 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_653
timestamp 1636986456
transform 1 0 64952 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_665
timestamp 18001
transform 1 0 66056 0 -1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_671
timestamp 18001
transform 1 0 66608 0 -1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_673
timestamp 1636986456
transform 1 0 66792 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_685
timestamp 1636986456
transform 1 0 67896 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_697
timestamp 1636986456
transform 1 0 69000 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_709
timestamp 1636986456
transform 1 0 70104 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_721
timestamp 18001
transform 1 0 71208 0 -1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_727
timestamp 18001
transform 1 0 71760 0 -1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_729
timestamp 1636986456
transform 1 0 71944 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_741
timestamp 1636986456
transform 1 0 73048 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_753
timestamp 1636986456
transform 1 0 74152 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_765
timestamp 1636986456
transform 1 0 75256 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_777
timestamp 18001
transform 1 0 76360 0 -1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_783
timestamp 18001
transform 1 0 76912 0 -1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_785
timestamp 1636986456
transform 1 0 77096 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_797
timestamp 1636986456
transform 1 0 78200 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_809
timestamp 1636986456
transform 1 0 79304 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_821
timestamp 1636986456
transform 1 0 80408 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_833
timestamp 18001
transform 1 0 81512 0 -1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_839
timestamp 18001
transform 1 0 82064 0 -1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_841
timestamp 1636986456
transform 1 0 82248 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_853
timestamp 1636986456
transform 1 0 83352 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_865
timestamp 1636986456
transform 1 0 84456 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_877
timestamp 1636986456
transform 1 0 85560 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_889
timestamp 18001
transform 1 0 86664 0 -1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_895
timestamp 18001
transform 1 0 87216 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_149_897
timestamp 18001
transform 1 0 87400 0 -1 86496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_149_905
timestamp 18001
transform 1 0 88136 0 -1 86496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_150_3
timestamp 1636986456
transform 1 0 5152 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_15
timestamp 1636986456
transform 1 0 6256 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_150_27
timestamp 18001
transform 1 0 7360 0 1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_29
timestamp 1636986456
transform 1 0 7544 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_41
timestamp 1636986456
transform 1 0 8648 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_53
timestamp 1636986456
transform 1 0 9752 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_65
timestamp 1636986456
transform 1 0 10856 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_77
timestamp 18001
transform 1 0 11960 0 1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_83
timestamp 18001
transform 1 0 12512 0 1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_85
timestamp 1636986456
transform 1 0 12696 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_97
timestamp 1636986456
transform 1 0 13800 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_109
timestamp 1636986456
transform 1 0 14904 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_121
timestamp 1636986456
transform 1 0 16008 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_133
timestamp 18001
transform 1 0 17112 0 1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_139
timestamp 18001
transform 1 0 17664 0 1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_141
timestamp 1636986456
transform 1 0 17848 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_153
timestamp 1636986456
transform 1 0 18952 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_165
timestamp 1636986456
transform 1 0 20056 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_177
timestamp 1636986456
transform 1 0 21160 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_189
timestamp 18001
transform 1 0 22264 0 1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_195
timestamp 18001
transform 1 0 22816 0 1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_197
timestamp 1636986456
transform 1 0 23000 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_209
timestamp 1636986456
transform 1 0 24104 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_221
timestamp 1636986456
transform 1 0 25208 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_233
timestamp 1636986456
transform 1 0 26312 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_245
timestamp 18001
transform 1 0 27416 0 1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_251
timestamp 18001
transform 1 0 27968 0 1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_253
timestamp 1636986456
transform 1 0 28152 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_265
timestamp 1636986456
transform 1 0 29256 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_277
timestamp 1636986456
transform 1 0 30360 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_289
timestamp 1636986456
transform 1 0 31464 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_301
timestamp 18001
transform 1 0 32568 0 1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_307
timestamp 18001
transform 1 0 33120 0 1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_309
timestamp 1636986456
transform 1 0 33304 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_321
timestamp 1636986456
transform 1 0 34408 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_333
timestamp 1636986456
transform 1 0 35512 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_150_345
timestamp 18001
transform 1 0 36616 0 1 86496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_150_353
timestamp 18001
transform 1 0 37352 0 1 86496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_150_359
timestamp 18001
transform 1 0 37904 0 1 86496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_150_363
timestamp 18001
transform 1 0 38272 0 1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_367
timestamp 1636986456
transform 1 0 38640 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_379
timestamp 1636986456
transform 1 0 39744 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_391
timestamp 1636986456
transform 1 0 40848 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_403
timestamp 1636986456
transform 1 0 41952 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_150_415
timestamp 18001
transform 1 0 43056 0 1 86496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_150_419
timestamp 18001
transform 1 0 43424 0 1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_421
timestamp 1636986456
transform 1 0 43608 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_433
timestamp 1636986456
transform 1 0 44712 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_445
timestamp 1636986456
transform 1 0 45816 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_457
timestamp 1636986456
transform 1 0 46920 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_469
timestamp 18001
transform 1 0 48024 0 1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_475
timestamp 18001
transform 1 0 48576 0 1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_477
timestamp 1636986456
transform 1 0 48760 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_489
timestamp 1636986456
transform 1 0 49864 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_501
timestamp 1636986456
transform 1 0 50968 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_513
timestamp 1636986456
transform 1 0 52072 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_525
timestamp 18001
transform 1 0 53176 0 1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_531
timestamp 18001
transform 1 0 53728 0 1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_533
timestamp 1636986456
transform 1 0 53912 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_545
timestamp 1636986456
transform 1 0 55016 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_557
timestamp 1636986456
transform 1 0 56120 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_569
timestamp 1636986456
transform 1 0 57224 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_581
timestamp 18001
transform 1 0 58328 0 1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_587
timestamp 18001
transform 1 0 58880 0 1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_589
timestamp 1636986456
transform 1 0 59064 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_601
timestamp 1636986456
transform 1 0 60168 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_613
timestamp 1636986456
transform 1 0 61272 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_625
timestamp 1636986456
transform 1 0 62376 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_637
timestamp 18001
transform 1 0 63480 0 1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_643
timestamp 18001
transform 1 0 64032 0 1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_645
timestamp 1636986456
transform 1 0 64216 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_657
timestamp 1636986456
transform 1 0 65320 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_669
timestamp 1636986456
transform 1 0 66424 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_681
timestamp 1636986456
transform 1 0 67528 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_693
timestamp 18001
transform 1 0 68632 0 1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_699
timestamp 18001
transform 1 0 69184 0 1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_701
timestamp 1636986456
transform 1 0 69368 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_713
timestamp 1636986456
transform 1 0 70472 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_725
timestamp 1636986456
transform 1 0 71576 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_737
timestamp 1636986456
transform 1 0 72680 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_749
timestamp 18001
transform 1 0 73784 0 1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_755
timestamp 18001
transform 1 0 74336 0 1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_757
timestamp 1636986456
transform 1 0 74520 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_769
timestamp 1636986456
transform 1 0 75624 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_781
timestamp 1636986456
transform 1 0 76728 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_793
timestamp 1636986456
transform 1 0 77832 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_805
timestamp 18001
transform 1 0 78936 0 1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_811
timestamp 18001
transform 1 0 79488 0 1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_813
timestamp 1636986456
transform 1 0 79672 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_825
timestamp 1636986456
transform 1 0 80776 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_837
timestamp 1636986456
transform 1 0 81880 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_849
timestamp 1636986456
transform 1 0 82984 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_861
timestamp 18001
transform 1 0 84088 0 1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_867
timestamp 18001
transform 1 0 84640 0 1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_869
timestamp 1636986456
transform 1 0 84824 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_881
timestamp 1636986456
transform 1 0 85928 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_893
timestamp 1636986456
transform 1 0 87032 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_150_905
timestamp 18001
transform 1 0 88136 0 1 86496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_151_3
timestamp 1636986456
transform 1 0 5152 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_15
timestamp 1636986456
transform 1 0 6256 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_151_27
timestamp 18001
transform 1 0 7360 0 -1 87584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_151_29
timestamp 1636986456
transform 1 0 7544 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_41
timestamp 1636986456
transform 1 0 8648 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_151_53
timestamp 18001
transform 1 0 9752 0 -1 87584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_151_57
timestamp 1636986456
transform 1 0 10120 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_69
timestamp 1636986456
transform 1 0 11224 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_151_81
timestamp 18001
transform 1 0 12328 0 -1 87584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_151_85
timestamp 1636986456
transform 1 0 12696 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_97
timestamp 1636986456
transform 1 0 13800 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_151_109
timestamp 18001
transform 1 0 14904 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_151_130
timestamp 18001
transform 1 0 16836 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_151_139
timestamp 18001
transform 1 0 17664 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_151_141
timestamp 18001
transform 1 0 17848 0 -1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_147
timestamp 18001
transform 1 0 18400 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_151_153
timestamp 18001
transform 1 0 18952 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_151_160
timestamp 18001
transform 1 0 19596 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_151_174
timestamp 18001
transform 1 0 20884 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_151_182
timestamp 18001
transform 1 0 21620 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_151_188
timestamp 18001
transform 1 0 22172 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_151_202
timestamp 18001
transform 1 0 23460 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_151_209
timestamp 18001
transform 1 0 24104 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_151_217
timestamp 18001
transform 1 0 24840 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_151_223
timestamp 18001
transform 1 0 25392 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_151_225
timestamp 18001
transform 1 0 25576 0 -1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_231
timestamp 18001
transform 1 0 26128 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_151_237
timestamp 18001
transform 1 0 26680 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_151_244
timestamp 18001
transform 1 0 27324 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_151_258
timestamp 18001
transform 1 0 28612 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_151_266
timestamp 18001
transform 1 0 29348 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_151_272
timestamp 18001
transform 1 0 29900 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_151_285
timestamp 18001
transform 1 0 31096 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_151_292
timestamp 18001
transform 1 0 31740 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_151_300
timestamp 18001
transform 1 0 32476 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_151_306
timestamp 18001
transform 1 0 33028 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_151_309
timestamp 18001
transform 1 0 33304 0 -1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_315
timestamp 18001
transform 1 0 33856 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_151_320
timestamp 18001
transform 1 0 34316 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_151_327
timestamp 18001
transform 1 0 34960 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_151_335
timestamp 18001
transform 1 0 35696 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_151_341
timestamp 18001
transform 1 0 36248 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_151_359
timestamp 18001
transform 1 0 37904 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_151_382
timestamp 18001
transform 1 0 40020 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_151_390
timestamp 18001
transform 1 0 40756 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_151_397
timestamp 18001
transform 1 0 41400 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_151_403
timestamp 18001
transform 1 0 41952 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_151_411
timestamp 18001
transform 1 0 42688 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_151_417
timestamp 18001
transform 1 0 43240 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_151_425
timestamp 18001
transform 1 0 43976 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_151_432
timestamp 18001
transform 1 0 44620 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_151_438
timestamp 18001
transform 1 0 45172 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_151_445
timestamp 18001
transform 1 0 45816 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_151_452
timestamp 18001
transform 1 0 46460 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_151_459
timestamp 18001
transform 1 0 47104 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_151_466
timestamp 18001
transform 1 0 47748 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_151_473
timestamp 18001
transform 1 0 48392 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_151_480
timestamp 18001
transform 1 0 49036 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_151_487
timestamp 18001
transform 1 0 49680 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_151_494
timestamp 18001
transform 1 0 50324 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_151_502
timestamp 18001
transform 1 0 51060 0 -1 87584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_151_505
timestamp 1636986456
transform 1 0 51336 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_151_517
timestamp 18001
transform 1 0 52440 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_151_537
timestamp 18001
transform 1 0 54280 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_151_545
timestamp 18001
transform 1 0 55016 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_151_553
timestamp 18001
transform 1 0 55752 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_151_559
timestamp 18001
transform 1 0 56304 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_151_561
timestamp 18001
transform 1 0 56488 0 -1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_567
timestamp 18001
transform 1 0 57040 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_151_573
timestamp 18001
transform 1 0 57592 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_151_580
timestamp 18001
transform 1 0 58236 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_151_594
timestamp 18001
transform 1 0 59524 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_151_602
timestamp 18001
transform 1 0 60260 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_151_608
timestamp 18001
transform 1 0 60812 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_151_615
timestamp 18001
transform 1 0 61456 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_151_617
timestamp 18001
transform 1 0 61640 0 -1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_623
timestamp 18001
transform 1 0 62192 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_151_629
timestamp 18001
transform 1 0 62744 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_151_637
timestamp 18001
transform 1 0 63480 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_151_643
timestamp 18001
transform 1 0 64032 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_151_645
timestamp 18001
transform 1 0 64216 0 -1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_651
timestamp 18001
transform 1 0 64768 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_151_657
timestamp 18001
transform 1 0 65320 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_151_664
timestamp 18001
transform 1 0 65964 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_151_678
timestamp 18001
transform 1 0 67252 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_151_686
timestamp 18001
transform 1 0 67988 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_151_691
timestamp 18001
transform 1 0 68448 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_151_698
timestamp 18001
transform 1 0 69092 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_151_701
timestamp 18001
transform 1 0 69368 0 -1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_707
timestamp 18001
transform 1 0 69920 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_151_712
timestamp 18001
transform 1 0 70380 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_151_720
timestamp 18001
transform 1 0 71116 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_151_726
timestamp 18001
transform 1 0 71668 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_151_729
timestamp 18001
transform 1 0 71944 0 -1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_735
timestamp 18001
transform 1 0 72496 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_151_740
timestamp 18001
transform 1 0 72956 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_151_747
timestamp 18001
transform 1 0 73600 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_151_755
timestamp 18001
transform 1 0 74336 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_151_761
timestamp 18001
transform 1 0 74888 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_151_769
timestamp 18001
transform 1 0 75624 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_151_775
timestamp 18001
transform 1 0 76176 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_151_782
timestamp 18001
transform 1 0 76820 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_151_785
timestamp 18001
transform 1 0 77096 0 -1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_791
timestamp 18001
transform 1 0 77648 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_151_796
timestamp 18001
transform 1 0 78108 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_151_804
timestamp 18001
transform 1 0 78844 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_151_810
timestamp 18001
transform 1 0 79396 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_151_813
timestamp 18001
transform 1 0 79672 0 -1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_819
timestamp 18001
transform 1 0 80224 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_151_824
timestamp 18001
transform 1 0 80684 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_151_831
timestamp 18001
transform 1 0 81328 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_151_839
timestamp 18001
transform 1 0 82064 0 -1 87584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_151_845
timestamp 1636986456
transform 1 0 82616 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_151_857
timestamp 18001
transform 1 0 83720 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_151_865
timestamp 18001
transform 1 0 84456 0 -1 87584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_151_869
timestamp 1636986456
transform 1 0 84824 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_881
timestamp 1636986456
transform 1 0 85928 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_151_893
timestamp 18001
transform 1 0 87032 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_151_897
timestamp 18001
transform 1 0 87400 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_151_905
timestamp 18001
transform 1 0 88136 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  fpga_232
timestamp 18001
transform -1 0 46460 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_233
timestamp 18001
transform -1 0 50324 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_234
timestamp 18001
transform -1 0 47748 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_235
timestamp 18001
transform -1 0 41952 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_236
timestamp 18001
transform -1 0 49036 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_237
timestamp 18001
transform 1 0 88044 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_238
timestamp 18001
transform 1 0 88044 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_239
timestamp 18001
transform -1 0 43240 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_240
timestamp 18001
transform -1 0 45172 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_241
timestamp 18001
transform -1 0 49680 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_242
timestamp 18001
transform 1 0 88044 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_243
timestamp 18001
transform 1 0 88044 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_244
timestamp 18001
transform -1 0 45816 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_245
timestamp 18001
transform 1 0 88044 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_246
timestamp 18001
transform -1 0 47104 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_247
timestamp 18001
transform -1 0 48392 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 18001
transform 1 0 5152 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  input2
timestamp 18001
transform -1 0 37536 0 -1 87584
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 18001
transform -1 0 88320 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 18001
transform 1 0 88044 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 18001
transform 1 0 88044 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 18001
transform 1 0 88044 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 18001
transform 1 0 88044 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 18001
transform -1 0 88320 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 18001
transform 1 0 88044 0 -1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 18001
transform -1 0 88320 0 1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 18001
transform 1 0 88044 0 1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 18001
transform 1 0 88044 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 18001
transform 1 0 88044 0 1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 18001
transform -1 0 88320 0 1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 18001
transform -1 0 88320 0 -1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input16
timestamp 18001
transform -1 0 88320 0 1 74528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input17
timestamp 18001
transform -1 0 88320 0 1 75616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input18
timestamp 18001
transform -1 0 87860 0 1 76704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 18001
transform 1 0 88044 0 1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 18001
transform 1 0 88044 0 -1 78880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 18001
transform 1 0 88044 0 1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 18001
transform 1 0 88044 0 1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input23
timestamp 18001
transform -1 0 88320 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 18001
transform 1 0 88044 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input25
timestamp 18001
transform -1 0 88320 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input26
timestamp 18001
transform -1 0 88320 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input27
timestamp 18001
transform -1 0 88320 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input28
timestamp 18001
transform -1 0 88320 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input29
timestamp 18001
transform -1 0 88320 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input30
timestamp 18001
transform -1 0 88320 0 -1 40800
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input31
timestamp 18001
transform 1 0 15272 0 -1 87584
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 18001
transform 1 0 26220 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input33
timestamp 18001
transform 1 0 26864 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 18001
transform 1 0 28152 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input35
timestamp 18001
transform -1 0 29716 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input36
timestamp 18001
transform 1 0 52624 0 -1 87584
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input37
timestamp 18001
transform -1 0 53820 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input38
timestamp 18001
transform -1 0 54832 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input39
timestamp 18001
transform -1 0 56120 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input40
timestamp 18001
transform -1 0 16468 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input41
timestamp 18001
transform -1 0 57408 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input42
timestamp 18001
transform 1 0 57776 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input43
timestamp 18001
transform -1 0 59340 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input44
timestamp 18001
transform -1 0 60628 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 18001
transform -1 0 61272 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input46
timestamp 18001
transform -1 0 62560 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 18001
transform 1 0 63572 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input48
timestamp 18001
transform -1 0 65136 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 18001
transform -1 0 65780 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input50
timestamp 18001
transform -1 0 67068 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input51
timestamp 18001
transform -1 0 17480 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input52
timestamp 18001
transform -1 0 18768 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input53
timestamp 18001
transform 1 0 19136 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input54
timestamp 18001
transform -1 0 20700 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input55
timestamp 18001
transform -1 0 21988 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input56
timestamp 18001
transform -1 0 23276 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 18001
transform -1 0 23920 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input58
timestamp 18001
transform -1 0 25208 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 18001
transform 1 0 30728 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 18001
transform 1 0 41676 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 18001
transform -1 0 42596 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 18001
transform 1 0 43608 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 18001
transform 1 0 44896 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 18001
transform 1 0 68080 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input65
timestamp 18001
transform 1 0 68724 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input66
timestamp 18001
transform -1 0 70288 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input67
timestamp 18001
transform -1 0 71576 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input68
timestamp 18001
transform 1 0 31372 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input69
timestamp 18001
transform -1 0 72864 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 18001
transform -1 0 73508 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input71
timestamp 18001
transform -1 0 74796 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input72
timestamp 18001
transform -1 0 76084 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input73
timestamp 18001
transform 1 0 76452 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input74
timestamp 18001
transform -1 0 78016 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input75
timestamp 18001
transform 1 0 79028 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input76
timestamp 18001
transform 1 0 80316 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input77
timestamp 18001
transform -1 0 81236 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input78
timestamp 18001
transform 1 0 88044 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input79
timestamp 18001
transform -1 0 32936 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input80
timestamp 18001
transform -1 0 34224 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input81
timestamp 18001
transform 1 0 34592 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input82
timestamp 18001
transform 1 0 35880 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input83
timestamp 18001
transform -1 0 37444 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input84
timestamp 18001
transform -1 0 38732 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input85
timestamp 18001
transform 1 0 39100 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input86
timestamp 18001
transform -1 0 40664 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input87
timestamp 18001
transform -1 0 5428 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input88
timestamp 18001
transform -1 0 5428 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input89
timestamp 18001
transform -1 0 5428 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input90
timestamp 18001
transform -1 0 5428 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input91
timestamp 18001
transform -1 0 5428 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input92
timestamp 18001
transform -1 0 5428 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input93
timestamp 18001
transform -1 0 5428 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input94
timestamp 18001
transform -1 0 5428 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input95
timestamp 18001
transform -1 0 5428 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input96
timestamp 18001
transform -1 0 5428 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input97
timestamp 18001
transform -1 0 5428 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input98
timestamp 18001
transform -1 0 5428 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input99
timestamp 18001
transform 1 0 5152 0 1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input100
timestamp 18001
transform -1 0 5428 0 1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input101
timestamp 18001
transform 1 0 5152 0 1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input102
timestamp 18001
transform 1 0 5152 0 1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input103
timestamp 18001
transform -1 0 5428 0 -1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input104
timestamp 18001
transform -1 0 5428 0 1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input105
timestamp 18001
transform -1 0 5428 0 1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input106
timestamp 18001
transform -1 0 5428 0 1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input107
timestamp 18001
transform -1 0 5428 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input108
timestamp 18001
transform -1 0 5428 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input109
timestamp 18001
transform -1 0 5428 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input110
timestamp 18001
transform -1 0 5428 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input111
timestamp 18001
transform 1 0 5152 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input112
timestamp 18001
transform -1 0 5428 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input113
timestamp 18001
transform 1 0 5152 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input114
timestamp 18001
transform 1 0 5152 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input115
timestamp 18001
transform -1 0 87860 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input116
timestamp 18001
transform -1 0 88320 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input117
timestamp 18001
transform -1 0 87860 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  input118
timestamp 18001
transform 1 0 38456 0 -1 87584
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_2  output119
timestamp 18001
transform 1 0 87952 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output120
timestamp 18001
transform 1 0 87952 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output121
timestamp 18001
transform 1 0 87952 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output122
timestamp 18001
transform 1 0 87952 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp 18001
transform 1 0 87952 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output124
timestamp 18001
transform 1 0 87952 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output125
timestamp 18001
transform 1 0 87952 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output126
timestamp 18001
transform 1 0 87952 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output127
timestamp 18001
transform 1 0 87952 0 1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output128
timestamp 18001
transform 1 0 87952 0 1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output129
timestamp 18001
transform 1 0 87952 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output130
timestamp 18001
transform 1 0 87952 0 1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output131
timestamp 18001
transform 1 0 87952 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output132
timestamp 18001
transform 1 0 87952 0 1 58208
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output133
timestamp 18001
transform 1 0 87952 0 1 59296
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output134
timestamp 18001
transform 1 0 87952 0 1 60384
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output135
timestamp 18001
transform 1 0 87952 0 1 61472
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output136
timestamp 18001
transform 1 0 87952 0 -1 62560
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output137
timestamp 18001
transform 1 0 87952 0 1 63648
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output138
timestamp 18001
transform 1 0 87952 0 1 64736
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp 18001
transform 1 0 87952 0 1 65824
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output140
timestamp 18001
transform 1 0 87952 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output141
timestamp 18001
transform 1 0 87952 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output142
timestamp 18001
transform 1 0 87952 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output143
timestamp 18001
transform 1 0 87952 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output144
timestamp 18001
transform 1 0 87952 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output145
timestamp 18001
transform 1 0 87952 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output146
timestamp 18001
transform 1 0 87952 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output147
timestamp 18001
transform 1 0 87952 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output148
timestamp 18001
transform 1 0 30728 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output149
timestamp 18001
transform -1 0 41400 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output150
timestamp 18001
transform -1 0 42688 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output151
timestamp 18001
transform 1 0 43608 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output152
timestamp 18001
transform -1 0 44620 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output153
timestamp 18001
transform 1 0 68080 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output154
timestamp 18001
transform -1 0 69092 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output155
timestamp 18001
transform 1 0 70012 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output156
timestamp 18001
transform 1 0 71300 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output157
timestamp 18001
transform -1 0 31740 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output158
timestamp 18001
transform 1 0 72588 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output159
timestamp 18001
transform -1 0 73600 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output160
timestamp 18001
transform 1 0 74520 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output161
timestamp 18001
transform 1 0 75808 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output162
timestamp 18001
transform -1 0 76820 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output163
timestamp 18001
transform 1 0 77740 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output164
timestamp 18001
transform 1 0 79028 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output165
timestamp 18001
transform 1 0 80316 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output166
timestamp 18001
transform -1 0 81328 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output167
timestamp 18001
transform 1 0 82248 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output168
timestamp 18001
transform 1 0 32660 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output169
timestamp 18001
transform 1 0 33948 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output170
timestamp 18001
transform -1 0 34960 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output171
timestamp 18001
transform 1 0 35880 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output172
timestamp 18001
transform 1 0 37536 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output173
timestamp 18001
transform 1 0 37996 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output174
timestamp 18001
transform 1 0 39468 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output175
timestamp 18001
transform 1 0 40388 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output176
timestamp 18001
transform 1 0 15272 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output177
timestamp 18001
transform 1 0 26220 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output178
timestamp 18001
transform -1 0 27232 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output179
timestamp 18001
transform 1 0 28152 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output180
timestamp 18001
transform 1 0 29440 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output181
timestamp 18001
transform 1 0 52624 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output182
timestamp 18001
transform -1 0 53636 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output183
timestamp 18001
transform 1 0 54556 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output184
timestamp 18001
transform 1 0 55844 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output185
timestamp 18001
transform -1 0 16284 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output186
timestamp 18001
transform 1 0 57132 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output187
timestamp 18001
transform -1 0 58144 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output188
timestamp 18001
transform 1 0 59064 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output189
timestamp 18001
transform 1 0 60352 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output190
timestamp 18001
transform -1 0 61364 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output191
timestamp 18001
transform 1 0 62284 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output192
timestamp 18001
transform 1 0 63572 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output193
timestamp 18001
transform 1 0 64860 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output194
timestamp 18001
transform -1 0 65872 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output195
timestamp 18001
transform 1 0 66792 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output196
timestamp 18001
transform 1 0 17204 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output197
timestamp 18001
transform 1 0 18492 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output198
timestamp 18001
transform -1 0 19504 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output199
timestamp 18001
transform 1 0 20424 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output200
timestamp 18001
transform 1 0 21712 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output201
timestamp 18001
transform 1 0 23000 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output202
timestamp 18001
transform -1 0 24012 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output203
timestamp 18001
transform 1 0 24932 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output204
timestamp 18001
transform -1 0 5520 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output205
timestamp 18001
transform -1 0 5520 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output206
timestamp 18001
transform -1 0 5520 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output207
timestamp 18001
transform -1 0 5520 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output208
timestamp 18001
transform -1 0 5520 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output209
timestamp 18001
transform -1 0 5520 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output210
timestamp 18001
transform -1 0 5520 0 -1 68000
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output211
timestamp 18001
transform -1 0 5520 0 1 69088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output212
timestamp 18001
transform -1 0 5520 0 1 70176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output213
timestamp 18001
transform -1 0 5520 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output214
timestamp 18001
transform -1 0 5520 0 1 71264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output215
timestamp 18001
transform -1 0 5520 0 1 72352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output216
timestamp 18001
transform -1 0 5520 0 -1 73440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output217
timestamp 18001
transform -1 0 5520 0 1 74528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output218
timestamp 18001
transform -1 0 5520 0 1 75616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output219
timestamp 18001
transform -1 0 5520 0 1 76704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output220
timestamp 18001
transform -1 0 5520 0 1 77792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output221
timestamp 18001
transform -1 0 5520 0 -1 78880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output222
timestamp 18001
transform -1 0 5520 0 1 79968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output223
timestamp 18001
transform -1 0 5520 0 1 81056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output224
timestamp 18001
transform -1 0 5520 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output225
timestamp 18001
transform -1 0 5520 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output226
timestamp 18001
transform -1 0 5520 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output227
timestamp 18001
transform -1 0 5520 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output228
timestamp 18001
transform -1 0 5520 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output229
timestamp 18001
transform -1 0 5520 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output230
timestamp 18001
transform -1 0 5520 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output231
timestamp 18001
transform -1 0 5520 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_152
timestamp 18001
transform 1 0 4876 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 18001
transform -1 0 88596 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_153
timestamp 18001
transform 1 0 4876 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 18001
transform -1 0 88596 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_154
timestamp 18001
transform 1 0 4876 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 18001
transform -1 0 88596 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_155
timestamp 18001
transform 1 0 4876 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 18001
transform -1 0 88596 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_156
timestamp 18001
transform 1 0 4876 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 18001
transform -1 0 88596 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_1_Left_303
timestamp 18001
transform 1 0 4876 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_1_Right_585
timestamp 18001
transform -1 0 7912 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_3_Left_304
timestamp 18001
transform 1 0 85284 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_3_Right_11
timestamp 18001
transform -1 0 88596 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_1_Left_157
timestamp 18001
transform 1 0 4876 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_1_Right_445
timestamp 18001
transform -1 0 7912 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_3_Left_305
timestamp 18001
transform 1 0 85284 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_3_Right_12
timestamp 18001
transform -1 0 88596 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_1_Left_158
timestamp 18001
transform 1 0 4876 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_1_Right_446
timestamp 18001
transform -1 0 7912 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_3_Left_306
timestamp 18001
transform 1 0 85284 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_3_Right_13
timestamp 18001
transform -1 0 88596 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_1_Left_159
timestamp 18001
transform 1 0 4876 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_1_Right_447
timestamp 18001
transform -1 0 7912 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_3_Left_307
timestamp 18001
transform 1 0 85284 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_3_Right_14
timestamp 18001
transform -1 0 88596 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_1_Left_160
timestamp 18001
transform 1 0 4876 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_1_Right_448
timestamp 18001
transform -1 0 7912 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_3_Left_308
timestamp 18001
transform 1 0 85284 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_3_Right_15
timestamp 18001
transform -1 0 88596 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_1_Left_161
timestamp 18001
transform 1 0 4876 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_1_Right_449
timestamp 18001
transform -1 0 7912 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_3_Left_309
timestamp 18001
transform 1 0 85284 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_3_Right_16
timestamp 18001
transform -1 0 88596 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_1_Left_162
timestamp 18001
transform 1 0 4876 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_1_Right_450
timestamp 18001
transform -1 0 7912 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_3_Left_310
timestamp 18001
transform 1 0 85284 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_3_Right_17
timestamp 18001
transform -1 0 88596 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_1_Left_163
timestamp 18001
transform 1 0 4876 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_1_Right_451
timestamp 18001
transform -1 0 7912 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_3_Left_311
timestamp 18001
transform 1 0 85284 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_3_Right_18
timestamp 18001
transform -1 0 88596 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_1_Left_164
timestamp 18001
transform 1 0 4876 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_1_Right_452
timestamp 18001
transform -1 0 7912 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_3_Left_312
timestamp 18001
transform 1 0 85284 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_3_Right_19
timestamp 18001
transform -1 0 88596 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_1_Left_165
timestamp 18001
transform 1 0 4876 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_1_Right_453
timestamp 18001
transform -1 0 7912 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_3_Left_313
timestamp 18001
transform 1 0 85284 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_3_Right_20
timestamp 18001
transform -1 0 88596 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_1_Left_166
timestamp 18001
transform 1 0 4876 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_1_Right_454
timestamp 18001
transform -1 0 7912 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_3_Left_314
timestamp 18001
transform 1 0 85284 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_3_Right_21
timestamp 18001
transform -1 0 88596 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_1_Left_167
timestamp 18001
transform 1 0 4876 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_1_Right_455
timestamp 18001
transform -1 0 7912 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_3_Left_315
timestamp 18001
transform 1 0 85284 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_3_Right_22
timestamp 18001
transform -1 0 88596 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_1_Left_168
timestamp 18001
transform 1 0 4876 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_1_Right_456
timestamp 18001
transform -1 0 7912 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_3_Left_316
timestamp 18001
transform 1 0 85284 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_3_Right_23
timestamp 18001
transform -1 0 88596 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_1_Left_169
timestamp 18001
transform 1 0 4876 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_1_Right_457
timestamp 18001
transform -1 0 7912 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_3_Left_317
timestamp 18001
transform 1 0 85284 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_3_Right_24
timestamp 18001
transform -1 0 88596 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_1_Left_170
timestamp 18001
transform 1 0 4876 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_1_Right_458
timestamp 18001
transform -1 0 7912 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_3_Left_318
timestamp 18001
transform 1 0 85284 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_3_Right_25
timestamp 18001
transform -1 0 88596 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_1_Left_171
timestamp 18001
transform 1 0 4876 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_1_Right_459
timestamp 18001
transform -1 0 7912 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_3_Left_319
timestamp 18001
transform 1 0 85284 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_3_Right_26
timestamp 18001
transform -1 0 88596 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_1_Left_172
timestamp 18001
transform 1 0 4876 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_1_Right_460
timestamp 18001
transform -1 0 7912 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_3_Left_320
timestamp 18001
transform 1 0 85284 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_3_Right_27
timestamp 18001
transform -1 0 88596 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_1_Left_173
timestamp 18001
transform 1 0 4876 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_1_Right_461
timestamp 18001
transform -1 0 7912 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_3_Left_321
timestamp 18001
transform 1 0 85284 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_3_Right_28
timestamp 18001
transform -1 0 88596 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_1_Left_174
timestamp 18001
transform 1 0 4876 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_1_Right_462
timestamp 18001
transform -1 0 7912 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_3_Left_322
timestamp 18001
transform 1 0 85284 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_3_Right_29
timestamp 18001
transform -1 0 88596 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_1_Left_175
timestamp 18001
transform 1 0 4876 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_1_Right_463
timestamp 18001
transform -1 0 7912 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_3_Left_323
timestamp 18001
transform 1 0 85284 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_3_Right_30
timestamp 18001
transform -1 0 88596 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_1_Left_176
timestamp 18001
transform 1 0 4876 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_1_Right_464
timestamp 18001
transform -1 0 7912 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_3_Left_324
timestamp 18001
transform 1 0 85284 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_3_Right_31
timestamp 18001
transform -1 0 88596 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_1_Left_177
timestamp 18001
transform 1 0 4876 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_1_Right_465
timestamp 18001
transform -1 0 7912 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_3_Left_325
timestamp 18001
transform 1 0 85284 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_3_Right_32
timestamp 18001
transform -1 0 88596 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_1_Left_178
timestamp 18001
transform 1 0 4876 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_1_Right_466
timestamp 18001
transform -1 0 7912 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_3_Left_326
timestamp 18001
transform 1 0 85284 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_3_Right_33
timestamp 18001
transform -1 0 88596 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_1_Left_179
timestamp 18001
transform 1 0 4876 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_1_Right_467
timestamp 18001
transform -1 0 7912 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_3_Left_327
timestamp 18001
transform 1 0 85284 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_3_Right_34
timestamp 18001
transform -1 0 88596 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_1_Left_180
timestamp 18001
transform 1 0 4876 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_1_Right_468
timestamp 18001
transform -1 0 7912 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_3_Left_328
timestamp 18001
transform 1 0 85284 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_3_Right_35
timestamp 18001
transform -1 0 88596 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_1_Left_181
timestamp 18001
transform 1 0 4876 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_1_Right_469
timestamp 18001
transform -1 0 7912 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_3_Left_329
timestamp 18001
transform 1 0 85284 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_3_Right_36
timestamp 18001
transform -1 0 88596 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_1_Left_182
timestamp 18001
transform 1 0 4876 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_1_Right_470
timestamp 18001
transform -1 0 7912 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_3_Left_330
timestamp 18001
transform 1 0 85284 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_3_Right_37
timestamp 18001
transform -1 0 88596 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_1_Left_183
timestamp 18001
transform 1 0 4876 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_1_Right_471
timestamp 18001
transform -1 0 7912 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_3_Left_331
timestamp 18001
transform 1 0 85284 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_3_Right_38
timestamp 18001
transform -1 0 88596 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_1_Left_184
timestamp 18001
transform 1 0 4876 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_1_Right_472
timestamp 18001
transform -1 0 7912 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_3_Left_332
timestamp 18001
transform 1 0 85284 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_3_Right_39
timestamp 18001
transform -1 0 88596 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_1_Left_185
timestamp 18001
transform 1 0 4876 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_1_Right_473
timestamp 18001
transform -1 0 7912 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_3_Left_333
timestamp 18001
transform 1 0 85284 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_3_Right_40
timestamp 18001
transform -1 0 88596 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_1_Left_186
timestamp 18001
transform 1 0 4876 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_1_Right_474
timestamp 18001
transform -1 0 7912 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_3_Left_334
timestamp 18001
transform 1 0 85284 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_3_Right_41
timestamp 18001
transform -1 0 88596 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_1_Left_187
timestamp 18001
transform 1 0 4876 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_1_Right_475
timestamp 18001
transform -1 0 7912 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_3_Left_335
timestamp 18001
transform 1 0 85284 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_3_Right_42
timestamp 18001
transform -1 0 88596 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_1_Left_188
timestamp 18001
transform 1 0 4876 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_1_Right_476
timestamp 18001
transform -1 0 7912 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_3_Left_336
timestamp 18001
transform 1 0 85284 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_3_Right_43
timestamp 18001
transform -1 0 88596 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_1_Left_189
timestamp 18001
transform 1 0 4876 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_1_Right_477
timestamp 18001
transform -1 0 7912 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_3_Left_337
timestamp 18001
transform 1 0 85284 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_3_Right_44
timestamp 18001
transform -1 0 88596 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_1_Left_190
timestamp 18001
transform 1 0 4876 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_1_Right_478
timestamp 18001
transform -1 0 7912 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_3_Left_338
timestamp 18001
transform 1 0 85284 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_3_Right_45
timestamp 18001
transform -1 0 88596 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_1_Left_191
timestamp 18001
transform 1 0 4876 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_1_Right_479
timestamp 18001
transform -1 0 7912 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_3_Left_339
timestamp 18001
transform 1 0 85284 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_3_Right_46
timestamp 18001
transform -1 0 88596 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_1_Left_192
timestamp 18001
transform 1 0 4876 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_1_Right_480
timestamp 18001
transform -1 0 7912 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_3_Left_340
timestamp 18001
transform 1 0 85284 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_3_Right_47
timestamp 18001
transform -1 0 88596 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_1_Left_193
timestamp 18001
transform 1 0 4876 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_1_Right_481
timestamp 18001
transform -1 0 7912 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_3_Left_341
timestamp 18001
transform 1 0 85284 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_3_Right_48
timestamp 18001
transform -1 0 88596 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_1_Left_194
timestamp 18001
transform 1 0 4876 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_1_Right_482
timestamp 18001
transform -1 0 7912 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_3_Left_342
timestamp 18001
transform 1 0 85284 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_3_Right_49
timestamp 18001
transform -1 0 88596 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_1_Left_195
timestamp 18001
transform 1 0 4876 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_1_Right_483
timestamp 18001
transform -1 0 7912 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_3_Left_343
timestamp 18001
transform 1 0 85284 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_3_Right_50
timestamp 18001
transform -1 0 88596 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_1_Left_196
timestamp 18001
transform 1 0 4876 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_1_Right_484
timestamp 18001
transform -1 0 7912 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_3_Left_344
timestamp 18001
transform 1 0 85284 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_3_Right_51
timestamp 18001
transform -1 0 88596 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_1_Left_197
timestamp 18001
transform 1 0 4876 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_1_Right_485
timestamp 18001
transform -1 0 7912 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_3_Left_345
timestamp 18001
transform 1 0 85284 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_3_Right_52
timestamp 18001
transform -1 0 88596 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_1_Left_198
timestamp 18001
transform 1 0 4876 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_1_Right_486
timestamp 18001
transform -1 0 7912 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_3_Left_346
timestamp 18001
transform 1 0 85284 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_3_Right_53
timestamp 18001
transform -1 0 88596 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_1_Left_199
timestamp 18001
transform 1 0 4876 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_1_Right_487
timestamp 18001
transform -1 0 7912 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_3_Left_347
timestamp 18001
transform 1 0 85284 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_3_Right_54
timestamp 18001
transform -1 0 88596 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_1_Left_200
timestamp 18001
transform 1 0 4876 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_1_Right_488
timestamp 18001
transform -1 0 7912 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_3_Left_348
timestamp 18001
transform 1 0 85284 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_3_Right_55
timestamp 18001
transform -1 0 88596 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_1_Left_201
timestamp 18001
transform 1 0 4876 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_1_Right_489
timestamp 18001
transform -1 0 7912 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_3_Left_349
timestamp 18001
transform 1 0 85284 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_3_Right_56
timestamp 18001
transform -1 0 88596 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_1_Left_202
timestamp 18001
transform 1 0 4876 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_1_Right_490
timestamp 18001
transform -1 0 7912 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_3_Left_350
timestamp 18001
transform 1 0 85284 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_3_Right_57
timestamp 18001
transform -1 0 88596 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_1_Left_203
timestamp 18001
transform 1 0 4876 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_1_Right_491
timestamp 18001
transform -1 0 7912 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_3_Left_351
timestamp 18001
transform 1 0 85284 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_3_Right_58
timestamp 18001
transform -1 0 88596 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_1_Left_204
timestamp 18001
transform 1 0 4876 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_1_Right_492
timestamp 18001
transform -1 0 7912 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_3_Left_352
timestamp 18001
transform 1 0 85284 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_3_Right_59
timestamp 18001
transform -1 0 88596 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_1_Left_205
timestamp 18001
transform 1 0 4876 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_1_Right_493
timestamp 18001
transform -1 0 7912 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_3_Left_353
timestamp 18001
transform 1 0 85284 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_3_Right_60
timestamp 18001
transform -1 0 88596 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_1_Left_206
timestamp 18001
transform 1 0 4876 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_1_Right_494
timestamp 18001
transform -1 0 7912 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_3_Left_354
timestamp 18001
transform 1 0 85284 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_3_Right_61
timestamp 18001
transform -1 0 88596 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_1_Left_207
timestamp 18001
transform 1 0 4876 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_1_Right_495
timestamp 18001
transform -1 0 7912 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_3_Left_355
timestamp 18001
transform 1 0 85284 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_3_Right_62
timestamp 18001
transform -1 0 88596 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_1_Left_208
timestamp 18001
transform 1 0 4876 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_1_Right_496
timestamp 18001
transform -1 0 7912 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_3_Left_356
timestamp 18001
transform 1 0 85284 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_3_Right_63
timestamp 18001
transform -1 0 88596 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_1_Left_209
timestamp 18001
transform 1 0 4876 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_1_Right_497
timestamp 18001
transform -1 0 7912 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_3_Left_357
timestamp 18001
transform 1 0 85284 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_3_Right_64
timestamp 18001
transform -1 0 88596 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_1_Left_210
timestamp 18001
transform 1 0 4876 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_1_Right_498
timestamp 18001
transform -1 0 7912 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_3_Left_358
timestamp 18001
transform 1 0 85284 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_3_Right_65
timestamp 18001
transform -1 0 88596 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_1_Left_211
timestamp 18001
transform 1 0 4876 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_1_Right_499
timestamp 18001
transform -1 0 7912 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_3_Left_359
timestamp 18001
transform 1 0 85284 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_3_Right_66
timestamp 18001
transform -1 0 88596 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_1_Left_212
timestamp 18001
transform 1 0 4876 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_1_Right_500
timestamp 18001
transform -1 0 7912 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_3_Left_360
timestamp 18001
transform 1 0 85284 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_3_Right_67
timestamp 18001
transform -1 0 88596 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_1_Left_213
timestamp 18001
transform 1 0 4876 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_1_Right_501
timestamp 18001
transform -1 0 7912 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_3_Left_361
timestamp 18001
transform 1 0 85284 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_3_Right_68
timestamp 18001
transform -1 0 88596 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_1_Left_214
timestamp 18001
transform 1 0 4876 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_1_Right_502
timestamp 18001
transform -1 0 7912 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_3_Left_362
timestamp 18001
transform 1 0 85284 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_3_Right_69
timestamp 18001
transform -1 0 88596 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_1_Left_215
timestamp 18001
transform 1 0 4876 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_1_Right_503
timestamp 18001
transform -1 0 7912 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_3_Left_363
timestamp 18001
transform 1 0 85284 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_3_Right_70
timestamp 18001
transform -1 0 88596 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_1_Left_216
timestamp 18001
transform 1 0 4876 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_1_Right_504
timestamp 18001
transform -1 0 7912 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_3_Left_364
timestamp 18001
transform 1 0 85284 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_3_Right_71
timestamp 18001
transform -1 0 88596 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_1_Left_217
timestamp 18001
transform 1 0 4876 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_1_Right_505
timestamp 18001
transform -1 0 7912 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_3_Left_365
timestamp 18001
transform 1 0 85284 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_3_Right_72
timestamp 18001
transform -1 0 88596 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_1_Left_218
timestamp 18001
transform 1 0 4876 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_1_Right_506
timestamp 18001
transform -1 0 7912 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_3_Left_366
timestamp 18001
transform 1 0 85284 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_3_Right_73
timestamp 18001
transform -1 0 88596 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_1_Left_219
timestamp 18001
transform 1 0 4876 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_1_Right_507
timestamp 18001
transform -1 0 7912 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_3_Left_367
timestamp 18001
transform 1 0 85284 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_3_Right_74
timestamp 18001
transform -1 0 88596 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_1_Left_220
timestamp 18001
transform 1 0 4876 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_1_Right_508
timestamp 18001
transform -1 0 7912 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_3_Left_368
timestamp 18001
transform 1 0 85284 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_3_Right_75
timestamp 18001
transform -1 0 88596 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_1_Left_221
timestamp 18001
transform 1 0 4876 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_1_Right_509
timestamp 18001
transform -1 0 7912 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_3_Left_369
timestamp 18001
transform 1 0 85284 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_3_Right_76
timestamp 18001
transform -1 0 88596 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_1_Left_222
timestamp 18001
transform 1 0 4876 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_1_Right_510
timestamp 18001
transform -1 0 7912 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_3_Left_370
timestamp 18001
transform 1 0 85284 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_3_Right_77
timestamp 18001
transform -1 0 88596 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_1_Left_223
timestamp 18001
transform 1 0 4876 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_1_Right_511
timestamp 18001
transform -1 0 7912 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_5_Left_371
timestamp 18001
transform 1 0 85284 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_5_Right_78
timestamp 18001
transform -1 0 88596 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_1_Left_224
timestamp 18001
transform 1 0 4876 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_1_Right_512
timestamp 18001
transform -1 0 7912 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_5_Left_372
timestamp 18001
transform 1 0 85284 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_5_Right_79
timestamp 18001
transform -1 0 88596 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_1_Left_225
timestamp 18001
transform 1 0 4876 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_1_Right_513
timestamp 18001
transform -1 0 7912 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_5_Left_373
timestamp 18001
transform 1 0 85284 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_5_Right_80
timestamp 18001
transform -1 0 88596 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_1_Left_226
timestamp 18001
transform 1 0 4876 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_1_Right_514
timestamp 18001
transform -1 0 7912 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_5_Left_374
timestamp 18001
transform 1 0 85284 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_5_Right_81
timestamp 18001
transform -1 0 88596 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_1_Left_227
timestamp 18001
transform 1 0 4876 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_1_Right_515
timestamp 18001
transform -1 0 7912 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_5_Left_375
timestamp 18001
transform 1 0 85284 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_5_Right_82
timestamp 18001
transform -1 0 88596 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_1_Left_228
timestamp 18001
transform 1 0 4876 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_1_Right_516
timestamp 18001
transform -1 0 7912 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_5_Left_376
timestamp 18001
transform 1 0 85284 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_5_Right_83
timestamp 18001
transform -1 0 88596 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_1_Left_229
timestamp 18001
transform 1 0 4876 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_1_Right_517
timestamp 18001
transform -1 0 7912 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_5_Left_377
timestamp 18001
transform 1 0 85284 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_5_Right_84
timestamp 18001
transform -1 0 88596 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_1_Left_230
timestamp 18001
transform 1 0 4876 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_1_Right_518
timestamp 18001
transform -1 0 7912 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_3_Left_378
timestamp 18001
transform 1 0 85284 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_3_Right_85
timestamp 18001
transform -1 0 88596 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_1_Left_231
timestamp 18001
transform 1 0 4876 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_1_Right_519
timestamp 18001
transform -1 0 7912 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_3_Left_379
timestamp 18001
transform 1 0 85284 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_3_Right_86
timestamp 18001
transform -1 0 88596 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_1_Left_232
timestamp 18001
transform 1 0 4876 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_1_Right_520
timestamp 18001
transform -1 0 7912 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_3_Left_380
timestamp 18001
transform 1 0 85284 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_3_Right_87
timestamp 18001
transform -1 0 88596 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_1_Left_233
timestamp 18001
transform 1 0 4876 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_1_Right_521
timestamp 18001
transform -1 0 7912 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_3_Left_381
timestamp 18001
transform 1 0 85284 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_3_Right_88
timestamp 18001
transform -1 0 88596 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_1_Left_234
timestamp 18001
transform 1 0 4876 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_1_Right_522
timestamp 18001
transform -1 0 7912 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_3_Left_382
timestamp 18001
transform 1 0 85284 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_3_Right_89
timestamp 18001
transform -1 0 88596 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_1_Left_235
timestamp 18001
transform 1 0 4876 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_1_Right_523
timestamp 18001
transform -1 0 7912 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_3_Left_383
timestamp 18001
transform 1 0 85284 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_3_Right_90
timestamp 18001
transform -1 0 88596 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_1_Left_236
timestamp 18001
transform 1 0 4876 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_1_Right_524
timestamp 18001
transform -1 0 7912 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_3_Left_384
timestamp 18001
transform 1 0 85284 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_3_Right_91
timestamp 18001
transform -1 0 88596 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_1_Left_237
timestamp 18001
transform 1 0 4876 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_1_Right_525
timestamp 18001
transform -1 0 7912 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_3_Left_385
timestamp 18001
transform 1 0 85284 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_3_Right_92
timestamp 18001
transform -1 0 88596 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_1_Left_238
timestamp 18001
transform 1 0 4876 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_1_Right_526
timestamp 18001
transform -1 0 7912 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_3_Left_386
timestamp 18001
transform 1 0 85284 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_3_Right_93
timestamp 18001
transform -1 0 88596 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_1_Left_239
timestamp 18001
transform 1 0 4876 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_1_Right_527
timestamp 18001
transform -1 0 7912 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_3_Left_387
timestamp 18001
transform 1 0 85284 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_3_Right_94
timestamp 18001
transform -1 0 88596 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_1_Left_240
timestamp 18001
transform 1 0 4876 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_1_Right_528
timestamp 18001
transform -1 0 7912 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_3_Left_388
timestamp 18001
transform 1 0 85284 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_3_Right_95
timestamp 18001
transform -1 0 88596 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_1_Left_241
timestamp 18001
transform 1 0 4876 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_1_Right_529
timestamp 18001
transform -1 0 7912 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_3_Left_389
timestamp 18001
transform 1 0 85284 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_3_Right_96
timestamp 18001
transform -1 0 88596 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_1_Left_242
timestamp 18001
transform 1 0 4876 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_1_Right_530
timestamp 18001
transform -1 0 7912 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_3_Left_390
timestamp 18001
transform 1 0 85284 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_3_Right_97
timestamp 18001
transform -1 0 88596 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_1_Left_243
timestamp 18001
transform 1 0 4876 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_1_Right_531
timestamp 18001
transform -1 0 7912 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_3_Left_391
timestamp 18001
transform 1 0 85284 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_3_Right_98
timestamp 18001
transform -1 0 88596 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_1_Left_244
timestamp 18001
transform 1 0 4876 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_1_Right_532
timestamp 18001
transform -1 0 7912 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_3_Left_392
timestamp 18001
transform 1 0 85284 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_3_Right_99
timestamp 18001
transform -1 0 88596 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_1_Left_245
timestamp 18001
transform 1 0 4876 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_1_Right_533
timestamp 18001
transform -1 0 7912 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_3_Left_393
timestamp 18001
transform 1 0 85284 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_3_Right_100
timestamp 18001
transform -1 0 88596 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_1_Left_246
timestamp 18001
transform 1 0 4876 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_1_Right_534
timestamp 18001
transform -1 0 7912 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_3_Left_394
timestamp 18001
transform 1 0 85284 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_3_Right_101
timestamp 18001
transform -1 0 88596 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_1_Left_247
timestamp 18001
transform 1 0 4876 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_1_Right_535
timestamp 18001
transform -1 0 7912 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_3_Left_395
timestamp 18001
transform 1 0 85284 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_3_Right_102
timestamp 18001
transform -1 0 88596 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_1_Left_248
timestamp 18001
transform 1 0 4876 0 -1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_1_Right_536
timestamp 18001
transform -1 0 7912 0 -1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_3_Left_396
timestamp 18001
transform 1 0 85284 0 -1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_3_Right_103
timestamp 18001
transform -1 0 88596 0 -1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_1_Left_249
timestamp 18001
transform 1 0 4876 0 1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_1_Right_537
timestamp 18001
transform -1 0 7912 0 1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_3_Left_397
timestamp 18001
transform 1 0 85284 0 1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_3_Right_104
timestamp 18001
transform -1 0 88596 0 1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_1_Left_250
timestamp 18001
transform 1 0 4876 0 -1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_1_Right_538
timestamp 18001
transform -1 0 7912 0 -1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_3_Left_398
timestamp 18001
transform 1 0 85284 0 -1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_3_Right_105
timestamp 18001
transform -1 0 88596 0 -1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_1_Left_251
timestamp 18001
transform 1 0 4876 0 1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_1_Right_539
timestamp 18001
transform -1 0 7912 0 1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_3_Left_399
timestamp 18001
transform 1 0 85284 0 1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_3_Right_106
timestamp 18001
transform -1 0 88596 0 1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_1_Left_252
timestamp 18001
transform 1 0 4876 0 -1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_1_Right_540
timestamp 18001
transform -1 0 7912 0 -1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_3_Left_400
timestamp 18001
transform 1 0 85284 0 -1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_3_Right_107
timestamp 18001
transform -1 0 88596 0 -1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_1_Left_253
timestamp 18001
transform 1 0 4876 0 1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_1_Right_541
timestamp 18001
transform -1 0 7912 0 1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_3_Left_401
timestamp 18001
transform 1 0 85284 0 1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_3_Right_108
timestamp 18001
transform -1 0 88596 0 1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_1_Left_254
timestamp 18001
transform 1 0 4876 0 -1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_1_Right_542
timestamp 18001
transform -1 0 7912 0 -1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_3_Left_402
timestamp 18001
transform 1 0 85284 0 -1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_3_Right_109
timestamp 18001
transform -1 0 88596 0 -1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_1_Left_255
timestamp 18001
transform 1 0 4876 0 1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_1_Right_543
timestamp 18001
transform -1 0 7912 0 1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_3_Left_403
timestamp 18001
transform 1 0 85284 0 1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_3_Right_110
timestamp 18001
transform -1 0 88596 0 1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_1_Left_256
timestamp 18001
transform 1 0 4876 0 -1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_1_Right_544
timestamp 18001
transform -1 0 7912 0 -1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_3_Left_404
timestamp 18001
transform 1 0 85284 0 -1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_3_Right_111
timestamp 18001
transform -1 0 88596 0 -1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_1_Left_257
timestamp 18001
transform 1 0 4876 0 1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_1_Right_545
timestamp 18001
transform -1 0 7912 0 1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_3_Left_405
timestamp 18001
transform 1 0 85284 0 1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_3_Right_112
timestamp 18001
transform -1 0 88596 0 1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_1_Left_258
timestamp 18001
transform 1 0 4876 0 -1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_1_Right_546
timestamp 18001
transform -1 0 7912 0 -1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_3_Left_406
timestamp 18001
transform 1 0 85284 0 -1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_3_Right_113
timestamp 18001
transform -1 0 88596 0 -1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_1_Left_259
timestamp 18001
transform 1 0 4876 0 1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_1_Right_547
timestamp 18001
transform -1 0 7912 0 1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_3_Left_407
timestamp 18001
transform 1 0 85284 0 1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_3_Right_114
timestamp 18001
transform -1 0 88596 0 1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_1_Left_260
timestamp 18001
transform 1 0 4876 0 -1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_1_Right_548
timestamp 18001
transform -1 0 7912 0 -1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_3_Left_408
timestamp 18001
transform 1 0 85284 0 -1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_3_Right_115
timestamp 18001
transform -1 0 88596 0 -1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_1_Left_261
timestamp 18001
transform 1 0 4876 0 1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_1_Right_549
timestamp 18001
transform -1 0 7912 0 1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_3_Left_409
timestamp 18001
transform 1 0 85284 0 1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_3_Right_116
timestamp 18001
transform -1 0 88596 0 1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_1_Left_262
timestamp 18001
transform 1 0 4876 0 -1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_1_Right_550
timestamp 18001
transform -1 0 7912 0 -1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_3_Left_410
timestamp 18001
transform 1 0 85284 0 -1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_3_Right_117
timestamp 18001
transform -1 0 88596 0 -1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_1_Left_263
timestamp 18001
transform 1 0 4876 0 1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_1_Right_551
timestamp 18001
transform -1 0 7912 0 1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_3_Left_411
timestamp 18001
transform 1 0 85284 0 1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_3_Right_118
timestamp 18001
transform -1 0 88596 0 1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_1_Left_264
timestamp 18001
transform 1 0 4876 0 -1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_1_Right_552
timestamp 18001
transform -1 0 7912 0 -1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_3_Left_412
timestamp 18001
transform 1 0 85284 0 -1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_3_Right_119
timestamp 18001
transform -1 0 88596 0 -1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_1_Left_265
timestamp 18001
transform 1 0 4876 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_1_Right_553
timestamp 18001
transform -1 0 7912 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_3_Left_413
timestamp 18001
transform 1 0 85284 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_3_Right_120
timestamp 18001
transform -1 0 88596 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_1_Left_266
timestamp 18001
transform 1 0 4876 0 -1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_1_Right_554
timestamp 18001
transform -1 0 7912 0 -1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_3_Left_414
timestamp 18001
transform 1 0 85284 0 -1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_3_Right_121
timestamp 18001
transform -1 0 88596 0 -1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_1_Left_267
timestamp 18001
transform 1 0 4876 0 1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_1_Right_555
timestamp 18001
transform -1 0 7912 0 1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_3_Left_415
timestamp 18001
transform 1 0 85284 0 1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_3_Right_122
timestamp 18001
transform -1 0 88596 0 1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_117_1_Left_268
timestamp 18001
transform 1 0 4876 0 -1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_117_1_Right_556
timestamp 18001
transform -1 0 7912 0 -1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_117_3_Left_416
timestamp 18001
transform 1 0 85284 0 -1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_117_3_Right_123
timestamp 18001
transform -1 0 88596 0 -1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_118_1_Left_269
timestamp 18001
transform 1 0 4876 0 1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_118_1_Right_557
timestamp 18001
transform -1 0 7912 0 1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_118_3_Left_417
timestamp 18001
transform 1 0 85284 0 1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_118_3_Right_124
timestamp 18001
transform -1 0 88596 0 1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_119_1_Left_270
timestamp 18001
transform 1 0 4876 0 -1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_119_1_Right_558
timestamp 18001
transform -1 0 7912 0 -1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_119_3_Left_418
timestamp 18001
transform 1 0 85284 0 -1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_119_3_Right_125
timestamp 18001
transform -1 0 88596 0 -1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_120_1_Left_271
timestamp 18001
transform 1 0 4876 0 1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_120_1_Right_559
timestamp 18001
transform -1 0 7912 0 1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_120_3_Left_419
timestamp 18001
transform 1 0 85284 0 1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_120_3_Right_126
timestamp 18001
transform -1 0 88596 0 1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_121_1_Left_272
timestamp 18001
transform 1 0 4876 0 -1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_121_1_Right_560
timestamp 18001
transform -1 0 7912 0 -1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_121_3_Left_420
timestamp 18001
transform 1 0 85284 0 -1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_121_3_Right_127
timestamp 18001
transform -1 0 88596 0 -1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_122_1_Left_273
timestamp 18001
transform 1 0 4876 0 1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_122_1_Right_561
timestamp 18001
transform -1 0 7912 0 1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_122_3_Left_421
timestamp 18001
transform 1 0 85284 0 1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_122_3_Right_128
timestamp 18001
transform -1 0 88596 0 1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_123_1_Left_274
timestamp 18001
transform 1 0 4876 0 -1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_123_1_Right_562
timestamp 18001
transform -1 0 7912 0 -1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_123_3_Left_422
timestamp 18001
transform 1 0 85284 0 -1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_123_3_Right_129
timestamp 18001
transform -1 0 88596 0 -1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_124_1_Left_275
timestamp 18001
transform 1 0 4876 0 1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_124_1_Right_563
timestamp 18001
transform -1 0 7912 0 1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_124_3_Left_423
timestamp 18001
transform 1 0 85284 0 1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_124_3_Right_130
timestamp 18001
transform -1 0 88596 0 1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_125_1_Left_276
timestamp 18001
transform 1 0 4876 0 -1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_125_1_Right_564
timestamp 18001
transform -1 0 7912 0 -1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_125_3_Left_424
timestamp 18001
transform 1 0 85284 0 -1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_125_3_Right_131
timestamp 18001
transform -1 0 88596 0 -1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_126_1_Left_277
timestamp 18001
transform 1 0 4876 0 1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_126_1_Right_565
timestamp 18001
transform -1 0 7912 0 1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_126_3_Left_425
timestamp 18001
transform 1 0 85284 0 1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_126_3_Right_132
timestamp 18001
transform -1 0 88596 0 1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_127_1_Left_278
timestamp 18001
transform 1 0 4876 0 -1 74528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_127_1_Right_566
timestamp 18001
transform -1 0 7912 0 -1 74528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_127_3_Left_426
timestamp 18001
transform 1 0 85284 0 -1 74528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_127_3_Right_133
timestamp 18001
transform -1 0 88596 0 -1 74528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_128_1_Left_279
timestamp 18001
transform 1 0 4876 0 1 74528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_128_1_Right_567
timestamp 18001
transform -1 0 7912 0 1 74528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_128_3_Left_427
timestamp 18001
transform 1 0 85284 0 1 74528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_128_3_Right_134
timestamp 18001
transform -1 0 88596 0 1 74528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_129_1_Left_280
timestamp 18001
transform 1 0 4876 0 -1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_129_1_Right_568
timestamp 18001
transform -1 0 7912 0 -1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_129_3_Left_428
timestamp 18001
transform 1 0 85284 0 -1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_129_3_Right_135
timestamp 18001
transform -1 0 88596 0 -1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_130_1_Left_281
timestamp 18001
transform 1 0 4876 0 1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_130_1_Right_569
timestamp 18001
transform -1 0 7912 0 1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_130_3_Left_429
timestamp 18001
transform 1 0 85284 0 1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_130_3_Right_136
timestamp 18001
transform -1 0 88596 0 1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_131_1_Left_282
timestamp 18001
transform 1 0 4876 0 -1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_131_1_Right_570
timestamp 18001
transform -1 0 7912 0 -1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_131_3_Left_430
timestamp 18001
transform 1 0 85284 0 -1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_131_3_Right_137
timestamp 18001
transform -1 0 88596 0 -1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_132_1_Left_283
timestamp 18001
transform 1 0 4876 0 1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_132_1_Right_571
timestamp 18001
transform -1 0 7912 0 1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_132_3_Left_431
timestamp 18001
transform 1 0 85284 0 1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_132_3_Right_138
timestamp 18001
transform -1 0 88596 0 1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_133_1_Left_284
timestamp 18001
transform 1 0 4876 0 -1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_133_1_Right_572
timestamp 18001
transform -1 0 7912 0 -1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_133_3_Left_432
timestamp 18001
transform 1 0 85284 0 -1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_133_3_Right_139
timestamp 18001
transform -1 0 88596 0 -1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_134_1_Left_285
timestamp 18001
transform 1 0 4876 0 1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_134_1_Right_573
timestamp 18001
transform -1 0 7912 0 1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_134_3_Left_433
timestamp 18001
transform 1 0 85284 0 1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_134_3_Right_140
timestamp 18001
transform -1 0 88596 0 1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_135_1_Left_286
timestamp 18001
transform 1 0 4876 0 -1 78880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_135_1_Right_574
timestamp 18001
transform -1 0 7912 0 -1 78880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_135_3_Left_434
timestamp 18001
transform 1 0 85284 0 -1 78880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_135_3_Right_141
timestamp 18001
transform -1 0 88596 0 -1 78880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_136_1_Left_287
timestamp 18001
transform 1 0 4876 0 1 78880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_136_1_Right_575
timestamp 18001
transform -1 0 7912 0 1 78880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_136_3_Left_435
timestamp 18001
transform 1 0 85284 0 1 78880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_136_3_Right_142
timestamp 18001
transform -1 0 88596 0 1 78880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_137_1_Left_288
timestamp 18001
transform 1 0 4876 0 -1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_137_1_Right_576
timestamp 18001
transform -1 0 7912 0 -1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_137_3_Left_436
timestamp 18001
transform 1 0 85284 0 -1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_137_3_Right_143
timestamp 18001
transform -1 0 88596 0 -1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_138_1_Left_289
timestamp 18001
transform 1 0 4876 0 1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_138_1_Right_577
timestamp 18001
transform -1 0 7912 0 1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_138_3_Left_437
timestamp 18001
transform 1 0 85284 0 1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_138_3_Right_144
timestamp 18001
transform -1 0 88596 0 1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_139_1_Left_290
timestamp 18001
transform 1 0 4876 0 -1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_139_1_Right_578
timestamp 18001
transform -1 0 7912 0 -1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_139_3_Left_438
timestamp 18001
transform 1 0 85284 0 -1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_139_3_Right_145
timestamp 18001
transform -1 0 88596 0 -1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_140_1_Left_291
timestamp 18001
transform 1 0 4876 0 1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_140_1_Right_579
timestamp 18001
transform -1 0 7912 0 1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_140_3_Left_439
timestamp 18001
transform 1 0 85284 0 1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_140_3_Right_146
timestamp 18001
transform -1 0 88596 0 1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_141_1_Left_292
timestamp 18001
transform 1 0 4876 0 -1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_141_1_Right_580
timestamp 18001
transform -1 0 7912 0 -1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_141_3_Left_440
timestamp 18001
transform 1 0 85284 0 -1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_141_3_Right_147
timestamp 18001
transform -1 0 88596 0 -1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_142_1_Left_293
timestamp 18001
transform 1 0 4876 0 1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_142_1_Right_581
timestamp 18001
transform -1 0 7912 0 1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_142_3_Left_441
timestamp 18001
transform 1 0 85284 0 1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_142_3_Right_148
timestamp 18001
transform -1 0 88596 0 1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_143_1_Left_294
timestamp 18001
transform 1 0 4876 0 -1 83232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_143_1_Right_582
timestamp 18001
transform -1 0 7912 0 -1 83232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_143_3_Left_442
timestamp 18001
transform 1 0 85284 0 -1 83232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_143_3_Right_149
timestamp 18001
transform -1 0 88596 0 -1 83232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_144_1_Left_295
timestamp 18001
transform 1 0 4876 0 1 83232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_144_1_Right_583
timestamp 18001
transform -1 0 7912 0 1 83232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_144_3_Left_443
timestamp 18001
transform 1 0 85284 0 1 83232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_144_3_Right_150
timestamp 18001
transform -1 0 88596 0 1 83232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_145_1_Left_296
timestamp 18001
transform 1 0 4876 0 -1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_145_1_Right_584
timestamp 18001
transform -1 0 7912 0 -1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_145_3_Left_444
timestamp 18001
transform 1 0 85284 0 -1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_145_3_Right_151
timestamp 18001
transform -1 0 88596 0 -1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_146_Left_297
timestamp 18001
transform 1 0 4876 0 1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_146_Right_5
timestamp 18001
transform -1 0 88596 0 1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_147_Left_298
timestamp 18001
transform 1 0 4876 0 -1 85408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_147_Right_6
timestamp 18001
transform -1 0 88596 0 -1 85408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_148_Left_299
timestamp 18001
transform 1 0 4876 0 1 85408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_148_Right_7
timestamp 18001
transform -1 0 88596 0 1 85408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_149_Left_300
timestamp 18001
transform 1 0 4876 0 -1 86496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_149_Right_8
timestamp 18001
transform -1 0 88596 0 -1 86496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_150_Left_301
timestamp 18001
transform 1 0 4876 0 1 86496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_150_Right_9
timestamp 18001
transform -1 0 88596 0 1 86496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_151_Left_302
timestamp 18001
transform 1 0 4876 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_151_Right_10
timestamp 18001
transform -1 0 88596 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_586
timestamp 18001
transform 1 0 7452 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_587
timestamp 18001
transform 1 0 10028 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_588
timestamp 18001
transform 1 0 12604 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_589
timestamp 18001
transform 1 0 15180 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_590
timestamp 18001
transform 1 0 17756 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_591
timestamp 18001
transform 1 0 20332 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_592
timestamp 18001
transform 1 0 22908 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_593
timestamp 18001
transform 1 0 25484 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_594
timestamp 18001
transform 1 0 28060 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_595
timestamp 18001
transform 1 0 30636 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_596
timestamp 18001
transform 1 0 33212 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_597
timestamp 18001
transform 1 0 35788 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_598
timestamp 18001
transform 1 0 38364 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_599
timestamp 18001
transform 1 0 40940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_600
timestamp 18001
transform 1 0 43516 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_601
timestamp 18001
transform 1 0 46092 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_602
timestamp 18001
transform 1 0 48668 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_603
timestamp 18001
transform 1 0 51244 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_604
timestamp 18001
transform 1 0 53820 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_605
timestamp 18001
transform 1 0 56396 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_606
timestamp 18001
transform 1 0 58972 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_607
timestamp 18001
transform 1 0 61548 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_608
timestamp 18001
transform 1 0 64124 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_609
timestamp 18001
transform 1 0 66700 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_610
timestamp 18001
transform 1 0 69276 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_611
timestamp 18001
transform 1 0 71852 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_612
timestamp 18001
transform 1 0 74428 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_613
timestamp 18001
transform 1 0 77004 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_614
timestamp 18001
transform 1 0 79580 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_615
timestamp 18001
transform 1 0 82156 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_616
timestamp 18001
transform 1 0 84732 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_617
timestamp 18001
transform 1 0 87308 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_618
timestamp 18001
transform 1 0 10028 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_619
timestamp 18001
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_620
timestamp 18001
transform 1 0 20332 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_621
timestamp 18001
transform 1 0 25484 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_622
timestamp 18001
transform 1 0 30636 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_623
timestamp 18001
transform 1 0 35788 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_624
timestamp 18001
transform 1 0 40940 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_625
timestamp 18001
transform 1 0 46092 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_626
timestamp 18001
transform 1 0 51244 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_627
timestamp 18001
transform 1 0 56396 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_628
timestamp 18001
transform 1 0 61548 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_629
timestamp 18001
transform 1 0 66700 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_630
timestamp 18001
transform 1 0 71852 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_631
timestamp 18001
transform 1 0 77004 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_632
timestamp 18001
transform 1 0 82156 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_633
timestamp 18001
transform 1 0 87308 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_634
timestamp 18001
transform 1 0 7452 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_635
timestamp 18001
transform 1 0 12604 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_636
timestamp 18001
transform 1 0 17756 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_637
timestamp 18001
transform 1 0 22908 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_638
timestamp 18001
transform 1 0 28060 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_639
timestamp 18001
transform 1 0 33212 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_640
timestamp 18001
transform 1 0 38364 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_641
timestamp 18001
transform 1 0 43516 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_642
timestamp 18001
transform 1 0 48668 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_643
timestamp 18001
transform 1 0 53820 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_644
timestamp 18001
transform 1 0 58972 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_645
timestamp 18001
transform 1 0 64124 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_646
timestamp 18001
transform 1 0 69276 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_647
timestamp 18001
transform 1 0 74428 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_648
timestamp 18001
transform 1 0 79580 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_649
timestamp 18001
transform 1 0 84732 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_650
timestamp 18001
transform 1 0 10028 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_651
timestamp 18001
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_652
timestamp 18001
transform 1 0 20332 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_653
timestamp 18001
transform 1 0 25484 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_654
timestamp 18001
transform 1 0 30636 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_655
timestamp 18001
transform 1 0 35788 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_656
timestamp 18001
transform 1 0 40940 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_657
timestamp 18001
transform 1 0 46092 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_658
timestamp 18001
transform 1 0 51244 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_659
timestamp 18001
transform 1 0 56396 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_660
timestamp 18001
transform 1 0 61548 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_661
timestamp 18001
transform 1 0 66700 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_662
timestamp 18001
transform 1 0 71852 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_663
timestamp 18001
transform 1 0 77004 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_664
timestamp 18001
transform 1 0 82156 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_665
timestamp 18001
transform 1 0 87308 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_666
timestamp 18001
transform 1 0 7452 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_667
timestamp 18001
transform 1 0 10028 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_668
timestamp 18001
transform 1 0 12604 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_669
timestamp 18001
transform 1 0 15180 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_670
timestamp 18001
transform 1 0 17756 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_671
timestamp 18001
transform 1 0 20332 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_672
timestamp 18001
transform 1 0 22908 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_673
timestamp 18001
transform 1 0 25484 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_674
timestamp 18001
transform 1 0 28060 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_675
timestamp 18001
transform 1 0 30636 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_676
timestamp 18001
transform 1 0 33212 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_677
timestamp 18001
transform 1 0 35788 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_678
timestamp 18001
transform 1 0 38364 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_679
timestamp 18001
transform 1 0 40940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_680
timestamp 18001
transform 1 0 43516 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_681
timestamp 18001
transform 1 0 46092 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_682
timestamp 18001
transform 1 0 48668 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_683
timestamp 18001
transform 1 0 51244 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_684
timestamp 18001
transform 1 0 53820 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_685
timestamp 18001
transform 1 0 56396 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_686
timestamp 18001
transform 1 0 58972 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_687
timestamp 18001
transform 1 0 61548 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_688
timestamp 18001
transform 1 0 64124 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_689
timestamp 18001
transform 1 0 66700 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_690
timestamp 18001
transform 1 0 69276 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_691
timestamp 18001
transform 1 0 71852 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_692
timestamp 18001
transform 1 0 74428 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_693
timestamp 18001
transform 1 0 77004 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_694
timestamp 18001
transform 1 0 79580 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_695
timestamp 18001
transform 1 0 82156 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_696
timestamp 18001
transform 1 0 84732 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_697
timestamp 18001
transform 1 0 87308 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1_698
timestamp 18001
transform 1 0 7452 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_3_896
timestamp 18001
transform 1 0 87860 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1_699
timestamp 18001
transform 1 0 7452 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_3_897
timestamp 18001
transform 1 0 87860 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_1_700
timestamp 18001
transform 1 0 7452 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_3_898
timestamp 18001
transform 1 0 87860 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_1_701
timestamp 18001
transform 1 0 7452 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_3_899
timestamp 18001
transform 1 0 87860 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_1_702
timestamp 18001
transform 1 0 7452 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_3_900
timestamp 18001
transform 1 0 87860 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_1_703
timestamp 18001
transform 1 0 7452 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_3_901
timestamp 18001
transform 1 0 87860 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_1_704
timestamp 18001
transform 1 0 7452 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_3_902
timestamp 18001
transform 1 0 87860 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_1_705
timestamp 18001
transform 1 0 7452 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_3_903
timestamp 18001
transform 1 0 87860 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_1_706
timestamp 18001
transform 1 0 7452 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_3_904
timestamp 18001
transform 1 0 87860 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_1_707
timestamp 18001
transform 1 0 7452 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_3_905
timestamp 18001
transform 1 0 87860 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_1_708
timestamp 18001
transform 1 0 7452 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_3_906
timestamp 18001
transform 1 0 87860 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_1_709
timestamp 18001
transform 1 0 7452 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_3_907
timestamp 18001
transform 1 0 87860 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_1_710
timestamp 18001
transform 1 0 7452 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_3_908
timestamp 18001
transform 1 0 87860 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_1_711
timestamp 18001
transform 1 0 7452 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_3_909
timestamp 18001
transform 1 0 87860 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_1_712
timestamp 18001
transform 1 0 7452 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_3_910
timestamp 18001
transform 1 0 87860 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_1_713
timestamp 18001
transform 1 0 7452 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_3_911
timestamp 18001
transform 1 0 87860 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_1_714
timestamp 18001
transform 1 0 7452 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_3_912
timestamp 18001
transform 1 0 87860 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_1_715
timestamp 18001
transform 1 0 7452 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_3_913
timestamp 18001
transform 1 0 87860 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_1_716
timestamp 18001
transform 1 0 7452 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_3_914
timestamp 18001
transform 1 0 87860 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_1_717
timestamp 18001
transform 1 0 7452 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_3_915
timestamp 18001
transform 1 0 87860 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_1_718
timestamp 18001
transform 1 0 7452 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_3_916
timestamp 18001
transform 1 0 87860 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_1_719
timestamp 18001
transform 1 0 7452 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_3_917
timestamp 18001
transform 1 0 87860 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_1_720
timestamp 18001
transform 1 0 7452 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_3_918
timestamp 18001
transform 1 0 87860 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_1_721
timestamp 18001
transform 1 0 7452 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_3_919
timestamp 18001
transform 1 0 87860 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_1_722
timestamp 18001
transform 1 0 7452 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_3_920
timestamp 18001
transform 1 0 87860 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_1_723
timestamp 18001
transform 1 0 7452 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_3_921
timestamp 18001
transform 1 0 87860 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_1_724
timestamp 18001
transform 1 0 7452 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_3_922
timestamp 18001
transform 1 0 87860 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1_725
timestamp 18001
transform 1 0 7452 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_3_923
timestamp 18001
transform 1 0 87860 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1_726
timestamp 18001
transform 1 0 7452 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_3_924
timestamp 18001
transform 1 0 87860 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1_727
timestamp 18001
transform 1 0 7452 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_3_925
timestamp 18001
transform 1 0 87860 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_1_728
timestamp 18001
transform 1 0 7452 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_3_926
timestamp 18001
transform 1 0 87860 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_1_729
timestamp 18001
transform 1 0 7452 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_3_927
timestamp 18001
transform 1 0 87860 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_1_730
timestamp 18001
transform 1 0 7452 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_3_928
timestamp 18001
transform 1 0 87860 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1_731
timestamp 18001
transform 1 0 7452 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_5_929
timestamp 18001
transform 1 0 87860 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1_732
timestamp 18001
transform 1 0 7452 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_5_930
timestamp 18001
transform 1 0 87860 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1_733
timestamp 18001
transform 1 0 7452 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_5_931
timestamp 18001
transform 1 0 87860 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1_734
timestamp 18001
transform 1 0 7452 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_5_932
timestamp 18001
transform 1 0 87860 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1_735
timestamp 18001
transform 1 0 7452 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_3_933
timestamp 18001
transform 1 0 87860 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1_736
timestamp 18001
transform 1 0 7452 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_3_934
timestamp 18001
transform 1 0 87860 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1_737
timestamp 18001
transform 1 0 7452 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_3_935
timestamp 18001
transform 1 0 87860 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1_738
timestamp 18001
transform 1 0 7452 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_3_936
timestamp 18001
transform 1 0 87860 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1_739
timestamp 18001
transform 1 0 7452 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_3_937
timestamp 18001
transform 1 0 87860 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1_740
timestamp 18001
transform 1 0 7452 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_3_938
timestamp 18001
transform 1 0 87860 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1_741
timestamp 18001
transform 1 0 7452 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_3_939
timestamp 18001
transform 1 0 87860 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1_742
timestamp 18001
transform 1 0 7452 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_3_940
timestamp 18001
transform 1 0 87860 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1_743
timestamp 18001
transform 1 0 7452 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_3_941
timestamp 18001
transform 1 0 87860 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1_744
timestamp 18001
transform 1 0 7452 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_3_942
timestamp 18001
transform 1 0 87860 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1_745
timestamp 18001
transform 1 0 7452 0 1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_3_943
timestamp 18001
transform 1 0 87860 0 1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_1_746
timestamp 18001
transform 1 0 7452 0 1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_3_944
timestamp 18001
transform 1 0 87860 0 1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_1_747
timestamp 18001
transform 1 0 7452 0 1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_3_945
timestamp 18001
transform 1 0 87860 0 1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_1_748
timestamp 18001
transform 1 0 7452 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_3_946
timestamp 18001
transform 1 0 87860 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_1_749
timestamp 18001
transform 1 0 7452 0 1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_3_947
timestamp 18001
transform 1 0 87860 0 1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_1_750
timestamp 18001
transform 1 0 7452 0 1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_3_948
timestamp 18001
transform 1 0 87860 0 1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_1_751
timestamp 18001
transform 1 0 7452 0 1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_3_949
timestamp 18001
transform 1 0 87860 0 1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_1_752
timestamp 18001
transform 1 0 7452 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_3_950
timestamp 18001
transform 1 0 87860 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_1_753
timestamp 18001
transform 1 0 7452 0 1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_3_951
timestamp 18001
transform 1 0 87860 0 1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1_754
timestamp 18001
transform 1 0 7452 0 1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_3_952
timestamp 18001
transform 1 0 87860 0 1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1_755
timestamp 18001
transform 1 0 7452 0 1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_3_953
timestamp 18001
transform 1 0 87860 0 1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1_756
timestamp 18001
transform 1 0 7452 0 1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_3_954
timestamp 18001
transform 1 0 87860 0 1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1_757
timestamp 18001
transform 1 0 7452 0 1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_3_955
timestamp 18001
transform 1 0 87860 0 1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1_758
timestamp 18001
transform 1 0 7452 0 1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_3_956
timestamp 18001
transform 1 0 87860 0 1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1_759
timestamp 18001
transform 1 0 7452 0 1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_3_957
timestamp 18001
transform 1 0 87860 0 1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1_760
timestamp 18001
transform 1 0 7452 0 1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_3_958
timestamp 18001
transform 1 0 87860 0 1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1_761
timestamp 18001
transform 1 0 7452 0 1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_3_959
timestamp 18001
transform 1 0 87860 0 1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1_762
timestamp 18001
transform 1 0 7452 0 1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_3_960
timestamp 18001
transform 1 0 87860 0 1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1_763
timestamp 18001
transform 1 0 7452 0 1 78880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_3_961
timestamp 18001
transform 1 0 87860 0 1 78880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1_764
timestamp 18001
transform 1 0 7452 0 1 79968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_3_962
timestamp 18001
transform 1 0 87860 0 1 79968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_140_1_765
timestamp 18001
transform 1 0 7452 0 1 81056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_140_3_963
timestamp 18001
transform 1 0 87860 0 1 81056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_142_1_766
timestamp 18001
transform 1 0 7452 0 1 82144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_142_3_964
timestamp 18001
transform 1 0 87860 0 1 82144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_144_1_767
timestamp 18001
transform 1 0 7452 0 1 83232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_144_3_965
timestamp 18001
transform 1 0 87860 0 1 83232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_768
timestamp 18001
transform 1 0 7452 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_769
timestamp 18001
transform 1 0 10028 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_770
timestamp 18001
transform 1 0 12604 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_771
timestamp 18001
transform 1 0 15180 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_772
timestamp 18001
transform 1 0 17756 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_773
timestamp 18001
transform 1 0 20332 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_774
timestamp 18001
transform 1 0 22908 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_775
timestamp 18001
transform 1 0 25484 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_776
timestamp 18001
transform 1 0 28060 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_777
timestamp 18001
transform 1 0 30636 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_778
timestamp 18001
transform 1 0 33212 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_779
timestamp 18001
transform 1 0 35788 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_780
timestamp 18001
transform 1 0 38364 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_781
timestamp 18001
transform 1 0 40940 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_782
timestamp 18001
transform 1 0 43516 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_783
timestamp 18001
transform 1 0 46092 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_784
timestamp 18001
transform 1 0 48668 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_785
timestamp 18001
transform 1 0 51244 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_786
timestamp 18001
transform 1 0 53820 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_787
timestamp 18001
transform 1 0 56396 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_788
timestamp 18001
transform 1 0 58972 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_789
timestamp 18001
transform 1 0 61548 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_790
timestamp 18001
transform 1 0 64124 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_791
timestamp 18001
transform 1 0 66700 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_792
timestamp 18001
transform 1 0 69276 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_793
timestamp 18001
transform 1 0 71852 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_794
timestamp 18001
transform 1 0 74428 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_795
timestamp 18001
transform 1 0 77004 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_796
timestamp 18001
transform 1 0 79580 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_797
timestamp 18001
transform 1 0 82156 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_798
timestamp 18001
transform 1 0 84732 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_799
timestamp 18001
transform 1 0 87308 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_800
timestamp 18001
transform 1 0 10028 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_801
timestamp 18001
transform 1 0 15180 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_802
timestamp 18001
transform 1 0 20332 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_803
timestamp 18001
transform 1 0 25484 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_804
timestamp 18001
transform 1 0 30636 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_805
timestamp 18001
transform 1 0 35788 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_806
timestamp 18001
transform 1 0 40940 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_807
timestamp 18001
transform 1 0 46092 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_808
timestamp 18001
transform 1 0 51244 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_809
timestamp 18001
transform 1 0 56396 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_810
timestamp 18001
transform 1 0 61548 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_811
timestamp 18001
transform 1 0 66700 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_812
timestamp 18001
transform 1 0 71852 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_813
timestamp 18001
transform 1 0 77004 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_814
timestamp 18001
transform 1 0 82156 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_815
timestamp 18001
transform 1 0 87308 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_816
timestamp 18001
transform 1 0 7452 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_817
timestamp 18001
transform 1 0 12604 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_818
timestamp 18001
transform 1 0 17756 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_819
timestamp 18001
transform 1 0 22908 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_820
timestamp 18001
transform 1 0 28060 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_821
timestamp 18001
transform 1 0 33212 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_822
timestamp 18001
transform 1 0 38364 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_823
timestamp 18001
transform 1 0 43516 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_824
timestamp 18001
transform 1 0 48668 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_825
timestamp 18001
transform 1 0 53820 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_826
timestamp 18001
transform 1 0 58972 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_827
timestamp 18001
transform 1 0 64124 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_828
timestamp 18001
transform 1 0 69276 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_829
timestamp 18001
transform 1 0 74428 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_830
timestamp 18001
transform 1 0 79580 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_831
timestamp 18001
transform 1 0 84732 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_832
timestamp 18001
transform 1 0 10028 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_833
timestamp 18001
transform 1 0 15180 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_834
timestamp 18001
transform 1 0 20332 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_835
timestamp 18001
transform 1 0 25484 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_836
timestamp 18001
transform 1 0 30636 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_837
timestamp 18001
transform 1 0 35788 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_838
timestamp 18001
transform 1 0 40940 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_839
timestamp 18001
transform 1 0 46092 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_840
timestamp 18001
transform 1 0 51244 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_841
timestamp 18001
transform 1 0 56396 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_842
timestamp 18001
transform 1 0 61548 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_843
timestamp 18001
transform 1 0 66700 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_844
timestamp 18001
transform 1 0 71852 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_845
timestamp 18001
transform 1 0 77004 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_846
timestamp 18001
transform 1 0 82156 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_847
timestamp 18001
transform 1 0 87308 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_848
timestamp 18001
transform 1 0 7452 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_849
timestamp 18001
transform 1 0 12604 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_850
timestamp 18001
transform 1 0 17756 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_851
timestamp 18001
transform 1 0 22908 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_852
timestamp 18001
transform 1 0 28060 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_853
timestamp 18001
transform 1 0 33212 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_854
timestamp 18001
transform 1 0 38364 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_855
timestamp 18001
transform 1 0 43516 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_856
timestamp 18001
transform 1 0 48668 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_857
timestamp 18001
transform 1 0 53820 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_858
timestamp 18001
transform 1 0 58972 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_859
timestamp 18001
transform 1 0 64124 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_860
timestamp 18001
transform 1 0 69276 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_861
timestamp 18001
transform 1 0 74428 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_862
timestamp 18001
transform 1 0 79580 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_863
timestamp 18001
transform 1 0 84732 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_864
timestamp 18001
transform 1 0 7452 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_865
timestamp 18001
transform 1 0 10028 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_866
timestamp 18001
transform 1 0 12604 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_867
timestamp 18001
transform 1 0 15180 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_868
timestamp 18001
transform 1 0 17756 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_869
timestamp 18001
transform 1 0 20332 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_870
timestamp 18001
transform 1 0 22908 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_871
timestamp 18001
transform 1 0 25484 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_872
timestamp 18001
transform 1 0 28060 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_873
timestamp 18001
transform 1 0 30636 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_874
timestamp 18001
transform 1 0 33212 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_875
timestamp 18001
transform 1 0 35788 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_876
timestamp 18001
transform 1 0 38364 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_877
timestamp 18001
transform 1 0 40940 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_878
timestamp 18001
transform 1 0 43516 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_879
timestamp 18001
transform 1 0 46092 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_880
timestamp 18001
transform 1 0 48668 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_881
timestamp 18001
transform 1 0 51244 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_882
timestamp 18001
transform 1 0 53820 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_883
timestamp 18001
transform 1 0 56396 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_884
timestamp 18001
transform 1 0 58972 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_885
timestamp 18001
transform 1 0 61548 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_886
timestamp 18001
transform 1 0 64124 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_887
timestamp 18001
transform 1 0 66700 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_888
timestamp 18001
transform 1 0 69276 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_889
timestamp 18001
transform 1 0 71852 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_890
timestamp 18001
transform 1 0 74428 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_891
timestamp 18001
transform 1 0 77004 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_892
timestamp 18001
transform 1 0 79580 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_893
timestamp 18001
transform 1 0 82156 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_894
timestamp 18001
transform 1 0 84732 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_895
timestamp 18001
transform 1 0 87308 0 -1 87584
box -38 -48 130 592
<< labels >>
flabel metal2 s 39726 88000 39782 88800 0 FreeSans 224 90 0 0 clk
port 0 nsew signal input
flabel metal3 s 3000 45168 3800 45288 0 FreeSans 480 0 0 0 config_data_in
port 1 nsew signal input
flabel metal3 s 89200 47208 90000 47328 0 FreeSans 480 0 0 0 config_data_out
port 2 nsew signal output
flabel metal2 s 36506 88000 36562 88800 0 FreeSans 224 90 0 0 config_en
port 3 nsew signal input
flabel metal3 s 89200 30208 90000 30328 0 FreeSans 480 0 0 0 io_east_in[0]
port 4 nsew signal input
flabel metal3 s 89200 41088 90000 41208 0 FreeSans 480 0 0 0 io_east_in[10]
port 5 nsew signal input
flabel metal3 s 89200 42448 90000 42568 0 FreeSans 480 0 0 0 io_east_in[11]
port 6 nsew signal input
flabel metal3 s 89200 43128 90000 43248 0 FreeSans 480 0 0 0 io_east_in[12]
port 7 nsew signal input
flabel metal3 s 89200 43808 90000 43928 0 FreeSans 480 0 0 0 io_east_in[13]
port 8 nsew signal input
flabel metal2 s 3018 3000 3074 3800 0 FreeSans 224 90 0 0 io_east_in[14]
port 9 nsew signal input
flabel metal2 s 3662 3000 3718 3800 0 FreeSans 224 90 0 0 io_east_in[15]
port 10 nsew signal input
flabel metal3 s 89200 66928 90000 67048 0 FreeSans 480 0 0 0 io_east_in[16]
port 11 nsew signal input
flabel metal3 s 89200 67608 90000 67728 0 FreeSans 480 0 0 0 io_east_in[17]
port 12 nsew signal input
flabel metal3 s 89200 68968 90000 69088 0 FreeSans 480 0 0 0 io_east_in[18]
port 13 nsew signal input
flabel metal3 s 89200 70328 90000 70448 0 FreeSans 480 0 0 0 io_east_in[19]
port 14 nsew signal input
flabel metal3 s 89200 31568 90000 31688 0 FreeSans 480 0 0 0 io_east_in[1]
port 15 nsew signal input
flabel metal3 s 89200 71008 90000 71128 0 FreeSans 480 0 0 0 io_east_in[20]
port 16 nsew signal input
flabel metal3 s 89200 72368 90000 72488 0 FreeSans 480 0 0 0 io_east_in[21]
port 17 nsew signal input
flabel metal3 s 89200 73048 90000 73168 0 FreeSans 480 0 0 0 io_east_in[22]
port 18 nsew signal input
flabel metal3 s 89200 74408 90000 74528 0 FreeSans 480 0 0 0 io_east_in[23]
port 19 nsew signal input
flabel metal3 s 89200 75768 90000 75888 0 FreeSans 480 0 0 0 io_east_in[24]
port 20 nsew signal input
flabel metal3 s 89200 76448 90000 76568 0 FreeSans 480 0 0 0 io_east_in[25]
port 21 nsew signal input
flabel metal3 s 89200 77808 90000 77928 0 FreeSans 480 0 0 0 io_east_in[26]
port 22 nsew signal input
flabel metal3 s 89200 78488 90000 78608 0 FreeSans 480 0 0 0 io_east_in[27]
port 23 nsew signal input
flabel metal3 s 89200 79848 90000 79968 0 FreeSans 480 0 0 0 io_east_in[28]
port 24 nsew signal input
flabel metal3 s 89200 81208 90000 81328 0 FreeSans 480 0 0 0 io_east_in[29]
port 25 nsew signal input
flabel metal3 s 89200 32248 90000 32368 0 FreeSans 480 0 0 0 io_east_in[2]
port 26 nsew signal input
flabel metal2 s 4306 3000 4362 3800 0 FreeSans 224 90 0 0 io_east_in[30]
port 27 nsew signal input
flabel metal2 s 4950 3000 5006 3800 0 FreeSans 224 90 0 0 io_east_in[31]
port 28 nsew signal input
flabel metal3 s 89200 33608 90000 33728 0 FreeSans 480 0 0 0 io_east_in[3]
port 29 nsew signal input
flabel metal3 s 89200 34968 90000 35088 0 FreeSans 480 0 0 0 io_east_in[4]
port 30 nsew signal input
flabel metal3 s 89200 35648 90000 35768 0 FreeSans 480 0 0 0 io_east_in[5]
port 31 nsew signal input
flabel metal3 s 89200 37008 90000 37128 0 FreeSans 480 0 0 0 io_east_in[6]
port 32 nsew signal input
flabel metal3 s 89200 37688 90000 37808 0 FreeSans 480 0 0 0 io_east_in[7]
port 33 nsew signal input
flabel metal3 s 89200 39048 90000 39168 0 FreeSans 480 0 0 0 io_east_in[8]
port 34 nsew signal input
flabel metal3 s 89200 40408 90000 40528 0 FreeSans 480 0 0 0 io_east_in[9]
port 35 nsew signal input
flabel metal3 s 89200 15248 90000 15368 0 FreeSans 480 0 0 0 io_east_out[0]
port 36 nsew signal output
flabel metal3 s 89200 26128 90000 26248 0 FreeSans 480 0 0 0 io_east_out[10]
port 37 nsew signal output
flabel metal3 s 89200 26808 90000 26928 0 FreeSans 480 0 0 0 io_east_out[11]
port 38 nsew signal output
flabel metal3 s 89200 28168 90000 28288 0 FreeSans 480 0 0 0 io_east_out[12]
port 39 nsew signal output
flabel metal3 s 89200 29528 90000 29648 0 FreeSans 480 0 0 0 io_east_out[13]
port 40 nsew signal output
flabel metal2 s 46166 88000 46222 88800 0 FreeSans 224 90 0 0 io_east_out[14]
port 41 nsew signal output
flabel metal2 s 50030 88000 50086 88800 0 FreeSans 224 90 0 0 io_east_out[15]
port 42 nsew signal output
flabel metal3 s 89200 51288 90000 51408 0 FreeSans 480 0 0 0 io_east_out[16]
port 43 nsew signal output
flabel metal3 s 89200 52648 90000 52768 0 FreeSans 480 0 0 0 io_east_out[17]
port 44 nsew signal output
flabel metal3 s 89200 54008 90000 54128 0 FreeSans 480 0 0 0 io_east_out[18]
port 45 nsew signal output
flabel metal3 s 89200 54688 90000 54808 0 FreeSans 480 0 0 0 io_east_out[19]
port 46 nsew signal output
flabel metal3 s 89200 15928 90000 16048 0 FreeSans 480 0 0 0 io_east_out[1]
port 47 nsew signal output
flabel metal3 s 89200 56048 90000 56168 0 FreeSans 480 0 0 0 io_east_out[20]
port 48 nsew signal output
flabel metal3 s 89200 56728 90000 56848 0 FreeSans 480 0 0 0 io_east_out[21]
port 49 nsew signal output
flabel metal3 s 89200 58088 90000 58208 0 FreeSans 480 0 0 0 io_east_out[22]
port 50 nsew signal output
flabel metal3 s 89200 59448 90000 59568 0 FreeSans 480 0 0 0 io_east_out[23]
port 51 nsew signal output
flabel metal3 s 89200 60128 90000 60248 0 FreeSans 480 0 0 0 io_east_out[24]
port 52 nsew signal output
flabel metal3 s 89200 61488 90000 61608 0 FreeSans 480 0 0 0 io_east_out[25]
port 53 nsew signal output
flabel metal3 s 89200 62168 90000 62288 0 FreeSans 480 0 0 0 io_east_out[26]
port 54 nsew signal output
flabel metal3 s 89200 63528 90000 63648 0 FreeSans 480 0 0 0 io_east_out[27]
port 55 nsew signal output
flabel metal3 s 89200 64888 90000 65008 0 FreeSans 480 0 0 0 io_east_out[28]
port 56 nsew signal output
flabel metal3 s 89200 65568 90000 65688 0 FreeSans 480 0 0 0 io_east_out[29]
port 57 nsew signal output
flabel metal3 s 89200 17288 90000 17408 0 FreeSans 480 0 0 0 io_east_out[2]
port 58 nsew signal output
flabel metal2 s 47454 88000 47510 88800 0 FreeSans 224 90 0 0 io_east_out[30]
port 59 nsew signal output
flabel metal2 s 41658 88000 41714 88800 0 FreeSans 224 90 0 0 io_east_out[31]
port 60 nsew signal output
flabel metal3 s 89200 18648 90000 18768 0 FreeSans 480 0 0 0 io_east_out[3]
port 61 nsew signal output
flabel metal3 s 89200 19328 90000 19448 0 FreeSans 480 0 0 0 io_east_out[4]
port 62 nsew signal output
flabel metal3 s 89200 20688 90000 20808 0 FreeSans 480 0 0 0 io_east_out[5]
port 63 nsew signal output
flabel metal3 s 89200 21368 90000 21488 0 FreeSans 480 0 0 0 io_east_out[6]
port 64 nsew signal output
flabel metal3 s 89200 22728 90000 22848 0 FreeSans 480 0 0 0 io_east_out[7]
port 65 nsew signal output
flabel metal3 s 89200 24088 90000 24208 0 FreeSans 480 0 0 0 io_east_out[8]
port 66 nsew signal output
flabel metal3 s 89200 24768 90000 24888 0 FreeSans 480 0 0 0 io_east_out[9]
port 67 nsew signal output
flabel metal2 s 15254 88000 15310 88800 0 FreeSans 224 90 0 0 io_north_in[0]
port 68 nsew signal input
flabel metal2 s 26202 88000 26258 88800 0 FreeSans 224 90 0 0 io_north_in[10]
port 69 nsew signal input
flabel metal2 s 26846 88000 26902 88800 0 FreeSans 224 90 0 0 io_north_in[11]
port 70 nsew signal input
flabel metal2 s 28134 88000 28190 88800 0 FreeSans 224 90 0 0 io_north_in[12]
port 71 nsew signal input
flabel metal2 s 29422 88000 29478 88800 0 FreeSans 224 90 0 0 io_north_in[13]
port 72 nsew signal input
flabel metal2 s 5594 3000 5650 3800 0 FreeSans 224 90 0 0 io_north_in[14]
port 73 nsew signal input
flabel metal2 s 6238 3000 6294 3800 0 FreeSans 224 90 0 0 io_north_in[15]
port 74 nsew signal input
flabel metal2 s 52606 88000 52662 88800 0 FreeSans 224 90 0 0 io_north_in[16]
port 75 nsew signal input
flabel metal2 s 53250 88000 53306 88800 0 FreeSans 224 90 0 0 io_north_in[17]
port 76 nsew signal input
flabel metal2 s 54538 88000 54594 88800 0 FreeSans 224 90 0 0 io_north_in[18]
port 77 nsew signal input
flabel metal2 s 55826 88000 55882 88800 0 FreeSans 224 90 0 0 io_north_in[19]
port 78 nsew signal input
flabel metal2 s 15898 88000 15954 88800 0 FreeSans 224 90 0 0 io_north_in[1]
port 79 nsew signal input
flabel metal2 s 57114 88000 57170 88800 0 FreeSans 224 90 0 0 io_north_in[20]
port 80 nsew signal input
flabel metal2 s 57758 88000 57814 88800 0 FreeSans 224 90 0 0 io_north_in[21]
port 81 nsew signal input
flabel metal2 s 59046 88000 59102 88800 0 FreeSans 224 90 0 0 io_north_in[22]
port 82 nsew signal input
flabel metal2 s 60334 88000 60390 88800 0 FreeSans 224 90 0 0 io_north_in[23]
port 83 nsew signal input
flabel metal2 s 60978 88000 61034 88800 0 FreeSans 224 90 0 0 io_north_in[24]
port 84 nsew signal input
flabel metal2 s 62266 88000 62322 88800 0 FreeSans 224 90 0 0 io_north_in[25]
port 85 nsew signal input
flabel metal2 s 63554 88000 63610 88800 0 FreeSans 224 90 0 0 io_north_in[26]
port 86 nsew signal input
flabel metal2 s 64842 88000 64898 88800 0 FreeSans 224 90 0 0 io_north_in[27]
port 87 nsew signal input
flabel metal2 s 65486 88000 65542 88800 0 FreeSans 224 90 0 0 io_north_in[28]
port 88 nsew signal input
flabel metal2 s 66774 88000 66830 88800 0 FreeSans 224 90 0 0 io_north_in[29]
port 89 nsew signal input
flabel metal2 s 17186 88000 17242 88800 0 FreeSans 224 90 0 0 io_north_in[2]
port 90 nsew signal input
flabel metal2 s 6882 3000 6938 3800 0 FreeSans 224 90 0 0 io_north_in[30]
port 91 nsew signal input
flabel metal2 s 7526 3000 7582 3800 0 FreeSans 224 90 0 0 io_north_in[31]
port 92 nsew signal input
flabel metal2 s 18474 88000 18530 88800 0 FreeSans 224 90 0 0 io_north_in[3]
port 93 nsew signal input
flabel metal2 s 19118 88000 19174 88800 0 FreeSans 224 90 0 0 io_north_in[4]
port 94 nsew signal input
flabel metal2 s 20406 88000 20462 88800 0 FreeSans 224 90 0 0 io_north_in[5]
port 95 nsew signal input
flabel metal2 s 21694 88000 21750 88800 0 FreeSans 224 90 0 0 io_north_in[6]
port 96 nsew signal input
flabel metal2 s 22982 88000 23038 88800 0 FreeSans 224 90 0 0 io_north_in[7]
port 97 nsew signal input
flabel metal2 s 23626 88000 23682 88800 0 FreeSans 224 90 0 0 io_north_in[8]
port 98 nsew signal input
flabel metal2 s 24914 88000 24970 88800 0 FreeSans 224 90 0 0 io_north_in[9]
port 99 nsew signal input
flabel metal2 s 30710 88000 30766 88800 0 FreeSans 224 90 0 0 io_north_out[0]
port 100 nsew signal output
flabel metal2 s 41014 88000 41070 88800 0 FreeSans 224 90 0 0 io_north_out[10]
port 101 nsew signal output
flabel metal2 s 42302 88000 42358 88800 0 FreeSans 224 90 0 0 io_north_out[11]
port 102 nsew signal output
flabel metal2 s 43590 88000 43646 88800 0 FreeSans 224 90 0 0 io_north_out[12]
port 103 nsew signal output
flabel metal2 s 44234 88000 44290 88800 0 FreeSans 224 90 0 0 io_north_out[13]
port 104 nsew signal output
flabel metal2 s 48742 88000 48798 88800 0 FreeSans 224 90 0 0 io_north_out[14]
port 105 nsew signal output
flabel metal3 s 89200 47888 90000 48008 0 FreeSans 480 0 0 0 io_north_out[15]
port 106 nsew signal output
flabel metal2 s 68062 88000 68118 88800 0 FreeSans 224 90 0 0 io_north_out[16]
port 107 nsew signal output
flabel metal2 s 68706 88000 68762 88800 0 FreeSans 224 90 0 0 io_north_out[17]
port 108 nsew signal output
flabel metal2 s 69994 88000 70050 88800 0 FreeSans 224 90 0 0 io_north_out[18]
port 109 nsew signal output
flabel metal2 s 71282 88000 71338 88800 0 FreeSans 224 90 0 0 io_north_out[19]
port 110 nsew signal output
flabel metal2 s 31354 88000 31410 88800 0 FreeSans 224 90 0 0 io_north_out[1]
port 111 nsew signal output
flabel metal2 s 72570 88000 72626 88800 0 FreeSans 224 90 0 0 io_north_out[20]
port 112 nsew signal output
flabel metal2 s 73214 88000 73270 88800 0 FreeSans 224 90 0 0 io_north_out[21]
port 113 nsew signal output
flabel metal2 s 74502 88000 74558 88800 0 FreeSans 224 90 0 0 io_north_out[22]
port 114 nsew signal output
flabel metal2 s 75790 88000 75846 88800 0 FreeSans 224 90 0 0 io_north_out[23]
port 115 nsew signal output
flabel metal2 s 76434 88000 76490 88800 0 FreeSans 224 90 0 0 io_north_out[24]
port 116 nsew signal output
flabel metal2 s 77722 88000 77778 88800 0 FreeSans 224 90 0 0 io_north_out[25]
port 117 nsew signal output
flabel metal2 s 79010 88000 79066 88800 0 FreeSans 224 90 0 0 io_north_out[26]
port 118 nsew signal output
flabel metal2 s 80298 88000 80354 88800 0 FreeSans 224 90 0 0 io_north_out[27]
port 119 nsew signal output
flabel metal2 s 80942 88000 80998 88800 0 FreeSans 224 90 0 0 io_north_out[28]
port 120 nsew signal output
flabel metal2 s 82230 88000 82286 88800 0 FreeSans 224 90 0 0 io_north_out[29]
port 121 nsew signal output
flabel metal2 s 32642 88000 32698 88800 0 FreeSans 224 90 0 0 io_north_out[2]
port 122 nsew signal output
flabel metal3 s 89200 44488 90000 44608 0 FreeSans 480 0 0 0 io_north_out[30]
port 123 nsew signal output
flabel metal2 s 42946 88000 43002 88800 0 FreeSans 224 90 0 0 io_north_out[31]
port 124 nsew signal output
flabel metal2 s 33930 88000 33986 88800 0 FreeSans 224 90 0 0 io_north_out[3]
port 125 nsew signal output
flabel metal2 s 34574 88000 34630 88800 0 FreeSans 224 90 0 0 io_north_out[4]
port 126 nsew signal output
flabel metal2 s 35862 88000 35918 88800 0 FreeSans 224 90 0 0 io_north_out[5]
port 127 nsew signal output
flabel metal2 s 37150 88000 37206 88800 0 FreeSans 224 90 0 0 io_north_out[6]
port 128 nsew signal output
flabel metal2 s 38438 88000 38494 88800 0 FreeSans 224 90 0 0 io_north_out[7]
port 129 nsew signal output
flabel metal2 s 39082 88000 39138 88800 0 FreeSans 224 90 0 0 io_north_out[8]
port 130 nsew signal output
flabel metal2 s 40370 88000 40426 88800 0 FreeSans 224 90 0 0 io_north_out[9]
port 131 nsew signal output
flabel metal2 s 30710 3000 30766 3800 0 FreeSans 224 90 0 0 io_south_in[0]
port 132 nsew signal input
flabel metal2 s 41658 3000 41714 3800 0 FreeSans 224 90 0 0 io_south_in[10]
port 133 nsew signal input
flabel metal2 s 42302 3000 42358 3800 0 FreeSans 224 90 0 0 io_south_in[11]
port 134 nsew signal input
flabel metal2 s 43590 3000 43646 3800 0 FreeSans 224 90 0 0 io_south_in[12]
port 135 nsew signal input
flabel metal2 s 44878 3000 44934 3800 0 FreeSans 224 90 0 0 io_south_in[13]
port 136 nsew signal input
flabel metal2 s 8170 3000 8226 3800 0 FreeSans 224 90 0 0 io_south_in[14]
port 137 nsew signal input
flabel metal2 s 8814 3000 8870 3800 0 FreeSans 224 90 0 0 io_south_in[15]
port 138 nsew signal input
flabel metal2 s 68062 3000 68118 3800 0 FreeSans 224 90 0 0 io_south_in[16]
port 139 nsew signal input
flabel metal2 s 68706 3000 68762 3800 0 FreeSans 224 90 0 0 io_south_in[17]
port 140 nsew signal input
flabel metal2 s 69994 3000 70050 3800 0 FreeSans 224 90 0 0 io_south_in[18]
port 141 nsew signal input
flabel metal2 s 71282 3000 71338 3800 0 FreeSans 224 90 0 0 io_south_in[19]
port 142 nsew signal input
flabel metal2 s 31354 3000 31410 3800 0 FreeSans 224 90 0 0 io_south_in[1]
port 143 nsew signal input
flabel metal2 s 72570 3000 72626 3800 0 FreeSans 224 90 0 0 io_south_in[20]
port 144 nsew signal input
flabel metal2 s 73214 3000 73270 3800 0 FreeSans 224 90 0 0 io_south_in[21]
port 145 nsew signal input
flabel metal2 s 74502 3000 74558 3800 0 FreeSans 224 90 0 0 io_south_in[22]
port 146 nsew signal input
flabel metal2 s 75790 3000 75846 3800 0 FreeSans 224 90 0 0 io_south_in[23]
port 147 nsew signal input
flabel metal2 s 76434 3000 76490 3800 0 FreeSans 224 90 0 0 io_south_in[24]
port 148 nsew signal input
flabel metal2 s 77722 3000 77778 3800 0 FreeSans 224 90 0 0 io_south_in[25]
port 149 nsew signal input
flabel metal2 s 79010 3000 79066 3800 0 FreeSans 224 90 0 0 io_south_in[26]
port 150 nsew signal input
flabel metal2 s 80298 3000 80354 3800 0 FreeSans 224 90 0 0 io_south_in[27]
port 151 nsew signal input
flabel metal2 s 80942 3000 80998 3800 0 FreeSans 224 90 0 0 io_south_in[28]
port 152 nsew signal input
flabel metal3 s 89200 10488 90000 10608 0 FreeSans 480 0 0 0 io_south_in[29]
port 153 nsew signal input
flabel metal2 s 32642 3000 32698 3800 0 FreeSans 224 90 0 0 io_south_in[2]
port 154 nsew signal input
flabel metal2 s 9458 3000 9514 3800 0 FreeSans 224 90 0 0 io_south_in[30]
port 155 nsew signal input
flabel metal2 s 10102 3000 10158 3800 0 FreeSans 224 90 0 0 io_south_in[31]
port 156 nsew signal input
flabel metal2 s 33930 3000 33986 3800 0 FreeSans 224 90 0 0 io_south_in[3]
port 157 nsew signal input
flabel metal2 s 34574 3000 34630 3800 0 FreeSans 224 90 0 0 io_south_in[4]
port 158 nsew signal input
flabel metal2 s 35862 3000 35918 3800 0 FreeSans 224 90 0 0 io_south_in[5]
port 159 nsew signal input
flabel metal2 s 37150 3000 37206 3800 0 FreeSans 224 90 0 0 io_south_in[6]
port 160 nsew signal input
flabel metal2 s 38438 3000 38494 3800 0 FreeSans 224 90 0 0 io_south_in[7]
port 161 nsew signal input
flabel metal2 s 39082 3000 39138 3800 0 FreeSans 224 90 0 0 io_south_in[8]
port 162 nsew signal input
flabel metal2 s 40370 3000 40426 3800 0 FreeSans 224 90 0 0 io_south_in[9]
port 163 nsew signal input
flabel metal2 s 15254 3000 15310 3800 0 FreeSans 224 90 0 0 io_south_out[0]
port 164 nsew signal output
flabel metal2 s 26202 3000 26258 3800 0 FreeSans 224 90 0 0 io_south_out[10]
port 165 nsew signal output
flabel metal2 s 26846 3000 26902 3800 0 FreeSans 224 90 0 0 io_south_out[11]
port 166 nsew signal output
flabel metal2 s 28134 3000 28190 3800 0 FreeSans 224 90 0 0 io_south_out[12]
port 167 nsew signal output
flabel metal2 s 29422 3000 29478 3800 0 FreeSans 224 90 0 0 io_south_out[13]
port 168 nsew signal output
flabel metal2 s 44878 88000 44934 88800 0 FreeSans 224 90 0 0 io_south_out[14]
port 169 nsew signal output
flabel metal2 s 49386 88000 49442 88800 0 FreeSans 224 90 0 0 io_south_out[15]
port 170 nsew signal output
flabel metal2 s 52606 3000 52662 3800 0 FreeSans 224 90 0 0 io_south_out[16]
port 171 nsew signal output
flabel metal2 s 53250 3000 53306 3800 0 FreeSans 224 90 0 0 io_south_out[17]
port 172 nsew signal output
flabel metal2 s 54538 3000 54594 3800 0 FreeSans 224 90 0 0 io_south_out[18]
port 173 nsew signal output
flabel metal2 s 55826 3000 55882 3800 0 FreeSans 224 90 0 0 io_south_out[19]
port 174 nsew signal output
flabel metal2 s 15898 3000 15954 3800 0 FreeSans 224 90 0 0 io_south_out[1]
port 175 nsew signal output
flabel metal2 s 57114 3000 57170 3800 0 FreeSans 224 90 0 0 io_south_out[20]
port 176 nsew signal output
flabel metal2 s 57758 3000 57814 3800 0 FreeSans 224 90 0 0 io_south_out[21]
port 177 nsew signal output
flabel metal2 s 59046 3000 59102 3800 0 FreeSans 224 90 0 0 io_south_out[22]
port 178 nsew signal output
flabel metal2 s 60334 3000 60390 3800 0 FreeSans 224 90 0 0 io_south_out[23]
port 179 nsew signal output
flabel metal2 s 60978 3000 61034 3800 0 FreeSans 224 90 0 0 io_south_out[24]
port 180 nsew signal output
flabel metal2 s 62266 3000 62322 3800 0 FreeSans 224 90 0 0 io_south_out[25]
port 181 nsew signal output
flabel metal2 s 63554 3000 63610 3800 0 FreeSans 224 90 0 0 io_south_out[26]
port 182 nsew signal output
flabel metal2 s 64842 3000 64898 3800 0 FreeSans 224 90 0 0 io_south_out[27]
port 183 nsew signal output
flabel metal2 s 65486 3000 65542 3800 0 FreeSans 224 90 0 0 io_south_out[28]
port 184 nsew signal output
flabel metal2 s 66774 3000 66830 3800 0 FreeSans 224 90 0 0 io_south_out[29]
port 185 nsew signal output
flabel metal2 s 17186 3000 17242 3800 0 FreeSans 224 90 0 0 io_south_out[2]
port 186 nsew signal output
flabel metal3 s 89200 45168 90000 45288 0 FreeSans 480 0 0 0 io_south_out[30]
port 187 nsew signal output
flabel metal3 s 89200 46528 90000 46648 0 FreeSans 480 0 0 0 io_south_out[31]
port 188 nsew signal output
flabel metal2 s 18474 3000 18530 3800 0 FreeSans 224 90 0 0 io_south_out[3]
port 189 nsew signal output
flabel metal2 s 19118 3000 19174 3800 0 FreeSans 224 90 0 0 io_south_out[4]
port 190 nsew signal output
flabel metal2 s 20406 3000 20462 3800 0 FreeSans 224 90 0 0 io_south_out[5]
port 191 nsew signal output
flabel metal2 s 21694 3000 21750 3800 0 FreeSans 224 90 0 0 io_south_out[6]
port 192 nsew signal output
flabel metal2 s 22982 3000 23038 3800 0 FreeSans 224 90 0 0 io_south_out[7]
port 193 nsew signal output
flabel metal2 s 23626 3000 23682 3800 0 FreeSans 224 90 0 0 io_south_out[8]
port 194 nsew signal output
flabel metal2 s 24914 3000 24970 3800 0 FreeSans 224 90 0 0 io_south_out[9]
port 195 nsew signal output
flabel metal3 s 3000 15248 3800 15368 0 FreeSans 480 0 0 0 io_west_in[0]
port 196 nsew signal input
flabel metal3 s 3000 26128 3800 26248 0 FreeSans 480 0 0 0 io_west_in[10]
port 197 nsew signal input
flabel metal3 s 3000 26808 3800 26928 0 FreeSans 480 0 0 0 io_west_in[11]
port 198 nsew signal input
flabel metal3 s 3000 28168 3800 28288 0 FreeSans 480 0 0 0 io_west_in[12]
port 199 nsew signal input
flabel metal3 s 3000 29528 3800 29648 0 FreeSans 480 0 0 0 io_west_in[13]
port 200 nsew signal input
flabel metal2 s 10746 3000 10802 3800 0 FreeSans 224 90 0 0 io_west_in[14]
port 201 nsew signal input
flabel metal2 s 11390 3000 11446 3800 0 FreeSans 224 90 0 0 io_west_in[15]
port 202 nsew signal input
flabel metal3 s 3000 51288 3800 51408 0 FreeSans 480 0 0 0 io_west_in[16]
port 203 nsew signal input
flabel metal3 s 3000 52648 3800 52768 0 FreeSans 480 0 0 0 io_west_in[17]
port 204 nsew signal input
flabel metal3 s 3000 54008 3800 54128 0 FreeSans 480 0 0 0 io_west_in[18]
port 205 nsew signal input
flabel metal3 s 3000 54688 3800 54808 0 FreeSans 480 0 0 0 io_west_in[19]
port 206 nsew signal input
flabel metal3 s 3000 15928 3800 16048 0 FreeSans 480 0 0 0 io_west_in[1]
port 207 nsew signal input
flabel metal3 s 3000 56048 3800 56168 0 FreeSans 480 0 0 0 io_west_in[20]
port 208 nsew signal input
flabel metal3 s 3000 56728 3800 56848 0 FreeSans 480 0 0 0 io_west_in[21]
port 209 nsew signal input
flabel metal3 s 3000 58088 3800 58208 0 FreeSans 480 0 0 0 io_west_in[22]
port 210 nsew signal input
flabel metal3 s 3000 59448 3800 59568 0 FreeSans 480 0 0 0 io_west_in[23]
port 211 nsew signal input
flabel metal3 s 3000 60128 3800 60248 0 FreeSans 480 0 0 0 io_west_in[24]
port 212 nsew signal input
flabel metal3 s 3000 61488 3800 61608 0 FreeSans 480 0 0 0 io_west_in[25]
port 213 nsew signal input
flabel metal3 s 3000 62168 3800 62288 0 FreeSans 480 0 0 0 io_west_in[26]
port 214 nsew signal input
flabel metal3 s 3000 63528 3800 63648 0 FreeSans 480 0 0 0 io_west_in[27]
port 215 nsew signal input
flabel metal3 s 3000 64888 3800 65008 0 FreeSans 480 0 0 0 io_west_in[28]
port 216 nsew signal input
flabel metal3 s 3000 65568 3800 65688 0 FreeSans 480 0 0 0 io_west_in[29]
port 217 nsew signal input
flabel metal3 s 3000 17288 3800 17408 0 FreeSans 480 0 0 0 io_west_in[2]
port 218 nsew signal input
flabel metal2 s 12034 3000 12090 3800 0 FreeSans 224 90 0 0 io_west_in[30]
port 219 nsew signal input
flabel metal2 s 12678 3000 12734 3800 0 FreeSans 224 90 0 0 io_west_in[31]
port 220 nsew signal input
flabel metal3 s 3000 18648 3800 18768 0 FreeSans 480 0 0 0 io_west_in[3]
port 221 nsew signal input
flabel metal3 s 3000 19328 3800 19448 0 FreeSans 480 0 0 0 io_west_in[4]
port 222 nsew signal input
flabel metal3 s 3000 20688 3800 20808 0 FreeSans 480 0 0 0 io_west_in[5]
port 223 nsew signal input
flabel metal3 s 3000 21368 3800 21488 0 FreeSans 480 0 0 0 io_west_in[6]
port 224 nsew signal input
flabel metal3 s 3000 22728 3800 22848 0 FreeSans 480 0 0 0 io_west_in[7]
port 225 nsew signal input
flabel metal3 s 3000 24088 3800 24208 0 FreeSans 480 0 0 0 io_west_in[8]
port 226 nsew signal input
flabel metal3 s 3000 24768 3800 24888 0 FreeSans 480 0 0 0 io_west_in[9]
port 227 nsew signal input
flabel metal3 s 3000 30208 3800 30328 0 FreeSans 480 0 0 0 io_west_out[0]
port 228 nsew signal output
flabel metal3 s 3000 41088 3800 41208 0 FreeSans 480 0 0 0 io_west_out[10]
port 229 nsew signal output
flabel metal3 s 3000 42448 3800 42568 0 FreeSans 480 0 0 0 io_west_out[11]
port 230 nsew signal output
flabel metal3 s 3000 43128 3800 43248 0 FreeSans 480 0 0 0 io_west_out[12]
port 231 nsew signal output
flabel metal3 s 3000 44488 3800 44608 0 FreeSans 480 0 0 0 io_west_out[13]
port 232 nsew signal output
flabel metal2 s 45522 88000 45578 88800 0 FreeSans 224 90 0 0 io_west_out[14]
port 233 nsew signal output
flabel metal3 s 89200 48568 90000 48688 0 FreeSans 480 0 0 0 io_west_out[15]
port 234 nsew signal output
flabel metal3 s 3000 66928 3800 67048 0 FreeSans 480 0 0 0 io_west_out[16]
port 235 nsew signal output
flabel metal3 s 3000 67608 3800 67728 0 FreeSans 480 0 0 0 io_west_out[17]
port 236 nsew signal output
flabel metal3 s 3000 68968 3800 69088 0 FreeSans 480 0 0 0 io_west_out[18]
port 237 nsew signal output
flabel metal3 s 3000 70328 3800 70448 0 FreeSans 480 0 0 0 io_west_out[19]
port 238 nsew signal output
flabel metal3 s 3000 31568 3800 31688 0 FreeSans 480 0 0 0 io_west_out[1]
port 239 nsew signal output
flabel metal3 s 3000 71008 3800 71128 0 FreeSans 480 0 0 0 io_west_out[20]
port 240 nsew signal output
flabel metal3 s 3000 72368 3800 72488 0 FreeSans 480 0 0 0 io_west_out[21]
port 241 nsew signal output
flabel metal3 s 3000 73048 3800 73168 0 FreeSans 480 0 0 0 io_west_out[22]
port 242 nsew signal output
flabel metal3 s 3000 74408 3800 74528 0 FreeSans 480 0 0 0 io_west_out[23]
port 243 nsew signal output
flabel metal3 s 3000 75768 3800 75888 0 FreeSans 480 0 0 0 io_west_out[24]
port 244 nsew signal output
flabel metal3 s 3000 76448 3800 76568 0 FreeSans 480 0 0 0 io_west_out[25]
port 245 nsew signal output
flabel metal3 s 3000 77808 3800 77928 0 FreeSans 480 0 0 0 io_west_out[26]
port 246 nsew signal output
flabel metal3 s 3000 78488 3800 78608 0 FreeSans 480 0 0 0 io_west_out[27]
port 247 nsew signal output
flabel metal3 s 3000 79848 3800 79968 0 FreeSans 480 0 0 0 io_west_out[28]
port 248 nsew signal output
flabel metal3 s 3000 81208 3800 81328 0 FreeSans 480 0 0 0 io_west_out[29]
port 249 nsew signal output
flabel metal3 s 3000 32248 3800 32368 0 FreeSans 480 0 0 0 io_west_out[2]
port 250 nsew signal output
flabel metal2 s 46810 88000 46866 88800 0 FreeSans 224 90 0 0 io_west_out[30]
port 251 nsew signal output
flabel metal2 s 48098 88000 48154 88800 0 FreeSans 224 90 0 0 io_west_out[31]
port 252 nsew signal output
flabel metal3 s 3000 33608 3800 33728 0 FreeSans 480 0 0 0 io_west_out[3]
port 253 nsew signal output
flabel metal3 s 3000 34968 3800 35088 0 FreeSans 480 0 0 0 io_west_out[4]
port 254 nsew signal output
flabel metal3 s 3000 35648 3800 35768 0 FreeSans 480 0 0 0 io_west_out[5]
port 255 nsew signal output
flabel metal3 s 3000 37008 3800 37128 0 FreeSans 480 0 0 0 io_west_out[6]
port 256 nsew signal output
flabel metal3 s 3000 37688 3800 37808 0 FreeSans 480 0 0 0 io_west_out[7]
port 257 nsew signal output
flabel metal3 s 3000 39048 3800 39168 0 FreeSans 480 0 0 0 io_west_out[8]
port 258 nsew signal output
flabel metal3 s 3000 40408 3800 40528 0 FreeSans 480 0 0 0 io_west_out[9]
port 259 nsew signal output
flabel metal3 s 89200 12528 90000 12648 0 FreeSans 480 0 0 0 le_clk
port 260 nsew signal input
flabel metal3 s 89200 13208 90000 13328 0 FreeSans 480 0 0 0 le_en
port 261 nsew signal input
flabel metal3 s 89200 14568 90000 14688 0 FreeSans 480 0 0 0 le_nrst
port 262 nsew signal input
flabel metal2 s 37794 88000 37850 88800 0 FreeSans 224 90 0 0 nrst
port 263 nsew signal input
flabel metal4 s 3356 3376 3676 89104 0 FreeSans 1920 90 0 0 vccd1
port 264 nsew power bidirectional
flabel metal5 s 3356 3376 90116 3696 0 FreeSans 2560 0 0 0 vccd1
port 264 nsew power bidirectional
flabel metal5 s 3356 88784 90116 89104 0 FreeSans 2560 0 0 0 vccd1
port 264 nsew power bidirectional
flabel metal4 s 89796 3376 90116 89104 0 FreeSans 1920 90 0 0 vccd1
port 264 nsew power bidirectional
flabel metal4 s 17716 2716 18036 10187 0 FreeSans 1920 90 0 0 vccd1
port 264 nsew power bidirectional
flabel metal4 s 17716 81029 18036 89764 0 FreeSans 1920 90 0 0 vccd1
port 264 nsew power bidirectional
flabel metal4 s 36116 2716 36436 10187 0 FreeSans 1920 90 0 0 vccd1
port 264 nsew power bidirectional
flabel metal4 s 36116 81029 36436 89764 0 FreeSans 1920 90 0 0 vccd1
port 264 nsew power bidirectional
flabel metal4 s 54516 2716 54836 10187 0 FreeSans 1920 90 0 0 vccd1
port 264 nsew power bidirectional
flabel metal4 s 54516 81029 54836 89764 0 FreeSans 1920 90 0 0 vccd1
port 264 nsew power bidirectional
flabel metal4 s 72916 2716 73236 10187 0 FreeSans 1920 90 0 0 vccd1
port 264 nsew power bidirectional
flabel metal4 s 72916 81029 73236 89764 0 FreeSans 1920 90 0 0 vccd1
port 264 nsew power bidirectional
flabel metal5 s 2696 17736 90776 18056 0 FreeSans 2560 0 0 0 vccd1
port 264 nsew power bidirectional
flabel metal5 s 2696 36136 90776 36456 0 FreeSans 2560 0 0 0 vccd1
port 264 nsew power bidirectional
flabel metal5 s 2696 54536 90776 54856 0 FreeSans 2560 0 0 0 vccd1
port 264 nsew power bidirectional
flabel metal5 s 2696 72936 90776 73256 0 FreeSans 2560 0 0 0 vccd1
port 264 nsew power bidirectional
flabel metal4 s 5876 7024 6196 84912 0 FreeSans 1920 90 0 0 vccd1
port 264 nsew power bidirectional
flabel metal4 s 86468 7024 86788 84912 0 FreeSans 1920 90 0 0 vccd1
port 264 nsew power bidirectional
flabel metal4 s 2696 2716 3016 89764 0 FreeSans 1920 90 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal5 s 2696 2716 90776 3036 0 FreeSans 2560 0 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal5 s 2696 89444 90776 89764 0 FreeSans 2560 0 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal4 s 90456 2716 90776 89764 0 FreeSans 1920 90 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal4 s 18376 2716 18696 10187 0 FreeSans 1920 90 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal4 s 18376 81029 18696 89764 0 FreeSans 1920 90 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal4 s 36776 2716 37096 10187 0 FreeSans 1920 90 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal4 s 36776 81029 37096 89764 0 FreeSans 1920 90 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal4 s 55176 2716 55496 10187 0 FreeSans 1920 90 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal4 s 55176 81029 55496 89764 0 FreeSans 1920 90 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal4 s 73576 2716 73896 10187 0 FreeSans 1920 90 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal4 s 73576 81029 73896 89764 0 FreeSans 1920 90 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal5 s 2696 18396 90776 18716 0 FreeSans 2560 0 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal5 s 2696 36796 90776 37116 0 FreeSans 2560 0 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal5 s 2696 55196 90776 55516 0 FreeSans 2560 0 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal5 s 2696 73596 90776 73916 0 FreeSans 2560 0 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal4 s 6612 7024 6932 84912 0 FreeSans 1920 90 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal4 s 87204 7024 87524 84912 0 FreeSans 1920 90 0 0 vssd1
port 265 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 3000 3000 90000 88800
<< end >>
