magic
tech sky130A
magscale 1 2
timestamp 1752714626
<< viali >>
rect 10892 87433 10926 87467
rect 15061 87433 15095 87467
rect 16993 87433 17027 87467
rect 18281 87433 18315 87467
rect 19569 87433 19603 87467
rect 21501 87433 21535 87467
rect 22789 87433 22823 87467
rect 23433 87433 23467 87467
rect 24721 87433 24755 87467
rect 26009 87433 26043 87467
rect 27297 87433 27331 87467
rect 29229 87433 29263 87467
rect 30948 87433 30982 87467
rect 31391 87433 31425 87467
rect 32788 87433 32822 87467
rect 34076 87433 34110 87467
rect 35364 87433 35398 87467
rect 36100 87433 36134 87467
rect 37296 87433 37330 87467
rect 37877 87433 37911 87467
rect 38225 87433 38259 87467
rect 39688 87433 39722 87467
rect 40516 87433 40550 87467
rect 40821 87433 40855 87467
rect 42339 87433 42373 87467
rect 43828 87433 43862 87467
rect 44271 87433 44305 87467
rect 52413 87433 52447 87467
rect 55633 87433 55667 87467
rect 56921 87433 56955 87467
rect 57565 87433 57599 87467
rect 60141 87433 60175 87467
rect 63361 87433 63395 87467
rect 64649 87433 64683 87467
rect 65293 87433 65327 87467
rect 68208 87433 68242 87467
rect 69588 87433 69622 87467
rect 70031 87433 70065 87467
rect 71428 87433 71462 87467
rect 72716 87433 72750 87467
rect 73251 87433 73285 87467
rect 74740 87433 74774 87467
rect 75936 87433 75970 87467
rect 77316 87433 77350 87467
rect 77759 87433 77793 87467
rect 79156 87433 79190 87467
rect 80444 87433 80478 87467
rect 80979 87433 81013 87467
rect 82468 87433 82502 87467
rect 10737 87331 10771 87365
rect 16395 87353 16429 87387
rect 16533 87365 16567 87399
rect 17177 87331 17211 87365
rect 18587 87333 18621 87367
rect 19875 87333 19909 87367
rect 20613 87333 20647 87367
rect 20765 87365 20799 87399
rect 21823 87353 21857 87387
rect 23203 87353 23237 87387
rect 23617 87331 23651 87365
rect 24905 87331 24939 87365
rect 26331 87353 26365 87387
rect 27619 87353 27653 87387
rect 28341 87333 28375 87367
rect 28493 87365 28527 87399
rect 29551 87353 29585 87387
rect 38473 87365 38507 87399
rect 41049 87365 41083 87399
rect 42937 87365 42971 87399
rect 44869 87365 44903 87399
rect 45513 87365 45547 87399
rect 46249 87365 46283 87399
rect 46801 87365 46835 87399
rect 47445 87365 47479 87399
rect 48089 87365 48123 87399
rect 48825 87365 48859 87399
rect 49377 87365 49411 87399
rect 50021 87365 50055 87399
rect 50665 87365 50699 87399
rect 30745 87331 30779 87365
rect 31560 87331 31594 87365
rect 32633 87331 32667 87365
rect 33873 87331 33907 87365
rect 35161 87331 35195 87365
rect 35945 87331 35979 87365
rect 37141 87331 37175 87365
rect 38061 87331 38095 87365
rect 39485 87331 39519 87365
rect 40361 87331 40395 87365
rect 42545 87331 42579 87365
rect 43673 87331 43707 87365
rect 44477 87331 44511 87365
rect 54099 87333 54133 87367
rect 54253 87365 54287 87399
rect 54805 87365 54839 87399
rect 54529 87331 54563 87365
rect 55955 87353 55989 87387
rect 57243 87353 57277 87387
rect 57749 87331 57783 87365
rect 59251 87333 59285 87367
rect 59405 87365 59439 87399
rect 60447 87333 60481 87367
rect 61829 87333 61863 87367
rect 61981 87365 62015 87399
rect 62533 87365 62567 87399
rect 62257 87331 62291 87365
rect 63683 87353 63717 87387
rect 64971 87353 65005 87387
rect 65477 87331 65511 87365
rect 66979 87333 67013 87367
rect 67133 87365 67167 87399
rect 68005 87331 68039 87365
rect 69433 87331 69467 87365
rect 70200 87331 70234 87365
rect 71273 87331 71307 87365
rect 72513 87331 72547 87365
rect 73420 87331 73454 87365
rect 74585 87331 74619 87365
rect 75733 87331 75767 87365
rect 77150 87331 77184 87365
rect 77928 87331 77962 87365
rect 79001 87331 79035 87365
rect 80289 87331 80323 87365
rect 81148 87331 81182 87365
rect 82313 87331 82347 87365
rect 15337 87297 15371 87331
rect 18419 87297 18453 87331
rect 19707 87297 19741 87331
rect 52597 87297 52631 87331
rect 60279 87297 60313 87331
rect 23019 87229 23053 87263
rect 27435 87229 27469 87263
rect 39073 87229 39107 87263
rect 39901 87229 39935 87263
rect 57059 87229 57093 87263
rect 62395 87229 62429 87263
rect 64787 87229 64821 87263
rect 15521 87161 15555 87195
rect 16211 87161 16245 87195
rect 17327 87161 17361 87195
rect 20443 87161 20477 87195
rect 21639 87161 21673 87195
rect 23777 87161 23811 87195
rect 25064 87161 25098 87195
rect 26147 87161 26181 87195
rect 28171 87161 28205 87195
rect 29367 87161 29401 87195
rect 41833 87161 41867 87195
rect 42109 87161 42143 87195
rect 52781 87161 52815 87195
rect 53931 87161 53965 87195
rect 54679 87161 54713 87195
rect 55771 87161 55805 87195
rect 57909 87161 57943 87195
rect 59083 87161 59117 87195
rect 61659 87161 61693 87195
rect 63499 87161 63533 87195
rect 65637 87161 65671 87195
rect 66811 87161 66845 87195
rect 41804 86889 41838 86923
rect 41603 86719 41637 86753
rect 31069 84713 31103 84747
rect 45421 84713 45455 84747
rect 12853 84645 12887 84679
rect 11749 84577 11783 84611
rect 45605 84577 45639 84611
rect 51401 84577 51435 84611
rect 30585 84509 30619 84543
rect 30885 84509 30919 84543
rect 41049 84509 41083 84543
rect 42753 84509 42787 84543
rect 42937 84509 42971 84543
rect 48089 84509 48123 84543
rect 10645 84441 10679 84475
rect 13957 84441 13991 84475
rect 29965 84441 29999 84475
rect 40821 84441 40855 84475
rect 45789 84441 45823 84475
rect 45973 84441 46007 84475
rect 49193 84441 49227 84475
rect 50297 84441 50331 84475
rect 88063 81381 88097 81415
rect 88265 81279 88299 81313
rect 87741 81245 87775 81279
rect 87741 80225 87775 80259
rect 5469 80191 5503 80225
rect 88265 80191 88299 80225
rect 5263 80089 5297 80123
rect 88063 80089 88097 80123
rect 5469 78627 5503 78661
rect 88265 78627 88299 78661
rect 87925 78593 87959 78627
rect 88063 78525 88097 78559
rect 5263 78457 5297 78491
rect 5469 78015 5503 78049
rect 88265 78015 88299 78049
rect 87741 77981 87775 78015
rect 5263 77913 5297 77947
rect 88063 77913 88097 77947
rect 87809 76961 87843 76995
rect 5469 76927 5503 76961
rect 5263 76825 5297 76859
rect 87557 76825 87591 76859
rect 88017 76825 88051 76859
rect 88063 75941 88097 75975
rect 87741 75873 87775 75907
rect 5469 75839 5503 75873
rect 88269 75839 88303 75873
rect 5263 75737 5297 75771
rect 5263 74853 5297 74887
rect 88063 74853 88097 74887
rect 87741 74785 87775 74819
rect 5469 74751 5503 74785
rect 88269 74751 88303 74785
rect 5469 73187 5503 73221
rect 88265 73187 88299 73221
rect 88063 73153 88097 73187
rect 87925 73085 87959 73119
rect 5263 73017 5297 73051
rect 5469 72575 5503 72609
rect 88063 72541 88097 72575
rect 88265 72569 88299 72603
rect 5263 72473 5297 72507
rect 87741 72473 87775 72507
rect 88063 71589 88097 71623
rect 5469 71487 5503 71521
rect 88265 71487 88299 71521
rect 87741 71453 87775 71487
rect 5263 71385 5297 71419
rect 88063 70501 88097 70535
rect 87741 70433 87775 70467
rect 5469 70399 5503 70433
rect 88233 70399 88267 70433
rect 5263 70297 5297 70331
rect 5469 69311 5503 69345
rect 88063 69277 88097 69311
rect 88265 69305 88299 69339
rect 5263 69209 5297 69243
rect 87741 69209 87775 69243
rect 87925 67781 87959 67815
rect 5469 67747 5503 67781
rect 88265 67747 88299 67781
rect 88063 67645 88097 67679
rect 5263 67577 5297 67611
rect 5469 67135 5503 67169
rect 88063 67101 88097 67135
rect 88265 67129 88299 67163
rect 5263 67033 5297 67067
rect 87741 67033 87775 67067
rect 5217 66047 5251 66081
rect 87969 66047 88003 66081
rect 5377 66013 5411 66047
rect 5493 65945 5527 65979
rect 88181 65945 88215 65979
rect 5217 64959 5251 64993
rect 87969 64959 88003 64993
rect 5377 64925 5411 64959
rect 5493 64857 5527 64891
rect 88181 64857 88215 64891
rect 7517 64585 7551 64619
rect 5377 63905 5411 63939
rect 5217 63871 5251 63905
rect 87969 63871 88003 63905
rect 5493 63837 5527 63871
rect 7401 63837 7435 63871
rect 6781 63769 6815 63803
rect 88181 63769 88215 63803
rect 7517 63225 7551 63259
rect 5377 62409 5411 62443
rect 88181 62341 88215 62375
rect 5171 62307 5205 62341
rect 87969 62307 88003 62341
rect 5493 62273 5527 62307
rect 5217 61695 5251 61729
rect 87969 61695 88003 61729
rect 5376 61661 5410 61695
rect 5493 61593 5527 61627
rect 88181 61593 88215 61627
rect 5217 60607 5251 60641
rect 87969 60607 88003 60641
rect 5376 60573 5410 60607
rect 5493 60505 5527 60539
rect 88181 60505 88215 60539
rect 5217 59519 5251 59553
rect 87969 59519 88003 59553
rect 5377 59485 5411 59519
rect 5493 59417 5527 59451
rect 88181 59417 88215 59451
rect 5217 58431 5251 58465
rect 88017 58431 88051 58465
rect 5493 58397 5527 58431
rect 5376 58329 5410 58363
rect 88181 58329 88215 58363
rect 5377 56969 5411 57003
rect 5171 56867 5205 56901
rect 88017 56867 88051 56901
rect 5493 56833 5527 56867
rect 88181 56833 88215 56867
rect 5493 56289 5527 56323
rect 5171 56255 5205 56289
rect 87969 56255 88003 56289
rect 5377 56221 5411 56255
rect 88181 56153 88215 56187
rect 5493 55201 5527 55235
rect 5171 55167 5205 55201
rect 87969 55167 88003 55201
rect 5377 55133 5411 55167
rect 88181 55065 88215 55099
rect 5493 54113 5527 54147
rect 5171 54079 5205 54113
rect 87969 54079 88003 54113
rect 5377 54045 5411 54079
rect 88181 54045 88215 54079
rect 5493 53025 5527 53059
rect 5171 52991 5205 53025
rect 87969 52991 88003 53025
rect 5377 52957 5411 52991
rect 88181 52889 88215 52923
rect 5377 51529 5411 51563
rect 5171 51427 5205 51461
rect 87969 51427 88003 51461
rect 5493 51393 5527 51427
rect 88181 51325 88215 51359
rect 85625 50713 85659 50747
rect 85625 49625 85659 49659
rect 88201 48605 88235 48639
rect 85625 48537 85659 48571
rect 88201 47993 88235 48027
rect 87969 47551 88003 47585
rect 88181 47449 88215 47483
rect 88201 46905 88235 46939
rect 88201 45817 88235 45851
rect 5376 45545 5410 45579
rect 7333 45545 7367 45579
rect 85809 45545 85843 45579
rect 7149 45477 7183 45511
rect 85993 45477 86027 45511
rect 5171 45375 5205 45409
rect 5493 45341 5527 45375
rect 86177 45341 86211 45375
rect 88201 45341 88235 45375
rect 85625 45273 85659 45307
rect 7517 45001 7551 45035
rect 5469 44899 5503 44933
rect 88265 44899 88299 44933
rect 87925 44865 87959 44899
rect 88063 44797 88097 44831
rect 5263 44729 5297 44763
rect 87741 44389 87775 44423
rect 5469 44287 5503 44321
rect 88265 44281 88299 44315
rect 5263 44185 5297 44219
rect 88063 44185 88097 44219
rect 5469 42723 5503 42757
rect 88265 42723 88299 42757
rect 87925 42689 87959 42723
rect 88063 42621 88097 42655
rect 5263 42553 5297 42587
rect 5263 41737 5297 41771
rect 88063 41737 88097 41771
rect 5469 41635 5503 41669
rect 88265 41635 88299 41669
rect 87925 41601 87959 41635
rect 5469 40547 5503 40581
rect 87925 40513 87959 40547
rect 88269 40513 88303 40547
rect 5263 40377 5297 40411
rect 88201 40105 88235 40139
rect 5469 39459 5503 39493
rect 88269 39459 88303 39493
rect 87833 39425 87867 39459
rect 88063 39357 88097 39391
rect 5263 39289 5297 39323
rect 5263 38949 5297 38983
rect 88063 38949 88097 38983
rect 5469 38847 5503 38881
rect 88269 38847 88303 38881
rect 87741 38813 87775 38847
rect 5469 37283 5503 37317
rect 88265 37283 88299 37317
rect 87925 37249 87959 37283
rect 88063 37181 88097 37215
rect 5263 37113 5297 37147
rect 5469 36195 5503 36229
rect 88265 36195 88299 36229
rect 87925 36161 87959 36195
rect 5263 36093 5297 36127
rect 88063 36093 88097 36127
rect 5469 35107 5503 35141
rect 88265 35107 88299 35141
rect 87925 35073 87959 35107
rect 88063 35005 88097 35039
rect 5263 34937 5297 34971
rect 87925 34121 87959 34155
rect 5469 34019 5503 34053
rect 88265 34019 88299 34053
rect 88063 33917 88097 33951
rect 5263 33849 5297 33883
rect 5263 33509 5297 33543
rect 87741 33509 87775 33543
rect 5469 33407 5503 33441
rect 88063 33373 88097 33407
rect 88265 33401 88299 33435
rect 5469 31843 5503 31877
rect 88265 31843 88299 31877
rect 87925 31809 87959 31843
rect 88063 31741 88097 31775
rect 5263 31673 5297 31707
rect 5469 30755 5503 30789
rect 88265 30755 88299 30789
rect 87925 30721 87959 30755
rect 88063 30653 88097 30687
rect 5263 30585 5297 30619
rect 5171 29667 5205 29701
rect 87969 29667 88003 29701
rect 5493 29633 5527 29667
rect 5377 29565 5411 29599
rect 88181 29497 88215 29531
rect 5171 28579 5205 28613
rect 87969 28579 88003 28613
rect 5493 28545 5527 28579
rect 5377 28477 5411 28511
rect 88181 28409 88215 28443
rect 5493 28069 5527 28103
rect 5217 27967 5251 28001
rect 87969 27967 88003 28001
rect 5377 27865 5411 27899
rect 88181 27865 88215 27899
rect 5171 26403 5205 26437
rect 87969 26403 88003 26437
rect 5493 26369 5527 26403
rect 5377 26301 5411 26335
rect 88181 26233 88215 26267
rect 5171 25315 5205 25349
rect 87969 25315 88003 25349
rect 5493 25281 5527 25315
rect 5376 25213 5410 25247
rect 88181 25145 88215 25179
rect 5171 24227 5205 24261
rect 87969 24227 88003 24261
rect 5493 24193 5527 24227
rect 5376 24125 5410 24159
rect 88181 24057 88215 24091
rect 5171 23139 5205 23173
rect 87969 23139 88003 23173
rect 5493 23105 5527 23139
rect 5377 23037 5411 23071
rect 88181 22969 88215 23003
rect 5493 22561 5527 22595
rect 5171 22527 5205 22561
rect 87969 22527 88003 22561
rect 5376 22493 5410 22527
rect 88181 22425 88215 22459
rect 5377 21065 5411 21099
rect 5217 20963 5251 20997
rect 87969 20963 88003 20997
rect 5493 20929 5527 20963
rect 88181 20929 88215 20963
rect 5171 19875 5205 19909
rect 87969 19875 88003 19909
rect 5493 19841 5527 19875
rect 5377 19773 5411 19807
rect 88181 19705 88215 19739
rect 5171 18787 5205 18821
rect 87969 18787 88003 18821
rect 5493 18753 5527 18787
rect 5377 18685 5411 18719
rect 88181 18617 88215 18651
rect 5171 17699 5205 17733
rect 87969 17699 88003 17733
rect 5493 17665 5527 17699
rect 5377 17597 5411 17631
rect 88181 17529 88215 17563
rect 5217 17087 5251 17121
rect 88017 17087 88051 17121
rect 5493 17053 5527 17087
rect 5377 16985 5411 17019
rect 88181 16985 88215 17019
rect 5217 15523 5251 15557
rect 87969 15523 88003 15557
rect 5493 15489 5527 15523
rect 5377 15421 5411 15455
rect 88181 15421 88215 15455
rect 88201 15013 88235 15047
rect 87465 14945 87499 14979
rect 87808 14911 87842 14945
rect 88017 14809 88051 14843
rect 85625 14265 85659 14299
rect 85625 13449 85659 13483
rect 87649 13381 87683 13415
rect 88226 13347 88260 13381
rect 87925 13313 87959 13347
rect 88201 12905 88235 12939
rect 87808 12735 87842 12769
rect 87465 12701 87499 12735
rect 88017 12701 88051 12735
rect 85625 12361 85659 12395
rect 88109 12361 88143 12395
rect 85625 11205 85659 11239
rect 87741 10593 87775 10627
rect 88265 10559 88299 10593
rect 88063 10457 88097 10491
rect 88265 10083 88299 10117
rect 87925 10049 87959 10083
rect 88063 9981 88097 10015
rect 45421 7465 45455 7499
rect 45973 7465 46007 7499
rect 45605 7397 45639 7431
rect 45789 7397 45823 7431
rect 30747 5289 30781 5323
rect 31504 5289 31538 5323
rect 33875 5289 33909 5323
rect 35163 5289 35197 5323
rect 35899 5289 35933 5323
rect 37095 5289 37129 5323
rect 38475 5289 38509 5323
rect 39232 5289 39266 5323
rect 41603 5289 41637 5323
rect 42891 5289 42925 5323
rect 43627 5289 43661 5323
rect 44823 5289 44857 5323
rect 68007 5289 68041 5323
rect 69387 5289 69421 5323
rect 71227 5289 71261 5323
rect 72515 5289 72549 5323
rect 73365 5289 73399 5323
rect 74539 5289 74573 5323
rect 75735 5289 75769 5323
rect 77115 5289 77149 5323
rect 78955 5289 78989 5323
rect 80243 5289 80277 5323
rect 32771 5221 32805 5255
rect 40499 5221 40533 5255
rect 70123 5221 70157 5255
rect 77851 5221 77885 5255
rect 15337 5119 15371 5153
rect 16104 5119 16138 5153
rect 17177 5119 17211 5153
rect 18417 5119 18451 5153
rect 19753 5119 19787 5153
rect 20489 5119 20523 5153
rect 21685 5119 21719 5153
rect 23065 5119 23099 5153
rect 23832 5119 23866 5153
rect 24905 5119 24939 5153
rect 26193 5119 26227 5153
rect 27481 5119 27515 5153
rect 28217 5119 28251 5153
rect 29413 5119 29447 5153
rect 30931 5093 30965 5127
rect 31345 5119 31379 5153
rect 32633 5119 32667 5153
rect 34059 5093 34093 5127
rect 35347 5093 35381 5127
rect 36083 5113 36117 5147
rect 36221 5085 36255 5119
rect 37279 5093 37313 5127
rect 38659 5093 38693 5127
rect 39073 5119 39107 5153
rect 40361 5119 40395 5153
rect 41787 5093 41821 5127
rect 43075 5093 43109 5127
rect 43797 5113 43831 5147
rect 43949 5085 43983 5119
rect 45007 5093 45041 5127
rect 52549 5119 52583 5153
rect 53929 5119 53963 5153
rect 54781 5119 54815 5153
rect 55817 5119 55851 5153
rect 57057 5119 57091 5153
rect 57964 5119 57998 5153
rect 59129 5119 59163 5153
rect 60277 5119 60311 5153
rect 61657 5119 61691 5153
rect 62472 5119 62506 5153
rect 63545 5119 63579 5153
rect 64785 5119 64819 5153
rect 65692 5119 65726 5153
rect 66857 5119 66891 5153
rect 68191 5093 68225 5127
rect 69555 5113 69589 5147
rect 69985 5119 70019 5153
rect 69709 5085 69743 5119
rect 70261 5085 70295 5119
rect 71411 5093 71445 5127
rect 72699 5093 72733 5127
rect 73205 5119 73239 5153
rect 74723 5113 74757 5147
rect 74861 5085 74895 5119
rect 75919 5093 75953 5127
rect 77283 5113 77317 5147
rect 77713 5119 77747 5153
rect 77437 5085 77471 5119
rect 77989 5085 78023 5119
rect 79139 5093 79173 5127
rect 80427 5093 80461 5127
rect 15492 5017 15526 5051
rect 15935 5017 15969 5051
rect 17332 5017 17366 5051
rect 18620 5017 18654 5051
rect 19908 5017 19942 5051
rect 20644 5017 20678 5051
rect 21840 5017 21874 5051
rect 23220 5017 23254 5051
rect 23663 5017 23697 5051
rect 25060 5017 25094 5051
rect 26348 5017 26382 5051
rect 27636 5017 27670 5051
rect 28372 5017 28406 5051
rect 29568 5017 29602 5051
rect 30517 5017 30551 5051
rect 31161 5017 31195 5051
rect 32449 5017 32483 5051
rect 33737 5017 33771 5051
rect 35025 5017 35059 5051
rect 36957 5017 36991 5051
rect 38245 5017 38279 5051
rect 38889 5017 38923 5051
rect 40177 5017 40211 5051
rect 41465 5017 41499 5051
rect 42753 5017 42787 5051
rect 44685 5017 44719 5051
rect 52752 5017 52786 5051
rect 54132 5017 54166 5051
rect 54575 5017 54609 5051
rect 55972 5017 56006 5051
rect 57260 5017 57294 5051
rect 57795 5017 57829 5051
rect 59284 5017 59318 5051
rect 60480 5017 60514 5051
rect 61860 5017 61894 5051
rect 62303 5017 62337 5051
rect 63700 5017 63734 5051
rect 64988 5017 65022 5051
rect 65523 5017 65557 5051
rect 67012 5017 67046 5051
rect 67869 5017 67903 5051
rect 71089 5017 71123 5051
rect 72377 5017 72411 5051
rect 73021 5017 73055 5051
rect 75597 5017 75631 5051
rect 78817 5017 78851 5051
rect 80105 5017 80139 5051
<< metal1 >>
rect 4876 87610 88596 87632
rect 4876 87558 18382 87610
rect 18434 87558 18446 87610
rect 18498 87558 18510 87610
rect 18562 87558 18574 87610
rect 18626 87558 18638 87610
rect 18690 87558 36782 87610
rect 36834 87558 36846 87610
rect 36898 87558 36910 87610
rect 36962 87558 36974 87610
rect 37026 87558 37038 87610
rect 37090 87558 55182 87610
rect 55234 87558 55246 87610
rect 55298 87558 55310 87610
rect 55362 87558 55374 87610
rect 55426 87558 55438 87610
rect 55490 87558 73582 87610
rect 73634 87558 73646 87610
rect 73698 87558 73710 87610
rect 73762 87558 73774 87610
rect 73826 87558 73838 87610
rect 73890 87558 88596 87610
rect 4876 87536 88596 87558
rect 10630 87424 10636 87476
rect 10688 87464 10694 87476
rect 10880 87467 10938 87473
rect 10880 87464 10892 87467
rect 10688 87436 10892 87464
rect 10688 87424 10694 87436
rect 10880 87433 10892 87436
rect 10926 87433 10938 87467
rect 10880 87427 10938 87433
rect 15049 87467 15107 87473
rect 15049 87433 15061 87467
rect 15095 87464 15107 87467
rect 15138 87464 15144 87476
rect 15095 87436 15144 87464
rect 15095 87433 15107 87436
rect 15049 87427 15107 87433
rect 15138 87424 15144 87436
rect 15196 87424 15202 87476
rect 16981 87467 17039 87473
rect 16981 87433 16993 87467
rect 17027 87464 17039 87467
rect 17070 87464 17076 87476
rect 17027 87436 17076 87464
rect 17027 87433 17039 87436
rect 16981 87427 17039 87433
rect 17070 87424 17076 87436
rect 17128 87424 17134 87476
rect 18266 87424 18272 87476
rect 18324 87424 18330 87476
rect 19557 87467 19615 87473
rect 19557 87433 19569 87467
rect 19603 87464 19615 87467
rect 19646 87464 19652 87476
rect 19603 87436 19652 87464
rect 19603 87433 19615 87436
rect 19557 87427 19615 87433
rect 19646 87424 19652 87436
rect 19704 87424 19710 87476
rect 21489 87467 21547 87473
rect 21489 87433 21501 87467
rect 21535 87464 21547 87467
rect 21578 87464 21584 87476
rect 21535 87436 21584 87464
rect 21535 87433 21547 87436
rect 21489 87427 21547 87433
rect 21578 87424 21584 87436
rect 21636 87424 21642 87476
rect 22777 87467 22835 87473
rect 22777 87433 22789 87467
rect 22823 87464 22835 87467
rect 22866 87464 22872 87476
rect 22823 87436 22872 87464
rect 22823 87433 22835 87436
rect 22777 87427 22835 87433
rect 22866 87424 22872 87436
rect 22924 87424 22930 87476
rect 23421 87467 23479 87473
rect 23421 87433 23433 87467
rect 23467 87464 23479 87467
rect 23510 87464 23516 87476
rect 23467 87436 23516 87464
rect 23467 87433 23479 87436
rect 23421 87427 23479 87433
rect 23510 87424 23516 87436
rect 23568 87424 23574 87476
rect 24709 87467 24767 87473
rect 24709 87433 24721 87467
rect 24755 87464 24767 87467
rect 24798 87464 24804 87476
rect 24755 87436 24804 87464
rect 24755 87433 24767 87436
rect 24709 87427 24767 87433
rect 24798 87424 24804 87436
rect 24856 87424 24862 87476
rect 25997 87467 26055 87473
rect 25997 87433 26009 87467
rect 26043 87464 26055 87467
rect 26086 87464 26092 87476
rect 26043 87436 26092 87464
rect 26043 87433 26055 87436
rect 25997 87427 26055 87433
rect 26086 87424 26092 87436
rect 26144 87424 26150 87476
rect 27285 87467 27343 87473
rect 27285 87433 27297 87467
rect 27331 87464 27343 87467
rect 27374 87464 27380 87476
rect 27331 87436 27380 87464
rect 27331 87433 27343 87436
rect 27285 87427 27343 87433
rect 27374 87424 27380 87436
rect 27432 87424 27438 87476
rect 29217 87467 29275 87473
rect 29217 87433 29229 87467
rect 29263 87464 29275 87467
rect 29306 87464 29312 87476
rect 29263 87436 29312 87464
rect 29263 87433 29275 87436
rect 29217 87427 29275 87433
rect 29306 87424 29312 87436
rect 29364 87424 29370 87476
rect 30594 87424 30600 87476
rect 30652 87464 30658 87476
rect 30936 87467 30994 87473
rect 30936 87464 30948 87467
rect 30652 87436 30948 87464
rect 30652 87424 30658 87436
rect 30936 87433 30948 87436
rect 30982 87433 30994 87467
rect 30936 87427 30994 87433
rect 31238 87424 31244 87476
rect 31296 87464 31302 87476
rect 31379 87467 31437 87473
rect 31379 87464 31391 87467
rect 31296 87436 31391 87464
rect 31296 87424 31302 87436
rect 31379 87433 31391 87436
rect 31425 87433 31437 87467
rect 31379 87427 31437 87433
rect 32526 87424 32532 87476
rect 32584 87464 32590 87476
rect 32776 87467 32834 87473
rect 32776 87464 32788 87467
rect 32584 87436 32788 87464
rect 32584 87424 32590 87436
rect 32776 87433 32788 87436
rect 32822 87433 32834 87467
rect 32776 87427 32834 87433
rect 33814 87424 33820 87476
rect 33872 87464 33878 87476
rect 34064 87467 34122 87473
rect 34064 87464 34076 87467
rect 33872 87436 34076 87464
rect 33872 87424 33878 87436
rect 34064 87433 34076 87436
rect 34110 87433 34122 87467
rect 34064 87427 34122 87433
rect 35102 87424 35108 87476
rect 35160 87464 35166 87476
rect 35352 87467 35410 87473
rect 35352 87464 35364 87467
rect 35160 87436 35364 87464
rect 35160 87424 35166 87436
rect 35352 87433 35364 87436
rect 35398 87433 35410 87467
rect 35352 87427 35410 87433
rect 35746 87424 35752 87476
rect 35804 87464 35810 87476
rect 36088 87467 36146 87473
rect 36088 87464 36100 87467
rect 35804 87436 36100 87464
rect 35804 87424 35810 87436
rect 36088 87433 36100 87436
rect 36134 87433 36146 87467
rect 36088 87427 36146 87433
rect 37126 87424 37132 87476
rect 37184 87464 37190 87476
rect 37284 87467 37342 87473
rect 37284 87464 37296 87467
rect 37184 87436 37296 87464
rect 37184 87424 37190 87436
rect 37284 87433 37296 87436
rect 37330 87433 37342 87467
rect 37284 87427 37342 87433
rect 37678 87424 37684 87476
rect 37736 87464 37742 87476
rect 37865 87467 37923 87473
rect 37865 87464 37877 87467
rect 37736 87436 37877 87464
rect 37736 87424 37742 87436
rect 37865 87433 37877 87436
rect 37911 87433 37923 87467
rect 37865 87427 37923 87433
rect 38213 87467 38271 87473
rect 38213 87433 38225 87467
rect 38259 87464 38271 87467
rect 38322 87464 38328 87476
rect 38259 87436 38328 87464
rect 38259 87433 38271 87436
rect 38213 87427 38271 87433
rect 10722 87322 10728 87374
rect 10780 87322 10786 87374
rect 15156 87328 15184 87424
rect 15782 87356 15788 87408
rect 15840 87396 15846 87408
rect 16521 87399 16579 87405
rect 15840 87384 16288 87396
rect 16383 87387 16441 87393
rect 16383 87384 16395 87387
rect 15840 87368 16395 87384
rect 15840 87356 15846 87368
rect 16260 87356 16395 87368
rect 16383 87353 16395 87356
rect 16429 87384 16441 87387
rect 16521 87384 16533 87399
rect 16429 87365 16533 87384
rect 16567 87365 16579 87399
rect 16429 87359 16579 87365
rect 17088 87362 17116 87424
rect 18284 87396 18312 87424
rect 19664 87396 19692 87424
rect 18284 87373 18588 87396
rect 19664 87373 19876 87396
rect 17165 87365 17223 87371
rect 18284 87368 18633 87373
rect 19664 87368 19921 87373
rect 17165 87362 17177 87365
rect 16429 87356 16564 87359
rect 16429 87353 16441 87356
rect 16383 87347 16441 87353
rect 15325 87331 15383 87337
rect 17088 87334 17177 87362
rect 15325 87328 15337 87331
rect 15156 87300 15337 87328
rect 15325 87297 15337 87300
rect 15371 87297 15383 87331
rect 17165 87331 17177 87334
rect 17211 87331 17223 87365
rect 18560 87367 18633 87368
rect 17165 87325 17223 87331
rect 15325 87291 15383 87297
rect 18266 87288 18272 87340
rect 18324 87328 18330 87340
rect 18407 87331 18465 87337
rect 18560 87336 18587 87367
rect 18407 87328 18419 87331
rect 18324 87300 18419 87328
rect 18324 87288 18330 87300
rect 18407 87297 18419 87300
rect 18453 87297 18465 87331
rect 18575 87333 18587 87336
rect 18621 87333 18633 87367
rect 19848 87367 19921 87368
rect 18575 87327 18633 87333
rect 18407 87291 18465 87297
rect 19554 87288 19560 87340
rect 19612 87328 19618 87340
rect 19695 87331 19753 87337
rect 19848 87336 19875 87367
rect 19695 87328 19707 87331
rect 19612 87300 19707 87328
rect 19612 87288 19618 87300
rect 19695 87297 19707 87300
rect 19741 87297 19753 87331
rect 19863 87333 19875 87336
rect 19909 87333 19921 87367
rect 20290 87356 20296 87408
rect 20348 87364 20354 87408
rect 20753 87399 20811 87405
rect 20601 87367 20659 87373
rect 20601 87364 20613 87367
rect 20348 87356 20613 87364
rect 20308 87336 20613 87356
rect 19863 87327 19921 87333
rect 20601 87333 20613 87336
rect 20647 87364 20659 87367
rect 20753 87365 20765 87399
rect 20799 87365 20811 87399
rect 20753 87364 20811 87365
rect 20647 87359 20811 87364
rect 21596 87384 21624 87424
rect 22884 87396 22912 87424
rect 21811 87387 21869 87393
rect 21811 87384 21823 87387
rect 20647 87336 20796 87359
rect 21596 87356 21823 87384
rect 21811 87353 21823 87356
rect 21857 87353 21869 87387
rect 22884 87384 23004 87396
rect 23191 87387 23249 87393
rect 23191 87384 23203 87387
rect 22884 87368 23203 87384
rect 22976 87356 23203 87368
rect 21811 87347 21869 87353
rect 23191 87353 23203 87356
rect 23237 87353 23249 87387
rect 23191 87347 23249 87353
rect 23528 87362 23556 87424
rect 23605 87365 23663 87371
rect 23605 87362 23617 87365
rect 20647 87333 20659 87336
rect 23528 87334 23617 87362
rect 20601 87327 20659 87333
rect 23605 87331 23617 87334
rect 23651 87331 23663 87365
rect 24816 87362 24844 87424
rect 26104 87384 26132 87424
rect 26319 87387 26377 87393
rect 26319 87384 26331 87387
rect 24893 87365 24951 87371
rect 24893 87362 24905 87365
rect 24816 87334 24905 87362
rect 23605 87325 23663 87331
rect 24893 87331 24905 87334
rect 24939 87331 24951 87365
rect 26104 87356 26331 87384
rect 26319 87353 26331 87356
rect 26365 87353 26377 87387
rect 27392 87384 27420 87424
rect 27607 87387 27665 87393
rect 27607 87384 27619 87387
rect 27392 87356 27619 87384
rect 26319 87347 26377 87353
rect 27607 87353 27619 87356
rect 27653 87353 27665 87387
rect 28018 87356 28024 87408
rect 28076 87364 28082 87408
rect 28481 87399 28539 87405
rect 28329 87367 28387 87373
rect 28329 87364 28341 87367
rect 28076 87356 28341 87364
rect 27607 87347 27665 87353
rect 28036 87336 28341 87356
rect 24893 87325 24951 87331
rect 28329 87333 28341 87336
rect 28375 87364 28387 87367
rect 28481 87365 28493 87399
rect 28527 87365 28539 87399
rect 28481 87364 28539 87365
rect 28375 87359 28539 87364
rect 29324 87384 29352 87424
rect 29539 87387 29597 87393
rect 29539 87384 29551 87387
rect 28375 87336 28524 87359
rect 29324 87356 29551 87384
rect 29539 87353 29551 87356
rect 29585 87353 29597 87387
rect 29539 87347 29597 87353
rect 28375 87333 28387 87336
rect 28329 87327 28387 87333
rect 30594 87322 30600 87374
rect 30652 87362 30658 87374
rect 30733 87365 30791 87371
rect 30733 87362 30745 87365
rect 30652 87334 30745 87362
rect 30652 87322 30658 87334
rect 30733 87331 30745 87334
rect 30779 87331 30791 87365
rect 30733 87325 30791 87331
rect 31514 87322 31520 87374
rect 31572 87371 31578 87374
rect 31572 87365 31606 87371
rect 31594 87331 31606 87365
rect 31572 87325 31606 87331
rect 31572 87322 31578 87325
rect 32618 87322 32624 87374
rect 32676 87322 32682 87374
rect 33722 87322 33728 87374
rect 33780 87362 33786 87374
rect 33861 87365 33919 87371
rect 33861 87362 33873 87365
rect 33780 87334 33873 87362
rect 33780 87322 33786 87334
rect 33861 87331 33873 87334
rect 33907 87331 33919 87365
rect 33861 87325 33919 87331
rect 34918 87322 34924 87374
rect 34976 87362 34982 87374
rect 35149 87365 35207 87371
rect 35149 87362 35161 87365
rect 34976 87334 35161 87362
rect 34976 87322 34982 87334
rect 35149 87331 35161 87334
rect 35195 87331 35207 87365
rect 35149 87325 35207 87331
rect 35930 87322 35936 87374
rect 35988 87322 35994 87374
rect 37126 87322 37132 87374
rect 37184 87322 37190 87374
rect 19695 87291 19753 87297
rect 22682 87220 22688 87272
rect 22740 87260 22746 87272
rect 23007 87263 23065 87269
rect 23007 87260 23019 87263
rect 22740 87232 23019 87260
rect 22740 87220 22746 87232
rect 23007 87229 23019 87232
rect 23053 87229 23065 87263
rect 23007 87223 23065 87229
rect 27098 87220 27104 87272
rect 27156 87260 27162 87272
rect 27423 87263 27481 87269
rect 27423 87260 27435 87263
rect 27156 87232 27435 87260
rect 27156 87220 27162 87232
rect 27423 87229 27435 87232
rect 27469 87229 27481 87263
rect 37880 87260 37908 87427
rect 38322 87424 38328 87436
rect 38380 87424 38386 87476
rect 38966 87424 38972 87476
rect 39024 87464 39030 87476
rect 39676 87467 39734 87473
rect 39676 87464 39688 87467
rect 39024 87436 39688 87464
rect 39024 87424 39030 87436
rect 39676 87433 39688 87436
rect 39722 87433 39734 87467
rect 39676 87427 39734 87433
rect 40254 87424 40260 87476
rect 40312 87464 40318 87476
rect 40504 87467 40562 87473
rect 40504 87464 40516 87467
rect 40312 87436 40516 87464
rect 40312 87424 40318 87436
rect 40504 87433 40516 87436
rect 40550 87433 40562 87467
rect 40504 87427 40562 87433
rect 40809 87467 40867 87473
rect 40809 87433 40821 87467
rect 40855 87464 40867 87467
rect 40898 87464 40904 87476
rect 40855 87436 40904 87464
rect 40855 87433 40867 87436
rect 40809 87427 40867 87433
rect 40898 87424 40904 87436
rect 40956 87424 40962 87476
rect 42186 87424 42192 87476
rect 42244 87464 42250 87476
rect 42327 87467 42385 87473
rect 42327 87464 42339 87467
rect 42244 87436 42339 87464
rect 42244 87424 42250 87436
rect 42327 87433 42339 87436
rect 42373 87433 42385 87467
rect 42327 87427 42385 87433
rect 43474 87424 43480 87476
rect 43532 87464 43538 87476
rect 43816 87467 43874 87473
rect 43816 87464 43828 87467
rect 43532 87436 43828 87464
rect 43532 87424 43538 87436
rect 43816 87433 43828 87436
rect 43862 87433 43874 87467
rect 43816 87427 43874 87433
rect 44118 87424 44124 87476
rect 44176 87464 44182 87476
rect 44259 87467 44317 87473
rect 44259 87464 44271 87467
rect 44176 87436 44271 87464
rect 44176 87424 44182 87436
rect 44259 87433 44271 87436
rect 44305 87433 44317 87467
rect 44259 87427 44317 87433
rect 52401 87467 52459 87473
rect 52401 87433 52413 87467
rect 52447 87464 52459 87467
rect 52490 87464 52496 87476
rect 52447 87436 52496 87464
rect 52447 87433 52459 87436
rect 52401 87427 52459 87433
rect 52490 87424 52496 87436
rect 52548 87424 52554 87476
rect 55621 87467 55679 87473
rect 55621 87433 55633 87467
rect 55667 87464 55679 87467
rect 55710 87464 55716 87476
rect 55667 87436 55716 87464
rect 55667 87433 55679 87436
rect 55621 87427 55679 87433
rect 55710 87424 55716 87436
rect 55768 87424 55774 87476
rect 56909 87467 56967 87473
rect 56909 87433 56921 87467
rect 56955 87464 56967 87467
rect 56998 87464 57004 87476
rect 56955 87436 57004 87464
rect 56955 87433 56967 87436
rect 56909 87427 56967 87433
rect 56998 87424 57004 87436
rect 57056 87424 57062 87476
rect 57553 87467 57611 87473
rect 57553 87433 57565 87467
rect 57599 87464 57611 87467
rect 57642 87464 57648 87476
rect 57599 87436 57648 87464
rect 57599 87433 57611 87436
rect 57553 87427 57611 87433
rect 57642 87424 57648 87436
rect 57700 87424 57706 87476
rect 60129 87467 60187 87473
rect 60129 87433 60141 87467
rect 60175 87464 60187 87467
rect 60218 87464 60224 87476
rect 60175 87436 60224 87464
rect 60175 87433 60187 87436
rect 60129 87427 60187 87433
rect 60218 87424 60224 87436
rect 60276 87424 60282 87476
rect 63349 87467 63407 87473
rect 63349 87433 63361 87467
rect 63395 87464 63407 87467
rect 63438 87464 63444 87476
rect 63395 87436 63444 87464
rect 63395 87433 63407 87436
rect 63349 87427 63407 87433
rect 63438 87424 63444 87436
rect 63496 87424 63502 87476
rect 64637 87467 64695 87473
rect 64637 87433 64649 87467
rect 64683 87464 64695 87467
rect 64726 87464 64732 87476
rect 64683 87436 64732 87464
rect 64683 87433 64695 87436
rect 64637 87427 64695 87433
rect 64726 87424 64732 87436
rect 64784 87424 64790 87476
rect 65281 87467 65339 87473
rect 65281 87433 65293 87467
rect 65327 87464 65339 87467
rect 65370 87464 65376 87476
rect 65327 87436 65376 87464
rect 65327 87433 65339 87436
rect 65281 87427 65339 87433
rect 65370 87424 65376 87436
rect 65428 87424 65434 87476
rect 67946 87424 67952 87476
rect 68004 87464 68010 87476
rect 68196 87467 68254 87473
rect 68196 87464 68208 87467
rect 68004 87436 68208 87464
rect 68004 87424 68010 87436
rect 68196 87433 68208 87436
rect 68242 87433 68254 87467
rect 68196 87427 68254 87433
rect 69234 87424 69240 87476
rect 69292 87464 69298 87476
rect 69576 87467 69634 87473
rect 69576 87464 69588 87467
rect 69292 87436 69588 87464
rect 69292 87424 69298 87436
rect 69576 87433 69588 87436
rect 69622 87433 69634 87467
rect 69576 87427 69634 87433
rect 69878 87424 69884 87476
rect 69936 87464 69942 87476
rect 70019 87467 70077 87473
rect 70019 87464 70031 87467
rect 69936 87436 70031 87464
rect 69936 87424 69942 87436
rect 70019 87433 70031 87436
rect 70065 87433 70077 87467
rect 70019 87427 70077 87433
rect 71166 87424 71172 87476
rect 71224 87464 71230 87476
rect 71416 87467 71474 87473
rect 71416 87464 71428 87467
rect 71224 87436 71428 87464
rect 71224 87424 71230 87436
rect 71416 87433 71428 87436
rect 71462 87433 71474 87467
rect 71416 87427 71474 87433
rect 72454 87424 72460 87476
rect 72512 87464 72518 87476
rect 72704 87467 72762 87473
rect 72704 87464 72716 87467
rect 72512 87436 72716 87464
rect 72512 87424 72518 87436
rect 72704 87433 72716 87436
rect 72750 87433 72762 87467
rect 72704 87427 72762 87433
rect 73098 87424 73104 87476
rect 73156 87464 73162 87476
rect 73239 87467 73297 87473
rect 73239 87464 73251 87467
rect 73156 87436 73251 87464
rect 73156 87424 73162 87436
rect 73239 87433 73251 87436
rect 73285 87433 73297 87467
rect 73239 87427 73297 87433
rect 74386 87424 74392 87476
rect 74444 87464 74450 87476
rect 74728 87467 74786 87473
rect 74728 87464 74740 87467
rect 74444 87436 74740 87464
rect 74444 87424 74450 87436
rect 74728 87433 74740 87436
rect 74774 87433 74786 87467
rect 74728 87427 74786 87433
rect 75674 87424 75680 87476
rect 75732 87464 75738 87476
rect 75924 87467 75982 87473
rect 75924 87464 75936 87467
rect 75732 87436 75936 87464
rect 75732 87424 75738 87436
rect 75924 87433 75936 87436
rect 75970 87433 75982 87467
rect 75924 87427 75982 87433
rect 76962 87424 76968 87476
rect 77020 87464 77026 87476
rect 77304 87467 77362 87473
rect 77304 87464 77316 87467
rect 77020 87436 77316 87464
rect 77020 87424 77026 87436
rect 77304 87433 77316 87436
rect 77350 87433 77362 87467
rect 77304 87427 77362 87433
rect 77606 87424 77612 87476
rect 77664 87464 77670 87476
rect 77747 87467 77805 87473
rect 77747 87464 77759 87467
rect 77664 87436 77759 87464
rect 77664 87424 77670 87436
rect 77747 87433 77759 87436
rect 77793 87433 77805 87467
rect 77747 87427 77805 87433
rect 78894 87424 78900 87476
rect 78952 87464 78958 87476
rect 79144 87467 79202 87473
rect 79144 87464 79156 87467
rect 78952 87436 79156 87464
rect 78952 87424 78958 87436
rect 79144 87433 79156 87436
rect 79190 87433 79202 87467
rect 79144 87427 79202 87433
rect 80182 87424 80188 87476
rect 80240 87464 80246 87476
rect 80432 87467 80490 87473
rect 80432 87464 80444 87467
rect 80240 87436 80444 87464
rect 80240 87424 80246 87436
rect 80432 87433 80444 87436
rect 80478 87433 80490 87467
rect 80432 87427 80490 87433
rect 80826 87424 80832 87476
rect 80884 87464 80890 87476
rect 80967 87467 81025 87473
rect 80967 87464 80979 87467
rect 80884 87436 80979 87464
rect 80884 87424 80890 87436
rect 80967 87433 80979 87436
rect 81013 87433 81025 87467
rect 80967 87427 81025 87433
rect 82114 87424 82120 87476
rect 82172 87464 82178 87476
rect 82456 87467 82514 87473
rect 82456 87464 82468 87467
rect 82172 87436 82468 87464
rect 82172 87424 82178 87436
rect 82456 87433 82468 87436
rect 82502 87433 82514 87467
rect 82456 87427 82514 87433
rect 38461 87399 38519 87405
rect 38461 87396 38473 87399
rect 38049 87365 38107 87371
rect 38049 87331 38061 87365
rect 38095 87362 38107 87365
rect 38138 87362 38144 87374
rect 38095 87334 38144 87362
rect 38095 87331 38107 87334
rect 38049 87325 38107 87331
rect 38138 87322 38144 87334
rect 38196 87322 38202 87374
rect 38248 87368 38473 87396
rect 38248 87260 38276 87368
rect 38461 87365 38473 87368
rect 38507 87365 38519 87399
rect 40916 87396 40944 87424
rect 41037 87399 41095 87405
rect 41037 87396 41049 87399
rect 38461 87359 38519 87365
rect 39242 87322 39248 87374
rect 39300 87362 39306 87374
rect 39473 87365 39531 87371
rect 39473 87362 39485 87365
rect 39300 87334 39485 87362
rect 39300 87322 39306 87334
rect 39473 87331 39485 87334
rect 39519 87331 39531 87365
rect 39473 87325 39531 87331
rect 40346 87322 40352 87374
rect 40404 87322 40410 87374
rect 40916 87368 41049 87396
rect 41037 87365 41049 87368
rect 41083 87365 41095 87399
rect 42554 87371 42560 87374
rect 41037 87359 41095 87365
rect 42533 87365 42560 87371
rect 42533 87331 42545 87365
rect 42533 87325 42560 87331
rect 42554 87322 42560 87325
rect 42612 87322 42618 87374
rect 42830 87356 42836 87408
rect 42888 87396 42894 87408
rect 42925 87399 42983 87405
rect 42925 87396 42937 87399
rect 42888 87368 42937 87396
rect 42888 87356 42894 87368
rect 42925 87365 42937 87368
rect 42971 87365 42983 87399
rect 42925 87359 42983 87365
rect 43658 87322 43664 87374
rect 43716 87322 43722 87374
rect 44465 87365 44523 87371
rect 44465 87331 44477 87365
rect 44511 87362 44523 87365
rect 44670 87362 44676 87374
rect 44511 87334 44676 87362
rect 44511 87331 44523 87334
rect 44465 87325 44523 87331
rect 44670 87322 44676 87334
rect 44728 87322 44734 87374
rect 44762 87356 44768 87408
rect 44820 87396 44826 87408
rect 44857 87399 44915 87405
rect 44857 87396 44869 87399
rect 44820 87368 44869 87396
rect 44820 87356 44826 87368
rect 44857 87365 44869 87368
rect 44903 87365 44915 87399
rect 44857 87359 44915 87365
rect 45406 87356 45412 87408
rect 45464 87396 45470 87408
rect 45501 87399 45559 87405
rect 45501 87396 45513 87399
rect 45464 87368 45513 87396
rect 45464 87356 45470 87368
rect 45501 87365 45513 87368
rect 45547 87365 45559 87399
rect 45501 87359 45559 87365
rect 46050 87356 46056 87408
rect 46108 87396 46114 87408
rect 46237 87399 46295 87405
rect 46237 87396 46249 87399
rect 46108 87368 46249 87396
rect 46108 87356 46114 87368
rect 46237 87365 46249 87368
rect 46283 87365 46295 87399
rect 46237 87359 46295 87365
rect 46694 87356 46700 87408
rect 46752 87396 46758 87408
rect 46789 87399 46847 87405
rect 46789 87396 46801 87399
rect 46752 87368 46801 87396
rect 46752 87356 46758 87368
rect 46789 87365 46801 87368
rect 46835 87365 46847 87399
rect 46789 87359 46847 87365
rect 47338 87356 47344 87408
rect 47396 87396 47402 87408
rect 47433 87399 47491 87405
rect 47433 87396 47445 87399
rect 47396 87368 47445 87396
rect 47396 87356 47402 87368
rect 47433 87365 47445 87368
rect 47479 87365 47491 87399
rect 47433 87359 47491 87365
rect 47982 87356 47988 87408
rect 48040 87396 48046 87408
rect 48077 87399 48135 87405
rect 48077 87396 48089 87399
rect 48040 87368 48089 87396
rect 48040 87356 48046 87368
rect 48077 87365 48089 87368
rect 48123 87365 48135 87399
rect 48077 87359 48135 87365
rect 48626 87356 48632 87408
rect 48684 87396 48690 87408
rect 48813 87399 48871 87405
rect 48813 87396 48825 87399
rect 48684 87368 48825 87396
rect 48684 87356 48690 87368
rect 48813 87365 48825 87368
rect 48859 87365 48871 87399
rect 48813 87359 48871 87365
rect 49270 87356 49276 87408
rect 49328 87396 49334 87408
rect 49365 87399 49423 87405
rect 49365 87396 49377 87399
rect 49328 87368 49377 87396
rect 49328 87356 49334 87368
rect 49365 87365 49377 87368
rect 49411 87365 49423 87399
rect 49365 87359 49423 87365
rect 49914 87356 49920 87408
rect 49972 87396 49978 87408
rect 50009 87399 50067 87405
rect 50009 87396 50021 87399
rect 49972 87368 50021 87396
rect 49972 87356 49978 87368
rect 50009 87365 50021 87368
rect 50055 87365 50067 87399
rect 50009 87359 50067 87365
rect 50558 87356 50564 87408
rect 50616 87396 50622 87408
rect 50653 87399 50711 87405
rect 50653 87396 50665 87399
rect 50616 87368 50665 87396
rect 50616 87356 50622 87368
rect 50653 87365 50665 87368
rect 50699 87365 50711 87399
rect 50653 87359 50711 87365
rect 52508 87328 52536 87424
rect 53778 87356 53784 87408
rect 53836 87364 53842 87408
rect 54241 87399 54299 87405
rect 54087 87367 54145 87373
rect 54087 87364 54099 87367
rect 53836 87356 54099 87364
rect 52585 87331 52643 87337
rect 53796 87336 54099 87356
rect 52585 87328 52597 87331
rect 52508 87300 52597 87328
rect 52585 87297 52597 87300
rect 52631 87297 52643 87331
rect 54087 87333 54099 87336
rect 54133 87364 54145 87367
rect 54241 87365 54253 87399
rect 54287 87365 54299 87399
rect 54793 87399 54851 87405
rect 54793 87396 54805 87399
rect 54241 87364 54299 87365
rect 54133 87359 54299 87364
rect 54133 87336 54284 87359
rect 54133 87333 54145 87336
rect 54087 87327 54145 87333
rect 54422 87322 54428 87374
rect 54480 87362 54486 87374
rect 54532 87371 54805 87396
rect 54517 87368 54805 87371
rect 54517 87365 54575 87368
rect 54517 87362 54529 87365
rect 54480 87334 54529 87362
rect 54480 87322 54486 87334
rect 54517 87331 54529 87334
rect 54563 87331 54575 87365
rect 54793 87365 54805 87368
rect 54839 87365 54851 87399
rect 54793 87359 54851 87365
rect 55728 87384 55756 87424
rect 55943 87387 56001 87393
rect 55943 87384 55955 87387
rect 55728 87356 55955 87384
rect 55943 87353 55955 87356
rect 55989 87353 56001 87387
rect 57016 87384 57044 87424
rect 57231 87387 57289 87393
rect 57231 87384 57243 87387
rect 57016 87356 57243 87384
rect 55943 87347 56001 87353
rect 57231 87353 57243 87356
rect 57277 87353 57289 87387
rect 57231 87347 57289 87353
rect 57660 87362 57688 87424
rect 57737 87365 57795 87371
rect 57737 87362 57749 87365
rect 57660 87334 57749 87362
rect 54517 87325 54575 87331
rect 57737 87331 57749 87334
rect 57783 87331 57795 87365
rect 58930 87356 58936 87408
rect 58988 87364 58994 87408
rect 59393 87399 59451 87405
rect 59239 87367 59297 87373
rect 59239 87364 59251 87367
rect 58988 87356 59251 87364
rect 58948 87336 59251 87356
rect 57737 87325 57795 87331
rect 59239 87333 59251 87336
rect 59285 87364 59297 87367
rect 59393 87365 59405 87399
rect 59439 87365 59451 87399
rect 60236 87396 60264 87424
rect 60236 87373 60448 87396
rect 60236 87368 60493 87373
rect 59393 87364 59451 87365
rect 59285 87359 59451 87364
rect 60420 87367 60493 87368
rect 59285 87336 59436 87359
rect 59285 87333 59297 87336
rect 59239 87327 59297 87333
rect 52585 87291 52643 87297
rect 60126 87288 60132 87340
rect 60184 87328 60190 87340
rect 60267 87331 60325 87337
rect 60420 87336 60447 87367
rect 60267 87328 60279 87331
rect 60184 87300 60279 87328
rect 60184 87288 60190 87300
rect 60267 87297 60279 87300
rect 60313 87297 60325 87331
rect 60435 87333 60447 87336
rect 60481 87333 60493 87367
rect 61506 87356 61512 87408
rect 61564 87364 61570 87408
rect 61969 87399 62027 87405
rect 61817 87367 61875 87373
rect 61817 87364 61829 87367
rect 61564 87356 61829 87364
rect 61524 87336 61829 87356
rect 60435 87327 60493 87333
rect 61817 87333 61829 87336
rect 61863 87364 61875 87367
rect 61969 87365 61981 87399
rect 62015 87365 62027 87399
rect 62521 87399 62579 87405
rect 62521 87396 62533 87399
rect 61969 87364 62027 87365
rect 61863 87359 62027 87364
rect 61863 87336 62012 87359
rect 61863 87333 61875 87336
rect 61817 87327 61875 87333
rect 62150 87322 62156 87374
rect 62208 87362 62214 87374
rect 62260 87371 62533 87396
rect 62245 87368 62533 87371
rect 62245 87365 62303 87368
rect 62245 87362 62257 87365
rect 62208 87334 62257 87362
rect 62208 87322 62214 87334
rect 62245 87331 62257 87334
rect 62291 87331 62303 87365
rect 62521 87365 62533 87368
rect 62567 87365 62579 87399
rect 62521 87359 62579 87365
rect 63456 87384 63484 87424
rect 63671 87387 63729 87393
rect 63671 87384 63683 87387
rect 63456 87356 63683 87384
rect 63671 87353 63683 87356
rect 63717 87353 63729 87387
rect 64744 87384 64772 87424
rect 64959 87387 65017 87393
rect 64959 87384 64971 87387
rect 64744 87356 64971 87384
rect 63671 87347 63729 87353
rect 64959 87353 64971 87356
rect 65005 87353 65017 87387
rect 64959 87347 65017 87353
rect 65388 87362 65416 87424
rect 65465 87365 65523 87371
rect 65465 87362 65477 87365
rect 65388 87334 65477 87362
rect 62245 87325 62303 87331
rect 65465 87331 65477 87334
rect 65511 87331 65523 87365
rect 66658 87356 66664 87408
rect 66716 87364 66722 87408
rect 67121 87399 67179 87405
rect 66967 87367 67025 87373
rect 66967 87364 66979 87367
rect 66716 87356 66979 87364
rect 66676 87336 66979 87356
rect 65465 87325 65523 87331
rect 66967 87333 66979 87336
rect 67013 87364 67025 87367
rect 67121 87365 67133 87399
rect 67167 87365 67179 87399
rect 67121 87364 67179 87365
rect 67013 87359 67179 87364
rect 67013 87336 67164 87359
rect 67013 87333 67025 87336
rect 66967 87327 67025 87333
rect 67854 87322 67860 87374
rect 67912 87362 67918 87374
rect 67993 87365 68051 87371
rect 67993 87362 68005 87365
rect 67912 87334 68005 87362
rect 67912 87322 67918 87334
rect 67993 87331 68005 87334
rect 68039 87331 68051 87365
rect 67993 87325 68051 87331
rect 69326 87322 69332 87374
rect 69384 87362 69390 87374
rect 69421 87365 69479 87371
rect 69421 87362 69433 87365
rect 69384 87334 69433 87362
rect 69384 87322 69390 87334
rect 69421 87331 69433 87334
rect 69467 87331 69479 87365
rect 69421 87325 69479 87331
rect 70062 87322 70068 87374
rect 70120 87362 70126 87374
rect 70188 87365 70246 87371
rect 70188 87362 70200 87365
rect 70120 87334 70200 87362
rect 70120 87322 70126 87334
rect 70188 87331 70200 87334
rect 70234 87331 70246 87365
rect 70188 87325 70246 87331
rect 71166 87322 71172 87374
rect 71224 87362 71230 87374
rect 71261 87365 71319 87371
rect 71261 87362 71273 87365
rect 71224 87334 71273 87362
rect 71224 87322 71230 87334
rect 71261 87331 71273 87334
rect 71307 87331 71319 87365
rect 71261 87325 71319 87331
rect 72270 87322 72276 87374
rect 72328 87362 72334 87374
rect 72501 87365 72559 87371
rect 72501 87362 72513 87365
rect 72328 87334 72513 87362
rect 72328 87322 72334 87334
rect 72501 87331 72513 87334
rect 72547 87331 72559 87365
rect 72501 87325 72559 87331
rect 73374 87322 73380 87374
rect 73432 87371 73438 87374
rect 73432 87365 73466 87371
rect 73454 87331 73466 87365
rect 73432 87325 73466 87331
rect 73432 87322 73438 87325
rect 74478 87322 74484 87374
rect 74536 87362 74542 87374
rect 74573 87365 74631 87371
rect 74573 87362 74585 87365
rect 74536 87334 74585 87362
rect 74536 87322 74542 87334
rect 74573 87331 74585 87334
rect 74619 87331 74631 87365
rect 74573 87325 74631 87331
rect 75582 87322 75588 87374
rect 75640 87362 75646 87374
rect 75721 87365 75779 87371
rect 75721 87362 75733 87365
rect 75640 87334 75733 87362
rect 75640 87322 75646 87334
rect 75721 87331 75733 87334
rect 75767 87331 75779 87365
rect 77138 87365 77196 87371
rect 77138 87362 77150 87365
rect 75721 87325 75779 87331
rect 60267 87291 60325 87297
rect 76686 87288 76692 87340
rect 76744 87328 76750 87340
rect 77072 87334 77150 87362
rect 77072 87328 77100 87334
rect 76744 87300 77100 87328
rect 77138 87331 77150 87334
rect 77184 87331 77196 87365
rect 77138 87325 77196 87331
rect 77790 87322 77796 87374
rect 77848 87362 77854 87374
rect 77916 87365 77974 87371
rect 77916 87362 77928 87365
rect 77848 87334 77928 87362
rect 77848 87322 77854 87334
rect 77916 87331 77928 87334
rect 77962 87331 77974 87365
rect 77916 87325 77974 87331
rect 78894 87322 78900 87374
rect 78952 87362 78958 87374
rect 78989 87365 79047 87371
rect 78989 87362 79001 87365
rect 78952 87334 79001 87362
rect 78952 87322 78958 87334
rect 78989 87331 79001 87334
rect 79035 87331 79047 87365
rect 78989 87325 79047 87331
rect 80274 87322 80280 87374
rect 80332 87322 80338 87374
rect 81102 87322 81108 87374
rect 81160 87371 81166 87374
rect 81160 87365 81194 87371
rect 81182 87331 81194 87365
rect 81160 87325 81194 87331
rect 81160 87322 81166 87325
rect 82206 87322 82212 87374
rect 82264 87362 82270 87374
rect 82301 87365 82359 87371
rect 82301 87362 82313 87365
rect 82264 87334 82313 87362
rect 82264 87322 82270 87334
rect 82301 87331 82313 87334
rect 82347 87331 82359 87365
rect 82301 87325 82359 87331
rect 76744 87288 76750 87300
rect 37880 87232 38276 87260
rect 27423 87223 27481 87229
rect 39058 87220 39064 87272
rect 39116 87260 39122 87272
rect 39889 87263 39947 87269
rect 39889 87260 39901 87263
rect 39116 87232 39901 87260
rect 39116 87220 39122 87232
rect 39889 87229 39901 87232
rect 39935 87229 39947 87263
rect 39889 87223 39947 87229
rect 56814 87220 56820 87272
rect 56872 87260 56878 87272
rect 57047 87263 57105 87269
rect 57047 87260 57059 87263
rect 56872 87232 57059 87260
rect 56872 87220 56878 87232
rect 57047 87229 57059 87232
rect 57093 87229 57105 87263
rect 57047 87223 57105 87229
rect 62334 87220 62340 87272
rect 62392 87269 62398 87272
rect 62392 87263 62441 87269
rect 62392 87229 62395 87263
rect 62429 87229 62441 87263
rect 62392 87223 62441 87229
rect 62392 87220 62398 87223
rect 64542 87220 64548 87272
rect 64600 87260 64606 87272
rect 64775 87263 64833 87269
rect 64775 87260 64787 87263
rect 64600 87232 64787 87260
rect 64600 87220 64606 87232
rect 64775 87229 64787 87232
rect 64821 87229 64833 87263
rect 64775 87223 64833 87229
rect 15506 87152 15512 87204
rect 15564 87152 15570 87204
rect 16058 87152 16064 87204
rect 16116 87192 16122 87204
rect 16199 87195 16257 87201
rect 16199 87192 16211 87195
rect 16116 87164 16211 87192
rect 16116 87152 16122 87164
rect 16199 87161 16211 87164
rect 16245 87161 16257 87195
rect 16199 87155 16257 87161
rect 17162 87152 17168 87204
rect 17220 87192 17226 87204
rect 20474 87201 20480 87204
rect 17315 87195 17373 87201
rect 17315 87192 17327 87195
rect 17220 87164 17327 87192
rect 17220 87152 17226 87164
rect 17315 87161 17327 87164
rect 17361 87161 17373 87195
rect 17315 87155 17373 87161
rect 20431 87195 20480 87201
rect 20431 87161 20443 87195
rect 20477 87161 20480 87195
rect 20431 87155 20480 87161
rect 20474 87152 20480 87155
rect 20532 87152 20538 87204
rect 21578 87152 21584 87204
rect 21636 87201 21642 87204
rect 23786 87201 23792 87204
rect 21636 87195 21685 87201
rect 21636 87161 21639 87195
rect 21673 87161 21685 87195
rect 21636 87155 21685 87161
rect 23765 87195 23792 87201
rect 23765 87161 23777 87195
rect 23765 87155 23792 87161
rect 21636 87152 21642 87155
rect 23786 87152 23792 87155
rect 23844 87152 23850 87204
rect 25074 87201 25080 87204
rect 25052 87195 25080 87201
rect 25052 87161 25064 87195
rect 25052 87155 25080 87161
rect 25074 87152 25080 87155
rect 25132 87152 25138 87204
rect 26086 87152 26092 87204
rect 26144 87201 26150 87204
rect 28202 87201 28208 87204
rect 26144 87195 26193 87201
rect 26144 87161 26147 87195
rect 26181 87161 26193 87195
rect 26144 87155 26193 87161
rect 28159 87195 28208 87201
rect 28159 87161 28171 87195
rect 28205 87161 28208 87195
rect 28159 87155 28208 87161
rect 26144 87152 26150 87155
rect 28202 87152 28208 87155
rect 28260 87152 28266 87204
rect 29306 87152 29312 87204
rect 29364 87201 29370 87204
rect 29364 87195 29413 87201
rect 29364 87161 29367 87195
rect 29401 87161 29413 87195
rect 29364 87155 29413 87161
rect 29364 87152 29370 87155
rect 41818 87152 41824 87204
rect 41876 87192 41882 87204
rect 42097 87195 42155 87201
rect 42097 87192 42109 87195
rect 41876 87164 42109 87192
rect 41876 87152 41882 87164
rect 42097 87161 42109 87164
rect 42143 87161 42155 87195
rect 42097 87155 42155 87161
rect 52674 87152 52680 87204
rect 52732 87192 52738 87204
rect 52769 87195 52827 87201
rect 52769 87192 52781 87195
rect 52732 87164 52781 87192
rect 52732 87152 52738 87164
rect 52769 87161 52781 87164
rect 52815 87161 52827 87195
rect 52769 87155 52827 87161
rect 53502 87152 53508 87204
rect 53560 87192 53566 87204
rect 53919 87195 53977 87201
rect 53919 87192 53931 87195
rect 53560 87164 53931 87192
rect 53560 87152 53566 87164
rect 53919 87161 53931 87164
rect 53965 87161 53977 87195
rect 53919 87155 53977 87161
rect 54422 87152 54428 87204
rect 54480 87192 54486 87204
rect 54667 87195 54725 87201
rect 54667 87192 54679 87195
rect 54480 87164 54679 87192
rect 54480 87152 54486 87164
rect 54667 87161 54679 87164
rect 54713 87161 54725 87195
rect 54667 87155 54725 87161
rect 55710 87152 55716 87204
rect 55768 87201 55774 87204
rect 57918 87201 57924 87204
rect 55768 87195 55817 87201
rect 55768 87161 55771 87195
rect 55805 87161 55817 87195
rect 55768 87155 55817 87161
rect 57897 87195 57924 87201
rect 57897 87161 57909 87195
rect 57897 87155 57924 87161
rect 55768 87152 55774 87155
rect 57918 87152 57924 87155
rect 57976 87152 57982 87204
rect 59022 87152 59028 87204
rect 59080 87201 59086 87204
rect 59080 87195 59129 87201
rect 59080 87161 59083 87195
rect 59117 87161 59129 87195
rect 59080 87155 59129 87161
rect 59080 87152 59086 87155
rect 61230 87152 61236 87204
rect 61288 87192 61294 87204
rect 61647 87195 61705 87201
rect 61647 87192 61659 87195
rect 61288 87164 61659 87192
rect 61288 87152 61294 87164
rect 61647 87161 61659 87164
rect 61693 87161 61705 87195
rect 61647 87155 61705 87161
rect 63438 87152 63444 87204
rect 63496 87201 63502 87204
rect 65646 87201 65652 87204
rect 63496 87195 63545 87201
rect 63496 87161 63499 87195
rect 63533 87161 63545 87195
rect 63496 87155 63545 87161
rect 65625 87195 65652 87201
rect 65625 87161 65637 87195
rect 65625 87155 65652 87161
rect 63496 87152 63502 87155
rect 65646 87152 65652 87155
rect 65704 87152 65710 87204
rect 66750 87152 66756 87204
rect 66808 87201 66814 87204
rect 66808 87195 66857 87201
rect 66808 87161 66811 87195
rect 66845 87161 66857 87195
rect 66808 87155 66857 87161
rect 66808 87152 66814 87155
rect 4876 87066 88596 87088
rect 4876 87014 17722 87066
rect 17774 87014 17786 87066
rect 17838 87014 17850 87066
rect 17902 87014 17914 87066
rect 17966 87014 17978 87066
rect 18030 87014 36122 87066
rect 36174 87014 36186 87066
rect 36238 87014 36250 87066
rect 36302 87014 36314 87066
rect 36366 87014 36378 87066
rect 36430 87014 54522 87066
rect 54574 87014 54586 87066
rect 54638 87014 54650 87066
rect 54702 87014 54714 87066
rect 54766 87014 54778 87066
rect 54830 87014 72922 87066
rect 72974 87014 72986 87066
rect 73038 87014 73050 87066
rect 73102 87014 73114 87066
rect 73166 87014 73178 87066
rect 73230 87014 88596 87066
rect 4876 86992 88596 87014
rect 41542 86880 41548 86932
rect 41600 86920 41606 86932
rect 41792 86923 41850 86929
rect 41792 86920 41804 86923
rect 41600 86892 41804 86920
rect 41600 86880 41606 86892
rect 41792 86889 41804 86892
rect 41838 86889 41850 86923
rect 41792 86883 41850 86889
rect 41450 86710 41456 86762
rect 41508 86750 41514 86762
rect 41591 86753 41649 86759
rect 41591 86750 41603 86753
rect 41508 86722 41603 86750
rect 41508 86710 41514 86722
rect 41591 86719 41603 86722
rect 41637 86719 41649 86753
rect 41591 86713 41649 86719
rect 4876 86522 88596 86544
rect 4876 86470 18382 86522
rect 18434 86470 18446 86522
rect 18498 86470 18510 86522
rect 18562 86470 18574 86522
rect 18626 86470 18638 86522
rect 18690 86470 36782 86522
rect 36834 86470 36846 86522
rect 36898 86470 36910 86522
rect 36962 86470 36974 86522
rect 37026 86470 37038 86522
rect 37090 86470 55182 86522
rect 55234 86470 55246 86522
rect 55298 86470 55310 86522
rect 55362 86470 55374 86522
rect 55426 86470 55438 86522
rect 55490 86470 73582 86522
rect 73634 86470 73646 86522
rect 73698 86470 73710 86522
rect 73762 86470 73774 86522
rect 73826 86470 73838 86522
rect 73890 86470 88596 86522
rect 4876 86448 88596 86470
rect 4876 85978 88596 86000
rect 4876 85926 17722 85978
rect 17774 85926 17786 85978
rect 17838 85926 17850 85978
rect 17902 85926 17914 85978
rect 17966 85926 17978 85978
rect 18030 85926 36122 85978
rect 36174 85926 36186 85978
rect 36238 85926 36250 85978
rect 36302 85926 36314 85978
rect 36366 85926 36378 85978
rect 36430 85926 54522 85978
rect 54574 85926 54586 85978
rect 54638 85926 54650 85978
rect 54702 85926 54714 85978
rect 54766 85926 54778 85978
rect 54830 85926 72922 85978
rect 72974 85926 72986 85978
rect 73038 85926 73050 85978
rect 73102 85926 73114 85978
rect 73166 85926 73178 85978
rect 73230 85926 88596 85978
rect 4876 85904 88596 85926
rect 4876 85434 88596 85456
rect 4876 85382 18382 85434
rect 18434 85382 18446 85434
rect 18498 85382 18510 85434
rect 18562 85382 18574 85434
rect 18626 85382 18638 85434
rect 18690 85382 36782 85434
rect 36834 85382 36846 85434
rect 36898 85382 36910 85434
rect 36962 85382 36974 85434
rect 37026 85382 37038 85434
rect 37090 85382 55182 85434
rect 55234 85382 55246 85434
rect 55298 85382 55310 85434
rect 55362 85382 55374 85434
rect 55426 85382 55438 85434
rect 55490 85382 73582 85434
rect 73634 85382 73646 85434
rect 73698 85382 73710 85434
rect 73762 85382 73774 85434
rect 73826 85382 73838 85434
rect 73890 85382 88596 85434
rect 4876 85360 88596 85382
rect 41818 84976 41824 85028
rect 41876 85016 41882 85028
rect 49086 85016 49092 85028
rect 41876 84988 49092 85016
rect 41876 84976 41882 84988
rect 49086 84976 49092 84988
rect 49144 84976 49150 85028
rect 4876 84890 88596 84912
rect 4876 84838 5954 84890
rect 6006 84838 6018 84890
rect 6070 84838 6082 84890
rect 6134 84838 6146 84890
rect 6198 84838 6210 84890
rect 6262 84838 17722 84890
rect 17774 84838 17786 84890
rect 17838 84838 17850 84890
rect 17902 84838 17914 84890
rect 17966 84838 17978 84890
rect 18030 84838 36122 84890
rect 36174 84838 36186 84890
rect 36238 84838 36250 84890
rect 36302 84838 36314 84890
rect 36366 84838 36378 84890
rect 36430 84838 54522 84890
rect 54574 84838 54586 84890
rect 54638 84838 54650 84890
rect 54702 84838 54714 84890
rect 54766 84838 54778 84890
rect 54830 84838 72922 84890
rect 72974 84838 72986 84890
rect 73038 84838 73050 84890
rect 73102 84838 73114 84890
rect 73166 84838 73178 84890
rect 73230 84838 86546 84890
rect 86598 84838 86610 84890
rect 86662 84838 86674 84890
rect 86726 84838 86738 84890
rect 86790 84838 86802 84890
rect 86854 84838 88596 84890
rect 4876 84816 88596 84838
rect 30686 84744 30692 84756
rect 27806 84716 30692 84744
rect 12746 84636 12752 84688
rect 12804 84676 12810 84688
rect 12841 84679 12899 84685
rect 12841 84676 12853 84679
rect 12804 84648 12853 84676
rect 12804 84636 12810 84648
rect 12841 84645 12853 84648
rect 12887 84676 12899 84679
rect 27806 84676 27834 84716
rect 30686 84704 30692 84716
rect 30744 84704 30750 84756
rect 31057 84747 31115 84753
rect 31057 84744 31069 84747
rect 30980 84716 31069 84744
rect 12887 84648 27834 84676
rect 12887 84645 12899 84648
rect 12841 84639 12899 84645
rect 11642 84568 11648 84620
rect 11700 84608 11706 84620
rect 11737 84611 11795 84617
rect 11737 84608 11749 84611
rect 11700 84580 11749 84608
rect 11700 84568 11706 84580
rect 11737 84577 11749 84580
rect 11783 84608 11795 84611
rect 30686 84608 30692 84620
rect 11783 84580 30692 84608
rect 11783 84577 11795 84580
rect 11737 84571 11795 84577
rect 30686 84568 30692 84580
rect 30744 84568 30750 84620
rect 30980 84608 31008 84716
rect 31057 84713 31069 84716
rect 31103 84744 31115 84747
rect 39610 84744 39616 84756
rect 31103 84716 39616 84744
rect 31103 84713 31115 84716
rect 31057 84707 31115 84713
rect 39610 84704 39616 84716
rect 39668 84704 39674 84756
rect 45409 84747 45467 84753
rect 45409 84713 45421 84747
rect 45455 84744 45467 84747
rect 46142 84744 46148 84756
rect 45455 84716 46148 84744
rect 45455 84713 45467 84716
rect 45409 84707 45467 84713
rect 46142 84704 46148 84716
rect 46200 84704 46206 84756
rect 31238 84636 31244 84688
rect 31296 84676 31302 84688
rect 39058 84676 39064 84688
rect 31296 84648 39064 84676
rect 31296 84636 31302 84648
rect 39058 84636 39064 84648
rect 39116 84676 39122 84688
rect 50190 84676 50196 84688
rect 39116 84648 50196 84676
rect 39116 84636 39122 84648
rect 50190 84636 50196 84648
rect 50248 84636 50254 84688
rect 30796 84580 31008 84608
rect 7410 84500 7416 84552
rect 7468 84540 7474 84552
rect 30573 84543 30631 84549
rect 7468 84512 29996 84540
rect 7468 84500 7474 84512
rect 10538 84432 10544 84484
rect 10596 84472 10602 84484
rect 10633 84475 10691 84481
rect 10633 84472 10645 84475
rect 10596 84444 10645 84472
rect 10596 84432 10602 84444
rect 10633 84441 10645 84444
rect 10679 84441 10691 84475
rect 10633 84435 10691 84441
rect 13850 84432 13856 84484
rect 13908 84472 13914 84484
rect 29968 84481 29996 84512
rect 30573 84509 30585 84543
rect 30619 84540 30631 84543
rect 30796 84540 30824 84580
rect 31146 84568 31152 84620
rect 31204 84608 31210 84620
rect 41818 84608 41824 84620
rect 31204 84580 41824 84608
rect 31204 84568 31210 84580
rect 41818 84568 41824 84580
rect 41876 84568 41882 84620
rect 45593 84611 45651 84617
rect 45593 84577 45605 84611
rect 45639 84608 45651 84611
rect 46050 84608 46056 84620
rect 45639 84580 46056 84608
rect 45639 84577 45651 84580
rect 45593 84571 45651 84577
rect 46050 84568 46056 84580
rect 46108 84568 46114 84620
rect 46142 84568 46148 84620
rect 46200 84608 46206 84620
rect 51294 84608 51300 84620
rect 46200 84580 51300 84608
rect 46200 84568 46206 84580
rect 51294 84568 51300 84580
rect 51352 84608 51358 84620
rect 51389 84611 51447 84617
rect 51389 84608 51401 84611
rect 51352 84580 51401 84608
rect 51352 84568 51358 84580
rect 51389 84577 51401 84580
rect 51435 84577 51447 84611
rect 51389 84571 51447 84577
rect 30619 84512 30824 84540
rect 30873 84543 30931 84549
rect 30619 84509 30631 84512
rect 30573 84503 30631 84509
rect 30873 84509 30885 84543
rect 30919 84540 30931 84543
rect 41037 84543 41095 84549
rect 41037 84540 41049 84543
rect 30919 84512 37494 84540
rect 30919 84509 30931 84512
rect 30873 84503 30931 84509
rect 13945 84475 14003 84481
rect 13945 84472 13957 84475
rect 13908 84444 13957 84472
rect 13908 84432 13914 84444
rect 13945 84441 13957 84444
rect 13991 84441 14003 84475
rect 13945 84435 14003 84441
rect 29953 84475 30011 84481
rect 29953 84441 29965 84475
rect 29999 84472 30011 84475
rect 30888 84472 30916 84503
rect 29999 84444 30916 84472
rect 37466 84472 37494 84512
rect 40824 84512 41049 84540
rect 40824 84481 40852 84512
rect 41037 84509 41049 84512
rect 41083 84509 41095 84543
rect 41037 84503 41095 84509
rect 42741 84543 42799 84549
rect 42741 84509 42753 84543
rect 42787 84540 42799 84543
rect 42925 84543 42983 84549
rect 42925 84540 42937 84543
rect 42787 84512 42937 84540
rect 42787 84509 42799 84512
rect 42741 84503 42799 84509
rect 42925 84509 42937 84512
rect 42971 84540 42983 84543
rect 47154 84540 47160 84552
rect 42971 84512 47160 84540
rect 42971 84509 42983 84512
rect 42925 84503 42983 84509
rect 47154 84500 47160 84512
rect 47212 84540 47218 84552
rect 48077 84543 48135 84549
rect 48077 84540 48089 84543
rect 47212 84512 48089 84540
rect 47212 84500 47218 84512
rect 48077 84509 48089 84512
rect 48123 84509 48135 84543
rect 48077 84503 48135 84509
rect 40809 84475 40867 84481
rect 40809 84472 40821 84475
rect 37466 84444 40821 84472
rect 29999 84441 30011 84444
rect 29953 84435 30011 84441
rect 40809 84441 40821 84444
rect 40855 84441 40867 84475
rect 40809 84435 40867 84441
rect 45777 84475 45835 84481
rect 45777 84441 45789 84475
rect 45823 84472 45835 84475
rect 45866 84472 45872 84484
rect 45823 84444 45872 84472
rect 45823 84441 45835 84444
rect 45777 84435 45835 84441
rect 45866 84432 45872 84444
rect 45924 84432 45930 84484
rect 45958 84432 45964 84484
rect 46016 84432 46022 84484
rect 49086 84432 49092 84484
rect 49144 84472 49150 84484
rect 49181 84475 49239 84481
rect 49181 84472 49193 84475
rect 49144 84444 49193 84472
rect 49144 84432 49150 84444
rect 49181 84441 49193 84444
rect 49227 84441 49239 84475
rect 49181 84435 49239 84441
rect 50190 84432 50196 84484
rect 50248 84472 50254 84484
rect 50285 84475 50343 84481
rect 50285 84472 50297 84475
rect 50248 84444 50297 84472
rect 50248 84432 50254 84444
rect 50285 84441 50297 84444
rect 50331 84441 50343 84475
rect 50285 84435 50343 84441
rect 4876 84346 88596 84368
rect 4876 84294 6690 84346
rect 6742 84294 6754 84346
rect 6806 84294 6818 84346
rect 6870 84294 6882 84346
rect 6934 84294 6946 84346
rect 6998 84294 18382 84346
rect 18434 84294 18446 84346
rect 18498 84294 18510 84346
rect 18562 84294 18574 84346
rect 18626 84294 18638 84346
rect 18690 84294 36782 84346
rect 36834 84294 36846 84346
rect 36898 84294 36910 84346
rect 36962 84294 36974 84346
rect 37026 84294 37038 84346
rect 37090 84294 55182 84346
rect 55234 84294 55246 84346
rect 55298 84294 55310 84346
rect 55362 84294 55374 84346
rect 55426 84294 55438 84346
rect 55490 84294 73582 84346
rect 73634 84294 73646 84346
rect 73698 84294 73710 84346
rect 73762 84294 73774 84346
rect 73826 84294 73838 84346
rect 73890 84294 87282 84346
rect 87334 84294 87346 84346
rect 87398 84294 87410 84346
rect 87462 84294 87474 84346
rect 87526 84294 87538 84346
rect 87590 84294 88596 84346
rect 4876 84272 88596 84294
rect 4876 83802 7912 83824
rect 4876 83750 5954 83802
rect 6006 83750 6018 83802
rect 6070 83750 6082 83802
rect 6134 83750 6146 83802
rect 6198 83750 6210 83802
rect 6262 83750 7912 83802
rect 4876 83728 7912 83750
rect 85284 83802 88596 83824
rect 85284 83750 86546 83802
rect 86598 83750 86610 83802
rect 86662 83750 86674 83802
rect 86726 83750 86738 83802
rect 86790 83750 86802 83802
rect 86854 83750 88596 83802
rect 85284 83728 88596 83750
rect 4876 83258 7912 83280
rect 4876 83206 6690 83258
rect 6742 83206 6754 83258
rect 6806 83206 6818 83258
rect 6870 83206 6882 83258
rect 6934 83206 6946 83258
rect 6998 83206 7912 83258
rect 4876 83184 7912 83206
rect 85284 83258 88596 83280
rect 85284 83206 87282 83258
rect 87334 83206 87346 83258
rect 87398 83206 87410 83258
rect 87462 83206 87474 83258
rect 87526 83206 87538 83258
rect 87590 83206 88596 83258
rect 85284 83184 88596 83206
rect 13850 83072 13856 83124
rect 13908 83112 13914 83124
rect 83310 83112 83316 83124
rect 13908 83084 83316 83112
rect 13908 83072 13914 83084
rect 83310 83072 83316 83084
rect 83368 83072 83374 83124
rect 47062 83004 47068 83056
rect 47120 83044 47126 83056
rect 47154 83044 47160 83056
rect 47120 83016 47160 83044
rect 47120 83004 47126 83016
rect 47154 83004 47160 83016
rect 47212 83044 47218 83056
rect 47982 83044 47988 83056
rect 47212 83016 47988 83044
rect 47212 83004 47218 83016
rect 47982 83004 47988 83016
rect 48040 83004 48046 83056
rect 4876 82714 7912 82736
rect 4876 82662 5954 82714
rect 6006 82662 6018 82714
rect 6070 82662 6082 82714
rect 6134 82662 6146 82714
rect 6198 82662 6210 82714
rect 6262 82662 7912 82714
rect 4876 82640 7912 82662
rect 85284 82714 88596 82736
rect 85284 82662 86546 82714
rect 86598 82662 86610 82714
rect 86662 82662 86674 82714
rect 86726 82662 86738 82714
rect 86790 82662 86802 82714
rect 86854 82662 88596 82714
rect 85284 82640 88596 82662
rect 14982 82392 14988 82444
rect 15040 82432 15046 82444
rect 15506 82432 15512 82444
rect 15040 82404 15512 82432
rect 15040 82392 15046 82404
rect 15506 82392 15512 82404
rect 15564 82392 15570 82444
rect 68942 82392 68948 82444
rect 69000 82432 69006 82444
rect 69326 82432 69332 82444
rect 69000 82404 69332 82432
rect 69000 82392 69006 82404
rect 69326 82392 69332 82404
rect 69384 82392 69390 82444
rect 7594 82324 7600 82376
rect 7652 82364 7658 82376
rect 11670 82364 11676 82376
rect 7652 82336 11676 82364
rect 7652 82324 7658 82336
rect 11670 82324 11676 82336
rect 11728 82324 11734 82376
rect 7226 82256 7232 82308
rect 7284 82296 7290 82308
rect 12774 82296 12780 82308
rect 7284 82268 12780 82296
rect 7284 82256 7290 82268
rect 12774 82256 12780 82268
rect 12832 82256 12838 82308
rect 4876 82170 7912 82192
rect 4876 82118 6690 82170
rect 6742 82118 6754 82170
rect 6806 82118 6818 82170
rect 6870 82118 6882 82170
rect 6934 82118 6946 82170
rect 6998 82118 7912 82170
rect 4876 82096 7912 82118
rect 85284 82170 88596 82192
rect 85284 82118 87282 82170
rect 87334 82118 87346 82170
rect 87398 82118 87410 82170
rect 87462 82118 87474 82170
rect 87526 82118 87538 82170
rect 87590 82118 88596 82170
rect 85284 82096 88596 82118
rect 7778 81712 7784 81764
rect 7836 81752 7842 81764
rect 9986 81752 9992 81764
rect 7836 81724 9992 81752
rect 7836 81712 7842 81724
rect 9986 81712 9992 81724
rect 10044 81712 10050 81764
rect 4876 81626 7912 81648
rect 4876 81574 5954 81626
rect 6006 81574 6018 81626
rect 6070 81574 6082 81626
rect 6134 81574 6146 81626
rect 6198 81574 6210 81626
rect 6262 81574 7912 81626
rect 4876 81552 7912 81574
rect 85284 81626 88596 81648
rect 85284 81574 86546 81626
rect 86598 81574 86610 81626
rect 86662 81574 86674 81626
rect 86726 81574 86738 81626
rect 86790 81574 86802 81626
rect 86854 81574 88596 81626
rect 85284 81552 88596 81574
rect 83494 81372 83500 81424
rect 83552 81412 83558 81424
rect 88051 81415 88109 81421
rect 88051 81412 88063 81415
rect 83552 81384 88063 81412
rect 83552 81372 83558 81384
rect 88051 81381 88063 81384
rect 88097 81381 88109 81415
rect 88051 81375 88109 81381
rect 88253 81313 88311 81319
rect 88253 81310 88265 81313
rect 87729 81279 87787 81285
rect 87729 81245 87741 81279
rect 87775 81276 87787 81279
rect 88112 81282 88265 81310
rect 88112 81276 88140 81282
rect 87775 81248 88140 81276
rect 88253 81279 88265 81282
rect 88299 81310 88311 81313
rect 88299 81296 88416 81310
rect 88299 81282 88376 81296
rect 88299 81279 88311 81282
rect 88253 81273 88311 81279
rect 87775 81245 87787 81248
rect 87729 81239 87787 81245
rect 88370 81244 88376 81282
rect 88428 81244 88434 81296
rect 4876 81082 7912 81104
rect 4876 81030 6690 81082
rect 6742 81030 6754 81082
rect 6806 81030 6818 81082
rect 6870 81030 6882 81082
rect 6934 81030 6946 81082
rect 6998 81030 7912 81082
rect 4876 81008 7912 81030
rect 85284 81082 88596 81104
rect 85284 81030 87282 81082
rect 87334 81030 87346 81082
rect 87398 81030 87410 81082
rect 87462 81030 87474 81082
rect 87526 81030 87538 81082
rect 87590 81030 88596 81082
rect 85284 81008 88596 81030
rect 4876 80538 7912 80560
rect 4876 80486 5954 80538
rect 6006 80486 6018 80538
rect 6070 80486 6082 80538
rect 6134 80486 6146 80538
rect 6198 80486 6210 80538
rect 6262 80486 7912 80538
rect 4876 80464 7912 80486
rect 85284 80538 88596 80560
rect 85284 80486 86546 80538
rect 86598 80486 86610 80538
rect 86662 80486 86674 80538
rect 86726 80486 86738 80538
rect 86790 80486 86802 80538
rect 86854 80486 88596 80538
rect 85284 80464 88596 80486
rect 87729 80259 87787 80265
rect 5457 80225 5515 80231
rect 5457 80191 5469 80225
rect 5503 80191 5515 80225
rect 87729 80225 87741 80259
rect 87775 80256 87787 80259
rect 87775 80234 88300 80256
rect 87775 80228 88284 80234
rect 87775 80225 87787 80228
rect 87729 80219 87787 80225
rect 88253 80225 88284 80228
rect 5457 80188 5515 80191
rect 7134 80188 7140 80200
rect 5457 80185 7140 80188
rect 5472 80160 7140 80185
rect 7134 80148 7140 80160
rect 7192 80148 7198 80200
rect 83494 80148 83500 80200
rect 83552 80188 83558 80200
rect 88253 80191 88265 80225
rect 83552 80160 88094 80188
rect 88253 80185 88284 80191
rect 88278 80182 88284 80185
rect 88336 80182 88342 80234
rect 83552 80148 83558 80160
rect 2902 80080 2908 80132
rect 2960 80120 2966 80132
rect 88066 80129 88094 80160
rect 5251 80123 5309 80129
rect 5251 80120 5263 80123
rect 2960 80092 5263 80120
rect 2960 80080 2966 80092
rect 5251 80089 5263 80092
rect 5297 80089 5309 80123
rect 5251 80083 5309 80089
rect 88051 80123 88109 80129
rect 88051 80089 88063 80123
rect 88097 80089 88109 80123
rect 88051 80083 88109 80089
rect 4876 79994 7912 80016
rect 4876 79942 6690 79994
rect 6742 79942 6754 79994
rect 6806 79942 6818 79994
rect 6870 79942 6882 79994
rect 6934 79942 6946 79994
rect 6998 79942 7912 79994
rect 4876 79920 7912 79942
rect 85284 79994 88596 80016
rect 85284 79942 87282 79994
rect 87334 79942 87346 79994
rect 87398 79942 87410 79994
rect 87462 79942 87474 79994
rect 87526 79942 87538 79994
rect 87590 79942 88596 79994
rect 85284 79920 88596 79942
rect 4876 79450 7912 79472
rect 4876 79398 5954 79450
rect 6006 79398 6018 79450
rect 6070 79398 6082 79450
rect 6134 79398 6146 79450
rect 6198 79398 6210 79450
rect 6262 79398 7912 79450
rect 4876 79376 7912 79398
rect 85284 79450 88596 79472
rect 85284 79398 86546 79450
rect 86598 79398 86610 79450
rect 86662 79398 86674 79450
rect 86726 79398 86738 79450
rect 86790 79398 86802 79450
rect 86854 79398 88596 79450
rect 85284 79376 88596 79398
rect 4876 78906 7912 78928
rect 4876 78854 6690 78906
rect 6742 78854 6754 78906
rect 6806 78854 6818 78906
rect 6870 78854 6882 78906
rect 6934 78854 6946 78906
rect 6998 78854 7912 78906
rect 4876 78832 7912 78854
rect 85284 78906 88596 78928
rect 85284 78854 87282 78906
rect 87334 78854 87346 78906
rect 87398 78854 87410 78906
rect 87462 78854 87474 78906
rect 87526 78854 87538 78906
rect 87590 78854 88596 78906
rect 85284 78832 88596 78854
rect 7134 78692 7140 78704
rect 5472 78667 7140 78692
rect 5457 78664 7140 78667
rect 5457 78661 5515 78664
rect 5457 78627 5469 78661
rect 5503 78627 5515 78661
rect 7134 78652 7140 78664
rect 7192 78652 7198 78704
rect 88278 78667 88284 78670
rect 88253 78661 88284 78667
rect 88253 78658 88265 78661
rect 87928 78633 88265 78658
rect 5457 78621 5515 78627
rect 87913 78630 88265 78633
rect 87913 78627 87971 78630
rect 87913 78593 87925 78627
rect 87959 78593 87971 78627
rect 88253 78627 88265 78630
rect 88253 78621 88284 78627
rect 88278 78618 88284 78621
rect 88336 78618 88342 78670
rect 87913 78587 87971 78593
rect 88002 78516 88008 78568
rect 88060 78565 88066 78568
rect 88060 78559 88109 78565
rect 88060 78525 88063 78559
rect 88097 78525 88109 78559
rect 88060 78519 88109 78525
rect 88060 78516 88066 78519
rect 2902 78448 2908 78500
rect 2960 78488 2966 78500
rect 5251 78491 5309 78497
rect 5251 78488 5263 78491
rect 2960 78460 5263 78488
rect 2960 78448 2966 78460
rect 5251 78457 5263 78460
rect 5297 78457 5309 78491
rect 5251 78451 5309 78457
rect 4876 78362 7912 78384
rect 4876 78310 5954 78362
rect 6006 78310 6018 78362
rect 6070 78310 6082 78362
rect 6134 78310 6146 78362
rect 6198 78310 6210 78362
rect 6262 78310 7912 78362
rect 4876 78288 7912 78310
rect 85284 78362 88596 78384
rect 85284 78310 86546 78362
rect 86598 78310 86610 78362
rect 86662 78310 86674 78362
rect 86726 78310 86738 78362
rect 86790 78310 86802 78362
rect 86854 78310 88596 78362
rect 85284 78288 88596 78310
rect 88278 78055 88284 78058
rect 5457 78049 5515 78055
rect 5457 78015 5469 78049
rect 5503 78015 5515 78049
rect 88253 78049 88284 78055
rect 88253 78046 88265 78049
rect 5457 78012 5515 78015
rect 7134 78012 7140 78024
rect 5457 78009 7140 78012
rect 5472 77984 7140 78009
rect 7134 77972 7140 77984
rect 7192 77972 7198 78024
rect 87729 78015 87787 78021
rect 87729 77981 87741 78015
rect 87775 78012 87787 78015
rect 88112 78018 88265 78046
rect 88112 78012 88140 78018
rect 87775 77984 88140 78012
rect 88253 78015 88265 78018
rect 88253 78009 88284 78015
rect 88278 78006 88284 78009
rect 88336 78006 88342 78058
rect 87775 77981 87787 77984
rect 87729 77975 87787 77981
rect 2902 77904 2908 77956
rect 2960 77944 2966 77956
rect 5251 77947 5309 77953
rect 5251 77944 5263 77947
rect 2960 77916 5263 77944
rect 2960 77904 2966 77916
rect 5251 77913 5263 77916
rect 5297 77913 5309 77947
rect 5251 77907 5309 77913
rect 87818 77904 87824 77956
rect 87876 77944 87882 77956
rect 88051 77947 88109 77953
rect 88051 77944 88063 77947
rect 87876 77916 88063 77944
rect 87876 77904 87882 77916
rect 88051 77913 88063 77916
rect 88097 77913 88109 77947
rect 88051 77907 88109 77913
rect 4876 77818 7912 77840
rect 4876 77766 6690 77818
rect 6742 77766 6754 77818
rect 6806 77766 6818 77818
rect 6870 77766 6882 77818
rect 6934 77766 6946 77818
rect 6998 77766 7912 77818
rect 4876 77744 7912 77766
rect 85284 77818 88596 77840
rect 85284 77766 87282 77818
rect 87334 77766 87346 77818
rect 87398 77766 87410 77818
rect 87462 77766 87474 77818
rect 87526 77766 87538 77818
rect 87590 77766 88596 77818
rect 85284 77744 88596 77766
rect 4876 77274 7912 77296
rect 4876 77222 5954 77274
rect 6006 77222 6018 77274
rect 6070 77222 6082 77274
rect 6134 77222 6146 77274
rect 6198 77222 6210 77274
rect 6262 77222 7912 77274
rect 4876 77200 7912 77222
rect 85284 77274 88596 77296
rect 85284 77222 86546 77274
rect 86598 77222 86610 77274
rect 86662 77222 86674 77274
rect 86726 77222 86738 77274
rect 86790 77222 86802 77274
rect 86854 77222 88596 77274
rect 85284 77200 88596 77222
rect 87797 76995 87855 77001
rect 5457 76961 5515 76967
rect 5457 76927 5469 76961
rect 5503 76927 5515 76961
rect 87797 76961 87809 76995
rect 87843 76992 87855 76995
rect 87843 76964 88048 76992
rect 87843 76961 87855 76964
rect 87797 76955 87855 76961
rect 5457 76924 5515 76927
rect 7134 76924 7140 76936
rect 5457 76921 7140 76924
rect 5472 76896 7140 76921
rect 7134 76884 7140 76896
rect 7192 76884 7198 76936
rect 88020 76868 88048 76964
rect 2718 76816 2724 76868
rect 2776 76856 2782 76868
rect 5251 76859 5309 76865
rect 5251 76856 5263 76859
rect 2776 76828 5263 76856
rect 2776 76816 2782 76828
rect 5251 76825 5263 76828
rect 5297 76825 5309 76859
rect 5251 76819 5309 76825
rect 86622 76816 86628 76868
rect 86680 76856 86686 76868
rect 87545 76859 87603 76865
rect 87545 76856 87557 76859
rect 86680 76828 87557 76856
rect 86680 76816 86686 76828
rect 87545 76825 87557 76828
rect 87591 76825 87603 76859
rect 87545 76819 87603 76825
rect 88002 76816 88008 76868
rect 88060 76816 88066 76868
rect 4876 76730 7912 76752
rect 4876 76678 6690 76730
rect 6742 76678 6754 76730
rect 6806 76678 6818 76730
rect 6870 76678 6882 76730
rect 6934 76678 6946 76730
rect 6998 76678 7912 76730
rect 4876 76656 7912 76678
rect 85284 76730 88596 76752
rect 85284 76678 87282 76730
rect 87334 76678 87346 76730
rect 87398 76678 87410 76730
rect 87462 76678 87474 76730
rect 87526 76678 87538 76730
rect 87590 76678 88596 76730
rect 85284 76656 88596 76678
rect 4876 76186 7912 76208
rect 4876 76134 5954 76186
rect 6006 76134 6018 76186
rect 6070 76134 6082 76186
rect 6134 76134 6146 76186
rect 6198 76134 6210 76186
rect 6262 76134 7912 76186
rect 4876 76112 7912 76134
rect 85284 76186 88596 76208
rect 85284 76134 86546 76186
rect 86598 76134 86610 76186
rect 86662 76134 86674 76186
rect 86726 76134 86738 76186
rect 86790 76134 86802 76186
rect 86854 76134 88596 76186
rect 85284 76112 88596 76134
rect 86898 75932 86904 75984
rect 86956 75972 86962 75984
rect 88051 75975 88109 75981
rect 88051 75972 88063 75975
rect 86956 75944 88063 75972
rect 86956 75932 86962 75944
rect 88051 75941 88063 75944
rect 88097 75941 88109 75975
rect 88051 75935 88109 75941
rect 87729 75907 87787 75913
rect 5457 75873 5515 75879
rect 5457 75839 5469 75873
rect 5503 75870 5515 75873
rect 87729 75873 87741 75907
rect 87775 75904 87787 75907
rect 87775 75876 88324 75904
rect 87775 75873 87787 75876
rect 5503 75842 5800 75870
rect 87729 75867 87787 75873
rect 88257 75873 88324 75876
rect 5503 75839 5515 75842
rect 5457 75833 5515 75839
rect 5772 75836 5800 75842
rect 7134 75836 7140 75848
rect 5772 75808 7140 75836
rect 7134 75796 7140 75808
rect 7192 75796 7198 75848
rect 88257 75839 88269 75873
rect 88303 75870 88324 75873
rect 88303 75848 88508 75870
rect 88303 75842 88468 75848
rect 88303 75839 88315 75842
rect 88257 75833 88315 75839
rect 88462 75796 88468 75842
rect 88520 75796 88526 75848
rect 2902 75728 2908 75780
rect 2960 75768 2966 75780
rect 5251 75771 5309 75777
rect 5251 75768 5263 75771
rect 2960 75740 5263 75768
rect 2960 75728 2966 75740
rect 5251 75737 5263 75740
rect 5297 75737 5309 75771
rect 5251 75731 5309 75737
rect 4876 75642 7912 75664
rect 4876 75590 6690 75642
rect 6742 75590 6754 75642
rect 6806 75590 6818 75642
rect 6870 75590 6882 75642
rect 6934 75590 6946 75642
rect 6998 75590 7912 75642
rect 4876 75568 7912 75590
rect 85284 75642 88596 75664
rect 85284 75590 87282 75642
rect 87334 75590 87346 75642
rect 87398 75590 87410 75642
rect 87462 75590 87474 75642
rect 87526 75590 87538 75642
rect 87590 75590 88596 75642
rect 85284 75568 88596 75590
rect 4876 75098 7912 75120
rect 4876 75046 5954 75098
rect 6006 75046 6018 75098
rect 6070 75046 6082 75098
rect 6134 75046 6146 75098
rect 6198 75046 6210 75098
rect 6262 75046 7912 75098
rect 4876 75024 7912 75046
rect 85284 75098 88596 75120
rect 85284 75046 86546 75098
rect 86598 75046 86610 75098
rect 86662 75046 86674 75098
rect 86726 75046 86738 75098
rect 86790 75046 86802 75098
rect 86854 75046 88596 75098
rect 85284 75024 88596 75046
rect 4374 74844 4380 74896
rect 4432 74884 4438 74896
rect 5251 74887 5309 74893
rect 5251 74884 5263 74887
rect 4432 74856 5263 74884
rect 4432 74844 4438 74856
rect 5251 74853 5263 74856
rect 5297 74853 5309 74887
rect 5251 74847 5309 74853
rect 84414 74844 84420 74896
rect 84472 74884 84478 74896
rect 88051 74887 88109 74893
rect 88051 74884 88063 74887
rect 84472 74856 88063 74884
rect 84472 74844 84478 74856
rect 88051 74853 88063 74856
rect 88097 74853 88109 74887
rect 88051 74847 88109 74853
rect 87729 74819 87787 74825
rect 5457 74785 5515 74791
rect 5457 74751 5469 74785
rect 5503 74782 5515 74785
rect 5662 74782 5668 74794
rect 5503 74754 5668 74782
rect 5503 74751 5515 74754
rect 5457 74745 5515 74751
rect 5662 74742 5668 74754
rect 5720 74742 5726 74794
rect 87729 74785 87741 74819
rect 87775 74816 87787 74819
rect 87775 74788 88140 74816
rect 87775 74785 87787 74788
rect 87729 74779 87787 74785
rect 88112 74782 88140 74788
rect 88257 74785 88315 74791
rect 88257 74782 88269 74785
rect 88112 74754 88269 74782
rect 88257 74751 88269 74754
rect 88303 74782 88315 74785
rect 88554 74782 88560 74828
rect 88303 74776 88560 74782
rect 88612 74776 88618 74828
rect 88303 74754 88600 74776
rect 88303 74751 88315 74754
rect 88257 74745 88315 74751
rect 4876 74554 7912 74576
rect 4876 74502 6690 74554
rect 6742 74502 6754 74554
rect 6806 74502 6818 74554
rect 6870 74502 6882 74554
rect 6934 74502 6946 74554
rect 6998 74502 7912 74554
rect 4876 74480 7912 74502
rect 85284 74554 88596 74576
rect 85284 74502 87282 74554
rect 87334 74502 87346 74554
rect 87398 74502 87410 74554
rect 87462 74502 87474 74554
rect 87526 74502 87538 74554
rect 87590 74502 88596 74554
rect 85284 74480 88596 74502
rect 4876 74010 7912 74032
rect 4876 73958 5954 74010
rect 6006 73958 6018 74010
rect 6070 73958 6082 74010
rect 6134 73958 6146 74010
rect 6198 73958 6210 74010
rect 6262 73958 7912 74010
rect 4876 73936 7912 73958
rect 85284 74010 88596 74032
rect 85284 73958 86546 74010
rect 86598 73958 86610 74010
rect 86662 73958 86674 74010
rect 86726 73958 86738 74010
rect 86790 73958 86802 74010
rect 86854 73958 88596 74010
rect 85284 73936 88596 73958
rect 4876 73466 7912 73488
rect 4876 73414 6690 73466
rect 6742 73414 6754 73466
rect 6806 73414 6818 73466
rect 6870 73414 6882 73466
rect 6934 73414 6946 73466
rect 6998 73414 7912 73466
rect 4876 73392 7912 73414
rect 85284 73466 88596 73488
rect 85284 73414 87282 73466
rect 87334 73414 87346 73466
rect 87398 73414 87410 73466
rect 87462 73414 87474 73466
rect 87526 73414 87538 73466
rect 87590 73414 88596 73466
rect 85284 73392 88596 73414
rect 7134 73252 7140 73264
rect 5457 73221 5515 73227
rect 5457 73187 5469 73221
rect 5503 73218 5515 73221
rect 5772 73224 7140 73252
rect 5772 73218 5800 73224
rect 5503 73190 5800 73218
rect 7134 73212 7140 73224
rect 7192 73212 7198 73264
rect 88278 73227 88284 73230
rect 88253 73221 88284 73227
rect 5503 73187 5515 73190
rect 5457 73181 5515 73187
rect 88002 73144 88008 73196
rect 88060 73193 88066 73196
rect 88060 73187 88109 73193
rect 88060 73153 88063 73187
rect 88097 73153 88109 73187
rect 88253 73187 88265 73221
rect 88253 73181 88284 73187
rect 88278 73178 88284 73181
rect 88336 73178 88342 73230
rect 88060 73147 88109 73153
rect 88060 73144 88066 73147
rect 87913 73119 87971 73125
rect 87913 73085 87925 73119
rect 87959 73116 87971 73119
rect 88296 73116 88324 73178
rect 87959 73088 88324 73116
rect 87959 73085 87971 73088
rect 87913 73079 87971 73085
rect 2902 73008 2908 73060
rect 2960 73048 2966 73060
rect 5251 73051 5309 73057
rect 5251 73048 5263 73051
rect 2960 73020 5263 73048
rect 2960 73008 2966 73020
rect 5251 73017 5263 73020
rect 5297 73017 5309 73051
rect 5251 73011 5309 73017
rect 4876 72922 7912 72944
rect 4876 72870 5954 72922
rect 6006 72870 6018 72922
rect 6070 72870 6082 72922
rect 6134 72870 6146 72922
rect 6198 72870 6210 72922
rect 6262 72870 7912 72922
rect 4876 72848 7912 72870
rect 85284 72922 88596 72944
rect 85284 72870 86546 72922
rect 86598 72870 86610 72922
rect 86662 72870 86674 72922
rect 86726 72870 86738 72922
rect 86790 72870 86802 72922
rect 86854 72870 88596 72922
rect 85284 72848 88596 72870
rect 5457 72609 5515 72615
rect 88278 72609 88284 72612
rect 5457 72575 5469 72609
rect 5503 72606 5515 72609
rect 5503 72578 5800 72606
rect 88253 72603 88284 72609
rect 5503 72575 5515 72578
rect 5457 72569 5515 72575
rect 5772 72572 5800 72578
rect 7134 72572 7140 72584
rect 5772 72544 7140 72572
rect 7134 72532 7140 72544
rect 7192 72532 7198 72584
rect 87174 72532 87180 72584
rect 87232 72572 87238 72584
rect 88051 72575 88109 72581
rect 88051 72572 88063 72575
rect 87232 72544 88063 72572
rect 87232 72532 87238 72544
rect 88051 72541 88063 72544
rect 88097 72541 88109 72575
rect 88253 72569 88265 72603
rect 88253 72563 88284 72569
rect 88278 72560 88284 72563
rect 88336 72560 88342 72612
rect 88051 72535 88109 72541
rect 2902 72464 2908 72516
rect 2960 72504 2966 72516
rect 5251 72507 5309 72513
rect 5251 72504 5263 72507
rect 2960 72476 5263 72504
rect 2960 72464 2966 72476
rect 5251 72473 5263 72476
rect 5297 72473 5309 72507
rect 5251 72467 5309 72473
rect 87729 72507 87787 72513
rect 87729 72473 87741 72507
rect 87775 72504 87787 72507
rect 88296 72504 88324 72560
rect 87775 72476 88324 72504
rect 87775 72473 87787 72476
rect 87729 72467 87787 72473
rect 4876 72378 7912 72400
rect 4876 72326 6690 72378
rect 6742 72326 6754 72378
rect 6806 72326 6818 72378
rect 6870 72326 6882 72378
rect 6934 72326 6946 72378
rect 6998 72326 7912 72378
rect 4876 72304 7912 72326
rect 85284 72378 88596 72400
rect 85284 72326 87282 72378
rect 87334 72326 87346 72378
rect 87398 72326 87410 72378
rect 87462 72326 87474 72378
rect 87526 72326 87538 72378
rect 87590 72326 88596 72378
rect 85284 72304 88596 72326
rect 4876 71834 7912 71856
rect 4876 71782 5954 71834
rect 6006 71782 6018 71834
rect 6070 71782 6082 71834
rect 6134 71782 6146 71834
rect 6198 71782 6210 71834
rect 6262 71782 7912 71834
rect 4876 71760 7912 71782
rect 85284 71834 88596 71856
rect 85284 71782 86546 71834
rect 86598 71782 86610 71834
rect 86662 71782 86674 71834
rect 86726 71782 86738 71834
rect 86790 71782 86802 71834
rect 86854 71782 88596 71834
rect 85284 71760 88596 71782
rect 86898 71580 86904 71632
rect 86956 71620 86962 71632
rect 88051 71623 88109 71629
rect 88051 71620 88063 71623
rect 86956 71592 88063 71620
rect 86956 71580 86962 71592
rect 88051 71589 88063 71592
rect 88097 71589 88109 71623
rect 88051 71583 88109 71589
rect 88278 71527 88284 71530
rect 5457 71521 5515 71527
rect 5457 71487 5469 71521
rect 5503 71518 5515 71521
rect 88253 71521 88284 71527
rect 88253 71518 88265 71521
rect 5503 71490 5800 71518
rect 5503 71487 5515 71490
rect 5457 71481 5515 71487
rect 5772 71484 5800 71490
rect 7134 71484 7140 71496
rect 5772 71456 7140 71484
rect 7134 71444 7140 71456
rect 7192 71444 7198 71496
rect 87729 71487 87787 71493
rect 87729 71453 87741 71487
rect 87775 71484 87787 71487
rect 88112 71490 88265 71518
rect 88112 71484 88140 71490
rect 87775 71456 88140 71484
rect 88253 71487 88265 71490
rect 88253 71481 88284 71487
rect 88278 71478 88284 71481
rect 88336 71478 88342 71530
rect 87775 71453 87787 71456
rect 87729 71447 87787 71453
rect 2718 71376 2724 71428
rect 2776 71416 2782 71428
rect 5251 71419 5309 71425
rect 5251 71416 5263 71419
rect 2776 71388 5263 71416
rect 2776 71376 2782 71388
rect 5251 71385 5263 71388
rect 5297 71385 5309 71419
rect 5251 71379 5309 71385
rect 4876 71290 7912 71312
rect 4876 71238 6690 71290
rect 6742 71238 6754 71290
rect 6806 71238 6818 71290
rect 6870 71238 6882 71290
rect 6934 71238 6946 71290
rect 6998 71238 7912 71290
rect 4876 71216 7912 71238
rect 85284 71290 88596 71312
rect 85284 71238 87282 71290
rect 87334 71238 87346 71290
rect 87398 71238 87410 71290
rect 87462 71238 87474 71290
rect 87526 71238 87538 71290
rect 87590 71238 88596 71290
rect 85284 71216 88596 71238
rect 4876 70746 7912 70768
rect 4876 70694 5954 70746
rect 6006 70694 6018 70746
rect 6070 70694 6082 70746
rect 6134 70694 6146 70746
rect 6198 70694 6210 70746
rect 6262 70694 7912 70746
rect 4876 70672 7912 70694
rect 85284 70746 88596 70768
rect 85284 70694 86546 70746
rect 86598 70694 86610 70746
rect 86662 70694 86674 70746
rect 86726 70694 86738 70746
rect 86790 70694 86802 70746
rect 86854 70694 88596 70746
rect 85284 70672 88596 70694
rect 86898 70492 86904 70544
rect 86956 70532 86962 70544
rect 88051 70535 88109 70541
rect 88051 70532 88063 70535
rect 86956 70504 88063 70532
rect 86956 70492 86962 70504
rect 88051 70501 88063 70504
rect 88097 70501 88109 70535
rect 88051 70495 88109 70501
rect 87729 70467 87787 70473
rect 5457 70433 5515 70439
rect 5457 70399 5469 70433
rect 5503 70430 5515 70433
rect 87729 70433 87741 70467
rect 87775 70464 87787 70467
rect 88186 70464 88192 70476
rect 87775 70436 88192 70464
rect 87775 70433 87787 70436
rect 5503 70402 5800 70430
rect 87729 70427 87787 70433
rect 88186 70424 88192 70436
rect 88244 70439 88250 70476
rect 88244 70433 88279 70439
rect 5503 70399 5515 70402
rect 5457 70393 5515 70399
rect 5772 70396 5800 70402
rect 7134 70396 7140 70408
rect 5772 70368 7140 70396
rect 7134 70356 7140 70368
rect 7192 70356 7198 70408
rect 88204 70402 88233 70424
rect 88221 70399 88233 70402
rect 88267 70399 88279 70433
rect 88221 70393 88279 70399
rect 2902 70288 2908 70340
rect 2960 70328 2966 70340
rect 5251 70331 5309 70337
rect 5251 70328 5263 70331
rect 2960 70300 5263 70328
rect 2960 70288 2966 70300
rect 5251 70297 5263 70300
rect 5297 70297 5309 70331
rect 5251 70291 5309 70297
rect 4876 70202 7912 70224
rect 4876 70150 6690 70202
rect 6742 70150 6754 70202
rect 6806 70150 6818 70202
rect 6870 70150 6882 70202
rect 6934 70150 6946 70202
rect 6998 70150 7912 70202
rect 4876 70128 7912 70150
rect 85284 70202 88596 70224
rect 85284 70150 87282 70202
rect 87334 70150 87346 70202
rect 87398 70150 87410 70202
rect 87462 70150 87474 70202
rect 87526 70150 87538 70202
rect 87590 70150 88596 70202
rect 85284 70128 88596 70150
rect 4876 69658 7912 69680
rect 4876 69606 5954 69658
rect 6006 69606 6018 69658
rect 6070 69606 6082 69658
rect 6134 69606 6146 69658
rect 6198 69606 6210 69658
rect 6262 69606 7912 69658
rect 4876 69584 7912 69606
rect 85284 69658 88596 69680
rect 85284 69606 86546 69658
rect 86598 69606 86610 69658
rect 86662 69606 86674 69658
rect 86726 69606 86738 69658
rect 86790 69606 86802 69658
rect 86854 69606 88596 69658
rect 85284 69584 88596 69606
rect 5457 69345 5515 69351
rect 5457 69311 5469 69345
rect 5503 69342 5515 69345
rect 5662 69342 5668 69354
rect 5503 69314 5668 69342
rect 5503 69311 5515 69314
rect 5457 69305 5515 69311
rect 5662 69302 5668 69314
rect 5720 69302 5726 69354
rect 88253 69339 88311 69345
rect 86898 69268 86904 69320
rect 86956 69308 86962 69320
rect 88051 69311 88109 69317
rect 88051 69308 88063 69311
rect 86956 69280 88063 69308
rect 86956 69268 86962 69280
rect 88051 69277 88063 69280
rect 88097 69277 88109 69311
rect 88253 69305 88265 69339
rect 88299 69336 88311 69339
rect 88299 69308 88416 69336
rect 88554 69308 88560 69320
rect 88299 69305 88311 69308
rect 88253 69299 88311 69305
rect 88051 69271 88109 69277
rect 88388 69280 88560 69308
rect 4374 69200 4380 69252
rect 4432 69240 4438 69252
rect 5251 69243 5309 69249
rect 5251 69240 5263 69243
rect 4432 69212 5263 69240
rect 4432 69200 4438 69212
rect 5251 69209 5263 69212
rect 5297 69209 5309 69243
rect 5251 69203 5309 69209
rect 87729 69243 87787 69249
rect 87729 69209 87741 69243
rect 87775 69240 87787 69243
rect 88388 69240 88416 69280
rect 88554 69268 88560 69280
rect 88612 69268 88618 69320
rect 87775 69212 88416 69240
rect 87775 69209 87787 69212
rect 87729 69203 87787 69209
rect 4876 69114 7912 69136
rect 4876 69062 6690 69114
rect 6742 69062 6754 69114
rect 6806 69062 6818 69114
rect 6870 69062 6882 69114
rect 6934 69062 6946 69114
rect 6998 69062 7912 69114
rect 4876 69040 7912 69062
rect 85284 69114 88596 69136
rect 85284 69062 87282 69114
rect 87334 69062 87346 69114
rect 87398 69062 87410 69114
rect 87462 69062 87474 69114
rect 87526 69062 87538 69114
rect 87590 69062 88596 69114
rect 85284 69040 88596 69062
rect 4876 68570 7912 68592
rect 4876 68518 5954 68570
rect 6006 68518 6018 68570
rect 6070 68518 6082 68570
rect 6134 68518 6146 68570
rect 6198 68518 6210 68570
rect 6262 68518 7912 68570
rect 4876 68496 7912 68518
rect 85284 68570 88596 68592
rect 85284 68518 86546 68570
rect 86598 68518 86610 68570
rect 86662 68518 86674 68570
rect 86726 68518 86738 68570
rect 86790 68518 86802 68570
rect 86854 68518 88596 68570
rect 85284 68496 88596 68518
rect 4876 68026 7912 68048
rect 4876 67974 6690 68026
rect 6742 67974 6754 68026
rect 6806 67974 6818 68026
rect 6870 67974 6882 68026
rect 6934 67974 6946 68026
rect 6998 67974 7912 68026
rect 4876 67952 7912 67974
rect 85284 68026 88596 68048
rect 85284 67974 87282 68026
rect 87334 67974 87346 68026
rect 87398 67974 87410 68026
rect 87462 67974 87474 68026
rect 87526 67974 87538 68026
rect 87590 67974 88596 68026
rect 85284 67952 88596 67974
rect 87913 67815 87971 67821
rect 5457 67781 5515 67787
rect 5457 67747 5469 67781
rect 5503 67778 5515 67781
rect 5662 67778 5668 67790
rect 5503 67750 5668 67778
rect 5503 67747 5515 67750
rect 5457 67741 5515 67747
rect 5662 67738 5668 67750
rect 5720 67738 5726 67790
rect 87913 67781 87925 67815
rect 87959 67812 87971 67815
rect 87959 67790 88324 67812
rect 87959 67784 88284 67790
rect 87959 67781 87971 67784
rect 87913 67775 87971 67781
rect 88253 67781 88284 67784
rect 88253 67747 88265 67781
rect 88253 67741 88284 67747
rect 88278 67738 88284 67741
rect 88336 67738 88342 67790
rect 84414 67636 84420 67688
rect 84472 67676 84478 67688
rect 88051 67679 88109 67685
rect 88051 67676 88063 67679
rect 84472 67648 88063 67676
rect 84472 67636 84478 67648
rect 88051 67645 88063 67648
rect 88097 67645 88109 67679
rect 88051 67639 88109 67645
rect 2902 67568 2908 67620
rect 2960 67608 2966 67620
rect 5251 67611 5309 67617
rect 5251 67608 5263 67611
rect 2960 67580 5263 67608
rect 2960 67568 2966 67580
rect 5251 67577 5263 67580
rect 5297 67577 5309 67611
rect 5251 67571 5309 67577
rect 4876 67482 7912 67504
rect 4876 67430 5954 67482
rect 6006 67430 6018 67482
rect 6070 67430 6082 67482
rect 6134 67430 6146 67482
rect 6198 67430 6210 67482
rect 6262 67430 7912 67482
rect 4876 67408 7912 67430
rect 85284 67482 88596 67504
rect 85284 67430 86546 67482
rect 86598 67430 86610 67482
rect 86662 67430 86674 67482
rect 86726 67430 86738 67482
rect 86790 67430 86802 67482
rect 86854 67430 88596 67482
rect 85284 67408 88596 67430
rect 5457 67169 5515 67175
rect 88278 67169 88284 67172
rect 5457 67135 5469 67169
rect 5503 67166 5515 67169
rect 5503 67138 5800 67166
rect 88253 67163 88284 67169
rect 5503 67135 5515 67138
rect 5457 67129 5515 67135
rect 5772 67132 5800 67138
rect 7134 67132 7140 67144
rect 5772 67104 7140 67132
rect 7134 67092 7140 67104
rect 7192 67092 7198 67144
rect 86898 67092 86904 67144
rect 86956 67132 86962 67144
rect 88051 67135 88109 67141
rect 88051 67132 88063 67135
rect 86956 67104 88063 67132
rect 86956 67092 86962 67104
rect 88051 67101 88063 67104
rect 88097 67101 88109 67135
rect 88253 67129 88265 67163
rect 88253 67123 88284 67129
rect 88278 67120 88284 67123
rect 88336 67120 88342 67172
rect 88051 67095 88109 67101
rect 2902 67024 2908 67076
rect 2960 67064 2966 67076
rect 5251 67067 5309 67073
rect 5251 67064 5263 67067
rect 2960 67036 5263 67064
rect 2960 67024 2966 67036
rect 5251 67033 5263 67036
rect 5297 67033 5309 67067
rect 5251 67027 5309 67033
rect 87729 67067 87787 67073
rect 87729 67033 87741 67067
rect 87775 67064 87787 67067
rect 88296 67064 88324 67120
rect 87775 67036 88324 67064
rect 87775 67033 87787 67036
rect 87729 67027 87787 67033
rect 4876 66938 7912 66960
rect 4876 66886 6690 66938
rect 6742 66886 6754 66938
rect 6806 66886 6818 66938
rect 6870 66886 6882 66938
rect 6934 66886 6946 66938
rect 6998 66886 7912 66938
rect 4876 66864 7912 66886
rect 85284 66938 88596 66960
rect 85284 66886 87282 66938
rect 87334 66886 87346 66938
rect 87398 66886 87410 66938
rect 87462 66886 87474 66938
rect 87526 66886 87538 66938
rect 87590 66886 88596 66938
rect 85284 66864 88596 66886
rect 4876 66394 7912 66416
rect 4876 66342 5954 66394
rect 6006 66342 6018 66394
rect 6070 66342 6082 66394
rect 6134 66342 6146 66394
rect 6198 66342 6210 66394
rect 6262 66342 7912 66394
rect 4876 66320 7912 66342
rect 85284 66394 88596 66416
rect 85284 66342 86546 66394
rect 86598 66342 86610 66394
rect 86662 66342 86674 66394
rect 86726 66342 86738 66394
rect 86790 66342 86802 66394
rect 86854 66342 88596 66394
rect 85284 66320 88596 66342
rect 5205 66081 5263 66087
rect 5205 66047 5217 66081
rect 5251 66047 5263 66081
rect 87957 66081 88015 66087
rect 87957 66078 87969 66081
rect 5205 66041 5263 66047
rect 5365 66047 5423 66053
rect 2902 65936 2908 65988
rect 2960 65976 2966 65988
rect 5220 65976 5248 66041
rect 5365 66013 5377 66047
rect 5411 66044 5423 66047
rect 7226 66044 7232 66056
rect 5411 66016 7232 66044
rect 5411 66013 5423 66016
rect 5365 66007 5423 66013
rect 7226 66004 7232 66016
rect 7284 66004 7290 66056
rect 87082 66004 87088 66056
rect 87140 66044 87146 66056
rect 87652 66050 87969 66078
rect 87652 66044 87680 66050
rect 87140 66016 87680 66044
rect 87957 66047 87969 66050
rect 88003 66047 88015 66081
rect 87957 66041 88015 66047
rect 87140 66004 87146 66016
rect 88186 65985 88192 65988
rect 5481 65979 5539 65985
rect 5481 65976 5493 65979
rect 2960 65948 5493 65976
rect 2960 65936 2966 65948
rect 5481 65945 5493 65948
rect 5527 65945 5539 65979
rect 5481 65939 5539 65945
rect 88169 65979 88192 65985
rect 88169 65945 88181 65979
rect 88169 65939 88192 65945
rect 88186 65936 88192 65939
rect 88244 65936 88250 65988
rect 4876 65850 7912 65872
rect 4876 65798 6690 65850
rect 6742 65798 6754 65850
rect 6806 65798 6818 65850
rect 6870 65798 6882 65850
rect 6934 65798 6946 65850
rect 6998 65798 7912 65850
rect 4876 65776 7912 65798
rect 85284 65850 88596 65872
rect 85284 65798 87282 65850
rect 87334 65798 87346 65850
rect 87398 65798 87410 65850
rect 87462 65798 87474 65850
rect 87526 65798 87538 65850
rect 87590 65798 88596 65850
rect 85284 65776 88596 65798
rect 4876 65306 7912 65328
rect 4876 65254 5954 65306
rect 6006 65254 6018 65306
rect 6070 65254 6082 65306
rect 6134 65254 6146 65306
rect 6198 65254 6210 65306
rect 6262 65254 7912 65306
rect 4876 65232 7912 65254
rect 85284 65306 88596 65328
rect 85284 65254 86546 65306
rect 86598 65254 86610 65306
rect 86662 65254 86674 65306
rect 86726 65254 86738 65306
rect 86790 65254 86802 65306
rect 86854 65254 88596 65306
rect 85284 65232 88596 65254
rect 5205 64993 5263 64999
rect 5205 64959 5217 64993
rect 5251 64959 5263 64993
rect 87957 64993 88015 64999
rect 87957 64990 87969 64993
rect 5205 64953 5263 64959
rect 5365 64959 5423 64965
rect 2902 64848 2908 64900
rect 2960 64888 2966 64900
rect 5220 64888 5248 64953
rect 5365 64925 5377 64959
rect 5411 64956 5423 64959
rect 7226 64956 7232 64968
rect 5411 64928 7232 64956
rect 5411 64925 5423 64928
rect 5365 64919 5423 64925
rect 7226 64916 7232 64928
rect 7284 64916 7290 64968
rect 87082 64916 87088 64968
rect 87140 64956 87146 64968
rect 87652 64962 87969 64990
rect 87652 64956 87680 64962
rect 87140 64928 87680 64956
rect 87957 64959 87969 64962
rect 88003 64959 88015 64993
rect 87957 64953 88015 64959
rect 87140 64916 87146 64928
rect 5481 64891 5539 64897
rect 5481 64888 5493 64891
rect 2960 64860 5493 64888
rect 2960 64848 2966 64860
rect 5481 64857 5493 64860
rect 5527 64857 5539 64891
rect 5481 64851 5539 64857
rect 88169 64891 88227 64897
rect 88169 64857 88181 64891
rect 88215 64888 88227 64891
rect 88370 64888 88376 64900
rect 88215 64860 88376 64888
rect 88215 64857 88227 64860
rect 88169 64851 88227 64857
rect 88370 64848 88376 64860
rect 88428 64848 88434 64900
rect 4876 64762 7912 64784
rect 4876 64710 6690 64762
rect 6742 64710 6754 64762
rect 6806 64710 6818 64762
rect 6870 64710 6882 64762
rect 6934 64710 6946 64762
rect 6998 64710 7912 64762
rect 4876 64688 7912 64710
rect 85284 64762 88596 64784
rect 85284 64710 87282 64762
rect 87334 64710 87346 64762
rect 87398 64710 87410 64762
rect 87462 64710 87474 64762
rect 87526 64710 87538 64762
rect 87590 64710 88596 64762
rect 85284 64688 88596 64710
rect 7410 64576 7416 64628
rect 7468 64616 7474 64628
rect 7505 64619 7563 64625
rect 7505 64616 7517 64619
rect 7468 64588 7517 64616
rect 7468 64576 7474 64588
rect 7505 64585 7517 64588
rect 7551 64585 7563 64619
rect 7505 64579 7563 64585
rect 4876 64218 7912 64240
rect 4876 64166 5954 64218
rect 6006 64166 6018 64218
rect 6070 64166 6082 64218
rect 6134 64166 6146 64218
rect 6198 64166 6210 64218
rect 6262 64166 7912 64218
rect 4876 64144 7912 64166
rect 85284 64218 88596 64240
rect 85284 64166 86546 64218
rect 86598 64166 86610 64218
rect 86662 64166 86674 64218
rect 86726 64166 86738 64218
rect 86790 64166 86802 64218
rect 86854 64166 88596 64218
rect 85284 64144 88596 64166
rect 5365 63939 5423 63945
rect 5202 63862 5208 63914
rect 5260 63868 5266 63914
rect 5365 63905 5377 63939
rect 5411 63936 5423 63939
rect 9618 63936 9624 63948
rect 5411 63908 9624 63936
rect 5411 63905 5423 63908
rect 5365 63899 5423 63905
rect 9618 63896 9624 63908
rect 9676 63896 9682 63948
rect 87957 63905 88015 63911
rect 87957 63902 87969 63905
rect 7410 63877 7416 63880
rect 5481 63871 5539 63877
rect 5481 63868 5493 63871
rect 5260 63862 5493 63868
rect 5220 63840 5493 63862
rect 5481 63837 5493 63840
rect 5527 63837 5539 63871
rect 5481 63831 5539 63837
rect 7389 63871 7416 63877
rect 7389 63837 7401 63871
rect 7389 63831 7416 63837
rect 7410 63828 7416 63831
rect 7468 63828 7474 63880
rect 84414 63828 84420 63880
rect 84472 63868 84478 63880
rect 87652 63874 87969 63902
rect 87652 63868 87680 63874
rect 84472 63840 87680 63868
rect 87957 63871 87969 63874
rect 88003 63871 88015 63905
rect 87957 63865 88015 63871
rect 84472 63828 84478 63840
rect 6769 63803 6827 63809
rect 6769 63769 6781 63803
rect 6815 63800 6827 63803
rect 7226 63800 7232 63812
rect 6815 63772 7232 63800
rect 6815 63769 6827 63772
rect 6769 63763 6827 63769
rect 7226 63760 7232 63772
rect 7284 63800 7290 63812
rect 7778 63800 7784 63812
rect 7284 63772 7784 63800
rect 7284 63760 7290 63772
rect 7778 63760 7784 63772
rect 7836 63760 7842 63812
rect 88169 63803 88227 63809
rect 88169 63769 88181 63803
rect 88215 63800 88227 63803
rect 88554 63800 88560 63812
rect 88215 63772 88560 63800
rect 88215 63769 88227 63772
rect 88169 63763 88227 63769
rect 88554 63760 88560 63772
rect 88612 63760 88618 63812
rect 4876 63674 7912 63696
rect 4876 63622 6690 63674
rect 6742 63622 6754 63674
rect 6806 63622 6818 63674
rect 6870 63622 6882 63674
rect 6934 63622 6946 63674
rect 6998 63622 7912 63674
rect 4876 63600 7912 63622
rect 85284 63674 88596 63696
rect 85284 63622 87282 63674
rect 87334 63622 87346 63674
rect 87398 63622 87410 63674
rect 87462 63622 87474 63674
rect 87526 63622 87538 63674
rect 87590 63622 88596 63674
rect 85284 63600 88596 63622
rect 7318 63216 7324 63268
rect 7376 63256 7382 63268
rect 7505 63259 7563 63265
rect 7505 63256 7517 63259
rect 7376 63228 7517 63256
rect 7376 63216 7382 63228
rect 7505 63225 7517 63228
rect 7551 63225 7563 63259
rect 7505 63219 7563 63225
rect 4876 63130 7912 63152
rect 4876 63078 5954 63130
rect 6006 63078 6018 63130
rect 6070 63078 6082 63130
rect 6134 63078 6146 63130
rect 6198 63078 6210 63130
rect 6262 63078 7912 63130
rect 4876 63056 7912 63078
rect 85284 63130 88596 63152
rect 85284 63078 86546 63130
rect 86598 63078 86610 63130
rect 86662 63078 86674 63130
rect 86726 63078 86738 63130
rect 86790 63078 86802 63130
rect 86854 63078 88596 63130
rect 85284 63056 88596 63078
rect 4876 62586 7912 62608
rect 4876 62534 6690 62586
rect 6742 62534 6754 62586
rect 6806 62534 6818 62586
rect 6870 62534 6882 62586
rect 6934 62534 6946 62586
rect 6998 62534 7912 62586
rect 4876 62512 7912 62534
rect 85284 62586 88596 62608
rect 85284 62534 87282 62586
rect 87334 62534 87346 62586
rect 87398 62534 87410 62586
rect 87462 62534 87474 62586
rect 87526 62534 87538 62586
rect 87590 62534 88596 62586
rect 85284 62512 88596 62534
rect 5365 62443 5423 62449
rect 5365 62409 5377 62443
rect 5411 62440 5423 62443
rect 7226 62440 7232 62452
rect 5411 62412 7232 62440
rect 5411 62409 5423 62412
rect 5365 62403 5423 62409
rect 7226 62400 7232 62412
rect 7284 62400 7290 62452
rect 4926 62298 4932 62350
rect 4984 62338 4990 62350
rect 5159 62341 5217 62347
rect 5159 62338 5171 62341
rect 4984 62310 5171 62338
rect 4984 62298 4990 62310
rect 5159 62307 5171 62310
rect 5205 62338 5217 62341
rect 5205 62313 5524 62338
rect 87082 62332 87088 62384
rect 87140 62372 87146 62384
rect 88169 62375 88227 62381
rect 87140 62344 87680 62372
rect 87140 62332 87146 62344
rect 87652 62338 87680 62344
rect 87957 62341 88015 62347
rect 87957 62338 87969 62341
rect 5205 62310 5539 62313
rect 87652 62310 87969 62338
rect 5205 62307 5217 62310
rect 5159 62301 5217 62307
rect 5481 62307 5539 62310
rect 5481 62273 5493 62307
rect 5527 62273 5539 62307
rect 87957 62307 87969 62310
rect 88003 62307 88015 62341
rect 88169 62341 88181 62375
rect 88215 62372 88227 62375
rect 88554 62372 88560 62384
rect 88215 62344 88560 62372
rect 88215 62341 88227 62344
rect 88169 62335 88227 62341
rect 88554 62332 88560 62344
rect 88612 62332 88618 62384
rect 87957 62301 88015 62307
rect 5481 62267 5539 62273
rect 4876 62042 7912 62064
rect 4876 61990 5954 62042
rect 6006 61990 6018 62042
rect 6070 61990 6082 62042
rect 6134 61990 6146 62042
rect 6198 61990 6210 62042
rect 6262 61990 7912 62042
rect 4876 61968 7912 61990
rect 85284 62042 88596 62064
rect 85284 61990 86546 62042
rect 86598 61990 86610 62042
rect 86662 61990 86674 62042
rect 86726 61990 86738 62042
rect 86790 61990 86802 62042
rect 86854 61990 88596 62042
rect 85284 61968 88596 61990
rect 5205 61729 5263 61735
rect 5205 61695 5217 61729
rect 5251 61695 5263 61729
rect 87957 61729 88015 61735
rect 87957 61726 87969 61729
rect 5205 61689 5263 61695
rect 5364 61695 5422 61701
rect 2902 61584 2908 61636
rect 2960 61624 2966 61636
rect 5220 61624 5248 61689
rect 5364 61661 5376 61695
rect 5410 61692 5422 61695
rect 7226 61692 7232 61704
rect 5410 61664 7232 61692
rect 5410 61661 5422 61664
rect 5364 61655 5422 61661
rect 7226 61652 7232 61664
rect 7284 61652 7290 61704
rect 87082 61652 87088 61704
rect 87140 61692 87146 61704
rect 87652 61698 87969 61726
rect 87652 61692 87680 61698
rect 87140 61664 87680 61692
rect 87957 61695 87969 61698
rect 88003 61695 88015 61729
rect 87957 61689 88015 61695
rect 87140 61652 87146 61664
rect 88186 61633 88192 61636
rect 5481 61627 5539 61633
rect 5481 61624 5493 61627
rect 2960 61596 5493 61624
rect 2960 61584 2966 61596
rect 5481 61593 5493 61596
rect 5527 61593 5539 61627
rect 5481 61587 5539 61593
rect 88169 61627 88192 61633
rect 88169 61593 88181 61627
rect 88169 61587 88192 61593
rect 88186 61584 88192 61587
rect 88244 61584 88250 61636
rect 4876 61498 7912 61520
rect 4876 61446 6690 61498
rect 6742 61446 6754 61498
rect 6806 61446 6818 61498
rect 6870 61446 6882 61498
rect 6934 61446 6946 61498
rect 6998 61446 7912 61498
rect 4876 61424 7912 61446
rect 85284 61498 88596 61520
rect 85284 61446 87282 61498
rect 87334 61446 87346 61498
rect 87398 61446 87410 61498
rect 87462 61446 87474 61498
rect 87526 61446 87538 61498
rect 87590 61446 88596 61498
rect 85284 61424 88596 61446
rect 4876 60954 7912 60976
rect 4876 60902 5954 60954
rect 6006 60902 6018 60954
rect 6070 60902 6082 60954
rect 6134 60902 6146 60954
rect 6198 60902 6210 60954
rect 6262 60902 7912 60954
rect 4876 60880 7912 60902
rect 85284 60954 88596 60976
rect 85284 60902 86546 60954
rect 86598 60902 86610 60954
rect 86662 60902 86674 60954
rect 86726 60902 86738 60954
rect 86790 60902 86802 60954
rect 86854 60902 88596 60954
rect 85284 60880 88596 60902
rect 5205 60641 5263 60647
rect 5205 60607 5217 60641
rect 5251 60607 5263 60641
rect 87957 60641 88015 60647
rect 87957 60638 87969 60641
rect 5205 60601 5263 60607
rect 5364 60607 5422 60613
rect 2902 60496 2908 60548
rect 2960 60536 2966 60548
rect 5220 60536 5248 60601
rect 5364 60573 5376 60607
rect 5410 60604 5422 60607
rect 7226 60604 7232 60616
rect 5410 60576 7232 60604
rect 5410 60573 5422 60576
rect 5364 60567 5422 60573
rect 7226 60564 7232 60576
rect 7284 60564 7290 60616
rect 87082 60564 87088 60616
rect 87140 60604 87146 60616
rect 87652 60610 87969 60638
rect 87652 60604 87680 60610
rect 87140 60576 87680 60604
rect 87957 60607 87969 60610
rect 88003 60607 88015 60641
rect 87957 60601 88015 60607
rect 87140 60564 87146 60576
rect 88186 60545 88192 60548
rect 5481 60539 5539 60545
rect 5481 60536 5493 60539
rect 2960 60508 5493 60536
rect 2960 60496 2966 60508
rect 5481 60505 5493 60508
rect 5527 60505 5539 60539
rect 5481 60499 5539 60505
rect 88169 60539 88192 60545
rect 88169 60505 88181 60539
rect 88169 60499 88192 60505
rect 88186 60496 88192 60499
rect 88244 60496 88250 60548
rect 4876 60410 7912 60432
rect 4876 60358 6690 60410
rect 6742 60358 6754 60410
rect 6806 60358 6818 60410
rect 6870 60358 6882 60410
rect 6934 60358 6946 60410
rect 6998 60358 7912 60410
rect 4876 60336 7912 60358
rect 85284 60410 88596 60432
rect 85284 60358 87282 60410
rect 87334 60358 87346 60410
rect 87398 60358 87410 60410
rect 87462 60358 87474 60410
rect 87526 60358 87538 60410
rect 87590 60358 88596 60410
rect 85284 60336 88596 60358
rect 4876 59866 7912 59888
rect 4876 59814 5954 59866
rect 6006 59814 6018 59866
rect 6070 59814 6082 59866
rect 6134 59814 6146 59866
rect 6198 59814 6210 59866
rect 6262 59814 7912 59866
rect 4876 59792 7912 59814
rect 85284 59866 88596 59888
rect 85284 59814 86546 59866
rect 86598 59814 86610 59866
rect 86662 59814 86674 59866
rect 86726 59814 86738 59866
rect 86790 59814 86802 59866
rect 86854 59814 88596 59866
rect 85284 59792 88596 59814
rect 5205 59553 5263 59559
rect 5205 59528 5217 59553
rect 5251 59528 5263 59553
rect 87957 59553 88015 59559
rect 87957 59550 87969 59553
rect 87652 59528 87969 59550
rect 5202 59476 5208 59528
rect 5260 59476 5266 59528
rect 5365 59519 5423 59525
rect 5365 59485 5377 59519
rect 5411 59516 5423 59519
rect 7226 59516 7232 59528
rect 5411 59488 7232 59516
rect 5411 59485 5423 59488
rect 5365 59479 5423 59485
rect 7226 59476 7232 59488
rect 7284 59476 7290 59528
rect 87634 59476 87640 59528
rect 87692 59522 87969 59528
rect 87692 59476 87698 59522
rect 87957 59519 87969 59522
rect 88003 59519 88015 59553
rect 87957 59513 88015 59519
rect 5220 59448 5248 59476
rect 5481 59451 5539 59457
rect 5481 59448 5493 59451
rect 5220 59420 5493 59448
rect 5481 59417 5493 59420
rect 5527 59417 5539 59451
rect 5481 59411 5539 59417
rect 88169 59451 88227 59457
rect 88169 59417 88181 59451
rect 88215 59448 88227 59451
rect 88370 59448 88376 59460
rect 88215 59420 88376 59448
rect 88215 59417 88227 59420
rect 88169 59411 88227 59417
rect 88370 59408 88376 59420
rect 88428 59408 88434 59460
rect 4876 59322 7912 59344
rect 4876 59270 6690 59322
rect 6742 59270 6754 59322
rect 6806 59270 6818 59322
rect 6870 59270 6882 59322
rect 6934 59270 6946 59322
rect 6998 59270 7912 59322
rect 4876 59248 7912 59270
rect 85284 59322 88596 59344
rect 85284 59270 87282 59322
rect 87334 59270 87346 59322
rect 87398 59270 87410 59322
rect 87462 59270 87474 59322
rect 87526 59270 87538 59322
rect 87590 59270 88596 59322
rect 85284 59248 88596 59270
rect 4876 58778 7912 58800
rect 4876 58726 5954 58778
rect 6006 58726 6018 58778
rect 6070 58726 6082 58778
rect 6134 58726 6146 58778
rect 6198 58726 6210 58778
rect 6262 58726 7912 58778
rect 4876 58704 7912 58726
rect 85284 58778 88596 58800
rect 85284 58726 86546 58778
rect 86598 58726 86610 58778
rect 86662 58726 86674 58778
rect 86726 58726 86738 58778
rect 86790 58726 86802 58778
rect 86854 58726 88596 58778
rect 85284 58704 88596 58726
rect 5202 58422 5208 58474
rect 5260 58428 5266 58474
rect 5481 58431 5539 58437
rect 5481 58428 5493 58431
rect 5260 58422 5493 58428
rect 5220 58400 5493 58422
rect 5481 58397 5493 58400
rect 5527 58397 5539 58431
rect 88002 58422 88008 58474
rect 88060 58422 88066 58474
rect 5481 58391 5539 58397
rect 5386 58369 5392 58372
rect 5364 58363 5392 58369
rect 5364 58329 5376 58363
rect 5364 58323 5392 58329
rect 5386 58320 5392 58323
rect 5444 58320 5450 58372
rect 88169 58363 88227 58369
rect 88169 58329 88181 58363
rect 88215 58360 88227 58363
rect 88554 58360 88560 58372
rect 88215 58332 88560 58360
rect 88215 58329 88227 58332
rect 88169 58323 88227 58329
rect 88554 58320 88560 58332
rect 88612 58320 88618 58372
rect 4876 58234 7912 58256
rect 4876 58182 6690 58234
rect 6742 58182 6754 58234
rect 6806 58182 6818 58234
rect 6870 58182 6882 58234
rect 6934 58182 6946 58234
rect 6998 58182 7912 58234
rect 4876 58160 7912 58182
rect 85284 58234 88596 58256
rect 85284 58182 87282 58234
rect 87334 58182 87346 58234
rect 87398 58182 87410 58234
rect 87462 58182 87474 58234
rect 87526 58182 87538 58234
rect 87590 58182 88596 58234
rect 85284 58160 88596 58182
rect 4876 57690 7912 57712
rect 4876 57638 5954 57690
rect 6006 57638 6018 57690
rect 6070 57638 6082 57690
rect 6134 57638 6146 57690
rect 6198 57638 6210 57690
rect 6262 57638 7912 57690
rect 4876 57616 7912 57638
rect 85284 57690 88596 57712
rect 85284 57638 86546 57690
rect 86598 57638 86610 57690
rect 86662 57638 86674 57690
rect 86726 57638 86738 57690
rect 86790 57638 86802 57690
rect 86854 57638 88596 57690
rect 85284 57616 88596 57638
rect 4876 57146 7912 57168
rect 4876 57094 6690 57146
rect 6742 57094 6754 57146
rect 6806 57094 6818 57146
rect 6870 57094 6882 57146
rect 6934 57094 6946 57146
rect 6998 57094 7912 57146
rect 4876 57072 7912 57094
rect 85284 57146 88596 57168
rect 85284 57094 87282 57146
rect 87334 57094 87346 57146
rect 87398 57094 87410 57146
rect 87462 57094 87474 57146
rect 87526 57094 87538 57146
rect 87590 57094 88596 57146
rect 85284 57072 88596 57094
rect 5365 57003 5423 57009
rect 5365 56969 5377 57003
rect 5411 57000 5423 57003
rect 7226 57000 7232 57012
rect 5411 56972 7232 57000
rect 5411 56969 5423 56972
rect 5365 56963 5423 56969
rect 7226 56960 7232 56972
rect 7284 56960 7290 57012
rect 4926 56858 4932 56910
rect 4984 56898 4990 56910
rect 5159 56901 5217 56907
rect 5159 56898 5171 56901
rect 4984 56870 5171 56898
rect 4984 56858 4990 56870
rect 5159 56867 5171 56870
rect 5205 56898 5217 56901
rect 5205 56873 5524 56898
rect 5205 56870 5539 56873
rect 5205 56867 5217 56870
rect 5159 56861 5217 56867
rect 5481 56867 5539 56870
rect 5481 56833 5493 56867
rect 5527 56833 5539 56867
rect 88002 56858 88008 56910
rect 88060 56858 88066 56910
rect 88169 56867 88227 56873
rect 5481 56827 5539 56833
rect 88169 56833 88181 56867
rect 88215 56864 88227 56867
rect 88830 56864 88836 56876
rect 88215 56836 88836 56864
rect 88215 56833 88227 56836
rect 88169 56827 88227 56833
rect 88830 56824 88836 56836
rect 88888 56824 88894 56876
rect 4876 56602 7912 56624
rect 4876 56550 5954 56602
rect 6006 56550 6018 56602
rect 6070 56550 6082 56602
rect 6134 56550 6146 56602
rect 6198 56550 6210 56602
rect 6262 56550 7912 56602
rect 4876 56528 7912 56550
rect 85284 56602 88596 56624
rect 85284 56550 86546 56602
rect 86598 56550 86610 56602
rect 86662 56550 86674 56602
rect 86726 56550 86738 56602
rect 86790 56550 86802 56602
rect 86854 56550 88596 56602
rect 85284 56528 88596 56550
rect 5481 56323 5539 56329
rect 5481 56320 5493 56323
rect 5174 56295 5493 56320
rect 5159 56292 5493 56295
rect 5159 56289 5217 56292
rect 2902 56212 2908 56264
rect 2960 56252 2966 56264
rect 5159 56255 5171 56289
rect 5205 56255 5217 56289
rect 5481 56289 5493 56292
rect 5527 56289 5539 56323
rect 5481 56283 5539 56289
rect 87957 56289 88015 56295
rect 87957 56286 87969 56289
rect 5159 56252 5217 56255
rect 2960 56249 5217 56252
rect 5365 56255 5423 56261
rect 2960 56224 5202 56249
rect 2960 56212 2966 56224
rect 5365 56221 5377 56255
rect 5411 56252 5423 56255
rect 7226 56252 7232 56264
rect 5411 56224 7232 56252
rect 5411 56221 5423 56224
rect 5365 56215 5423 56221
rect 7226 56212 7232 56224
rect 7284 56212 7290 56264
rect 87082 56212 87088 56264
rect 87140 56252 87146 56264
rect 87652 56258 87969 56286
rect 87652 56252 87680 56258
rect 87140 56224 87680 56252
rect 87957 56255 87969 56258
rect 88003 56255 88015 56289
rect 87957 56249 88015 56255
rect 87140 56212 87146 56224
rect 88186 56193 88192 56196
rect 88169 56187 88192 56193
rect 88169 56153 88181 56187
rect 88169 56147 88192 56153
rect 88186 56144 88192 56147
rect 88244 56144 88250 56196
rect 4876 56058 7912 56080
rect 4876 56006 6690 56058
rect 6742 56006 6754 56058
rect 6806 56006 6818 56058
rect 6870 56006 6882 56058
rect 6934 56006 6946 56058
rect 6998 56006 7912 56058
rect 4876 55984 7912 56006
rect 85284 56058 88596 56080
rect 85284 56006 87282 56058
rect 87334 56006 87346 56058
rect 87398 56006 87410 56058
rect 87462 56006 87474 56058
rect 87526 56006 87538 56058
rect 87590 56006 88596 56058
rect 85284 55984 88596 56006
rect 4876 55514 7912 55536
rect 4876 55462 5954 55514
rect 6006 55462 6018 55514
rect 6070 55462 6082 55514
rect 6134 55462 6146 55514
rect 6198 55462 6210 55514
rect 6262 55462 7912 55514
rect 4876 55440 7912 55462
rect 85284 55514 88596 55536
rect 85284 55462 86546 55514
rect 86598 55462 86610 55514
rect 86662 55462 86674 55514
rect 86726 55462 86738 55514
rect 86790 55462 86802 55514
rect 86854 55462 88596 55514
rect 85284 55440 88596 55462
rect 5481 55235 5539 55241
rect 5481 55232 5493 55235
rect 5174 55207 5493 55232
rect 5159 55204 5493 55207
rect 5159 55201 5217 55204
rect 2902 55124 2908 55176
rect 2960 55164 2966 55176
rect 5159 55167 5171 55201
rect 5205 55167 5217 55201
rect 5481 55201 5493 55204
rect 5527 55201 5539 55235
rect 5481 55195 5539 55201
rect 87957 55201 88015 55207
rect 87957 55198 87969 55201
rect 5159 55164 5217 55167
rect 2960 55161 5217 55164
rect 5365 55167 5423 55173
rect 2960 55136 5202 55161
rect 2960 55124 2966 55136
rect 5365 55133 5377 55167
rect 5411 55164 5423 55167
rect 7226 55164 7232 55176
rect 5411 55136 7232 55164
rect 5411 55133 5423 55136
rect 5365 55127 5423 55133
rect 7226 55124 7232 55136
rect 7284 55124 7290 55176
rect 87082 55124 87088 55176
rect 87140 55164 87146 55176
rect 87652 55170 87969 55198
rect 87652 55164 87680 55170
rect 87140 55136 87680 55164
rect 87957 55167 87969 55170
rect 88003 55167 88015 55201
rect 87957 55161 88015 55167
rect 87140 55124 87146 55136
rect 88186 55105 88192 55108
rect 88169 55099 88192 55105
rect 88169 55065 88181 55099
rect 88169 55059 88192 55065
rect 88186 55056 88192 55059
rect 88244 55056 88250 55108
rect 4876 54970 7912 54992
rect 4876 54918 6690 54970
rect 6742 54918 6754 54970
rect 6806 54918 6818 54970
rect 6870 54918 6882 54970
rect 6934 54918 6946 54970
rect 6998 54918 7912 54970
rect 4876 54896 7912 54918
rect 85284 54970 88596 54992
rect 85284 54918 87282 54970
rect 87334 54918 87346 54970
rect 87398 54918 87410 54970
rect 87462 54918 87474 54970
rect 87526 54918 87538 54970
rect 87590 54918 88596 54970
rect 85284 54896 88596 54918
rect 4876 54426 7912 54448
rect 4876 54374 5954 54426
rect 6006 54374 6018 54426
rect 6070 54374 6082 54426
rect 6134 54374 6146 54426
rect 6198 54374 6210 54426
rect 6262 54374 7912 54426
rect 4876 54352 7912 54374
rect 85284 54426 88596 54448
rect 85284 54374 86546 54426
rect 86598 54374 86610 54426
rect 86662 54374 86674 54426
rect 86726 54374 86738 54426
rect 86790 54374 86802 54426
rect 86854 54374 88596 54426
rect 85284 54352 88596 54374
rect 5481 54147 5539 54153
rect 5481 54144 5493 54147
rect 5174 54119 5493 54144
rect 5159 54116 5493 54119
rect 5159 54113 5217 54116
rect 5159 54088 5171 54113
rect 5110 54036 5116 54088
rect 5168 54079 5171 54088
rect 5205 54079 5217 54113
rect 5481 54113 5493 54116
rect 5527 54113 5539 54147
rect 5481 54107 5539 54113
rect 87957 54113 88015 54119
rect 87957 54110 87969 54113
rect 5168 54073 5217 54079
rect 5365 54079 5423 54085
rect 5168 54048 5202 54073
rect 5168 54036 5174 54048
rect 5365 54045 5377 54079
rect 5411 54076 5423 54079
rect 5662 54076 5668 54088
rect 5411 54048 5668 54076
rect 5411 54045 5423 54048
rect 5365 54039 5423 54045
rect 5662 54036 5668 54048
rect 5720 54036 5726 54088
rect 84414 54036 84420 54088
rect 84472 54076 84478 54088
rect 87652 54082 87969 54110
rect 87652 54076 87680 54082
rect 84472 54048 87680 54076
rect 87957 54079 87969 54082
rect 88003 54079 88015 54113
rect 87957 54073 88015 54079
rect 88169 54079 88227 54085
rect 84472 54036 84478 54048
rect 88169 54045 88181 54079
rect 88215 54076 88227 54079
rect 88646 54076 88652 54088
rect 88215 54048 88652 54076
rect 88215 54045 88227 54048
rect 88169 54039 88227 54045
rect 88646 54036 88652 54048
rect 88704 54036 88710 54088
rect 4876 53882 7912 53904
rect 4876 53830 6690 53882
rect 6742 53830 6754 53882
rect 6806 53830 6818 53882
rect 6870 53830 6882 53882
rect 6934 53830 6946 53882
rect 6998 53830 7912 53882
rect 4876 53808 7912 53830
rect 85284 53882 88596 53904
rect 85284 53830 87282 53882
rect 87334 53830 87346 53882
rect 87398 53830 87410 53882
rect 87462 53830 87474 53882
rect 87526 53830 87538 53882
rect 87590 53830 88596 53882
rect 85284 53808 88596 53830
rect 4876 53338 7912 53360
rect 4876 53286 5954 53338
rect 6006 53286 6018 53338
rect 6070 53286 6082 53338
rect 6134 53286 6146 53338
rect 6198 53286 6210 53338
rect 6262 53286 7912 53338
rect 4876 53264 7912 53286
rect 85284 53338 88596 53360
rect 85284 53286 86546 53338
rect 86598 53286 86610 53338
rect 86662 53286 86674 53338
rect 86726 53286 86738 53338
rect 86790 53286 86802 53338
rect 86854 53286 88596 53338
rect 85284 53264 88596 53286
rect 5481 53059 5539 53065
rect 5481 53056 5493 53059
rect 5174 53031 5493 53056
rect 5159 53028 5493 53031
rect 5159 53025 5217 53028
rect 2902 52948 2908 53000
rect 2960 52988 2966 53000
rect 5159 52991 5171 53025
rect 5205 52991 5217 53025
rect 5481 53025 5493 53028
rect 5527 53025 5539 53059
rect 5481 53019 5539 53025
rect 87957 53025 88015 53031
rect 87957 53022 87969 53025
rect 5159 52988 5217 52991
rect 2960 52985 5217 52988
rect 5365 52991 5423 52997
rect 2960 52960 5202 52985
rect 2960 52948 2966 52960
rect 5365 52957 5377 52991
rect 5411 52988 5423 52991
rect 7226 52988 7232 53000
rect 5411 52960 7232 52988
rect 5411 52957 5423 52960
rect 5365 52951 5423 52957
rect 7226 52948 7232 52960
rect 7284 52948 7290 53000
rect 87082 52948 87088 53000
rect 87140 52988 87146 53000
rect 87652 52994 87969 53022
rect 87652 52988 87680 52994
rect 87140 52960 87680 52988
rect 87957 52991 87969 52994
rect 88003 52991 88015 53025
rect 87957 52985 88015 52991
rect 87140 52948 87146 52960
rect 88169 52923 88227 52929
rect 88169 52889 88181 52923
rect 88215 52920 88227 52923
rect 88278 52920 88284 52932
rect 88215 52892 88284 52920
rect 88215 52889 88227 52892
rect 88169 52883 88227 52889
rect 88278 52880 88284 52892
rect 88336 52880 88342 52932
rect 4876 52794 7912 52816
rect 4876 52742 6690 52794
rect 6742 52742 6754 52794
rect 6806 52742 6818 52794
rect 6870 52742 6882 52794
rect 6934 52742 6946 52794
rect 6998 52742 7912 52794
rect 4876 52720 7912 52742
rect 85284 52794 88596 52816
rect 85284 52742 87282 52794
rect 87334 52742 87346 52794
rect 87398 52742 87410 52794
rect 87462 52742 87474 52794
rect 87526 52742 87538 52794
rect 87590 52742 88596 52794
rect 85284 52720 88596 52742
rect 4876 52250 7912 52272
rect 4876 52198 5954 52250
rect 6006 52198 6018 52250
rect 6070 52198 6082 52250
rect 6134 52198 6146 52250
rect 6198 52198 6210 52250
rect 6262 52198 7912 52250
rect 4876 52176 7912 52198
rect 85284 52250 88596 52272
rect 85284 52198 86546 52250
rect 86598 52198 86610 52250
rect 86662 52198 86674 52250
rect 86726 52198 86738 52250
rect 86790 52198 86802 52250
rect 86854 52198 88596 52250
rect 85284 52176 88596 52198
rect 4876 51706 7912 51728
rect 4876 51654 6690 51706
rect 6742 51654 6754 51706
rect 6806 51654 6818 51706
rect 6870 51654 6882 51706
rect 6934 51654 6946 51706
rect 6998 51654 7912 51706
rect 4876 51632 7912 51654
rect 85284 51706 88596 51728
rect 85284 51654 87282 51706
rect 87334 51654 87346 51706
rect 87398 51654 87410 51706
rect 87462 51654 87474 51706
rect 87526 51654 87538 51706
rect 87590 51654 88596 51706
rect 85284 51632 88596 51654
rect 5365 51563 5423 51569
rect 5365 51529 5377 51563
rect 5411 51560 5423 51563
rect 7226 51560 7232 51572
rect 5411 51532 7232 51560
rect 5411 51529 5423 51532
rect 5365 51523 5423 51529
rect 7226 51520 7232 51532
rect 7284 51520 7290 51572
rect 5159 51461 5217 51467
rect 2902 51384 2908 51436
rect 2960 51424 2966 51436
rect 5159 51427 5171 51461
rect 5205 51427 5217 51461
rect 85794 51452 85800 51504
rect 85852 51492 85858 51504
rect 85852 51467 88000 51492
rect 85852 51464 88015 51467
rect 85852 51452 85858 51464
rect 87957 51461 88015 51464
rect 5159 51424 5217 51427
rect 5481 51427 5539 51433
rect 5481 51424 5493 51427
rect 2960 51396 5493 51424
rect 2960 51384 2966 51396
rect 5481 51393 5493 51396
rect 5527 51393 5539 51427
rect 87957 51427 87969 51461
rect 88003 51427 88015 51461
rect 87957 51421 88015 51427
rect 5481 51387 5539 51393
rect 88186 51365 88192 51368
rect 88169 51359 88192 51365
rect 88169 51325 88181 51359
rect 88169 51319 88192 51325
rect 88186 51316 88192 51319
rect 88244 51316 88250 51368
rect 4876 51162 7912 51184
rect 4876 51110 5954 51162
rect 6006 51110 6018 51162
rect 6070 51110 6082 51162
rect 6134 51110 6146 51162
rect 6198 51110 6210 51162
rect 6262 51110 7912 51162
rect 4876 51088 7912 51110
rect 85284 51162 88596 51184
rect 85284 51110 86546 51162
rect 86598 51110 86610 51162
rect 86662 51110 86674 51162
rect 86726 51110 86738 51162
rect 86790 51110 86802 51162
rect 86854 51110 88596 51162
rect 85284 51088 88596 51110
rect 85426 50704 85432 50756
rect 85484 50744 85490 50756
rect 85613 50747 85671 50753
rect 85613 50744 85625 50747
rect 85484 50716 85625 50744
rect 85484 50704 85490 50716
rect 85613 50713 85625 50716
rect 85659 50713 85671 50747
rect 85613 50707 85671 50713
rect 4876 50618 7912 50640
rect 4876 50566 6690 50618
rect 6742 50566 6754 50618
rect 6806 50566 6818 50618
rect 6870 50566 6882 50618
rect 6934 50566 6946 50618
rect 6998 50566 7912 50618
rect 4876 50544 7912 50566
rect 85284 50618 88596 50640
rect 85284 50566 87282 50618
rect 87334 50566 87346 50618
rect 87398 50566 87410 50618
rect 87462 50566 87474 50618
rect 87526 50566 87538 50618
rect 87590 50566 88596 50618
rect 85284 50544 88596 50566
rect 4876 50074 7912 50096
rect 4876 50022 5954 50074
rect 6006 50022 6018 50074
rect 6070 50022 6082 50074
rect 6134 50022 6146 50074
rect 6198 50022 6210 50074
rect 6262 50022 7912 50074
rect 4876 50000 7912 50022
rect 85284 50074 88596 50096
rect 85284 50022 86546 50074
rect 86598 50022 86610 50074
rect 86662 50022 86674 50074
rect 86726 50022 86738 50074
rect 86790 50022 86802 50074
rect 86854 50022 88596 50074
rect 85284 50000 88596 50022
rect 85518 49616 85524 49668
rect 85576 49656 85582 49668
rect 85613 49659 85671 49665
rect 85613 49656 85625 49659
rect 85576 49628 85625 49656
rect 85576 49616 85582 49628
rect 85613 49625 85625 49628
rect 85659 49625 85671 49659
rect 85613 49619 85671 49625
rect 4876 49530 7912 49552
rect 4876 49478 6690 49530
rect 6742 49478 6754 49530
rect 6806 49478 6818 49530
rect 6870 49478 6882 49530
rect 6934 49478 6946 49530
rect 6998 49478 7912 49530
rect 4876 49456 7912 49478
rect 85284 49530 88596 49552
rect 85284 49478 87282 49530
rect 87334 49478 87346 49530
rect 87398 49478 87410 49530
rect 87462 49478 87474 49530
rect 87526 49478 87538 49530
rect 87590 49478 88596 49530
rect 85284 49456 88596 49478
rect 4876 48986 7912 49008
rect 4876 48934 5954 48986
rect 6006 48934 6018 48986
rect 6070 48934 6082 48986
rect 6134 48934 6146 48986
rect 6198 48934 6210 48986
rect 6262 48934 7912 48986
rect 4876 48912 7912 48934
rect 85284 48986 88596 49008
rect 85284 48934 86546 48986
rect 86598 48934 86610 48986
rect 86662 48934 86674 48986
rect 86726 48934 86738 48986
rect 86790 48934 86802 48986
rect 86854 48934 88596 48986
rect 85284 48912 88596 48934
rect 88186 48596 88192 48648
rect 88244 48596 88250 48648
rect 85334 48528 85340 48580
rect 85392 48568 85398 48580
rect 85613 48571 85671 48577
rect 85613 48568 85625 48571
rect 85392 48540 85625 48568
rect 85392 48528 85398 48540
rect 85613 48537 85625 48540
rect 85659 48537 85671 48571
rect 85613 48531 85671 48537
rect 4876 48442 7912 48464
rect 4876 48390 6690 48442
rect 6742 48390 6754 48442
rect 6806 48390 6818 48442
rect 6870 48390 6882 48442
rect 6934 48390 6946 48442
rect 6998 48390 7912 48442
rect 4876 48368 7912 48390
rect 85284 48442 88596 48464
rect 85284 48390 87282 48442
rect 87334 48390 87346 48442
rect 87398 48390 87410 48442
rect 87462 48390 87474 48442
rect 87526 48390 87538 48442
rect 87590 48390 88596 48442
rect 85284 48368 88596 48390
rect 88186 47984 88192 48036
rect 88244 47984 88250 48036
rect 4876 47898 7912 47920
rect 4876 47846 5954 47898
rect 6006 47846 6018 47898
rect 6070 47846 6082 47898
rect 6134 47846 6146 47898
rect 6198 47846 6210 47898
rect 6262 47846 7912 47898
rect 4876 47824 7912 47846
rect 85284 47898 88596 47920
rect 85284 47846 86546 47898
rect 86598 47846 86610 47898
rect 86662 47846 86674 47898
rect 86726 47846 86738 47898
rect 86790 47846 86802 47898
rect 86854 47846 88596 47898
rect 85284 47824 88596 47846
rect 87957 47585 88015 47591
rect 85794 47508 85800 47560
rect 85852 47548 85858 47560
rect 87957 47551 87969 47585
rect 88003 47551 88015 47585
rect 87957 47548 88015 47551
rect 85852 47545 88015 47548
rect 85852 47520 88000 47545
rect 85852 47508 85858 47520
rect 88186 47489 88192 47492
rect 88169 47483 88192 47489
rect 88169 47449 88181 47483
rect 88169 47443 88192 47449
rect 88186 47440 88192 47443
rect 88244 47440 88250 47492
rect 4876 47354 7912 47376
rect 4876 47302 6690 47354
rect 6742 47302 6754 47354
rect 6806 47302 6818 47354
rect 6870 47302 6882 47354
rect 6934 47302 6946 47354
rect 6998 47302 7912 47354
rect 4876 47280 7912 47302
rect 85284 47354 88596 47376
rect 85284 47302 87282 47354
rect 87334 47302 87346 47354
rect 87398 47302 87410 47354
rect 87462 47302 87474 47354
rect 87526 47302 87538 47354
rect 87590 47302 88596 47354
rect 85284 47280 88596 47302
rect 88186 46896 88192 46948
rect 88244 46896 88250 46948
rect 4876 46810 7912 46832
rect 4876 46758 5954 46810
rect 6006 46758 6018 46810
rect 6070 46758 6082 46810
rect 6134 46758 6146 46810
rect 6198 46758 6210 46810
rect 6262 46758 7912 46810
rect 4876 46736 7912 46758
rect 85284 46810 88596 46832
rect 85284 46758 86546 46810
rect 86598 46758 86610 46810
rect 86662 46758 86674 46810
rect 86726 46758 86738 46810
rect 86790 46758 86802 46810
rect 86854 46758 88596 46810
rect 85284 46736 88596 46758
rect 4876 46266 7912 46288
rect 4876 46214 6690 46266
rect 6742 46214 6754 46266
rect 6806 46214 6818 46266
rect 6870 46214 6882 46266
rect 6934 46214 6946 46266
rect 6998 46214 7912 46266
rect 4876 46192 7912 46214
rect 85284 46266 88596 46288
rect 85284 46214 87282 46266
rect 87334 46214 87346 46266
rect 87398 46214 87410 46266
rect 87462 46214 87474 46266
rect 87526 46214 87538 46266
rect 87590 46214 88596 46266
rect 85284 46192 88596 46214
rect 5386 45876 5392 45928
rect 5444 45916 5450 45928
rect 13878 45916 13884 45928
rect 5444 45888 13884 45916
rect 5444 45876 5450 45888
rect 13878 45876 13884 45888
rect 13936 45876 13942 45928
rect 46418 45876 46424 45928
rect 46476 45916 46482 45928
rect 51278 45916 51284 45928
rect 46476 45888 51284 45916
rect 46476 45876 46482 45888
rect 51278 45876 51284 45888
rect 51336 45916 51342 45928
rect 85794 45916 85800 45928
rect 51336 45888 85800 45916
rect 51336 45876 51342 45888
rect 85794 45876 85800 45888
rect 85852 45876 85858 45928
rect 88186 45808 88192 45860
rect 88244 45808 88250 45860
rect 4876 45722 7912 45744
rect 4876 45670 5954 45722
rect 6006 45670 6018 45722
rect 6070 45670 6082 45722
rect 6134 45670 6146 45722
rect 6198 45670 6210 45722
rect 6262 45670 7912 45722
rect 4876 45648 7912 45670
rect 85284 45722 88596 45744
rect 85284 45670 86546 45722
rect 86598 45670 86610 45722
rect 86662 45670 86674 45722
rect 86726 45670 86738 45722
rect 86790 45670 86802 45722
rect 86854 45670 88596 45722
rect 85284 45648 88596 45670
rect 5386 45585 5392 45588
rect 5364 45579 5392 45585
rect 5364 45545 5376 45579
rect 5364 45539 5392 45545
rect 5386 45536 5392 45539
rect 5444 45536 5450 45588
rect 7318 45536 7324 45588
rect 7376 45576 7382 45588
rect 9986 45576 9992 45588
rect 7376 45548 9992 45576
rect 7376 45536 7382 45548
rect 9986 45536 9992 45548
rect 10044 45536 10050 45588
rect 85794 45536 85800 45588
rect 85852 45536 85858 45588
rect 7134 45468 7140 45520
rect 7192 45468 7198 45520
rect 85978 45468 85984 45520
rect 86036 45468 86042 45520
rect 5159 45409 5217 45415
rect 5159 45406 5171 45409
rect 2902 45332 2908 45384
rect 2960 45372 2966 45384
rect 4852 45378 5171 45406
rect 4852 45372 4880 45378
rect 2960 45344 4880 45372
rect 5159 45375 5171 45378
rect 5205 45406 5217 45409
rect 5205 45381 5524 45406
rect 5205 45378 5539 45381
rect 5205 45375 5217 45378
rect 5159 45369 5217 45375
rect 5481 45375 5539 45378
rect 2960 45332 2966 45344
rect 5481 45341 5493 45375
rect 5527 45341 5539 45375
rect 5481 45335 5539 45341
rect 86162 45332 86168 45384
rect 86220 45332 86226 45384
rect 88186 45332 88192 45384
rect 88244 45332 88250 45384
rect 85610 45264 85616 45316
rect 85668 45264 85674 45316
rect 4876 45178 7912 45200
rect 4876 45126 6690 45178
rect 6742 45126 6754 45178
rect 6806 45126 6818 45178
rect 6870 45126 6882 45178
rect 6934 45126 6946 45178
rect 6998 45126 7912 45178
rect 4876 45104 7912 45126
rect 85284 45178 88596 45200
rect 85284 45126 87282 45178
rect 87334 45126 87346 45178
rect 87398 45126 87410 45178
rect 87462 45126 87474 45178
rect 87526 45126 87538 45178
rect 87590 45126 88596 45178
rect 85284 45104 88596 45126
rect 7502 44992 7508 45044
rect 7560 44992 7566 45044
rect 88278 44939 88284 44942
rect 5457 44933 5515 44939
rect 5457 44899 5469 44933
rect 5503 44899 5515 44933
rect 88253 44933 88284 44939
rect 5457 44896 5515 44899
rect 7134 44896 7140 44908
rect 5457 44893 7140 44896
rect 5472 44868 7140 44893
rect 7134 44856 7140 44868
rect 7192 44856 7198 44908
rect 87913 44899 87971 44905
rect 87913 44865 87925 44899
rect 87959 44896 87971 44899
rect 88253 44899 88265 44933
rect 88253 44896 88284 44899
rect 87959 44890 88284 44896
rect 88336 44890 88342 44942
rect 87959 44868 88296 44890
rect 87959 44865 87971 44868
rect 87913 44859 87971 44865
rect 87174 44788 87180 44840
rect 87232 44828 87238 44840
rect 88051 44831 88109 44837
rect 88051 44828 88063 44831
rect 87232 44800 88063 44828
rect 87232 44788 87238 44800
rect 88051 44797 88063 44800
rect 88097 44797 88109 44831
rect 88051 44791 88109 44797
rect 2902 44720 2908 44772
rect 2960 44760 2966 44772
rect 5251 44763 5309 44769
rect 5251 44760 5263 44763
rect 2960 44732 5263 44760
rect 2960 44720 2966 44732
rect 5251 44729 5263 44732
rect 5297 44729 5309 44763
rect 5251 44723 5309 44729
rect 4876 44634 7912 44656
rect 4876 44582 5954 44634
rect 6006 44582 6018 44634
rect 6070 44582 6082 44634
rect 6134 44582 6146 44634
rect 6198 44582 6210 44634
rect 6262 44582 7912 44634
rect 4876 44560 7912 44582
rect 85284 44634 88596 44656
rect 85284 44582 86546 44634
rect 86598 44582 86610 44634
rect 86662 44582 86674 44634
rect 86726 44582 86738 44634
rect 86790 44582 86802 44634
rect 86854 44582 88596 44634
rect 85284 44560 88596 44582
rect 87729 44423 87787 44429
rect 87729 44389 87741 44423
rect 87775 44420 87787 44423
rect 87775 44392 88296 44420
rect 87775 44389 87787 44392
rect 87729 44383 87787 44389
rect 5457 44321 5515 44327
rect 88268 44324 88296 44392
rect 88268 44321 88284 44324
rect 5457 44287 5469 44321
rect 5503 44287 5515 44321
rect 88253 44315 88284 44321
rect 5457 44284 5515 44287
rect 8146 44284 8152 44296
rect 5457 44281 8152 44284
rect 5472 44256 8152 44281
rect 8146 44244 8152 44256
rect 8204 44244 8210 44296
rect 85794 44244 85800 44296
rect 85852 44284 85858 44296
rect 85852 44256 88094 44284
rect 88253 44281 88265 44315
rect 88253 44275 88284 44281
rect 88278 44272 88284 44275
rect 88336 44272 88342 44324
rect 85852 44244 85858 44256
rect 2718 44176 2724 44228
rect 2776 44216 2782 44228
rect 88066 44225 88094 44256
rect 5251 44219 5309 44225
rect 5251 44216 5263 44219
rect 2776 44188 5263 44216
rect 2776 44176 2782 44188
rect 5251 44185 5263 44188
rect 5297 44185 5309 44219
rect 5251 44179 5309 44185
rect 88051 44219 88109 44225
rect 88051 44185 88063 44219
rect 88097 44185 88109 44219
rect 88051 44179 88109 44185
rect 4876 44090 7912 44112
rect 4876 44038 6690 44090
rect 6742 44038 6754 44090
rect 6806 44038 6818 44090
rect 6870 44038 6882 44090
rect 6934 44038 6946 44090
rect 6998 44038 7912 44090
rect 4876 44016 7912 44038
rect 85284 44090 88596 44112
rect 85284 44038 87282 44090
rect 87334 44038 87346 44090
rect 87398 44038 87410 44090
rect 87462 44038 87474 44090
rect 87526 44038 87538 44090
rect 87590 44038 88596 44090
rect 85284 44016 88596 44038
rect 4876 43546 7912 43568
rect 4876 43494 5954 43546
rect 6006 43494 6018 43546
rect 6070 43494 6082 43546
rect 6134 43494 6146 43546
rect 6198 43494 6210 43546
rect 6262 43494 7912 43546
rect 4876 43472 7912 43494
rect 85284 43546 88596 43568
rect 85284 43494 86546 43546
rect 86598 43494 86610 43546
rect 86662 43494 86674 43546
rect 86726 43494 86738 43546
rect 86790 43494 86802 43546
rect 86854 43494 88596 43546
rect 85284 43472 88596 43494
rect 4876 43002 7912 43024
rect 4876 42950 6690 43002
rect 6742 42950 6754 43002
rect 6806 42950 6818 43002
rect 6870 42950 6882 43002
rect 6934 42950 6946 43002
rect 6998 42950 7912 43002
rect 4876 42928 7912 42950
rect 85284 43002 88596 43024
rect 85284 42950 87282 43002
rect 87334 42950 87346 43002
rect 87398 42950 87410 43002
rect 87462 42950 87474 43002
rect 87526 42950 87538 43002
rect 87590 42950 88596 43002
rect 85284 42928 88596 42950
rect 88278 42763 88284 42766
rect 5457 42757 5515 42763
rect 5457 42723 5469 42757
rect 5503 42723 5515 42757
rect 88253 42757 88284 42763
rect 88253 42754 88265 42757
rect 5457 42720 5515 42723
rect 7134 42720 7140 42732
rect 5457 42717 7140 42720
rect 5472 42692 7140 42717
rect 7134 42680 7140 42692
rect 7192 42680 7198 42732
rect 87913 42723 87971 42729
rect 87913 42689 87925 42723
rect 87959 42720 87971 42723
rect 88250 42723 88265 42754
rect 88250 42720 88284 42723
rect 87959 42714 88284 42720
rect 88336 42714 88342 42766
rect 87959 42692 88278 42714
rect 87959 42689 87971 42692
rect 87913 42683 87971 42689
rect 86346 42612 86352 42664
rect 86404 42652 86410 42664
rect 88051 42655 88109 42661
rect 88051 42652 88063 42655
rect 86404 42624 88063 42652
rect 86404 42612 86410 42624
rect 88051 42621 88063 42624
rect 88097 42621 88109 42655
rect 88051 42615 88109 42621
rect 2902 42544 2908 42596
rect 2960 42584 2966 42596
rect 5251 42587 5309 42593
rect 5251 42584 5263 42587
rect 2960 42556 5263 42584
rect 2960 42544 2966 42556
rect 5251 42553 5263 42556
rect 5297 42553 5309 42587
rect 5251 42547 5309 42553
rect 4876 42458 7912 42480
rect 4876 42406 5954 42458
rect 6006 42406 6018 42458
rect 6070 42406 6082 42458
rect 6134 42406 6146 42458
rect 6198 42406 6210 42458
rect 6262 42406 7912 42458
rect 4876 42384 7912 42406
rect 85284 42458 88596 42480
rect 85284 42406 86546 42458
rect 86598 42406 86610 42458
rect 86662 42406 86674 42458
rect 86726 42406 86738 42458
rect 86790 42406 86802 42458
rect 86854 42406 88596 42458
rect 85284 42384 88596 42406
rect 4876 41914 7912 41936
rect 4876 41862 6690 41914
rect 6742 41862 6754 41914
rect 6806 41862 6818 41914
rect 6870 41862 6882 41914
rect 6934 41862 6946 41914
rect 6998 41862 7912 41914
rect 4876 41840 7912 41862
rect 85284 41914 88596 41936
rect 85284 41862 87282 41914
rect 87334 41862 87346 41914
rect 87398 41862 87410 41914
rect 87462 41862 87474 41914
rect 87526 41862 87538 41914
rect 87590 41862 88596 41914
rect 85284 41840 88596 41862
rect 4374 41728 4380 41780
rect 4432 41768 4438 41780
rect 5251 41771 5309 41777
rect 5251 41768 5263 41771
rect 4432 41740 5263 41768
rect 4432 41728 4438 41740
rect 5251 41737 5263 41740
rect 5297 41737 5309 41771
rect 5251 41731 5309 41737
rect 87174 41728 87180 41780
rect 87232 41768 87238 41780
rect 88051 41771 88109 41777
rect 88051 41768 88063 41771
rect 87232 41740 88063 41768
rect 87232 41728 87238 41740
rect 88051 41737 88063 41740
rect 88097 41737 88109 41771
rect 88051 41731 88109 41737
rect 5457 41669 5515 41675
rect 5457 41635 5469 41669
rect 5503 41666 5515 41669
rect 5662 41666 5668 41678
rect 5503 41638 5668 41666
rect 5503 41635 5515 41638
rect 5457 41629 5515 41635
rect 5662 41626 5668 41638
rect 5720 41626 5726 41678
rect 88278 41675 88284 41678
rect 88253 41669 88284 41675
rect 88253 41666 88265 41669
rect 87913 41635 87971 41641
rect 87913 41601 87925 41635
rect 87959 41632 87971 41635
rect 88250 41635 88265 41666
rect 88250 41632 88284 41635
rect 87959 41626 88284 41632
rect 88336 41626 88342 41678
rect 87959 41604 88278 41626
rect 87959 41601 87971 41604
rect 87913 41595 87971 41601
rect 4876 41370 7912 41392
rect 4876 41318 5954 41370
rect 6006 41318 6018 41370
rect 6070 41318 6082 41370
rect 6134 41318 6146 41370
rect 6198 41318 6210 41370
rect 6262 41318 7912 41370
rect 4876 41296 7912 41318
rect 85284 41370 88596 41392
rect 85284 41318 86546 41370
rect 86598 41318 86610 41370
rect 86662 41318 86674 41370
rect 86726 41318 86738 41370
rect 86790 41318 86802 41370
rect 86854 41318 88596 41370
rect 85284 41296 88596 41318
rect 4876 40826 7912 40848
rect 4876 40774 6690 40826
rect 6742 40774 6754 40826
rect 6806 40774 6818 40826
rect 6870 40774 6882 40826
rect 6934 40774 6946 40826
rect 6998 40774 7912 40826
rect 4876 40752 7912 40774
rect 85284 40826 88596 40848
rect 85284 40774 87282 40826
rect 87334 40774 87346 40826
rect 87398 40774 87410 40826
rect 87462 40774 87474 40826
rect 87526 40774 87538 40826
rect 87590 40774 88596 40826
rect 85284 40752 88596 40774
rect 5457 40581 5515 40587
rect 5457 40547 5469 40581
rect 5503 40547 5515 40581
rect 5457 40544 5515 40547
rect 7134 40544 7140 40556
rect 5457 40541 7140 40544
rect 5472 40516 7140 40541
rect 7134 40504 7140 40516
rect 7192 40504 7198 40556
rect 87910 40504 87916 40556
rect 87968 40504 87974 40556
rect 88278 40553 88284 40556
rect 88257 40547 88284 40553
rect 88257 40513 88269 40547
rect 88257 40507 88284 40513
rect 88278 40504 88284 40507
rect 88336 40504 88342 40556
rect 2902 40368 2908 40420
rect 2960 40408 2966 40420
rect 5251 40411 5309 40417
rect 5251 40408 5263 40411
rect 2960 40380 5263 40408
rect 2960 40368 2966 40380
rect 5251 40377 5263 40380
rect 5297 40377 5309 40411
rect 5251 40371 5309 40377
rect 4876 40282 7912 40304
rect 4876 40230 5954 40282
rect 6006 40230 6018 40282
rect 6070 40230 6082 40282
rect 6134 40230 6146 40282
rect 6198 40230 6210 40282
rect 6262 40230 7912 40282
rect 4876 40208 7912 40230
rect 85284 40282 88596 40304
rect 85284 40230 86546 40282
rect 86598 40230 86610 40282
rect 86662 40230 86674 40282
rect 86726 40230 86738 40282
rect 86790 40230 86802 40282
rect 86854 40230 88596 40282
rect 85284 40208 88596 40230
rect 88189 40139 88247 40145
rect 88189 40105 88201 40139
rect 88235 40136 88247 40139
rect 88278 40136 88284 40148
rect 88235 40108 88284 40136
rect 88235 40105 88247 40108
rect 88189 40099 88247 40105
rect 88278 40096 88284 40108
rect 88336 40096 88342 40148
rect 4876 39738 7912 39760
rect 4876 39686 6690 39738
rect 6742 39686 6754 39738
rect 6806 39686 6818 39738
rect 6870 39686 6882 39738
rect 6934 39686 6946 39738
rect 6998 39686 7912 39738
rect 4876 39664 7912 39686
rect 85284 39738 88596 39760
rect 85284 39686 87282 39738
rect 87334 39686 87346 39738
rect 87398 39686 87410 39738
rect 87462 39686 87474 39738
rect 87526 39686 87538 39738
rect 87590 39686 88596 39738
rect 85284 39664 88596 39686
rect 88278 39499 88284 39502
rect 5457 39493 5515 39499
rect 5457 39459 5469 39493
rect 5503 39459 5515 39493
rect 88257 39493 88284 39499
rect 88257 39490 88269 39493
rect 5457 39456 5515 39459
rect 7134 39456 7140 39468
rect 5457 39453 7140 39456
rect 5472 39428 7140 39453
rect 7134 39416 7140 39428
rect 7192 39416 7198 39468
rect 87821 39459 87879 39465
rect 87821 39425 87833 39459
rect 87867 39456 87879 39459
rect 88250 39459 88269 39490
rect 88250 39456 88284 39459
rect 87867 39450 88284 39456
rect 88336 39450 88342 39502
rect 87867 39428 88278 39450
rect 87867 39425 87879 39428
rect 87821 39419 87879 39425
rect 87174 39348 87180 39400
rect 87232 39388 87238 39400
rect 88051 39391 88109 39397
rect 88051 39388 88063 39391
rect 87232 39360 88063 39388
rect 87232 39348 87238 39360
rect 88051 39357 88063 39360
rect 88097 39357 88109 39391
rect 88051 39351 88109 39357
rect 2902 39280 2908 39332
rect 2960 39320 2966 39332
rect 5251 39323 5309 39329
rect 5251 39320 5263 39323
rect 2960 39292 5263 39320
rect 2960 39280 2966 39292
rect 5251 39289 5263 39292
rect 5297 39289 5309 39323
rect 5251 39283 5309 39289
rect 4876 39194 7912 39216
rect 4876 39142 5954 39194
rect 6006 39142 6018 39194
rect 6070 39142 6082 39194
rect 6134 39142 6146 39194
rect 6198 39142 6210 39194
rect 6262 39142 7912 39194
rect 4876 39120 7912 39142
rect 85284 39194 88596 39216
rect 85284 39142 86546 39194
rect 86598 39142 86610 39194
rect 86662 39142 86674 39194
rect 86726 39142 86738 39194
rect 86790 39142 86802 39194
rect 86854 39142 88596 39194
rect 85284 39120 88596 39142
rect 4374 38940 4380 38992
rect 4432 38980 4438 38992
rect 5251 38983 5309 38989
rect 5251 38980 5263 38983
rect 4432 38952 5263 38980
rect 4432 38940 4438 38952
rect 5251 38949 5263 38952
rect 5297 38949 5309 38983
rect 5251 38943 5309 38949
rect 84414 38940 84420 38992
rect 84472 38980 84478 38992
rect 88051 38983 88109 38989
rect 88051 38980 88063 38983
rect 84472 38952 88063 38980
rect 84472 38940 84478 38952
rect 88051 38949 88063 38952
rect 88097 38949 88109 38983
rect 88051 38943 88109 38949
rect 88278 38887 88284 38890
rect 5457 38881 5515 38887
rect 5457 38847 5469 38881
rect 5503 38847 5515 38881
rect 88257 38881 88284 38887
rect 88257 38878 88269 38881
rect 5457 38844 5515 38847
rect 7778 38844 7784 38856
rect 5457 38841 7784 38844
rect 5472 38816 7784 38841
rect 7778 38804 7784 38816
rect 7836 38804 7842 38856
rect 87729 38847 87787 38853
rect 87729 38813 87741 38847
rect 87775 38844 87787 38847
rect 88250 38847 88269 38878
rect 88250 38844 88284 38847
rect 87775 38838 88284 38844
rect 88336 38838 88342 38890
rect 87775 38816 88278 38838
rect 87775 38813 87787 38816
rect 87729 38807 87787 38813
rect 4876 38650 7912 38672
rect 4876 38598 6690 38650
rect 6742 38598 6754 38650
rect 6806 38598 6818 38650
rect 6870 38598 6882 38650
rect 6934 38598 6946 38650
rect 6998 38598 7912 38650
rect 4876 38576 7912 38598
rect 85284 38650 88596 38672
rect 85284 38598 87282 38650
rect 87334 38598 87346 38650
rect 87398 38598 87410 38650
rect 87462 38598 87474 38650
rect 87526 38598 87538 38650
rect 87590 38598 88596 38650
rect 85284 38576 88596 38598
rect 4876 38106 7912 38128
rect 4876 38054 5954 38106
rect 6006 38054 6018 38106
rect 6070 38054 6082 38106
rect 6134 38054 6146 38106
rect 6198 38054 6210 38106
rect 6262 38054 7912 38106
rect 4876 38032 7912 38054
rect 85284 38106 88596 38128
rect 85284 38054 86546 38106
rect 86598 38054 86610 38106
rect 86662 38054 86674 38106
rect 86726 38054 86738 38106
rect 86790 38054 86802 38106
rect 86854 38054 88596 38106
rect 85284 38032 88596 38054
rect 4876 37562 7912 37584
rect 4876 37510 6690 37562
rect 6742 37510 6754 37562
rect 6806 37510 6818 37562
rect 6870 37510 6882 37562
rect 6934 37510 6946 37562
rect 6998 37510 7912 37562
rect 4876 37488 7912 37510
rect 85284 37562 88596 37584
rect 85284 37510 87282 37562
rect 87334 37510 87346 37562
rect 87398 37510 87410 37562
rect 87462 37510 87474 37562
rect 87526 37510 87538 37562
rect 87590 37510 88596 37562
rect 85284 37488 88596 37510
rect 88278 37323 88284 37326
rect 5457 37317 5515 37323
rect 5457 37283 5469 37317
rect 5503 37314 5515 37317
rect 88253 37317 88284 37323
rect 88253 37314 88265 37317
rect 5503 37286 5800 37314
rect 5503 37283 5515 37286
rect 5457 37277 5515 37283
rect 5772 37280 5800 37286
rect 7226 37280 7232 37292
rect 5772 37252 7232 37280
rect 7226 37240 7232 37252
rect 7284 37240 7290 37292
rect 87928 37289 88265 37314
rect 87913 37286 88265 37289
rect 87913 37283 87971 37286
rect 87913 37249 87925 37283
rect 87959 37249 87971 37283
rect 88253 37283 88265 37286
rect 88253 37277 88284 37283
rect 88278 37274 88284 37277
rect 88336 37274 88342 37326
rect 87913 37243 87971 37249
rect 86346 37172 86352 37224
rect 86404 37212 86410 37224
rect 88051 37215 88109 37221
rect 88051 37212 88063 37215
rect 86404 37184 88063 37212
rect 86404 37172 86410 37184
rect 88051 37181 88063 37184
rect 88097 37181 88109 37215
rect 88051 37175 88109 37181
rect 2902 37104 2908 37156
rect 2960 37144 2966 37156
rect 5251 37147 5309 37153
rect 5251 37144 5263 37147
rect 2960 37116 5263 37144
rect 2960 37104 2966 37116
rect 5251 37113 5263 37116
rect 5297 37113 5309 37147
rect 5251 37107 5309 37113
rect 4876 37018 7912 37040
rect 4876 36966 5954 37018
rect 6006 36966 6018 37018
rect 6070 36966 6082 37018
rect 6134 36966 6146 37018
rect 6198 36966 6210 37018
rect 6262 36966 7912 37018
rect 4876 36944 7912 36966
rect 85284 37018 88596 37040
rect 85284 36966 86546 37018
rect 86598 36966 86610 37018
rect 86662 36966 86674 37018
rect 86726 36966 86738 37018
rect 86790 36966 86802 37018
rect 86854 36966 88596 37018
rect 85284 36944 88596 36966
rect 4876 36474 7912 36496
rect 4876 36422 6690 36474
rect 6742 36422 6754 36474
rect 6806 36422 6818 36474
rect 6870 36422 6882 36474
rect 6934 36422 6946 36474
rect 6998 36422 7912 36474
rect 4876 36400 7912 36422
rect 85284 36474 88596 36496
rect 85284 36422 87282 36474
rect 87334 36422 87346 36474
rect 87398 36422 87410 36474
rect 87462 36422 87474 36474
rect 87526 36422 87538 36474
rect 87590 36422 88596 36474
rect 85284 36400 88596 36422
rect 5457 36229 5515 36235
rect 5457 36195 5469 36229
rect 5503 36226 5515 36229
rect 5662 36226 5668 36238
rect 5503 36198 5668 36226
rect 5503 36195 5515 36198
rect 5457 36189 5515 36195
rect 5662 36186 5668 36198
rect 5720 36186 5726 36238
rect 88253 36229 88311 36235
rect 88253 36226 88265 36229
rect 87928 36201 88265 36226
rect 87913 36198 88265 36201
rect 87913 36195 87971 36198
rect 87913 36161 87925 36195
rect 87959 36161 87971 36195
rect 88253 36195 88265 36198
rect 88299 36226 88311 36229
rect 88299 36204 88600 36226
rect 88299 36198 88560 36204
rect 88299 36195 88311 36198
rect 88253 36189 88311 36195
rect 87913 36155 87971 36161
rect 88554 36152 88560 36198
rect 88612 36152 88618 36204
rect 4374 36084 4380 36136
rect 4432 36124 4438 36136
rect 5251 36127 5309 36133
rect 5251 36124 5263 36127
rect 4432 36096 5263 36124
rect 4432 36084 4438 36096
rect 5251 36093 5263 36096
rect 5297 36093 5309 36127
rect 5251 36087 5309 36093
rect 84414 36084 84420 36136
rect 84472 36124 84478 36136
rect 88051 36127 88109 36133
rect 88051 36124 88063 36127
rect 84472 36096 88063 36124
rect 84472 36084 84478 36096
rect 88051 36093 88063 36096
rect 88097 36093 88109 36127
rect 88051 36087 88109 36093
rect 4876 35930 7912 35952
rect 4876 35878 5954 35930
rect 6006 35878 6018 35930
rect 6070 35878 6082 35930
rect 6134 35878 6146 35930
rect 6198 35878 6210 35930
rect 6262 35878 7912 35930
rect 4876 35856 7912 35878
rect 85284 35930 88596 35952
rect 85284 35878 86546 35930
rect 86598 35878 86610 35930
rect 86662 35878 86674 35930
rect 86726 35878 86738 35930
rect 86790 35878 86802 35930
rect 86854 35878 88596 35930
rect 85284 35856 88596 35878
rect 4876 35386 7912 35408
rect 4876 35334 6690 35386
rect 6742 35334 6754 35386
rect 6806 35334 6818 35386
rect 6870 35334 6882 35386
rect 6934 35334 6946 35386
rect 6998 35334 7912 35386
rect 4876 35312 7912 35334
rect 85284 35386 88596 35408
rect 85284 35334 87282 35386
rect 87334 35334 87346 35386
rect 87398 35334 87410 35386
rect 87462 35334 87474 35386
rect 87526 35334 87538 35386
rect 87590 35334 88596 35386
rect 85284 35312 88596 35334
rect 88278 35147 88284 35150
rect 5457 35141 5515 35147
rect 5457 35107 5469 35141
rect 5503 35138 5515 35141
rect 88253 35141 88284 35147
rect 88253 35138 88265 35141
rect 5503 35110 5800 35138
rect 5503 35107 5515 35110
rect 5457 35101 5515 35107
rect 5772 35104 5800 35110
rect 7226 35104 7232 35116
rect 5772 35076 7232 35104
rect 7226 35064 7232 35076
rect 7284 35064 7290 35116
rect 87928 35113 88265 35138
rect 87913 35110 88265 35113
rect 87913 35107 87971 35110
rect 87913 35073 87925 35107
rect 87959 35073 87971 35107
rect 88253 35107 88265 35110
rect 88253 35101 88284 35107
rect 88278 35098 88284 35101
rect 88336 35098 88342 35150
rect 87913 35067 87971 35073
rect 86346 34996 86352 35048
rect 86404 35036 86410 35048
rect 88051 35039 88109 35045
rect 88051 35036 88063 35039
rect 86404 35008 88063 35036
rect 86404 34996 86410 35008
rect 88051 35005 88063 35008
rect 88097 35005 88109 35039
rect 88051 34999 88109 35005
rect 2902 34928 2908 34980
rect 2960 34968 2966 34980
rect 5251 34971 5309 34977
rect 5251 34968 5263 34971
rect 2960 34940 5263 34968
rect 2960 34928 2966 34940
rect 5251 34937 5263 34940
rect 5297 34937 5309 34971
rect 5251 34931 5309 34937
rect 4876 34842 7912 34864
rect 4876 34790 5954 34842
rect 6006 34790 6018 34842
rect 6070 34790 6082 34842
rect 6134 34790 6146 34842
rect 6198 34790 6210 34842
rect 6262 34790 7912 34842
rect 4876 34768 7912 34790
rect 85284 34842 88596 34864
rect 85284 34790 86546 34842
rect 86598 34790 86610 34842
rect 86662 34790 86674 34842
rect 86726 34790 86738 34842
rect 86790 34790 86802 34842
rect 86854 34790 88596 34842
rect 85284 34768 88596 34790
rect 4876 34298 7912 34320
rect 4876 34246 6690 34298
rect 6742 34246 6754 34298
rect 6806 34246 6818 34298
rect 6870 34246 6882 34298
rect 6934 34246 6946 34298
rect 6998 34246 7912 34298
rect 4876 34224 7912 34246
rect 85284 34298 88596 34320
rect 85284 34246 87282 34298
rect 87334 34246 87346 34298
rect 87398 34246 87410 34298
rect 87462 34246 87474 34298
rect 87526 34246 87538 34298
rect 87590 34246 88596 34298
rect 85284 34224 88596 34246
rect 87913 34155 87971 34161
rect 87913 34121 87925 34155
rect 87959 34152 87971 34155
rect 87959 34124 88324 34152
rect 87959 34121 87971 34124
rect 87913 34115 87971 34121
rect 88296 34062 88324 34124
rect 88278 34059 88284 34062
rect 5457 34053 5515 34059
rect 5457 34019 5469 34053
rect 5503 34050 5515 34053
rect 88253 34053 88284 34059
rect 5503 34022 5800 34050
rect 5503 34019 5515 34022
rect 5457 34013 5515 34019
rect 5772 34016 5800 34022
rect 7226 34016 7232 34028
rect 5772 33988 7232 34016
rect 7226 33976 7232 33988
rect 7284 33976 7290 34028
rect 88253 34019 88265 34053
rect 88253 34013 88284 34019
rect 88278 34010 88284 34013
rect 88336 34010 88342 34062
rect 86346 33908 86352 33960
rect 86404 33948 86410 33960
rect 88051 33951 88109 33957
rect 88051 33948 88063 33951
rect 86404 33920 88063 33948
rect 86404 33908 86410 33920
rect 88051 33917 88063 33920
rect 88097 33917 88109 33951
rect 88051 33911 88109 33917
rect 2902 33840 2908 33892
rect 2960 33880 2966 33892
rect 5251 33883 5309 33889
rect 5251 33880 5263 33883
rect 2960 33852 5263 33880
rect 2960 33840 2966 33852
rect 5251 33849 5263 33852
rect 5297 33849 5309 33883
rect 5251 33843 5309 33849
rect 4876 33754 7912 33776
rect 4876 33702 5954 33754
rect 6006 33702 6018 33754
rect 6070 33702 6082 33754
rect 6134 33702 6146 33754
rect 6198 33702 6210 33754
rect 6262 33702 7912 33754
rect 4876 33680 7912 33702
rect 85284 33754 88596 33776
rect 85284 33702 86546 33754
rect 86598 33702 86610 33754
rect 86662 33702 86674 33754
rect 86726 33702 86738 33754
rect 86790 33702 86802 33754
rect 86854 33702 88596 33754
rect 85284 33680 88596 33702
rect 4374 33500 4380 33552
rect 4432 33540 4438 33552
rect 5251 33543 5309 33549
rect 5251 33540 5263 33543
rect 4432 33512 5263 33540
rect 4432 33500 4438 33512
rect 5251 33509 5263 33512
rect 5297 33509 5309 33543
rect 5251 33503 5309 33509
rect 87729 33543 87787 33549
rect 87729 33509 87741 33543
rect 87775 33540 87787 33543
rect 87775 33512 88324 33540
rect 87775 33509 87787 33512
rect 87729 33503 87787 33509
rect 5457 33441 5515 33447
rect 5457 33407 5469 33441
rect 5503 33438 5515 33441
rect 5662 33438 5668 33450
rect 5503 33410 5668 33438
rect 5503 33407 5515 33410
rect 5457 33401 5515 33407
rect 5662 33398 5668 33410
rect 5720 33398 5726 33450
rect 88296 33441 88324 33512
rect 88253 33435 88324 33441
rect 84414 33364 84420 33416
rect 84472 33404 84478 33416
rect 88051 33407 88109 33413
rect 88051 33404 88063 33407
rect 84472 33376 88063 33404
rect 84472 33364 84478 33376
rect 88051 33373 88063 33376
rect 88097 33373 88109 33407
rect 88253 33401 88265 33435
rect 88299 33432 88324 33435
rect 88299 33416 88600 33432
rect 88299 33404 88560 33416
rect 88299 33401 88311 33404
rect 88253 33395 88311 33401
rect 88051 33367 88109 33373
rect 88554 33364 88560 33404
rect 88612 33364 88618 33416
rect 4876 33210 7912 33232
rect 4876 33158 6690 33210
rect 6742 33158 6754 33210
rect 6806 33158 6818 33210
rect 6870 33158 6882 33210
rect 6934 33158 6946 33210
rect 6998 33158 7912 33210
rect 4876 33136 7912 33158
rect 85284 33210 88596 33232
rect 85284 33158 87282 33210
rect 87334 33158 87346 33210
rect 87398 33158 87410 33210
rect 87462 33158 87474 33210
rect 87526 33158 87538 33210
rect 87590 33158 88596 33210
rect 85284 33136 88596 33158
rect 4876 32666 7912 32688
rect 4876 32614 5954 32666
rect 6006 32614 6018 32666
rect 6070 32614 6082 32666
rect 6134 32614 6146 32666
rect 6198 32614 6210 32666
rect 6262 32614 7912 32666
rect 4876 32592 7912 32614
rect 85284 32666 88596 32688
rect 85284 32614 86546 32666
rect 86598 32614 86610 32666
rect 86662 32614 86674 32666
rect 86726 32614 86738 32666
rect 86790 32614 86802 32666
rect 86854 32614 88596 32666
rect 85284 32592 88596 32614
rect 4876 32122 7912 32144
rect 4876 32070 6690 32122
rect 6742 32070 6754 32122
rect 6806 32070 6818 32122
rect 6870 32070 6882 32122
rect 6934 32070 6946 32122
rect 6998 32070 7912 32122
rect 4876 32048 7912 32070
rect 85284 32122 88596 32144
rect 85284 32070 87282 32122
rect 87334 32070 87346 32122
rect 87398 32070 87410 32122
rect 87462 32070 87474 32122
rect 87526 32070 87538 32122
rect 87590 32070 88596 32122
rect 85284 32048 88596 32070
rect 88278 31883 88284 31886
rect 5457 31877 5515 31883
rect 5457 31843 5469 31877
rect 5503 31874 5515 31877
rect 88253 31877 88284 31883
rect 88253 31874 88265 31877
rect 5503 31846 5800 31874
rect 5503 31843 5515 31846
rect 5457 31837 5515 31843
rect 5772 31840 5800 31846
rect 7226 31840 7232 31852
rect 5772 31812 7232 31840
rect 7226 31800 7232 31812
rect 7284 31800 7290 31852
rect 87913 31843 87971 31849
rect 87913 31809 87925 31843
rect 87959 31840 87971 31843
rect 88112 31846 88265 31874
rect 88112 31840 88140 31846
rect 87959 31812 88140 31840
rect 88253 31843 88265 31846
rect 88253 31837 88284 31843
rect 88278 31834 88284 31837
rect 88336 31834 88342 31886
rect 87959 31809 87971 31812
rect 87913 31803 87971 31809
rect 86346 31732 86352 31784
rect 86404 31772 86410 31784
rect 88051 31775 88109 31781
rect 88051 31772 88063 31775
rect 86404 31744 88063 31772
rect 86404 31732 86410 31744
rect 88051 31741 88063 31744
rect 88097 31741 88109 31775
rect 88051 31735 88109 31741
rect 2902 31664 2908 31716
rect 2960 31704 2966 31716
rect 5251 31707 5309 31713
rect 5251 31704 5263 31707
rect 2960 31676 5263 31704
rect 2960 31664 2966 31676
rect 5251 31673 5263 31676
rect 5297 31673 5309 31707
rect 5251 31667 5309 31673
rect 4876 31578 7912 31600
rect 4876 31526 5954 31578
rect 6006 31526 6018 31578
rect 6070 31526 6082 31578
rect 6134 31526 6146 31578
rect 6198 31526 6210 31578
rect 6262 31526 7912 31578
rect 4876 31504 7912 31526
rect 85284 31578 88596 31600
rect 85284 31526 86546 31578
rect 86598 31526 86610 31578
rect 86662 31526 86674 31578
rect 86726 31526 86738 31578
rect 86790 31526 86802 31578
rect 86854 31526 88596 31578
rect 85284 31504 88596 31526
rect 4876 31034 7912 31056
rect 4876 30982 6690 31034
rect 6742 30982 6754 31034
rect 6806 30982 6818 31034
rect 6870 30982 6882 31034
rect 6934 30982 6946 31034
rect 6998 30982 7912 31034
rect 4876 30960 7912 30982
rect 85284 31034 88596 31056
rect 85284 30982 87282 31034
rect 87334 30982 87346 31034
rect 87398 30982 87410 31034
rect 87462 30982 87474 31034
rect 87526 30982 87538 31034
rect 87590 30982 88596 31034
rect 85284 30960 88596 30982
rect 5457 30789 5515 30795
rect 5457 30755 5469 30789
rect 5503 30786 5515 30789
rect 5662 30786 5668 30798
rect 5503 30758 5668 30786
rect 5503 30755 5515 30758
rect 5457 30749 5515 30755
rect 5662 30746 5668 30758
rect 5720 30746 5726 30798
rect 88253 30789 88311 30795
rect 88253 30786 88265 30789
rect 87928 30761 88265 30786
rect 87913 30758 88265 30761
rect 87913 30755 87971 30758
rect 87913 30721 87925 30755
rect 87959 30721 87971 30755
rect 88253 30755 88265 30758
rect 88299 30786 88311 30789
rect 88299 30764 88600 30786
rect 88299 30758 88560 30764
rect 88299 30755 88311 30758
rect 88253 30749 88311 30755
rect 87913 30715 87971 30721
rect 88554 30712 88560 30758
rect 88612 30712 88618 30764
rect 88051 30687 88109 30693
rect 88051 30684 88063 30687
rect 85766 30656 88063 30684
rect 4374 30576 4380 30628
rect 4432 30616 4438 30628
rect 5251 30619 5309 30625
rect 5251 30616 5263 30619
rect 4432 30588 5263 30616
rect 4432 30576 4438 30588
rect 5251 30585 5263 30588
rect 5297 30585 5309 30619
rect 5251 30579 5309 30585
rect 84414 30576 84420 30628
rect 84472 30616 84478 30628
rect 85766 30616 85794 30656
rect 88051 30653 88063 30656
rect 88097 30653 88109 30687
rect 88051 30647 88109 30653
rect 84472 30588 85794 30616
rect 84472 30576 84478 30588
rect 4876 30490 7912 30512
rect 4876 30438 5954 30490
rect 6006 30438 6018 30490
rect 6070 30438 6082 30490
rect 6134 30438 6146 30490
rect 6198 30438 6210 30490
rect 6262 30438 7912 30490
rect 4876 30416 7912 30438
rect 85284 30490 88596 30512
rect 85284 30438 86546 30490
rect 86598 30438 86610 30490
rect 86662 30438 86674 30490
rect 86726 30438 86738 30490
rect 86790 30438 86802 30490
rect 86854 30438 88596 30490
rect 85284 30416 88596 30438
rect 4876 29946 7912 29968
rect 4876 29894 6690 29946
rect 6742 29894 6754 29946
rect 6806 29894 6818 29946
rect 6870 29894 6882 29946
rect 6934 29894 6946 29946
rect 6998 29894 7912 29946
rect 4876 29872 7912 29894
rect 85284 29946 88596 29968
rect 85284 29894 87282 29946
rect 87334 29894 87346 29946
rect 87398 29894 87410 29946
rect 87462 29894 87474 29946
rect 87526 29894 87538 29946
rect 87590 29894 88596 29946
rect 85284 29872 88596 29894
rect 5159 29701 5217 29707
rect 5159 29698 5171 29701
rect 2902 29624 2908 29676
rect 2960 29664 2966 29676
rect 4852 29670 5171 29698
rect 4852 29664 4880 29670
rect 2960 29636 4880 29664
rect 5159 29667 5171 29670
rect 5205 29698 5217 29701
rect 87957 29701 88015 29707
rect 87957 29698 87969 29701
rect 5205 29673 5524 29698
rect 5205 29670 5539 29673
rect 5205 29667 5217 29670
rect 5159 29661 5217 29667
rect 5481 29667 5539 29670
rect 2960 29624 2966 29636
rect 5481 29633 5493 29667
rect 5527 29633 5539 29667
rect 5481 29627 5539 29633
rect 86346 29624 86352 29676
rect 86404 29664 86410 29676
rect 87652 29670 87969 29698
rect 87652 29664 87680 29670
rect 86404 29636 87680 29664
rect 87957 29667 87969 29670
rect 88003 29667 88015 29701
rect 87957 29661 88015 29667
rect 86404 29624 86410 29636
rect 5365 29599 5423 29605
rect 5365 29565 5377 29599
rect 5411 29596 5423 29599
rect 7226 29596 7232 29608
rect 5411 29568 7232 29596
rect 5411 29565 5423 29568
rect 5365 29559 5423 29565
rect 7226 29556 7232 29568
rect 7284 29556 7290 29608
rect 88169 29531 88227 29537
rect 88169 29497 88181 29531
rect 88215 29528 88227 29531
rect 88278 29528 88284 29540
rect 88215 29500 88284 29528
rect 88215 29497 88227 29500
rect 88169 29491 88227 29497
rect 88278 29488 88284 29500
rect 88336 29488 88342 29540
rect 4876 29402 7912 29424
rect 4876 29350 5954 29402
rect 6006 29350 6018 29402
rect 6070 29350 6082 29402
rect 6134 29350 6146 29402
rect 6198 29350 6210 29402
rect 6262 29350 7912 29402
rect 4876 29328 7912 29350
rect 85284 29402 88596 29424
rect 85284 29350 86546 29402
rect 86598 29350 86610 29402
rect 86662 29350 86674 29402
rect 86726 29350 86738 29402
rect 86790 29350 86802 29402
rect 86854 29350 88596 29402
rect 85284 29328 88596 29350
rect 4876 28858 7912 28880
rect 4876 28806 6690 28858
rect 6742 28806 6754 28858
rect 6806 28806 6818 28858
rect 6870 28806 6882 28858
rect 6934 28806 6946 28858
rect 6998 28806 7912 28858
rect 4876 28784 7912 28806
rect 85284 28858 88596 28880
rect 85284 28806 87282 28858
rect 87334 28806 87346 28858
rect 87398 28806 87410 28858
rect 87462 28806 87474 28858
rect 87526 28806 87538 28858
rect 87590 28806 88596 28858
rect 85284 28784 88596 28806
rect 5159 28613 5217 28619
rect 5159 28610 5171 28613
rect 2902 28536 2908 28588
rect 2960 28576 2966 28588
rect 4852 28582 5171 28610
rect 4852 28576 4880 28582
rect 2960 28548 4880 28576
rect 5159 28579 5171 28582
rect 5205 28610 5217 28613
rect 87957 28613 88015 28619
rect 87957 28610 87969 28613
rect 5205 28585 5524 28610
rect 5205 28582 5539 28585
rect 5205 28579 5217 28582
rect 5159 28573 5217 28579
rect 5481 28579 5539 28582
rect 2960 28536 2966 28548
rect 5481 28545 5493 28579
rect 5527 28545 5539 28579
rect 5481 28539 5539 28545
rect 86346 28536 86352 28588
rect 86404 28576 86410 28588
rect 87652 28582 87969 28610
rect 87652 28576 87680 28582
rect 86404 28548 87680 28576
rect 87957 28579 87969 28582
rect 88003 28579 88015 28613
rect 87957 28573 88015 28579
rect 86404 28536 86410 28548
rect 5365 28511 5423 28517
rect 5365 28477 5377 28511
rect 5411 28508 5423 28511
rect 7226 28508 7232 28520
rect 5411 28480 7232 28508
rect 5411 28477 5423 28480
rect 5365 28471 5423 28477
rect 7226 28468 7232 28480
rect 7284 28468 7290 28520
rect 88186 28449 88192 28452
rect 88169 28443 88192 28449
rect 88169 28409 88181 28443
rect 88169 28403 88192 28409
rect 88186 28400 88192 28403
rect 88244 28400 88250 28452
rect 4876 28314 7912 28336
rect 4876 28262 5954 28314
rect 6006 28262 6018 28314
rect 6070 28262 6082 28314
rect 6134 28262 6146 28314
rect 6198 28262 6210 28314
rect 6262 28262 7912 28314
rect 4876 28240 7912 28262
rect 85284 28314 88596 28336
rect 85284 28262 86546 28314
rect 86598 28262 86610 28314
rect 86662 28262 86674 28314
rect 86726 28262 86738 28314
rect 86790 28262 86802 28314
rect 86854 28262 88596 28314
rect 85284 28240 88596 28262
rect 5110 28060 5116 28112
rect 5168 28100 5174 28112
rect 5481 28103 5539 28109
rect 5481 28100 5493 28103
rect 5168 28072 5493 28100
rect 5168 28060 5174 28072
rect 5481 28069 5493 28072
rect 5527 28069 5539 28103
rect 5481 28063 5539 28069
rect 5128 27998 5156 28060
rect 5205 28001 5263 28007
rect 5205 27998 5217 28001
rect 5128 27970 5217 27998
rect 5205 27967 5217 27970
rect 5251 27967 5263 28001
rect 87957 28001 88015 28007
rect 87957 27998 87969 28001
rect 5205 27961 5263 27967
rect 85242 27924 85248 27976
rect 85300 27964 85306 27976
rect 87652 27970 87969 27998
rect 87652 27964 87680 27970
rect 85300 27936 87680 27964
rect 87957 27967 87969 27970
rect 88003 27967 88015 28001
rect 87957 27961 88015 27967
rect 85300 27924 85306 27936
rect 5386 27905 5392 27908
rect 5365 27899 5392 27905
rect 5365 27865 5377 27899
rect 5365 27859 5392 27865
rect 5386 27856 5392 27859
rect 5444 27856 5450 27908
rect 88169 27899 88227 27905
rect 88169 27865 88181 27899
rect 88215 27896 88227 27899
rect 88922 27896 88928 27908
rect 88215 27868 88928 27896
rect 88215 27865 88227 27868
rect 88169 27859 88227 27865
rect 88922 27856 88928 27868
rect 88980 27856 88986 27908
rect 4876 27770 7912 27792
rect 4876 27718 6690 27770
rect 6742 27718 6754 27770
rect 6806 27718 6818 27770
rect 6870 27718 6882 27770
rect 6934 27718 6946 27770
rect 6998 27718 7912 27770
rect 4876 27696 7912 27718
rect 85284 27770 88596 27792
rect 85284 27718 87282 27770
rect 87334 27718 87346 27770
rect 87398 27718 87410 27770
rect 87462 27718 87474 27770
rect 87526 27718 87538 27770
rect 87590 27718 88596 27770
rect 85284 27696 88596 27718
rect 4876 27226 7912 27248
rect 4876 27174 5954 27226
rect 6006 27174 6018 27226
rect 6070 27174 6082 27226
rect 6134 27174 6146 27226
rect 6198 27174 6210 27226
rect 6262 27174 7912 27226
rect 4876 27152 7912 27174
rect 85284 27226 88596 27248
rect 85284 27174 86546 27226
rect 86598 27174 86610 27226
rect 86662 27174 86674 27226
rect 86726 27174 86738 27226
rect 86790 27174 86802 27226
rect 86854 27174 88596 27226
rect 85284 27152 88596 27174
rect 4876 26682 7912 26704
rect 4876 26630 6690 26682
rect 6742 26630 6754 26682
rect 6806 26630 6818 26682
rect 6870 26630 6882 26682
rect 6934 26630 6946 26682
rect 6998 26630 7912 26682
rect 4876 26608 7912 26630
rect 85284 26682 88596 26704
rect 85284 26630 87282 26682
rect 87334 26630 87346 26682
rect 87398 26630 87410 26682
rect 87462 26630 87474 26682
rect 87526 26630 87538 26682
rect 87590 26630 88596 26682
rect 85284 26608 88596 26630
rect 5159 26437 5217 26443
rect 2902 26360 2908 26412
rect 2960 26400 2966 26412
rect 5159 26403 5171 26437
rect 5205 26403 5217 26437
rect 5159 26400 5217 26403
rect 5481 26403 5539 26409
rect 5481 26400 5493 26403
rect 2960 26372 5493 26400
rect 2960 26360 2966 26372
rect 5481 26369 5493 26372
rect 5527 26369 5539 26403
rect 87726 26394 87732 26446
rect 87784 26434 87790 26446
rect 87957 26437 88015 26443
rect 87957 26434 87969 26437
rect 87784 26406 87969 26434
rect 87784 26394 87790 26406
rect 87957 26403 87969 26406
rect 88003 26403 88015 26437
rect 87957 26397 88015 26403
rect 5481 26363 5539 26369
rect 5365 26335 5423 26341
rect 5365 26301 5377 26335
rect 5411 26332 5423 26335
rect 7134 26332 7140 26344
rect 5411 26304 7140 26332
rect 5411 26301 5423 26304
rect 5365 26295 5423 26301
rect 7134 26292 7140 26304
rect 7192 26292 7198 26344
rect 88186 26273 88192 26276
rect 88169 26267 88192 26273
rect 88169 26233 88181 26267
rect 88169 26227 88192 26233
rect 88186 26224 88192 26227
rect 88244 26224 88250 26276
rect 4876 26138 7912 26160
rect 4876 26086 5954 26138
rect 6006 26086 6018 26138
rect 6070 26086 6082 26138
rect 6134 26086 6146 26138
rect 6198 26086 6210 26138
rect 6262 26086 7912 26138
rect 4876 26064 7912 26086
rect 85284 26138 88596 26160
rect 85284 26086 86546 26138
rect 86598 26086 86610 26138
rect 86662 26086 86674 26138
rect 86726 26086 86738 26138
rect 86790 26086 86802 26138
rect 86854 26086 88596 26138
rect 85284 26064 88596 26086
rect 4876 25594 7912 25616
rect 4876 25542 6690 25594
rect 6742 25542 6754 25594
rect 6806 25542 6818 25594
rect 6870 25542 6882 25594
rect 6934 25542 6946 25594
rect 6998 25542 7912 25594
rect 4876 25520 7912 25542
rect 85284 25594 88596 25616
rect 85284 25542 87282 25594
rect 87334 25542 87346 25594
rect 87398 25542 87410 25594
rect 87462 25542 87474 25594
rect 87526 25542 87538 25594
rect 87590 25542 88596 25594
rect 85284 25520 88596 25542
rect 4926 25306 4932 25358
rect 4984 25346 4990 25358
rect 5159 25349 5217 25355
rect 5159 25346 5171 25349
rect 4984 25318 5171 25346
rect 4984 25306 4990 25318
rect 5159 25315 5171 25318
rect 5205 25346 5217 25349
rect 5205 25321 5524 25346
rect 5205 25318 5539 25321
rect 5205 25315 5217 25318
rect 5159 25309 5217 25315
rect 5481 25315 5539 25318
rect 5481 25281 5493 25315
rect 5527 25281 5539 25315
rect 87726 25306 87732 25358
rect 87784 25346 87790 25358
rect 87957 25349 88015 25355
rect 87957 25346 87969 25349
rect 87784 25318 87969 25346
rect 87784 25306 87790 25318
rect 87957 25315 87969 25318
rect 88003 25315 88015 25349
rect 87957 25309 88015 25315
rect 5481 25275 5539 25281
rect 5364 25247 5422 25253
rect 5364 25213 5376 25247
rect 5410 25244 5422 25247
rect 7134 25244 7140 25256
rect 5410 25216 7140 25244
rect 5410 25213 5422 25216
rect 5364 25207 5422 25213
rect 7134 25204 7140 25216
rect 7192 25204 7198 25256
rect 88169 25179 88227 25185
rect 88169 25145 88181 25179
rect 88215 25176 88227 25179
rect 88554 25176 88560 25188
rect 88215 25148 88560 25176
rect 88215 25145 88227 25148
rect 88169 25139 88227 25145
rect 88554 25136 88560 25148
rect 88612 25136 88618 25188
rect 4876 25050 7912 25072
rect 4876 24998 5954 25050
rect 6006 24998 6018 25050
rect 6070 24998 6082 25050
rect 6134 24998 6146 25050
rect 6198 24998 6210 25050
rect 6262 24998 7912 25050
rect 4876 24976 7912 24998
rect 85284 25050 88596 25072
rect 85284 24998 86546 25050
rect 86598 24998 86610 25050
rect 86662 24998 86674 25050
rect 86726 24998 86738 25050
rect 86790 24998 86802 25050
rect 86854 24998 88596 25050
rect 85284 24976 88596 24998
rect 4876 24506 7912 24528
rect 4876 24454 6690 24506
rect 6742 24454 6754 24506
rect 6806 24454 6818 24506
rect 6870 24454 6882 24506
rect 6934 24454 6946 24506
rect 6998 24454 7912 24506
rect 4876 24432 7912 24454
rect 85284 24506 88596 24528
rect 85284 24454 87282 24506
rect 87334 24454 87346 24506
rect 87398 24454 87410 24506
rect 87462 24454 87474 24506
rect 87526 24454 87538 24506
rect 87590 24454 88596 24506
rect 85284 24432 88596 24454
rect 5159 24261 5217 24267
rect 2902 24184 2908 24236
rect 2960 24224 2966 24236
rect 5159 24227 5171 24261
rect 5205 24227 5217 24261
rect 5159 24224 5217 24227
rect 5481 24227 5539 24233
rect 5481 24224 5493 24227
rect 2960 24196 5493 24224
rect 2960 24184 2966 24196
rect 5481 24193 5493 24196
rect 5527 24193 5539 24227
rect 87726 24218 87732 24270
rect 87784 24258 87790 24270
rect 87957 24261 88015 24267
rect 87957 24258 87969 24261
rect 87784 24230 87969 24258
rect 87784 24218 87790 24230
rect 87957 24227 87969 24230
rect 88003 24227 88015 24261
rect 87957 24221 88015 24227
rect 5481 24187 5539 24193
rect 5364 24159 5422 24165
rect 5364 24125 5376 24159
rect 5410 24156 5422 24159
rect 7134 24156 7140 24168
rect 5410 24128 7140 24156
rect 5410 24125 5422 24128
rect 5364 24119 5422 24125
rect 7134 24116 7140 24128
rect 7192 24116 7198 24168
rect 88169 24091 88227 24097
rect 88169 24057 88181 24091
rect 88215 24088 88227 24091
rect 88278 24088 88284 24100
rect 88215 24060 88284 24088
rect 88215 24057 88227 24060
rect 88169 24051 88227 24057
rect 88278 24048 88284 24060
rect 88336 24048 88342 24100
rect 4876 23962 7912 23984
rect 4876 23910 5954 23962
rect 6006 23910 6018 23962
rect 6070 23910 6082 23962
rect 6134 23910 6146 23962
rect 6198 23910 6210 23962
rect 6262 23910 7912 23962
rect 4876 23888 7912 23910
rect 85284 23962 88596 23984
rect 85284 23910 86546 23962
rect 86598 23910 86610 23962
rect 86662 23910 86674 23962
rect 86726 23910 86738 23962
rect 86790 23910 86802 23962
rect 86854 23910 88596 23962
rect 85284 23888 88596 23910
rect 4876 23418 7912 23440
rect 4876 23366 6690 23418
rect 6742 23366 6754 23418
rect 6806 23366 6818 23418
rect 6870 23366 6882 23418
rect 6934 23366 6946 23418
rect 6998 23366 7912 23418
rect 4876 23344 7912 23366
rect 85284 23418 88596 23440
rect 85284 23366 87282 23418
rect 87334 23366 87346 23418
rect 87398 23366 87410 23418
rect 87462 23366 87474 23418
rect 87526 23366 87538 23418
rect 87590 23366 88596 23418
rect 85284 23344 88596 23366
rect 5159 23173 5217 23179
rect 2902 23096 2908 23148
rect 2960 23136 2966 23148
rect 5159 23139 5171 23173
rect 5205 23139 5217 23173
rect 87957 23173 88015 23179
rect 5159 23136 5217 23139
rect 5481 23139 5539 23145
rect 5481 23136 5493 23139
rect 2960 23108 5493 23136
rect 2960 23096 2966 23108
rect 5481 23105 5493 23108
rect 5527 23105 5539 23139
rect 5481 23099 5539 23105
rect 86346 23096 86352 23148
rect 86404 23136 86410 23148
rect 87957 23139 87969 23173
rect 88003 23139 88015 23173
rect 87957 23136 88015 23139
rect 86404 23133 88015 23136
rect 86404 23108 88000 23133
rect 86404 23096 86410 23108
rect 5365 23071 5423 23077
rect 5365 23037 5377 23071
rect 5411 23068 5423 23071
rect 7134 23068 7140 23080
rect 5411 23040 7140 23068
rect 5411 23037 5423 23040
rect 5365 23031 5423 23037
rect 7134 23028 7140 23040
rect 7192 23028 7198 23080
rect 88169 23003 88227 23009
rect 88169 22969 88181 23003
rect 88215 23000 88227 23003
rect 88278 23000 88284 23012
rect 88215 22972 88284 23000
rect 88215 22969 88227 22972
rect 88169 22963 88227 22969
rect 88278 22960 88284 22972
rect 88336 22960 88342 23012
rect 4876 22874 7912 22896
rect 4876 22822 5954 22874
rect 6006 22822 6018 22874
rect 6070 22822 6082 22874
rect 6134 22822 6146 22874
rect 6198 22822 6210 22874
rect 6262 22822 7912 22874
rect 4876 22800 7912 22822
rect 85284 22874 88596 22896
rect 85284 22822 86546 22874
rect 86598 22822 86610 22874
rect 86662 22822 86674 22874
rect 86726 22822 86738 22874
rect 86790 22822 86802 22874
rect 86854 22822 88596 22874
rect 85284 22800 88596 22822
rect 5481 22595 5539 22601
rect 5481 22592 5493 22595
rect 4926 22518 4932 22570
rect 4984 22558 4990 22570
rect 5174 22567 5493 22592
rect 5159 22564 5493 22567
rect 5159 22561 5217 22564
rect 5159 22558 5171 22561
rect 4984 22530 5171 22558
rect 4984 22518 4990 22530
rect 5159 22527 5171 22530
rect 5205 22527 5217 22561
rect 5481 22561 5493 22564
rect 5527 22561 5539 22595
rect 5481 22555 5539 22561
rect 87957 22561 88015 22567
rect 5159 22521 5217 22527
rect 5364 22527 5422 22533
rect 5364 22493 5376 22527
rect 5410 22524 5422 22527
rect 9158 22524 9164 22536
rect 5410 22496 9164 22524
rect 5410 22493 5422 22496
rect 5364 22487 5422 22493
rect 9158 22484 9164 22496
rect 9216 22484 9222 22536
rect 84414 22484 84420 22536
rect 84472 22524 84478 22536
rect 87957 22527 87969 22561
rect 88003 22527 88015 22561
rect 87957 22524 88015 22527
rect 84472 22521 88015 22524
rect 84472 22496 88000 22521
rect 84472 22484 84478 22496
rect 88169 22459 88227 22465
rect 88169 22425 88181 22459
rect 88215 22456 88227 22459
rect 88554 22456 88560 22468
rect 88215 22428 88560 22456
rect 88215 22425 88227 22428
rect 88169 22419 88227 22425
rect 88554 22416 88560 22428
rect 88612 22416 88618 22468
rect 4876 22330 7912 22352
rect 4876 22278 6690 22330
rect 6742 22278 6754 22330
rect 6806 22278 6818 22330
rect 6870 22278 6882 22330
rect 6934 22278 6946 22330
rect 6998 22278 7912 22330
rect 4876 22256 7912 22278
rect 85284 22330 88596 22352
rect 85284 22278 87282 22330
rect 87334 22278 87346 22330
rect 87398 22278 87410 22330
rect 87462 22278 87474 22330
rect 87526 22278 87538 22330
rect 87590 22278 88596 22330
rect 85284 22256 88596 22278
rect 4876 21786 7912 21808
rect 4876 21734 5954 21786
rect 6006 21734 6018 21786
rect 6070 21734 6082 21786
rect 6134 21734 6146 21786
rect 6198 21734 6210 21786
rect 6262 21734 7912 21786
rect 4876 21712 7912 21734
rect 85284 21786 88596 21808
rect 85284 21734 86546 21786
rect 86598 21734 86610 21786
rect 86662 21734 86674 21786
rect 86726 21734 86738 21786
rect 86790 21734 86802 21786
rect 86854 21734 88596 21786
rect 85284 21712 88596 21734
rect 4876 21242 7912 21264
rect 4876 21190 6690 21242
rect 6742 21190 6754 21242
rect 6806 21190 6818 21242
rect 6870 21190 6882 21242
rect 6934 21190 6946 21242
rect 6998 21190 7912 21242
rect 4876 21168 7912 21190
rect 85284 21242 88596 21264
rect 85284 21190 87282 21242
rect 87334 21190 87346 21242
rect 87398 21190 87410 21242
rect 87462 21190 87474 21242
rect 87526 21190 87538 21242
rect 87590 21190 88596 21242
rect 85284 21168 88596 21190
rect 5365 21099 5423 21105
rect 5365 21065 5377 21099
rect 5411 21096 5423 21099
rect 9250 21096 9256 21108
rect 5411 21068 9256 21096
rect 5411 21065 5423 21068
rect 5365 21059 5423 21065
rect 9250 21056 9256 21068
rect 9308 21056 9314 21108
rect 5202 20954 5208 21006
rect 5260 20960 5266 21006
rect 87957 20997 88015 21003
rect 5481 20963 5539 20969
rect 5481 20960 5493 20963
rect 5260 20954 5493 20960
rect 5220 20932 5493 20954
rect 5481 20929 5493 20932
rect 5527 20929 5539 20963
rect 5481 20923 5539 20929
rect 84414 20920 84420 20972
rect 84472 20960 84478 20972
rect 87957 20963 87969 20997
rect 88003 20963 88015 20997
rect 87957 20960 88015 20963
rect 84472 20957 88015 20960
rect 88169 20963 88227 20969
rect 84472 20932 88000 20957
rect 84472 20920 84478 20932
rect 88169 20929 88181 20963
rect 88215 20960 88227 20963
rect 88554 20960 88560 20972
rect 88215 20932 88560 20960
rect 88215 20929 88227 20932
rect 88169 20923 88227 20929
rect 88554 20920 88560 20932
rect 88612 20920 88618 20972
rect 4876 20698 7912 20720
rect 4876 20646 5954 20698
rect 6006 20646 6018 20698
rect 6070 20646 6082 20698
rect 6134 20646 6146 20698
rect 6198 20646 6210 20698
rect 6262 20646 7912 20698
rect 4876 20624 7912 20646
rect 85284 20698 88596 20720
rect 85284 20646 86546 20698
rect 86598 20646 86610 20698
rect 86662 20646 86674 20698
rect 86726 20646 86738 20698
rect 86790 20646 86802 20698
rect 86854 20646 88596 20698
rect 85284 20624 88596 20646
rect 4876 20154 7912 20176
rect 4876 20102 6690 20154
rect 6742 20102 6754 20154
rect 6806 20102 6818 20154
rect 6870 20102 6882 20154
rect 6934 20102 6946 20154
rect 6998 20102 7912 20154
rect 4876 20080 7912 20102
rect 85284 20154 88596 20176
rect 85284 20102 87282 20154
rect 87334 20102 87346 20154
rect 87398 20102 87410 20154
rect 87462 20102 87474 20154
rect 87526 20102 87538 20154
rect 87590 20102 88596 20154
rect 85284 20080 88596 20102
rect 4926 19866 4932 19918
rect 4984 19906 4990 19918
rect 5159 19909 5217 19915
rect 5159 19906 5171 19909
rect 4984 19878 5171 19906
rect 4984 19866 4990 19878
rect 5159 19875 5171 19878
rect 5205 19906 5217 19909
rect 5205 19881 5524 19906
rect 5205 19878 5539 19881
rect 5205 19875 5217 19878
rect 5159 19869 5217 19875
rect 5481 19875 5539 19878
rect 5481 19841 5493 19875
rect 5527 19841 5539 19875
rect 87726 19866 87732 19918
rect 87784 19906 87790 19918
rect 87957 19909 88015 19915
rect 87957 19906 87969 19909
rect 87784 19878 87969 19906
rect 87784 19866 87790 19878
rect 87957 19875 87969 19878
rect 88003 19875 88015 19909
rect 87957 19869 88015 19875
rect 5481 19835 5539 19841
rect 5365 19807 5423 19813
rect 5365 19773 5377 19807
rect 5411 19804 5423 19807
rect 7134 19804 7140 19816
rect 5411 19776 7140 19804
rect 5411 19773 5423 19776
rect 5365 19767 5423 19773
rect 7134 19764 7140 19776
rect 7192 19764 7198 19816
rect 88169 19739 88227 19745
rect 88169 19705 88181 19739
rect 88215 19736 88227 19739
rect 88554 19736 88560 19748
rect 88215 19708 88560 19736
rect 88215 19705 88227 19708
rect 88169 19699 88227 19705
rect 88554 19696 88560 19708
rect 88612 19696 88618 19748
rect 4876 19610 7912 19632
rect 4876 19558 5954 19610
rect 6006 19558 6018 19610
rect 6070 19558 6082 19610
rect 6134 19558 6146 19610
rect 6198 19558 6210 19610
rect 6262 19558 7912 19610
rect 4876 19536 7912 19558
rect 85284 19610 88596 19632
rect 85284 19558 86546 19610
rect 86598 19558 86610 19610
rect 86662 19558 86674 19610
rect 86726 19558 86738 19610
rect 86790 19558 86802 19610
rect 86854 19558 88596 19610
rect 85284 19536 88596 19558
rect 4876 19066 7912 19088
rect 4876 19014 6690 19066
rect 6742 19014 6754 19066
rect 6806 19014 6818 19066
rect 6870 19014 6882 19066
rect 6934 19014 6946 19066
rect 6998 19014 7912 19066
rect 4876 18992 7912 19014
rect 85284 19066 88596 19088
rect 85284 19014 87282 19066
rect 87334 19014 87346 19066
rect 87398 19014 87410 19066
rect 87462 19014 87474 19066
rect 87526 19014 87538 19066
rect 87590 19014 88596 19066
rect 85284 18992 88596 19014
rect 5159 18821 5217 18827
rect 2902 18744 2908 18796
rect 2960 18784 2966 18796
rect 5159 18787 5171 18821
rect 5205 18787 5217 18821
rect 5159 18784 5217 18787
rect 5481 18787 5539 18793
rect 5481 18784 5493 18787
rect 2960 18756 5493 18784
rect 2960 18744 2966 18756
rect 5481 18753 5493 18756
rect 5527 18753 5539 18787
rect 87726 18778 87732 18830
rect 87784 18818 87790 18830
rect 87957 18821 88015 18827
rect 87957 18818 87969 18821
rect 87784 18790 87969 18818
rect 87784 18778 87790 18790
rect 87957 18787 87969 18790
rect 88003 18787 88015 18821
rect 87957 18781 88015 18787
rect 5481 18747 5539 18753
rect 5365 18719 5423 18725
rect 5365 18685 5377 18719
rect 5411 18716 5423 18719
rect 7134 18716 7140 18728
rect 5411 18688 7140 18716
rect 5411 18685 5423 18688
rect 5365 18679 5423 18685
rect 7134 18676 7140 18688
rect 7192 18676 7198 18728
rect 88169 18651 88227 18657
rect 88169 18617 88181 18651
rect 88215 18648 88227 18651
rect 88278 18648 88284 18660
rect 88215 18620 88284 18648
rect 88215 18617 88227 18620
rect 88169 18611 88227 18617
rect 88278 18608 88284 18620
rect 88336 18608 88342 18660
rect 4876 18522 7912 18544
rect 4876 18470 5954 18522
rect 6006 18470 6018 18522
rect 6070 18470 6082 18522
rect 6134 18470 6146 18522
rect 6198 18470 6210 18522
rect 6262 18470 7912 18522
rect 4876 18448 7912 18470
rect 85284 18522 88596 18544
rect 85284 18470 86546 18522
rect 86598 18470 86610 18522
rect 86662 18470 86674 18522
rect 86726 18470 86738 18522
rect 86790 18470 86802 18522
rect 86854 18470 88596 18522
rect 85284 18448 88596 18470
rect 4876 17978 7912 18000
rect 4876 17926 6690 17978
rect 6742 17926 6754 17978
rect 6806 17926 6818 17978
rect 6870 17926 6882 17978
rect 6934 17926 6946 17978
rect 6998 17926 7912 17978
rect 4876 17904 7912 17926
rect 85284 17978 88596 18000
rect 85284 17926 87282 17978
rect 87334 17926 87346 17978
rect 87398 17926 87410 17978
rect 87462 17926 87474 17978
rect 87526 17926 87538 17978
rect 87590 17926 88596 17978
rect 85284 17904 88596 17926
rect 5159 17733 5217 17739
rect 5159 17730 5171 17733
rect 2902 17656 2908 17708
rect 2960 17696 2966 17708
rect 4852 17702 5171 17730
rect 4852 17696 4880 17702
rect 2960 17668 4880 17696
rect 5159 17699 5171 17702
rect 5205 17730 5217 17733
rect 87957 17733 88015 17739
rect 87957 17730 87969 17733
rect 5205 17705 5524 17730
rect 5205 17702 5539 17705
rect 5205 17699 5217 17702
rect 5159 17693 5217 17699
rect 5481 17699 5539 17702
rect 2960 17656 2966 17668
rect 5481 17665 5493 17699
rect 5527 17665 5539 17699
rect 5481 17659 5539 17665
rect 86346 17656 86352 17708
rect 86404 17696 86410 17708
rect 87652 17702 87969 17730
rect 87652 17696 87680 17702
rect 86404 17668 87680 17696
rect 87957 17699 87969 17702
rect 88003 17699 88015 17733
rect 87957 17693 88015 17699
rect 86404 17656 86410 17668
rect 5365 17631 5423 17637
rect 5365 17597 5377 17631
rect 5411 17628 5423 17631
rect 7226 17628 7232 17640
rect 5411 17600 7232 17628
rect 5411 17597 5423 17600
rect 5365 17591 5423 17597
rect 7226 17588 7232 17600
rect 7284 17588 7290 17640
rect 88186 17569 88192 17572
rect 88169 17563 88192 17569
rect 88169 17529 88181 17563
rect 88169 17523 88192 17529
rect 88186 17520 88192 17523
rect 88244 17520 88250 17572
rect 4876 17434 7912 17456
rect 4876 17382 5954 17434
rect 6006 17382 6018 17434
rect 6070 17382 6082 17434
rect 6134 17382 6146 17434
rect 6198 17382 6210 17434
rect 6262 17382 7912 17434
rect 4876 17360 7912 17382
rect 85284 17434 88596 17456
rect 85284 17382 86546 17434
rect 86598 17382 86610 17434
rect 86662 17382 86674 17434
rect 86726 17382 86738 17434
rect 86790 17382 86802 17434
rect 86854 17382 88596 17434
rect 85284 17360 88596 17382
rect 5202 17078 5208 17130
rect 5260 17084 5266 17130
rect 5481 17087 5539 17093
rect 5481 17084 5493 17087
rect 5260 17078 5493 17084
rect 5220 17056 5493 17078
rect 5481 17053 5493 17056
rect 5527 17053 5539 17087
rect 88002 17078 88008 17130
rect 88060 17078 88066 17130
rect 5481 17047 5539 17053
rect 5386 17025 5392 17028
rect 5365 17019 5392 17025
rect 5365 16985 5377 17019
rect 5365 16979 5392 16985
rect 5386 16976 5392 16979
rect 5444 16976 5450 17028
rect 88169 17019 88227 17025
rect 88169 16985 88181 17019
rect 88215 17016 88227 17019
rect 88554 17016 88560 17028
rect 88215 16988 88560 17016
rect 88215 16985 88227 16988
rect 88169 16979 88227 16985
rect 88554 16976 88560 16988
rect 88612 16976 88618 17028
rect 4876 16890 7912 16912
rect 4876 16838 6690 16890
rect 6742 16838 6754 16890
rect 6806 16838 6818 16890
rect 6870 16838 6882 16890
rect 6934 16838 6946 16890
rect 6998 16838 7912 16890
rect 4876 16816 7912 16838
rect 85284 16890 88596 16912
rect 85284 16838 87282 16890
rect 87334 16838 87346 16890
rect 87398 16838 87410 16890
rect 87462 16838 87474 16890
rect 87526 16838 87538 16890
rect 87590 16838 88596 16890
rect 85284 16816 88596 16838
rect 4876 16346 7912 16368
rect 4876 16294 5954 16346
rect 6006 16294 6018 16346
rect 6070 16294 6082 16346
rect 6134 16294 6146 16346
rect 6198 16294 6210 16346
rect 6262 16294 7912 16346
rect 4876 16272 7912 16294
rect 85284 16346 88596 16368
rect 85284 16294 86546 16346
rect 86598 16294 86610 16346
rect 86662 16294 86674 16346
rect 86726 16294 86738 16346
rect 86790 16294 86802 16346
rect 86854 16294 88596 16346
rect 85284 16272 88596 16294
rect 4876 15802 7912 15824
rect 4876 15750 6690 15802
rect 6742 15750 6754 15802
rect 6806 15750 6818 15802
rect 6870 15750 6882 15802
rect 6934 15750 6946 15802
rect 6998 15750 7912 15802
rect 4876 15728 7912 15750
rect 85284 15802 88596 15824
rect 85284 15750 87282 15802
rect 87334 15750 87346 15802
rect 87398 15750 87410 15802
rect 87462 15750 87474 15802
rect 87526 15750 87538 15802
rect 87590 15750 88596 15802
rect 85284 15728 88596 15750
rect 5202 15514 5208 15566
rect 5260 15520 5266 15566
rect 87957 15557 88015 15563
rect 87957 15554 87969 15557
rect 5481 15523 5539 15529
rect 5481 15520 5493 15523
rect 5260 15514 5493 15520
rect 5220 15492 5493 15514
rect 5481 15489 5493 15492
rect 5527 15489 5539 15523
rect 5481 15483 5539 15489
rect 84414 15480 84420 15532
rect 84472 15520 84478 15532
rect 87836 15526 87969 15554
rect 87836 15520 87864 15526
rect 84472 15492 87864 15520
rect 87957 15523 87969 15526
rect 88003 15523 88015 15557
rect 87957 15517 88015 15523
rect 84472 15480 84478 15492
rect 5365 15455 5423 15461
rect 5365 15421 5377 15455
rect 5411 15452 5423 15455
rect 5662 15452 5668 15464
rect 5411 15424 5668 15452
rect 5411 15421 5423 15424
rect 5365 15415 5423 15421
rect 5662 15412 5668 15424
rect 5720 15412 5726 15464
rect 88169 15455 88227 15461
rect 88169 15421 88181 15455
rect 88215 15452 88227 15455
rect 88554 15452 88560 15464
rect 88215 15424 88560 15452
rect 88215 15421 88227 15424
rect 88169 15415 88227 15421
rect 88554 15412 88560 15424
rect 88612 15412 88618 15464
rect 4876 15258 7912 15280
rect 4876 15206 5954 15258
rect 6006 15206 6018 15258
rect 6070 15206 6082 15258
rect 6134 15206 6146 15258
rect 6198 15206 6210 15258
rect 6262 15206 7912 15258
rect 4876 15184 7912 15206
rect 85284 15258 88596 15280
rect 85284 15206 86546 15258
rect 86598 15206 86610 15258
rect 86662 15206 86674 15258
rect 86726 15206 86738 15258
rect 86790 15206 86802 15258
rect 86854 15206 88596 15258
rect 85284 15184 88596 15206
rect 88189 15047 88247 15053
rect 88189 15044 88201 15047
rect 87468 15016 88201 15044
rect 85426 14936 85432 14988
rect 85484 14976 85490 14988
rect 85610 14976 85616 14988
rect 85484 14948 85616 14976
rect 85484 14936 85490 14948
rect 85610 14936 85616 14948
rect 85668 14976 85674 14988
rect 87468 14985 87496 15016
rect 88189 15013 88201 15016
rect 88235 15013 88247 15047
rect 88189 15007 88247 15013
rect 87453 14979 87511 14985
rect 87453 14976 87465 14979
rect 85668 14948 87465 14976
rect 85668 14936 85674 14948
rect 87453 14945 87465 14948
rect 87499 14945 87511 14979
rect 87453 14939 87511 14945
rect 87796 14945 87854 14951
rect 87796 14911 87808 14945
rect 87842 14942 87854 14945
rect 87842 14914 88048 14942
rect 87842 14911 87854 14914
rect 87796 14905 87854 14911
rect 88020 14852 88048 14914
rect 88002 14800 88008 14852
rect 88060 14800 88066 14852
rect 4876 14714 7912 14736
rect 4876 14662 6690 14714
rect 6742 14662 6754 14714
rect 6806 14662 6818 14714
rect 6870 14662 6882 14714
rect 6934 14662 6946 14714
rect 6998 14662 7912 14714
rect 4876 14640 7912 14662
rect 85284 14714 88596 14736
rect 85284 14662 87282 14714
rect 87334 14662 87346 14714
rect 87398 14662 87410 14714
rect 87462 14662 87474 14714
rect 87526 14662 87538 14714
rect 87590 14662 88596 14714
rect 85284 14640 88596 14662
rect 83678 14256 83684 14308
rect 83736 14296 83742 14308
rect 85610 14296 85616 14308
rect 83736 14268 85616 14296
rect 83736 14256 83742 14268
rect 85610 14256 85616 14268
rect 85668 14256 85674 14308
rect 4876 14170 7912 14192
rect 4876 14118 5954 14170
rect 6006 14118 6018 14170
rect 6070 14118 6082 14170
rect 6134 14118 6146 14170
rect 6198 14118 6210 14170
rect 6262 14118 7912 14170
rect 4876 14096 7912 14118
rect 85284 14170 88596 14192
rect 85284 14118 86546 14170
rect 86598 14118 86610 14170
rect 86662 14118 86674 14170
rect 86726 14118 86738 14170
rect 86790 14118 86802 14170
rect 86854 14118 88596 14170
rect 85284 14096 88596 14118
rect 4876 13626 7912 13648
rect 4876 13574 6690 13626
rect 6742 13574 6754 13626
rect 6806 13574 6818 13626
rect 6870 13574 6882 13626
rect 6934 13574 6946 13626
rect 6998 13574 7912 13626
rect 4876 13552 7912 13574
rect 85284 13626 88596 13648
rect 85284 13574 87282 13626
rect 87334 13574 87346 13626
rect 87398 13574 87410 13626
rect 87462 13574 87474 13626
rect 87526 13574 87538 13626
rect 87590 13574 88596 13626
rect 85284 13552 88596 13574
rect 83494 13440 83500 13492
rect 83552 13480 83558 13492
rect 85518 13480 85524 13492
rect 83552 13452 85524 13480
rect 83552 13440 83558 13452
rect 85518 13440 85524 13452
rect 85576 13480 85582 13492
rect 85613 13483 85671 13489
rect 85613 13480 85625 13483
rect 85576 13452 85625 13480
rect 85576 13440 85582 13452
rect 85613 13449 85625 13452
rect 85659 13480 85671 13483
rect 85659 13452 85794 13480
rect 85659 13449 85671 13452
rect 85613 13443 85671 13449
rect 85766 13344 85794 13452
rect 87637 13415 87695 13421
rect 87637 13381 87649 13415
rect 87683 13412 87695 13415
rect 87683 13384 88140 13412
rect 87683 13381 87695 13384
rect 87637 13375 87695 13381
rect 88112 13378 88140 13384
rect 88186 13378 88192 13390
rect 88244 13387 88250 13390
rect 88244 13381 88272 13387
rect 87910 13344 87916 13356
rect 85766 13316 87916 13344
rect 87910 13304 87916 13316
rect 87968 13304 87974 13356
rect 88112 13350 88192 13378
rect 88186 13338 88192 13350
rect 88260 13347 88272 13381
rect 88244 13341 88272 13347
rect 88244 13338 88250 13341
rect 4876 13082 7912 13104
rect 4876 13030 5954 13082
rect 6006 13030 6018 13082
rect 6070 13030 6082 13082
rect 6134 13030 6146 13082
rect 6198 13030 6210 13082
rect 6262 13030 7912 13082
rect 4876 13008 7912 13030
rect 85284 13082 88596 13104
rect 85284 13030 86546 13082
rect 86598 13030 86610 13082
rect 86662 13030 86674 13082
rect 86726 13030 86738 13082
rect 86790 13030 86802 13082
rect 86854 13030 88596 13082
rect 85284 13008 88596 13030
rect 87910 12896 87916 12948
rect 87968 12936 87974 12948
rect 88189 12939 88247 12945
rect 88189 12936 88201 12939
rect 87968 12908 88201 12936
rect 87968 12896 87974 12908
rect 88189 12905 88201 12908
rect 88235 12905 88247 12939
rect 88189 12899 88247 12905
rect 87796 12769 87854 12775
rect 87174 12692 87180 12744
rect 87232 12732 87238 12744
rect 87453 12735 87511 12741
rect 87453 12732 87465 12735
rect 87232 12704 87465 12732
rect 87232 12692 87238 12704
rect 87453 12701 87465 12704
rect 87499 12701 87511 12735
rect 87796 12735 87808 12769
rect 87842 12766 87854 12769
rect 87842 12741 88048 12766
rect 87842 12738 88063 12741
rect 87842 12735 87854 12738
rect 87796 12729 87854 12735
rect 88005 12735 88063 12738
rect 87453 12695 87511 12701
rect 88005 12701 88017 12735
rect 88051 12732 88063 12735
rect 88554 12732 88560 12744
rect 88051 12704 88560 12732
rect 88051 12701 88063 12704
rect 88005 12695 88063 12701
rect 88554 12692 88560 12704
rect 88612 12692 88618 12744
rect 4876 12538 7912 12560
rect 4876 12486 6690 12538
rect 6742 12486 6754 12538
rect 6806 12486 6818 12538
rect 6870 12486 6882 12538
rect 6934 12486 6946 12538
rect 6998 12486 7912 12538
rect 4876 12464 7912 12486
rect 85284 12538 88596 12560
rect 85284 12486 87282 12538
rect 87334 12486 87346 12538
rect 87398 12486 87410 12538
rect 87462 12486 87474 12538
rect 87526 12486 87538 12538
rect 87590 12486 88596 12538
rect 85284 12464 88596 12486
rect 83494 12352 83500 12404
rect 83552 12392 83558 12404
rect 85334 12392 85340 12404
rect 83552 12364 85340 12392
rect 83552 12352 83558 12364
rect 85334 12352 85340 12364
rect 85392 12392 85398 12404
rect 85613 12395 85671 12401
rect 85613 12392 85625 12395
rect 85392 12364 85625 12392
rect 85392 12352 85398 12364
rect 85613 12361 85625 12364
rect 85659 12392 85671 12395
rect 87174 12392 87180 12404
rect 85659 12364 87180 12392
rect 85659 12361 85671 12364
rect 85613 12355 85671 12361
rect 87174 12352 87180 12364
rect 87232 12392 87238 12404
rect 88097 12395 88155 12401
rect 88097 12392 88109 12395
rect 87232 12364 88109 12392
rect 87232 12352 87238 12364
rect 88097 12361 88109 12364
rect 88143 12361 88155 12395
rect 88097 12355 88155 12361
rect 4876 11994 7912 12016
rect 4876 11942 5954 11994
rect 6006 11942 6018 11994
rect 6070 11942 6082 11994
rect 6134 11942 6146 11994
rect 6198 11942 6210 11994
rect 6262 11942 7912 11994
rect 4876 11920 7912 11942
rect 85284 11994 88596 12016
rect 85284 11942 86546 11994
rect 86598 11942 86610 11994
rect 86662 11942 86674 11994
rect 86726 11942 86738 11994
rect 86790 11942 86802 11994
rect 86854 11942 88596 11994
rect 85284 11920 88596 11942
rect 83402 11740 83408 11792
rect 83460 11780 83466 11792
rect 83678 11780 83684 11792
rect 83460 11752 83684 11780
rect 83460 11740 83466 11752
rect 83678 11740 83684 11752
rect 83736 11740 83742 11792
rect 4876 11450 7912 11472
rect 4876 11398 6690 11450
rect 6742 11398 6754 11450
rect 6806 11398 6818 11450
rect 6870 11398 6882 11450
rect 6934 11398 6946 11450
rect 6998 11398 7912 11450
rect 4876 11376 7912 11398
rect 85284 11450 88596 11472
rect 85284 11398 87282 11450
rect 87334 11398 87346 11450
rect 87398 11398 87410 11450
rect 87462 11398 87474 11450
rect 87526 11398 87538 11450
rect 87590 11398 88596 11450
rect 85284 11376 88596 11398
rect 83310 11196 83316 11248
rect 83368 11236 83374 11248
rect 85613 11239 85671 11245
rect 85613 11236 85625 11239
rect 83368 11208 85625 11236
rect 83368 11196 83374 11208
rect 85613 11205 85625 11208
rect 85659 11205 85671 11239
rect 85613 11199 85671 11205
rect 4876 10906 7912 10928
rect 4876 10854 5954 10906
rect 6006 10854 6018 10906
rect 6070 10854 6082 10906
rect 6134 10854 6146 10906
rect 6198 10854 6210 10906
rect 6262 10854 7912 10906
rect 4876 10832 7912 10854
rect 85284 10906 88596 10928
rect 85284 10854 86546 10906
rect 86598 10854 86610 10906
rect 86662 10854 86674 10906
rect 86726 10854 86738 10906
rect 86790 10854 86802 10906
rect 86854 10854 88596 10906
rect 85284 10832 88596 10854
rect 87729 10627 87787 10633
rect 87729 10593 87741 10627
rect 87775 10624 87787 10627
rect 87775 10596 88140 10624
rect 87775 10593 87787 10596
rect 87729 10587 87787 10593
rect 88112 10564 88140 10596
rect 88253 10593 88311 10599
rect 88253 10564 88265 10593
rect 88112 10559 88265 10564
rect 88299 10590 88311 10593
rect 88299 10576 88416 10590
rect 88299 10562 88376 10576
rect 88299 10559 88324 10562
rect 83972 10528 87864 10556
rect 88112 10536 88324 10559
rect 83972 10420 84000 10528
rect 87836 10488 87864 10528
rect 88370 10524 88376 10562
rect 88428 10524 88434 10576
rect 88051 10491 88109 10497
rect 88051 10488 88063 10491
rect 87836 10460 88063 10488
rect 88051 10457 88063 10460
rect 88097 10457 88109 10491
rect 88051 10451 88109 10457
rect 82500 10392 84000 10420
rect 4876 10362 7912 10384
rect 4876 10310 6690 10362
rect 6742 10310 6754 10362
rect 6806 10310 6818 10362
rect 6870 10310 6882 10362
rect 6934 10310 6946 10362
rect 6998 10310 7912 10362
rect 4876 10288 7912 10310
rect 82500 10228 82528 10392
rect 85284 10362 88596 10384
rect 85284 10310 87282 10362
rect 87334 10310 87346 10362
rect 87398 10310 87410 10362
rect 87462 10310 87474 10362
rect 87526 10310 87538 10362
rect 87590 10310 88596 10362
rect 85284 10288 88596 10310
rect 45590 10176 45596 10228
rect 45648 10216 45654 10228
rect 46050 10216 46056 10228
rect 45648 10188 46056 10216
rect 45648 10176 45654 10188
rect 46050 10176 46056 10188
rect 46108 10176 46114 10228
rect 82482 10176 82488 10228
rect 82540 10176 82546 10228
rect 88253 10117 88311 10123
rect 88253 10114 88265 10117
rect 87913 10083 87971 10089
rect 87913 10049 87925 10083
rect 87959 10080 87971 10083
rect 88112 10086 88265 10114
rect 88112 10080 88140 10086
rect 87959 10052 88140 10080
rect 88253 10083 88265 10086
rect 88299 10114 88311 10117
rect 88299 10086 88508 10114
rect 88299 10083 88311 10086
rect 88253 10077 88311 10083
rect 88480 10080 88508 10086
rect 88554 10080 88560 10092
rect 88480 10052 88560 10080
rect 87959 10049 87971 10052
rect 87913 10043 87971 10049
rect 88554 10040 88560 10052
rect 88612 10040 88618 10092
rect 81378 9972 81384 10024
rect 81436 10012 81442 10024
rect 88051 10015 88109 10021
rect 88051 10012 88063 10015
rect 81436 9984 88063 10012
rect 81436 9972 81442 9984
rect 88051 9981 88063 9984
rect 88097 9981 88109 10015
rect 88051 9975 88109 9981
rect 4876 9818 7912 9840
rect 4876 9766 5954 9818
rect 6006 9766 6018 9818
rect 6070 9766 6082 9818
rect 6134 9766 6146 9818
rect 6198 9766 6210 9818
rect 6262 9766 7912 9818
rect 4876 9744 7912 9766
rect 85284 9818 88596 9840
rect 85284 9766 86546 9818
rect 86598 9766 86610 9818
rect 86662 9766 86674 9818
rect 86726 9766 86738 9818
rect 86790 9766 86802 9818
rect 86854 9766 88596 9818
rect 85284 9744 88596 9766
rect 4876 9274 7912 9296
rect 4876 9222 6690 9274
rect 6742 9222 6754 9274
rect 6806 9222 6818 9274
rect 6870 9222 6882 9274
rect 6934 9222 6946 9274
rect 6998 9222 7912 9274
rect 4876 9200 7912 9222
rect 85284 9274 88596 9296
rect 85284 9222 87282 9274
rect 87334 9222 87346 9274
rect 87398 9222 87410 9274
rect 87462 9222 87474 9274
rect 87526 9222 87538 9274
rect 87590 9222 88596 9274
rect 85284 9200 88596 9222
rect 4876 8730 7912 8752
rect 4876 8678 5954 8730
rect 6006 8678 6018 8730
rect 6070 8678 6082 8730
rect 6134 8678 6146 8730
rect 6198 8678 6210 8730
rect 6262 8678 7912 8730
rect 4876 8656 7912 8678
rect 85284 8730 88596 8752
rect 85284 8678 86546 8730
rect 86598 8678 86610 8730
rect 86662 8678 86674 8730
rect 86726 8678 86738 8730
rect 86790 8678 86802 8730
rect 86854 8678 88596 8730
rect 85284 8656 88596 8678
rect 4876 8186 7912 8208
rect 4876 8134 6690 8186
rect 6742 8134 6754 8186
rect 6806 8134 6818 8186
rect 6870 8134 6882 8186
rect 6934 8134 6946 8186
rect 6998 8134 7912 8186
rect 4876 8112 7912 8134
rect 85284 8186 88596 8208
rect 85284 8134 87282 8186
rect 87334 8134 87346 8186
rect 87398 8134 87410 8186
rect 87462 8134 87474 8186
rect 87526 8134 87538 8186
rect 87590 8134 88596 8186
rect 85284 8112 88596 8134
rect 4876 7642 88596 7664
rect 4876 7590 5954 7642
rect 6006 7590 6018 7642
rect 6070 7590 6082 7642
rect 6134 7590 6146 7642
rect 6198 7590 6210 7642
rect 6262 7590 17722 7642
rect 17774 7590 17786 7642
rect 17838 7590 17850 7642
rect 17902 7590 17914 7642
rect 17966 7590 17978 7642
rect 18030 7590 36122 7642
rect 36174 7590 36186 7642
rect 36238 7590 36250 7642
rect 36302 7590 36314 7642
rect 36366 7590 36378 7642
rect 36430 7590 54522 7642
rect 54574 7590 54586 7642
rect 54638 7590 54650 7642
rect 54702 7590 54714 7642
rect 54766 7590 54778 7642
rect 54830 7590 72922 7642
rect 72974 7590 72986 7642
rect 73038 7590 73050 7642
rect 73102 7590 73114 7642
rect 73166 7590 73178 7642
rect 73230 7590 86546 7642
rect 86598 7590 86610 7642
rect 86662 7590 86674 7642
rect 86726 7590 86738 7642
rect 86790 7590 86802 7642
rect 86854 7590 88596 7642
rect 4876 7568 88596 7590
rect 45409 7499 45467 7505
rect 45409 7465 45421 7499
rect 45455 7496 45467 7499
rect 45682 7496 45688 7508
rect 45455 7468 45688 7496
rect 45455 7465 45467 7468
rect 45409 7459 45467 7465
rect 45682 7456 45688 7468
rect 45740 7456 45746 7508
rect 45958 7456 45964 7508
rect 46016 7456 46022 7508
rect 45590 7388 45596 7440
rect 45648 7388 45654 7440
rect 45777 7431 45835 7437
rect 45777 7397 45789 7431
rect 45823 7428 45835 7431
rect 46050 7428 46056 7440
rect 45823 7400 46056 7428
rect 45823 7397 45835 7400
rect 45777 7391 45835 7397
rect 46050 7388 46056 7400
rect 46108 7428 46114 7440
rect 46108 7400 47154 7428
rect 46108 7388 46114 7400
rect 47126 7360 47154 7400
rect 83494 7360 83500 7372
rect 47126 7332 83500 7360
rect 83494 7320 83500 7332
rect 83552 7320 83558 7372
rect 45958 7252 45964 7304
rect 46016 7292 46022 7304
rect 83402 7292 83408 7304
rect 46016 7264 83408 7292
rect 46016 7252 46022 7264
rect 83402 7252 83408 7264
rect 83460 7252 83466 7304
rect 45590 7184 45596 7236
rect 45648 7224 45654 7236
rect 83586 7224 83592 7236
rect 45648 7196 83592 7224
rect 45648 7184 45654 7196
rect 83586 7184 83592 7196
rect 83644 7184 83650 7236
rect 4876 7098 88596 7120
rect 4876 7046 6690 7098
rect 6742 7046 6754 7098
rect 6806 7046 6818 7098
rect 6870 7046 6882 7098
rect 6934 7046 6946 7098
rect 6998 7046 18382 7098
rect 18434 7046 18446 7098
rect 18498 7046 18510 7098
rect 18562 7046 18574 7098
rect 18626 7046 18638 7098
rect 18690 7046 36782 7098
rect 36834 7046 36846 7098
rect 36898 7046 36910 7098
rect 36962 7046 36974 7098
rect 37026 7046 37038 7098
rect 37090 7046 55182 7098
rect 55234 7046 55246 7098
rect 55298 7046 55310 7098
rect 55362 7046 55374 7098
rect 55426 7046 55438 7098
rect 55490 7046 73582 7098
rect 73634 7046 73646 7098
rect 73698 7046 73710 7098
rect 73762 7046 73774 7098
rect 73826 7046 73838 7098
rect 73890 7046 87282 7098
rect 87334 7046 87346 7098
rect 87398 7046 87410 7098
rect 87462 7046 87474 7098
rect 87526 7046 87538 7098
rect 87590 7046 88596 7098
rect 4876 7024 88596 7046
rect 4876 6554 88596 6576
rect 4876 6502 17722 6554
rect 17774 6502 17786 6554
rect 17838 6502 17850 6554
rect 17902 6502 17914 6554
rect 17966 6502 17978 6554
rect 18030 6502 36122 6554
rect 36174 6502 36186 6554
rect 36238 6502 36250 6554
rect 36302 6502 36314 6554
rect 36366 6502 36378 6554
rect 36430 6502 54522 6554
rect 54574 6502 54586 6554
rect 54638 6502 54650 6554
rect 54702 6502 54714 6554
rect 54766 6502 54778 6554
rect 54830 6502 72922 6554
rect 72974 6502 72986 6554
rect 73038 6502 73050 6554
rect 73102 6502 73114 6554
rect 73166 6502 73178 6554
rect 73230 6502 88596 6554
rect 4876 6480 88596 6502
rect 4876 6010 88596 6032
rect 4876 5958 18382 6010
rect 18434 5958 18446 6010
rect 18498 5958 18510 6010
rect 18562 5958 18574 6010
rect 18626 5958 18638 6010
rect 18690 5958 36782 6010
rect 36834 5958 36846 6010
rect 36898 5958 36910 6010
rect 36962 5958 36974 6010
rect 37026 5958 37038 6010
rect 37090 5958 55182 6010
rect 55234 5958 55246 6010
rect 55298 5958 55310 6010
rect 55362 5958 55374 6010
rect 55426 5958 55438 6010
rect 55490 5958 73582 6010
rect 73634 5958 73646 6010
rect 73698 5958 73710 6010
rect 73762 5958 73774 6010
rect 73826 5958 73838 6010
rect 73890 5958 88596 6010
rect 4876 5936 88596 5958
rect 4876 5466 88596 5488
rect 4876 5414 17722 5466
rect 17774 5414 17786 5466
rect 17838 5414 17850 5466
rect 17902 5414 17914 5466
rect 17966 5414 17978 5466
rect 18030 5414 36122 5466
rect 36174 5414 36186 5466
rect 36238 5414 36250 5466
rect 36302 5414 36314 5466
rect 36366 5414 36378 5466
rect 36430 5414 54522 5466
rect 54574 5414 54586 5466
rect 54638 5414 54650 5466
rect 54702 5414 54714 5466
rect 54766 5414 54778 5466
rect 54830 5414 72922 5466
rect 72974 5414 72986 5466
rect 73038 5414 73050 5466
rect 73102 5414 73114 5466
rect 73166 5414 73178 5466
rect 73230 5414 88596 5466
rect 4876 5392 88596 5414
rect 30686 5280 30692 5332
rect 30744 5329 30750 5332
rect 31514 5329 31520 5332
rect 30744 5323 30793 5329
rect 30744 5289 30747 5323
rect 30781 5289 30793 5323
rect 30744 5283 30793 5289
rect 31492 5323 31520 5329
rect 31492 5289 31504 5323
rect 31492 5283 31520 5289
rect 30744 5280 30750 5283
rect 31514 5280 31520 5283
rect 31572 5280 31578 5332
rect 33814 5280 33820 5332
rect 33872 5329 33878 5332
rect 33872 5323 33921 5329
rect 33872 5289 33875 5323
rect 33909 5289 33921 5323
rect 33872 5283 33921 5289
rect 33872 5280 33878 5283
rect 35102 5280 35108 5332
rect 35160 5329 35166 5332
rect 35930 5329 35936 5332
rect 35160 5323 35209 5329
rect 35160 5289 35163 5323
rect 35197 5289 35209 5323
rect 35160 5283 35209 5289
rect 35887 5323 35936 5329
rect 35887 5289 35899 5323
rect 35933 5289 35936 5323
rect 35887 5283 35936 5289
rect 35160 5280 35166 5283
rect 35930 5280 35936 5283
rect 35988 5280 35994 5332
rect 37126 5329 37132 5332
rect 37083 5323 37132 5329
rect 37083 5289 37095 5323
rect 37129 5289 37132 5323
rect 37083 5283 37132 5289
rect 37126 5280 37132 5283
rect 37184 5280 37190 5332
rect 38414 5280 38420 5332
rect 38472 5329 38478 5332
rect 39242 5329 39248 5332
rect 38472 5323 38521 5329
rect 38472 5289 38475 5323
rect 38509 5289 38521 5323
rect 38472 5283 38521 5289
rect 39220 5323 39248 5329
rect 39220 5289 39232 5323
rect 39220 5283 39248 5289
rect 38472 5280 38478 5283
rect 39242 5280 39248 5283
rect 39300 5280 39306 5332
rect 41634 5329 41640 5332
rect 41591 5323 41640 5329
rect 41591 5289 41603 5323
rect 41637 5289 41640 5323
rect 41591 5283 41640 5289
rect 41634 5280 41640 5283
rect 41692 5280 41698 5332
rect 42830 5280 42836 5332
rect 42888 5329 42894 5332
rect 43658 5329 43664 5332
rect 42888 5323 42937 5329
rect 42888 5289 42891 5323
rect 42925 5289 42937 5323
rect 42888 5283 42937 5289
rect 43615 5323 43664 5329
rect 43615 5289 43627 5323
rect 43661 5289 43664 5323
rect 43615 5283 43664 5289
rect 42888 5280 42894 5283
rect 43658 5280 43664 5283
rect 43716 5280 43722 5332
rect 44762 5280 44768 5332
rect 44820 5329 44826 5332
rect 44820 5323 44869 5329
rect 44820 5289 44823 5323
rect 44857 5289 44869 5323
rect 44820 5283 44869 5289
rect 44820 5280 44826 5283
rect 67854 5280 67860 5332
rect 67912 5320 67918 5332
rect 67995 5323 68053 5329
rect 67995 5320 68007 5323
rect 67912 5292 68007 5320
rect 67912 5280 67918 5292
rect 67995 5289 68007 5292
rect 68041 5289 68053 5323
rect 67995 5283 68053 5289
rect 69326 5280 69332 5332
rect 69384 5329 69390 5332
rect 69384 5323 69433 5329
rect 69384 5289 69387 5323
rect 69421 5289 69433 5323
rect 69384 5283 69433 5289
rect 69384 5280 69390 5283
rect 71166 5280 71172 5332
rect 71224 5329 71230 5332
rect 71224 5323 71273 5329
rect 71224 5289 71227 5323
rect 71261 5289 71273 5323
rect 71224 5283 71273 5289
rect 71224 5280 71230 5283
rect 72270 5280 72276 5332
rect 72328 5320 72334 5332
rect 73374 5329 73380 5332
rect 72503 5323 72561 5329
rect 72503 5320 72515 5323
rect 72328 5292 72515 5320
rect 72328 5280 72334 5292
rect 72503 5289 72515 5292
rect 72549 5289 72561 5323
rect 72503 5283 72561 5289
rect 73353 5323 73380 5329
rect 73353 5289 73365 5323
rect 73353 5283 73380 5289
rect 73374 5280 73380 5283
rect 73432 5280 73438 5332
rect 74478 5280 74484 5332
rect 74536 5329 74542 5332
rect 74536 5323 74585 5329
rect 74536 5289 74539 5323
rect 74573 5289 74585 5323
rect 74536 5283 74585 5289
rect 74536 5280 74542 5283
rect 75582 5280 75588 5332
rect 75640 5320 75646 5332
rect 75723 5323 75781 5329
rect 75723 5320 75735 5323
rect 75640 5292 75735 5320
rect 75640 5280 75646 5292
rect 75723 5289 75735 5292
rect 75769 5289 75781 5323
rect 75723 5283 75781 5289
rect 76686 5280 76692 5332
rect 76744 5320 76750 5332
rect 77103 5323 77161 5329
rect 77103 5320 77115 5323
rect 76744 5292 77115 5320
rect 76744 5280 76750 5292
rect 77103 5289 77115 5292
rect 77149 5289 77161 5323
rect 77103 5283 77161 5289
rect 78894 5280 78900 5332
rect 78952 5329 78958 5332
rect 80274 5329 80280 5332
rect 78952 5323 79001 5329
rect 78952 5289 78955 5323
rect 78989 5289 79001 5323
rect 78952 5283 79001 5289
rect 80231 5323 80280 5329
rect 80231 5289 80243 5323
rect 80277 5289 80280 5323
rect 80231 5283 80280 5289
rect 78952 5280 78958 5283
rect 80274 5280 80280 5283
rect 80332 5280 80338 5332
rect 32710 5212 32716 5264
rect 32768 5261 32774 5264
rect 32768 5255 32817 5261
rect 32768 5221 32771 5255
rect 32805 5221 32817 5255
rect 32768 5215 32817 5221
rect 32768 5212 32774 5215
rect 40438 5212 40444 5264
rect 40496 5261 40502 5264
rect 40496 5255 40545 5261
rect 40496 5221 40499 5255
rect 40533 5221 40545 5255
rect 40496 5215 40545 5221
rect 40496 5212 40502 5215
rect 70062 5212 70068 5264
rect 70120 5261 70126 5264
rect 70120 5255 70169 5261
rect 70120 5221 70123 5255
rect 70157 5221 70169 5255
rect 70120 5215 70169 5221
rect 70120 5212 70126 5215
rect 77790 5212 77796 5264
rect 77848 5261 77854 5264
rect 77848 5255 77897 5261
rect 77848 5221 77851 5255
rect 77885 5221 77897 5255
rect 77848 5215 77897 5221
rect 77848 5212 77854 5215
rect 15230 5110 15236 5162
rect 15288 5150 15294 5162
rect 15325 5153 15383 5159
rect 15325 5150 15337 5153
rect 15288 5122 15337 5150
rect 15288 5110 15294 5122
rect 15325 5119 15337 5122
rect 15371 5119 15383 5153
rect 15325 5113 15383 5119
rect 16058 5110 16064 5162
rect 16116 5159 16122 5162
rect 16116 5153 16150 5159
rect 16138 5119 16150 5153
rect 16116 5113 16150 5119
rect 16116 5110 16122 5113
rect 17162 5110 17168 5162
rect 17220 5110 17226 5162
rect 18266 5110 18272 5162
rect 18324 5150 18330 5162
rect 18405 5153 18463 5159
rect 18405 5150 18417 5153
rect 18324 5122 18417 5150
rect 18324 5110 18330 5122
rect 18405 5119 18417 5122
rect 18451 5119 18463 5153
rect 18405 5113 18463 5119
rect 19646 5110 19652 5162
rect 19704 5150 19710 5162
rect 19741 5153 19799 5159
rect 19741 5150 19753 5153
rect 19704 5122 19753 5150
rect 19704 5110 19710 5122
rect 19741 5119 19753 5122
rect 19787 5119 19799 5153
rect 19741 5113 19799 5119
rect 20474 5110 20480 5162
rect 20532 5110 20538 5162
rect 21578 5110 21584 5162
rect 21636 5150 21642 5162
rect 21673 5153 21731 5159
rect 21673 5150 21685 5153
rect 21636 5122 21685 5150
rect 21636 5110 21642 5122
rect 21673 5119 21685 5122
rect 21719 5119 21731 5153
rect 21673 5113 21731 5119
rect 22958 5110 22964 5162
rect 23016 5150 23022 5162
rect 23053 5153 23111 5159
rect 23053 5150 23065 5153
rect 23016 5122 23065 5150
rect 23016 5110 23022 5122
rect 23053 5119 23065 5122
rect 23099 5119 23111 5153
rect 23053 5113 23111 5119
rect 23786 5110 23792 5162
rect 23844 5159 23850 5162
rect 23844 5153 23878 5159
rect 23866 5119 23878 5153
rect 23844 5113 23878 5119
rect 23844 5110 23850 5113
rect 24890 5110 24896 5162
rect 24948 5110 24954 5162
rect 26086 5110 26092 5162
rect 26144 5150 26150 5162
rect 26181 5153 26239 5159
rect 26181 5150 26193 5153
rect 26144 5122 26193 5150
rect 26144 5110 26150 5122
rect 26181 5119 26193 5122
rect 26227 5119 26239 5153
rect 26181 5113 26239 5119
rect 27374 5110 27380 5162
rect 27432 5150 27438 5162
rect 27469 5153 27527 5159
rect 27469 5150 27481 5153
rect 27432 5122 27481 5150
rect 27432 5110 27438 5122
rect 27469 5119 27481 5122
rect 27515 5119 27527 5153
rect 27469 5113 27527 5119
rect 28202 5110 28208 5162
rect 28260 5110 28266 5162
rect 29306 5110 29312 5162
rect 29364 5150 29370 5162
rect 29401 5153 29459 5159
rect 29401 5150 29413 5153
rect 29364 5122 29413 5150
rect 29364 5110 29370 5122
rect 29401 5119 29413 5122
rect 29447 5119 29459 5153
rect 31333 5153 31391 5159
rect 31333 5150 31345 5153
rect 30919 5127 30977 5133
rect 30919 5124 30931 5127
rect 29401 5113 29459 5119
rect 30704 5116 30931 5124
rect 30612 5096 30931 5116
rect 30612 5088 30732 5096
rect 30919 5093 30931 5096
rect 30965 5093 30977 5127
rect 30612 5060 30640 5088
rect 30919 5087 30977 5093
rect 31256 5122 31345 5150
rect 31256 5060 31284 5122
rect 31333 5119 31345 5122
rect 31379 5119 31391 5153
rect 32621 5153 32679 5159
rect 39061 5153 39119 5159
rect 32621 5150 32633 5153
rect 31333 5113 31391 5119
rect 32544 5122 32633 5150
rect 32544 5060 32572 5122
rect 32621 5119 32633 5122
rect 32667 5119 32679 5153
rect 36071 5147 36129 5153
rect 39061 5150 39073 5153
rect 36071 5144 36083 5147
rect 34047 5127 34105 5133
rect 34047 5124 34059 5127
rect 32621 5113 32679 5119
rect 33832 5096 34059 5124
rect 33832 5060 33860 5096
rect 34047 5093 34059 5096
rect 34093 5093 34105 5127
rect 35335 5127 35393 5133
rect 35764 5128 36083 5144
rect 35335 5124 35347 5127
rect 34047 5087 34105 5093
rect 35120 5096 35347 5124
rect 35120 5060 35148 5096
rect 35335 5093 35347 5096
rect 35381 5093 35393 5127
rect 35335 5087 35393 5093
rect 35746 5076 35752 5128
rect 35804 5116 36083 5128
rect 35804 5076 35810 5116
rect 36071 5113 36083 5116
rect 36117 5144 36129 5147
rect 36117 5125 36252 5144
rect 37267 5127 37325 5133
rect 36117 5119 36267 5125
rect 37267 5124 37279 5127
rect 36117 5116 36221 5119
rect 36117 5113 36129 5116
rect 36071 5107 36129 5113
rect 36209 5085 36221 5116
rect 36255 5085 36267 5119
rect 36209 5079 36267 5085
rect 37144 5096 37279 5124
rect 37144 5060 37172 5096
rect 37267 5093 37279 5096
rect 37313 5093 37325 5127
rect 38647 5127 38705 5133
rect 38647 5124 38659 5127
rect 38432 5116 38659 5124
rect 37267 5087 37325 5093
rect 38340 5096 38659 5116
rect 38340 5088 38460 5096
rect 38647 5093 38659 5096
rect 38693 5093 38705 5127
rect 38340 5060 38368 5088
rect 38647 5087 38705 5093
rect 38984 5122 39073 5150
rect 38984 5060 39012 5122
rect 39061 5119 39073 5122
rect 39107 5119 39119 5153
rect 40349 5153 40407 5159
rect 40349 5150 40361 5153
rect 39061 5113 39119 5119
rect 40272 5122 40361 5150
rect 40272 5060 40300 5122
rect 40349 5119 40361 5122
rect 40395 5119 40407 5153
rect 43785 5147 43843 5153
rect 43785 5144 43797 5147
rect 41775 5127 41833 5133
rect 41775 5124 41787 5127
rect 40349 5113 40407 5119
rect 41560 5096 41787 5124
rect 41560 5060 41588 5096
rect 41775 5093 41787 5096
rect 41821 5093 41833 5127
rect 43063 5127 43121 5133
rect 43492 5128 43797 5144
rect 43063 5124 43075 5127
rect 41775 5087 41833 5093
rect 42848 5096 43075 5124
rect 42848 5060 42876 5096
rect 43063 5093 43075 5096
rect 43109 5093 43121 5127
rect 43063 5087 43121 5093
rect 43474 5076 43480 5128
rect 43532 5116 43797 5128
rect 43532 5076 43538 5116
rect 43785 5113 43797 5116
rect 43831 5144 43843 5147
rect 43831 5125 43980 5144
rect 44995 5127 45053 5133
rect 43831 5119 43995 5125
rect 44995 5124 45007 5127
rect 43831 5116 43949 5119
rect 43831 5113 43843 5116
rect 43785 5107 43843 5113
rect 43937 5085 43949 5116
rect 43983 5085 43995 5119
rect 43937 5079 43995 5085
rect 44780 5096 45007 5124
rect 44780 5060 44808 5096
rect 44995 5093 45007 5096
rect 45041 5093 45053 5127
rect 52398 5110 52404 5162
rect 52456 5150 52462 5162
rect 52537 5153 52595 5159
rect 52537 5150 52549 5153
rect 52456 5122 52549 5150
rect 52456 5110 52462 5122
rect 52537 5119 52549 5122
rect 52583 5119 52595 5153
rect 52537 5113 52595 5119
rect 53686 5110 53692 5162
rect 53744 5150 53750 5162
rect 53917 5153 53975 5159
rect 53917 5150 53929 5153
rect 53744 5122 53929 5150
rect 53744 5110 53750 5122
rect 53917 5119 53929 5122
rect 53963 5119 53975 5153
rect 53917 5113 53975 5119
rect 54769 5153 54827 5159
rect 54769 5119 54781 5153
rect 54815 5150 54827 5153
rect 54882 5150 54888 5162
rect 54815 5122 54888 5150
rect 54815 5119 54827 5122
rect 54769 5113 54827 5119
rect 54882 5110 54888 5122
rect 54940 5110 54946 5162
rect 55710 5110 55716 5162
rect 55768 5150 55774 5162
rect 55805 5153 55863 5159
rect 55805 5150 55817 5153
rect 55768 5122 55817 5150
rect 55768 5110 55774 5122
rect 55805 5119 55817 5122
rect 55851 5119 55863 5153
rect 55805 5113 55863 5119
rect 56814 5110 56820 5162
rect 56872 5150 56878 5162
rect 57045 5153 57103 5159
rect 57045 5150 57057 5153
rect 56872 5122 57057 5150
rect 56872 5110 56878 5122
rect 57045 5119 57057 5122
rect 57091 5119 57103 5153
rect 57045 5113 57103 5119
rect 57918 5110 57924 5162
rect 57976 5159 57982 5162
rect 57976 5153 58010 5159
rect 57998 5119 58010 5153
rect 57976 5113 58010 5119
rect 57976 5110 57982 5113
rect 59022 5110 59028 5162
rect 59080 5150 59086 5162
rect 59117 5153 59175 5159
rect 59117 5150 59129 5153
rect 59080 5122 59129 5150
rect 59080 5110 59086 5122
rect 59117 5119 59129 5122
rect 59163 5119 59175 5153
rect 59117 5113 59175 5119
rect 60126 5110 60132 5162
rect 60184 5150 60190 5162
rect 60265 5153 60323 5159
rect 60265 5150 60277 5153
rect 60184 5122 60277 5150
rect 60184 5110 60190 5122
rect 60265 5119 60277 5122
rect 60311 5119 60323 5153
rect 60265 5113 60323 5119
rect 61414 5110 61420 5162
rect 61472 5150 61478 5162
rect 61645 5153 61703 5159
rect 61645 5150 61657 5153
rect 61472 5122 61657 5150
rect 61472 5110 61478 5122
rect 61645 5119 61657 5122
rect 61691 5119 61703 5153
rect 61645 5113 61703 5119
rect 62334 5110 62340 5162
rect 62392 5150 62398 5162
rect 62460 5153 62518 5159
rect 62460 5150 62472 5153
rect 62392 5122 62472 5150
rect 62392 5110 62398 5122
rect 62460 5119 62472 5122
rect 62506 5119 62518 5153
rect 62460 5113 62518 5119
rect 63438 5110 63444 5162
rect 63496 5150 63502 5162
rect 63533 5153 63591 5159
rect 63533 5150 63545 5153
rect 63496 5122 63545 5150
rect 63496 5110 63502 5122
rect 63533 5119 63545 5122
rect 63579 5119 63591 5153
rect 63533 5113 63591 5119
rect 64542 5110 64548 5162
rect 64600 5150 64606 5162
rect 64773 5153 64831 5159
rect 64773 5150 64785 5153
rect 64600 5122 64785 5150
rect 64600 5110 64606 5122
rect 64773 5119 64785 5122
rect 64819 5119 64831 5153
rect 64773 5113 64831 5119
rect 65646 5110 65652 5162
rect 65704 5159 65710 5162
rect 65704 5153 65738 5159
rect 65726 5119 65738 5153
rect 65704 5113 65738 5119
rect 65704 5110 65710 5113
rect 66750 5110 66756 5162
rect 66808 5150 66814 5162
rect 66845 5153 66903 5159
rect 66845 5150 66857 5153
rect 66808 5122 66857 5150
rect 66808 5110 66814 5122
rect 66845 5119 66857 5122
rect 66891 5119 66903 5153
rect 69543 5147 69601 5153
rect 69543 5144 69555 5147
rect 68179 5127 68237 5133
rect 69252 5128 69555 5144
rect 68179 5124 68191 5127
rect 66845 5113 66903 5119
rect 44995 5087 45053 5093
rect 67964 5096 68191 5124
rect 67964 5060 67992 5096
rect 68179 5093 68191 5096
rect 68225 5093 68237 5127
rect 68179 5087 68237 5093
rect 69234 5076 69240 5128
rect 69292 5116 69555 5128
rect 69292 5076 69298 5116
rect 69543 5113 69555 5116
rect 69589 5144 69601 5147
rect 69589 5125 69740 5144
rect 69589 5119 69755 5125
rect 69589 5116 69709 5119
rect 69589 5113 69601 5116
rect 69543 5107 69601 5113
rect 69697 5085 69709 5116
rect 69743 5085 69755 5119
rect 69878 5110 69884 5162
rect 69936 5150 69942 5162
rect 69973 5153 70031 5159
rect 69973 5150 69985 5153
rect 69936 5122 69985 5150
rect 69936 5110 69942 5122
rect 69973 5119 69985 5122
rect 70019 5150 70031 5153
rect 73193 5153 73251 5159
rect 73193 5150 73205 5153
rect 70019 5125 70292 5150
rect 71399 5127 71457 5133
rect 70019 5122 70307 5125
rect 71399 5124 71411 5127
rect 70019 5119 70031 5122
rect 69973 5113 70031 5119
rect 70249 5119 70307 5122
rect 69697 5079 69755 5085
rect 70249 5085 70261 5119
rect 70295 5085 70307 5119
rect 70249 5079 70307 5085
rect 71184 5096 71411 5124
rect 71184 5060 71212 5096
rect 71399 5093 71411 5096
rect 71445 5093 71457 5127
rect 72687 5127 72745 5133
rect 72687 5124 72699 5127
rect 71399 5087 71457 5093
rect 72472 5096 72699 5124
rect 72472 5060 72500 5096
rect 72687 5093 72699 5096
rect 72733 5093 72745 5127
rect 72687 5087 72745 5093
rect 73116 5122 73205 5150
rect 73116 5060 73144 5122
rect 73193 5119 73205 5122
rect 73239 5119 73251 5153
rect 74711 5147 74769 5153
rect 74711 5144 74723 5147
rect 74404 5128 74723 5144
rect 73193 5113 73251 5119
rect 74386 5076 74392 5128
rect 74444 5116 74723 5128
rect 74444 5076 74450 5116
rect 74711 5113 74723 5116
rect 74757 5144 74769 5147
rect 77271 5147 77329 5153
rect 77271 5144 77283 5147
rect 74757 5125 74892 5144
rect 75907 5127 75965 5133
rect 76980 5128 77283 5144
rect 74757 5119 74907 5125
rect 75907 5124 75919 5127
rect 74757 5116 74861 5119
rect 74757 5113 74769 5116
rect 74711 5107 74769 5113
rect 74849 5085 74861 5116
rect 74895 5085 74907 5119
rect 74849 5079 74907 5085
rect 75692 5096 75919 5124
rect 75692 5060 75720 5096
rect 75907 5093 75919 5096
rect 75953 5093 75965 5127
rect 75907 5087 75965 5093
rect 76962 5076 76968 5128
rect 77020 5116 77283 5128
rect 77020 5076 77026 5116
rect 77271 5113 77283 5116
rect 77317 5144 77329 5147
rect 77317 5125 77468 5144
rect 77317 5119 77483 5125
rect 77317 5116 77437 5119
rect 77317 5113 77329 5116
rect 77271 5107 77329 5113
rect 77425 5085 77437 5116
rect 77471 5085 77483 5119
rect 77606 5110 77612 5162
rect 77664 5150 77670 5162
rect 77701 5153 77759 5159
rect 77701 5150 77713 5153
rect 77664 5122 77713 5150
rect 77664 5110 77670 5122
rect 77701 5119 77713 5122
rect 77747 5150 77759 5153
rect 77747 5125 78020 5150
rect 79127 5127 79185 5133
rect 77747 5122 78035 5125
rect 79127 5124 79139 5127
rect 77747 5119 77759 5122
rect 77701 5113 77759 5119
rect 77977 5119 78035 5122
rect 77425 5079 77483 5085
rect 77977 5085 77989 5119
rect 78023 5085 78035 5119
rect 77977 5079 78035 5085
rect 78912 5096 79139 5124
rect 78912 5060 78940 5096
rect 79127 5093 79139 5096
rect 79173 5093 79185 5127
rect 80415 5127 80473 5133
rect 80415 5124 80427 5127
rect 79127 5087 79185 5093
rect 80200 5096 80427 5124
rect 80200 5060 80228 5096
rect 80415 5093 80427 5096
rect 80461 5093 80473 5127
rect 80415 5087 80473 5093
rect 15138 5008 15144 5060
rect 15196 5048 15202 5060
rect 15480 5051 15538 5057
rect 15480 5048 15492 5051
rect 15196 5020 15492 5048
rect 15196 5008 15202 5020
rect 15480 5017 15492 5020
rect 15526 5017 15538 5051
rect 15480 5011 15538 5017
rect 15782 5008 15788 5060
rect 15840 5048 15846 5060
rect 15923 5051 15981 5057
rect 15923 5048 15935 5051
rect 15840 5020 15935 5048
rect 15840 5008 15846 5020
rect 15923 5017 15935 5020
rect 15969 5017 15981 5051
rect 15923 5011 15981 5017
rect 17070 5008 17076 5060
rect 17128 5048 17134 5060
rect 17320 5051 17378 5057
rect 17320 5048 17332 5051
rect 17128 5020 17332 5048
rect 17128 5008 17134 5020
rect 17320 5017 17332 5020
rect 17366 5017 17378 5051
rect 17320 5011 17378 5017
rect 18266 5008 18272 5060
rect 18324 5048 18330 5060
rect 18608 5051 18666 5057
rect 18608 5048 18620 5051
rect 18324 5020 18620 5048
rect 18324 5008 18330 5020
rect 18608 5017 18620 5020
rect 18654 5017 18666 5051
rect 18608 5011 18666 5017
rect 19646 5008 19652 5060
rect 19704 5048 19710 5060
rect 19896 5051 19954 5057
rect 19896 5048 19908 5051
rect 19704 5020 19908 5048
rect 19704 5008 19710 5020
rect 19896 5017 19908 5020
rect 19942 5017 19954 5051
rect 19896 5011 19954 5017
rect 20290 5008 20296 5060
rect 20348 5048 20354 5060
rect 20632 5051 20690 5057
rect 20632 5048 20644 5051
rect 20348 5020 20644 5048
rect 20348 5008 20354 5020
rect 20632 5017 20644 5020
rect 20678 5017 20690 5051
rect 20632 5011 20690 5017
rect 21578 5008 21584 5060
rect 21636 5048 21642 5060
rect 21828 5051 21886 5057
rect 21828 5048 21840 5051
rect 21636 5020 21840 5048
rect 21636 5008 21642 5020
rect 21828 5017 21840 5020
rect 21874 5017 21886 5051
rect 21828 5011 21886 5017
rect 22866 5008 22872 5060
rect 22924 5048 22930 5060
rect 23208 5051 23266 5057
rect 23208 5048 23220 5051
rect 22924 5020 23220 5048
rect 22924 5008 22930 5020
rect 23208 5017 23220 5020
rect 23254 5017 23266 5051
rect 23208 5011 23266 5017
rect 23510 5008 23516 5060
rect 23568 5048 23574 5060
rect 23651 5051 23709 5057
rect 23651 5048 23663 5051
rect 23568 5020 23663 5048
rect 23568 5008 23574 5020
rect 23651 5017 23663 5020
rect 23697 5017 23709 5051
rect 23651 5011 23709 5017
rect 24798 5008 24804 5060
rect 24856 5048 24862 5060
rect 25048 5051 25106 5057
rect 25048 5048 25060 5051
rect 24856 5020 25060 5048
rect 24856 5008 24862 5020
rect 25048 5017 25060 5020
rect 25094 5017 25106 5051
rect 25048 5011 25106 5017
rect 26086 5008 26092 5060
rect 26144 5048 26150 5060
rect 26336 5051 26394 5057
rect 26336 5048 26348 5051
rect 26144 5020 26348 5048
rect 26144 5008 26150 5020
rect 26336 5017 26348 5020
rect 26382 5017 26394 5051
rect 26336 5011 26394 5017
rect 27374 5008 27380 5060
rect 27432 5048 27438 5060
rect 27624 5051 27682 5057
rect 27624 5048 27636 5051
rect 27432 5020 27636 5048
rect 27432 5008 27438 5020
rect 27624 5017 27636 5020
rect 27670 5017 27682 5051
rect 27624 5011 27682 5017
rect 28018 5008 28024 5060
rect 28076 5048 28082 5060
rect 28360 5051 28418 5057
rect 28360 5048 28372 5051
rect 28076 5020 28372 5048
rect 28076 5008 28082 5020
rect 28360 5017 28372 5020
rect 28406 5017 28418 5051
rect 28360 5011 28418 5017
rect 29306 5008 29312 5060
rect 29364 5048 29370 5060
rect 29556 5051 29614 5057
rect 29556 5048 29568 5051
rect 29364 5020 29568 5048
rect 29364 5008 29370 5020
rect 29556 5017 29568 5020
rect 29602 5017 29614 5051
rect 29556 5011 29614 5017
rect 30505 5051 30563 5057
rect 30505 5017 30517 5051
rect 30551 5048 30563 5051
rect 30594 5048 30600 5060
rect 30551 5020 30600 5048
rect 30551 5017 30563 5020
rect 30505 5011 30563 5017
rect 30594 5008 30600 5020
rect 30652 5008 30658 5060
rect 31149 5051 31207 5057
rect 31149 5017 31161 5051
rect 31195 5048 31207 5051
rect 31238 5048 31244 5060
rect 31195 5020 31244 5048
rect 31195 5017 31207 5020
rect 31149 5011 31207 5017
rect 31238 5008 31244 5020
rect 31296 5008 31302 5060
rect 32437 5051 32495 5057
rect 32437 5017 32449 5051
rect 32483 5048 32495 5051
rect 32526 5048 32532 5060
rect 32483 5020 32532 5048
rect 32483 5017 32495 5020
rect 32437 5011 32495 5017
rect 32526 5008 32532 5020
rect 32584 5008 32590 5060
rect 33725 5051 33783 5057
rect 33725 5017 33737 5051
rect 33771 5048 33783 5051
rect 33814 5048 33820 5060
rect 33771 5020 33820 5048
rect 33771 5017 33783 5020
rect 33725 5011 33783 5017
rect 33814 5008 33820 5020
rect 33872 5008 33878 5060
rect 35013 5051 35071 5057
rect 35013 5017 35025 5051
rect 35059 5048 35071 5051
rect 35102 5048 35108 5060
rect 35059 5020 35108 5048
rect 35059 5017 35071 5020
rect 35013 5011 35071 5017
rect 35102 5008 35108 5020
rect 35160 5008 35166 5060
rect 36945 5051 37003 5057
rect 36945 5017 36957 5051
rect 36991 5048 37003 5051
rect 37126 5048 37132 5060
rect 36991 5020 37132 5048
rect 36991 5017 37003 5020
rect 36945 5011 37003 5017
rect 37126 5008 37132 5020
rect 37184 5008 37190 5060
rect 38233 5051 38291 5057
rect 38233 5017 38245 5051
rect 38279 5048 38291 5051
rect 38322 5048 38328 5060
rect 38279 5020 38328 5048
rect 38279 5017 38291 5020
rect 38233 5011 38291 5017
rect 38322 5008 38328 5020
rect 38380 5008 38386 5060
rect 38877 5051 38935 5057
rect 38877 5017 38889 5051
rect 38923 5048 38935 5051
rect 38966 5048 38972 5060
rect 38923 5020 38972 5048
rect 38923 5017 38935 5020
rect 38877 5011 38935 5017
rect 38966 5008 38972 5020
rect 39024 5008 39030 5060
rect 40165 5051 40223 5057
rect 40165 5017 40177 5051
rect 40211 5048 40223 5051
rect 40254 5048 40260 5060
rect 40211 5020 40260 5048
rect 40211 5017 40223 5020
rect 40165 5011 40223 5017
rect 40254 5008 40260 5020
rect 40312 5008 40318 5060
rect 41453 5051 41511 5057
rect 41453 5017 41465 5051
rect 41499 5048 41511 5051
rect 41542 5048 41548 5060
rect 41499 5020 41548 5048
rect 41499 5017 41511 5020
rect 41453 5011 41511 5017
rect 41542 5008 41548 5020
rect 41600 5008 41606 5060
rect 42741 5051 42799 5057
rect 42741 5017 42753 5051
rect 42787 5048 42799 5051
rect 42830 5048 42836 5060
rect 42787 5020 42836 5048
rect 42787 5017 42799 5020
rect 42741 5011 42799 5017
rect 42830 5008 42836 5020
rect 42888 5008 42894 5060
rect 44673 5051 44731 5057
rect 44673 5017 44685 5051
rect 44719 5048 44731 5051
rect 44762 5048 44768 5060
rect 44719 5020 44768 5048
rect 44719 5017 44731 5020
rect 44673 5011 44731 5017
rect 44762 5008 44768 5020
rect 44820 5008 44826 5060
rect 52490 5008 52496 5060
rect 52548 5048 52554 5060
rect 52740 5051 52798 5057
rect 52740 5048 52752 5051
rect 52548 5020 52752 5048
rect 52548 5008 52554 5020
rect 52740 5017 52752 5020
rect 52786 5017 52798 5051
rect 52740 5011 52798 5017
rect 53778 5008 53784 5060
rect 53836 5048 53842 5060
rect 54120 5051 54178 5057
rect 54120 5048 54132 5051
rect 53836 5020 54132 5048
rect 53836 5008 53842 5020
rect 54120 5017 54132 5020
rect 54166 5017 54178 5051
rect 54120 5011 54178 5017
rect 54422 5008 54428 5060
rect 54480 5048 54486 5060
rect 54563 5051 54621 5057
rect 54563 5048 54575 5051
rect 54480 5020 54575 5048
rect 54480 5008 54486 5020
rect 54563 5017 54575 5020
rect 54609 5017 54621 5051
rect 54563 5011 54621 5017
rect 55710 5008 55716 5060
rect 55768 5048 55774 5060
rect 55960 5051 56018 5057
rect 55960 5048 55972 5051
rect 55768 5020 55972 5048
rect 55768 5008 55774 5020
rect 55960 5017 55972 5020
rect 56006 5017 56018 5051
rect 55960 5011 56018 5017
rect 56998 5008 57004 5060
rect 57056 5048 57062 5060
rect 57248 5051 57306 5057
rect 57248 5048 57260 5051
rect 57056 5020 57260 5048
rect 57056 5008 57062 5020
rect 57248 5017 57260 5020
rect 57294 5017 57306 5051
rect 57248 5011 57306 5017
rect 57642 5008 57648 5060
rect 57700 5048 57706 5060
rect 57783 5051 57841 5057
rect 57783 5048 57795 5051
rect 57700 5020 57795 5048
rect 57700 5008 57706 5020
rect 57783 5017 57795 5020
rect 57829 5017 57841 5051
rect 57783 5011 57841 5017
rect 58930 5008 58936 5060
rect 58988 5048 58994 5060
rect 59272 5051 59330 5057
rect 59272 5048 59284 5051
rect 58988 5020 59284 5048
rect 58988 5008 58994 5020
rect 59272 5017 59284 5020
rect 59318 5017 59330 5051
rect 59272 5011 59330 5017
rect 60218 5008 60224 5060
rect 60276 5048 60282 5060
rect 60468 5051 60526 5057
rect 60468 5048 60480 5051
rect 60276 5020 60480 5048
rect 60276 5008 60282 5020
rect 60468 5017 60480 5020
rect 60514 5017 60526 5051
rect 60468 5011 60526 5017
rect 61506 5008 61512 5060
rect 61564 5048 61570 5060
rect 61848 5051 61906 5057
rect 61848 5048 61860 5051
rect 61564 5020 61860 5048
rect 61564 5008 61570 5020
rect 61848 5017 61860 5020
rect 61894 5017 61906 5051
rect 61848 5011 61906 5017
rect 62150 5008 62156 5060
rect 62208 5048 62214 5060
rect 62291 5051 62349 5057
rect 62291 5048 62303 5051
rect 62208 5020 62303 5048
rect 62208 5008 62214 5020
rect 62291 5017 62303 5020
rect 62337 5017 62349 5051
rect 62291 5011 62349 5017
rect 63438 5008 63444 5060
rect 63496 5048 63502 5060
rect 63688 5051 63746 5057
rect 63688 5048 63700 5051
rect 63496 5020 63700 5048
rect 63496 5008 63502 5020
rect 63688 5017 63700 5020
rect 63734 5017 63746 5051
rect 63688 5011 63746 5017
rect 64726 5008 64732 5060
rect 64784 5048 64790 5060
rect 64976 5051 65034 5057
rect 64976 5048 64988 5051
rect 64784 5020 64988 5048
rect 64784 5008 64790 5020
rect 64976 5017 64988 5020
rect 65022 5017 65034 5051
rect 64976 5011 65034 5017
rect 65370 5008 65376 5060
rect 65428 5048 65434 5060
rect 65511 5051 65569 5057
rect 65511 5048 65523 5051
rect 65428 5020 65523 5048
rect 65428 5008 65434 5020
rect 65511 5017 65523 5020
rect 65557 5017 65569 5051
rect 65511 5011 65569 5017
rect 66658 5008 66664 5060
rect 66716 5048 66722 5060
rect 67000 5051 67058 5057
rect 67000 5048 67012 5051
rect 66716 5020 67012 5048
rect 66716 5008 66722 5020
rect 67000 5017 67012 5020
rect 67046 5017 67058 5051
rect 67000 5011 67058 5017
rect 67857 5051 67915 5057
rect 67857 5017 67869 5051
rect 67903 5048 67915 5051
rect 67946 5048 67952 5060
rect 67903 5020 67952 5048
rect 67903 5017 67915 5020
rect 67857 5011 67915 5017
rect 67946 5008 67952 5020
rect 68004 5008 68010 5060
rect 71077 5051 71135 5057
rect 71077 5017 71089 5051
rect 71123 5048 71135 5051
rect 71166 5048 71172 5060
rect 71123 5020 71172 5048
rect 71123 5017 71135 5020
rect 71077 5011 71135 5017
rect 71166 5008 71172 5020
rect 71224 5008 71230 5060
rect 72365 5051 72423 5057
rect 72365 5017 72377 5051
rect 72411 5048 72423 5051
rect 72454 5048 72460 5060
rect 72411 5020 72460 5048
rect 72411 5017 72423 5020
rect 72365 5011 72423 5017
rect 72454 5008 72460 5020
rect 72512 5008 72518 5060
rect 73009 5051 73067 5057
rect 73009 5017 73021 5051
rect 73055 5048 73067 5051
rect 73098 5048 73104 5060
rect 73055 5020 73104 5048
rect 73055 5017 73067 5020
rect 73009 5011 73067 5017
rect 73098 5008 73104 5020
rect 73156 5008 73162 5060
rect 75585 5051 75643 5057
rect 75585 5017 75597 5051
rect 75631 5048 75643 5051
rect 75674 5048 75680 5060
rect 75631 5020 75680 5048
rect 75631 5017 75643 5020
rect 75585 5011 75643 5017
rect 75674 5008 75680 5020
rect 75732 5008 75738 5060
rect 78805 5051 78863 5057
rect 78805 5017 78817 5051
rect 78851 5048 78863 5051
rect 78894 5048 78900 5060
rect 78851 5020 78900 5048
rect 78851 5017 78863 5020
rect 78805 5011 78863 5017
rect 78894 5008 78900 5020
rect 78952 5008 78958 5060
rect 80093 5051 80151 5057
rect 80093 5017 80105 5051
rect 80139 5048 80151 5051
rect 80182 5048 80188 5060
rect 80139 5020 80188 5048
rect 80139 5017 80151 5020
rect 80093 5011 80151 5017
rect 80182 5008 80188 5020
rect 80240 5008 80246 5060
rect 4876 4922 88596 4944
rect 4876 4870 18382 4922
rect 18434 4870 18446 4922
rect 18498 4870 18510 4922
rect 18562 4870 18574 4922
rect 18626 4870 18638 4922
rect 18690 4870 36782 4922
rect 36834 4870 36846 4922
rect 36898 4870 36910 4922
rect 36962 4870 36974 4922
rect 37026 4870 37038 4922
rect 37090 4870 55182 4922
rect 55234 4870 55246 4922
rect 55298 4870 55310 4922
rect 55362 4870 55374 4922
rect 55426 4870 55438 4922
rect 55490 4870 73582 4922
rect 73634 4870 73646 4922
rect 73698 4870 73710 4922
rect 73762 4870 73774 4922
rect 73826 4870 73838 4922
rect 73890 4870 88596 4922
rect 4876 4848 88596 4870
<< via1 >>
rect 18382 87558 18434 87610
rect 18446 87558 18498 87610
rect 18510 87558 18562 87610
rect 18574 87558 18626 87610
rect 18638 87558 18690 87610
rect 36782 87558 36834 87610
rect 36846 87558 36898 87610
rect 36910 87558 36962 87610
rect 36974 87558 37026 87610
rect 37038 87558 37090 87610
rect 55182 87558 55234 87610
rect 55246 87558 55298 87610
rect 55310 87558 55362 87610
rect 55374 87558 55426 87610
rect 55438 87558 55490 87610
rect 73582 87558 73634 87610
rect 73646 87558 73698 87610
rect 73710 87558 73762 87610
rect 73774 87558 73826 87610
rect 73838 87558 73890 87610
rect 10636 87424 10688 87476
rect 15144 87424 15196 87476
rect 17076 87424 17128 87476
rect 18272 87467 18324 87476
rect 18272 87433 18281 87467
rect 18281 87433 18315 87467
rect 18315 87433 18324 87467
rect 18272 87424 18324 87433
rect 19652 87424 19704 87476
rect 21584 87424 21636 87476
rect 22872 87424 22924 87476
rect 23516 87424 23568 87476
rect 24804 87424 24856 87476
rect 26092 87424 26144 87476
rect 27380 87424 27432 87476
rect 29312 87424 29364 87476
rect 30600 87424 30652 87476
rect 31244 87424 31296 87476
rect 32532 87424 32584 87476
rect 33820 87424 33872 87476
rect 35108 87424 35160 87476
rect 35752 87424 35804 87476
rect 37132 87424 37184 87476
rect 37684 87424 37736 87476
rect 10728 87365 10780 87374
rect 10728 87331 10737 87365
rect 10737 87331 10771 87365
rect 10771 87331 10780 87365
rect 10728 87322 10780 87331
rect 15788 87356 15840 87408
rect 18272 87288 18324 87340
rect 19560 87288 19612 87340
rect 20296 87356 20348 87408
rect 28024 87356 28076 87408
rect 30600 87322 30652 87374
rect 31520 87365 31572 87374
rect 31520 87331 31560 87365
rect 31560 87331 31572 87365
rect 31520 87322 31572 87331
rect 32624 87365 32676 87374
rect 32624 87331 32633 87365
rect 32633 87331 32667 87365
rect 32667 87331 32676 87365
rect 32624 87322 32676 87331
rect 33728 87322 33780 87374
rect 34924 87322 34976 87374
rect 35936 87365 35988 87374
rect 35936 87331 35945 87365
rect 35945 87331 35979 87365
rect 35979 87331 35988 87365
rect 35936 87322 35988 87331
rect 37132 87365 37184 87374
rect 37132 87331 37141 87365
rect 37141 87331 37175 87365
rect 37175 87331 37184 87365
rect 37132 87322 37184 87331
rect 22688 87220 22740 87272
rect 27104 87220 27156 87272
rect 38328 87424 38380 87476
rect 38972 87424 39024 87476
rect 40260 87424 40312 87476
rect 40904 87424 40956 87476
rect 42192 87424 42244 87476
rect 43480 87424 43532 87476
rect 44124 87424 44176 87476
rect 52496 87424 52548 87476
rect 55716 87424 55768 87476
rect 57004 87424 57056 87476
rect 57648 87424 57700 87476
rect 60224 87424 60276 87476
rect 63444 87424 63496 87476
rect 64732 87424 64784 87476
rect 65376 87424 65428 87476
rect 67952 87424 68004 87476
rect 69240 87424 69292 87476
rect 69884 87424 69936 87476
rect 71172 87424 71224 87476
rect 72460 87424 72512 87476
rect 73104 87424 73156 87476
rect 74392 87424 74444 87476
rect 75680 87424 75732 87476
rect 76968 87424 77020 87476
rect 77612 87424 77664 87476
rect 78900 87424 78952 87476
rect 80188 87424 80240 87476
rect 80832 87424 80884 87476
rect 82120 87424 82172 87476
rect 38144 87322 38196 87374
rect 39248 87322 39300 87374
rect 40352 87365 40404 87374
rect 40352 87331 40361 87365
rect 40361 87331 40395 87365
rect 40395 87331 40404 87365
rect 40352 87322 40404 87331
rect 42560 87365 42612 87374
rect 42560 87331 42579 87365
rect 42579 87331 42612 87365
rect 42560 87322 42612 87331
rect 42836 87356 42888 87408
rect 43664 87365 43716 87374
rect 43664 87331 43673 87365
rect 43673 87331 43707 87365
rect 43707 87331 43716 87365
rect 43664 87322 43716 87331
rect 44676 87322 44728 87374
rect 44768 87356 44820 87408
rect 45412 87356 45464 87408
rect 46056 87356 46108 87408
rect 46700 87356 46752 87408
rect 47344 87356 47396 87408
rect 47988 87356 48040 87408
rect 48632 87356 48684 87408
rect 49276 87356 49328 87408
rect 49920 87356 49972 87408
rect 50564 87356 50616 87408
rect 53784 87356 53836 87408
rect 54428 87322 54480 87374
rect 58936 87356 58988 87408
rect 60132 87288 60184 87340
rect 61512 87356 61564 87408
rect 62156 87322 62208 87374
rect 66664 87356 66716 87408
rect 67860 87322 67912 87374
rect 69332 87322 69384 87374
rect 70068 87322 70120 87374
rect 71172 87322 71224 87374
rect 72276 87322 72328 87374
rect 73380 87365 73432 87374
rect 73380 87331 73420 87365
rect 73420 87331 73432 87365
rect 73380 87322 73432 87331
rect 74484 87322 74536 87374
rect 75588 87322 75640 87374
rect 76692 87288 76744 87340
rect 77796 87322 77848 87374
rect 78900 87322 78952 87374
rect 80280 87365 80332 87374
rect 80280 87331 80289 87365
rect 80289 87331 80323 87365
rect 80323 87331 80332 87365
rect 80280 87322 80332 87331
rect 81108 87365 81160 87374
rect 81108 87331 81148 87365
rect 81148 87331 81160 87365
rect 81108 87322 81160 87331
rect 82212 87322 82264 87374
rect 39064 87263 39116 87272
rect 39064 87229 39073 87263
rect 39073 87229 39107 87263
rect 39107 87229 39116 87263
rect 39064 87220 39116 87229
rect 56820 87220 56872 87272
rect 62340 87220 62392 87272
rect 64548 87220 64600 87272
rect 15512 87195 15564 87204
rect 15512 87161 15521 87195
rect 15521 87161 15555 87195
rect 15555 87161 15564 87195
rect 15512 87152 15564 87161
rect 16064 87152 16116 87204
rect 17168 87152 17220 87204
rect 20480 87152 20532 87204
rect 21584 87152 21636 87204
rect 23792 87195 23844 87204
rect 23792 87161 23811 87195
rect 23811 87161 23844 87195
rect 23792 87152 23844 87161
rect 25080 87195 25132 87204
rect 25080 87161 25098 87195
rect 25098 87161 25132 87195
rect 25080 87152 25132 87161
rect 26092 87152 26144 87204
rect 28208 87152 28260 87204
rect 29312 87152 29364 87204
rect 41824 87195 41876 87204
rect 41824 87161 41833 87195
rect 41833 87161 41867 87195
rect 41867 87161 41876 87195
rect 41824 87152 41876 87161
rect 52680 87152 52732 87204
rect 53508 87152 53560 87204
rect 54428 87152 54480 87204
rect 55716 87152 55768 87204
rect 57924 87195 57976 87204
rect 57924 87161 57943 87195
rect 57943 87161 57976 87195
rect 57924 87152 57976 87161
rect 59028 87152 59080 87204
rect 61236 87152 61288 87204
rect 63444 87152 63496 87204
rect 65652 87195 65704 87204
rect 65652 87161 65671 87195
rect 65671 87161 65704 87195
rect 65652 87152 65704 87161
rect 66756 87152 66808 87204
rect 17722 87014 17774 87066
rect 17786 87014 17838 87066
rect 17850 87014 17902 87066
rect 17914 87014 17966 87066
rect 17978 87014 18030 87066
rect 36122 87014 36174 87066
rect 36186 87014 36238 87066
rect 36250 87014 36302 87066
rect 36314 87014 36366 87066
rect 36378 87014 36430 87066
rect 54522 87014 54574 87066
rect 54586 87014 54638 87066
rect 54650 87014 54702 87066
rect 54714 87014 54766 87066
rect 54778 87014 54830 87066
rect 72922 87014 72974 87066
rect 72986 87014 73038 87066
rect 73050 87014 73102 87066
rect 73114 87014 73166 87066
rect 73178 87014 73230 87066
rect 41548 86880 41600 86932
rect 41456 86710 41508 86762
rect 18382 86470 18434 86522
rect 18446 86470 18498 86522
rect 18510 86470 18562 86522
rect 18574 86470 18626 86522
rect 18638 86470 18690 86522
rect 36782 86470 36834 86522
rect 36846 86470 36898 86522
rect 36910 86470 36962 86522
rect 36974 86470 37026 86522
rect 37038 86470 37090 86522
rect 55182 86470 55234 86522
rect 55246 86470 55298 86522
rect 55310 86470 55362 86522
rect 55374 86470 55426 86522
rect 55438 86470 55490 86522
rect 73582 86470 73634 86522
rect 73646 86470 73698 86522
rect 73710 86470 73762 86522
rect 73774 86470 73826 86522
rect 73838 86470 73890 86522
rect 17722 85926 17774 85978
rect 17786 85926 17838 85978
rect 17850 85926 17902 85978
rect 17914 85926 17966 85978
rect 17978 85926 18030 85978
rect 36122 85926 36174 85978
rect 36186 85926 36238 85978
rect 36250 85926 36302 85978
rect 36314 85926 36366 85978
rect 36378 85926 36430 85978
rect 54522 85926 54574 85978
rect 54586 85926 54638 85978
rect 54650 85926 54702 85978
rect 54714 85926 54766 85978
rect 54778 85926 54830 85978
rect 72922 85926 72974 85978
rect 72986 85926 73038 85978
rect 73050 85926 73102 85978
rect 73114 85926 73166 85978
rect 73178 85926 73230 85978
rect 18382 85382 18434 85434
rect 18446 85382 18498 85434
rect 18510 85382 18562 85434
rect 18574 85382 18626 85434
rect 18638 85382 18690 85434
rect 36782 85382 36834 85434
rect 36846 85382 36898 85434
rect 36910 85382 36962 85434
rect 36974 85382 37026 85434
rect 37038 85382 37090 85434
rect 55182 85382 55234 85434
rect 55246 85382 55298 85434
rect 55310 85382 55362 85434
rect 55374 85382 55426 85434
rect 55438 85382 55490 85434
rect 73582 85382 73634 85434
rect 73646 85382 73698 85434
rect 73710 85382 73762 85434
rect 73774 85382 73826 85434
rect 73838 85382 73890 85434
rect 41824 84976 41876 85028
rect 49092 84976 49144 85028
rect 5954 84838 6006 84890
rect 6018 84838 6070 84890
rect 6082 84838 6134 84890
rect 6146 84838 6198 84890
rect 6210 84838 6262 84890
rect 17722 84838 17774 84890
rect 17786 84838 17838 84890
rect 17850 84838 17902 84890
rect 17914 84838 17966 84890
rect 17978 84838 18030 84890
rect 36122 84838 36174 84890
rect 36186 84838 36238 84890
rect 36250 84838 36302 84890
rect 36314 84838 36366 84890
rect 36378 84838 36430 84890
rect 54522 84838 54574 84890
rect 54586 84838 54638 84890
rect 54650 84838 54702 84890
rect 54714 84838 54766 84890
rect 54778 84838 54830 84890
rect 72922 84838 72974 84890
rect 72986 84838 73038 84890
rect 73050 84838 73102 84890
rect 73114 84838 73166 84890
rect 73178 84838 73230 84890
rect 86546 84838 86598 84890
rect 86610 84838 86662 84890
rect 86674 84838 86726 84890
rect 86738 84838 86790 84890
rect 86802 84838 86854 84890
rect 12752 84636 12804 84688
rect 30692 84704 30744 84756
rect 11648 84568 11700 84620
rect 30692 84568 30744 84620
rect 39616 84704 39668 84756
rect 46148 84704 46200 84756
rect 31244 84636 31296 84688
rect 39064 84636 39116 84688
rect 50196 84636 50248 84688
rect 7416 84500 7468 84552
rect 10544 84432 10596 84484
rect 13856 84432 13908 84484
rect 31152 84568 31204 84620
rect 41824 84568 41876 84620
rect 46056 84568 46108 84620
rect 46148 84568 46200 84620
rect 51300 84568 51352 84620
rect 47160 84500 47212 84552
rect 45872 84432 45924 84484
rect 45964 84475 46016 84484
rect 45964 84441 45973 84475
rect 45973 84441 46007 84475
rect 46007 84441 46016 84475
rect 45964 84432 46016 84441
rect 49092 84432 49144 84484
rect 50196 84432 50248 84484
rect 6690 84294 6742 84346
rect 6754 84294 6806 84346
rect 6818 84294 6870 84346
rect 6882 84294 6934 84346
rect 6946 84294 6998 84346
rect 18382 84294 18434 84346
rect 18446 84294 18498 84346
rect 18510 84294 18562 84346
rect 18574 84294 18626 84346
rect 18638 84294 18690 84346
rect 36782 84294 36834 84346
rect 36846 84294 36898 84346
rect 36910 84294 36962 84346
rect 36974 84294 37026 84346
rect 37038 84294 37090 84346
rect 55182 84294 55234 84346
rect 55246 84294 55298 84346
rect 55310 84294 55362 84346
rect 55374 84294 55426 84346
rect 55438 84294 55490 84346
rect 73582 84294 73634 84346
rect 73646 84294 73698 84346
rect 73710 84294 73762 84346
rect 73774 84294 73826 84346
rect 73838 84294 73890 84346
rect 87282 84294 87334 84346
rect 87346 84294 87398 84346
rect 87410 84294 87462 84346
rect 87474 84294 87526 84346
rect 87538 84294 87590 84346
rect 5954 83750 6006 83802
rect 6018 83750 6070 83802
rect 6082 83750 6134 83802
rect 6146 83750 6198 83802
rect 6210 83750 6262 83802
rect 86546 83750 86598 83802
rect 86610 83750 86662 83802
rect 86674 83750 86726 83802
rect 86738 83750 86790 83802
rect 86802 83750 86854 83802
rect 6690 83206 6742 83258
rect 6754 83206 6806 83258
rect 6818 83206 6870 83258
rect 6882 83206 6934 83258
rect 6946 83206 6998 83258
rect 87282 83206 87334 83258
rect 87346 83206 87398 83258
rect 87410 83206 87462 83258
rect 87474 83206 87526 83258
rect 87538 83206 87590 83258
rect 13856 83072 13908 83124
rect 83316 83072 83368 83124
rect 47068 83004 47120 83056
rect 47160 83004 47212 83056
rect 47988 83004 48040 83056
rect 5954 82662 6006 82714
rect 6018 82662 6070 82714
rect 6082 82662 6134 82714
rect 6146 82662 6198 82714
rect 6210 82662 6262 82714
rect 86546 82662 86598 82714
rect 86610 82662 86662 82714
rect 86674 82662 86726 82714
rect 86738 82662 86790 82714
rect 86802 82662 86854 82714
rect 14988 82392 15040 82444
rect 15512 82392 15564 82444
rect 68948 82392 69000 82444
rect 69332 82392 69384 82444
rect 7600 82324 7652 82376
rect 11676 82324 11728 82376
rect 7232 82256 7284 82308
rect 12780 82256 12832 82308
rect 6690 82118 6742 82170
rect 6754 82118 6806 82170
rect 6818 82118 6870 82170
rect 6882 82118 6934 82170
rect 6946 82118 6998 82170
rect 87282 82118 87334 82170
rect 87346 82118 87398 82170
rect 87410 82118 87462 82170
rect 87474 82118 87526 82170
rect 87538 82118 87590 82170
rect 7784 81712 7836 81764
rect 9992 81712 10044 81764
rect 5954 81574 6006 81626
rect 6018 81574 6070 81626
rect 6082 81574 6134 81626
rect 6146 81574 6198 81626
rect 6210 81574 6262 81626
rect 86546 81574 86598 81626
rect 86610 81574 86662 81626
rect 86674 81574 86726 81626
rect 86738 81574 86790 81626
rect 86802 81574 86854 81626
rect 83500 81372 83552 81424
rect 88376 81244 88428 81296
rect 6690 81030 6742 81082
rect 6754 81030 6806 81082
rect 6818 81030 6870 81082
rect 6882 81030 6934 81082
rect 6946 81030 6998 81082
rect 87282 81030 87334 81082
rect 87346 81030 87398 81082
rect 87410 81030 87462 81082
rect 87474 81030 87526 81082
rect 87538 81030 87590 81082
rect 5954 80486 6006 80538
rect 6018 80486 6070 80538
rect 6082 80486 6134 80538
rect 6146 80486 6198 80538
rect 6210 80486 6262 80538
rect 86546 80486 86598 80538
rect 86610 80486 86662 80538
rect 86674 80486 86726 80538
rect 86738 80486 86790 80538
rect 86802 80486 86854 80538
rect 88284 80225 88336 80234
rect 7140 80148 7192 80200
rect 83500 80148 83552 80200
rect 88284 80191 88299 80225
rect 88299 80191 88336 80225
rect 88284 80182 88336 80191
rect 2908 80080 2960 80132
rect 6690 79942 6742 79994
rect 6754 79942 6806 79994
rect 6818 79942 6870 79994
rect 6882 79942 6934 79994
rect 6946 79942 6998 79994
rect 87282 79942 87334 79994
rect 87346 79942 87398 79994
rect 87410 79942 87462 79994
rect 87474 79942 87526 79994
rect 87538 79942 87590 79994
rect 5954 79398 6006 79450
rect 6018 79398 6070 79450
rect 6082 79398 6134 79450
rect 6146 79398 6198 79450
rect 6210 79398 6262 79450
rect 86546 79398 86598 79450
rect 86610 79398 86662 79450
rect 86674 79398 86726 79450
rect 86738 79398 86790 79450
rect 86802 79398 86854 79450
rect 6690 78854 6742 78906
rect 6754 78854 6806 78906
rect 6818 78854 6870 78906
rect 6882 78854 6934 78906
rect 6946 78854 6998 78906
rect 87282 78854 87334 78906
rect 87346 78854 87398 78906
rect 87410 78854 87462 78906
rect 87474 78854 87526 78906
rect 87538 78854 87590 78906
rect 7140 78652 7192 78704
rect 88284 78661 88336 78670
rect 88284 78627 88299 78661
rect 88299 78627 88336 78661
rect 88284 78618 88336 78627
rect 88008 78516 88060 78568
rect 2908 78448 2960 78500
rect 5954 78310 6006 78362
rect 6018 78310 6070 78362
rect 6082 78310 6134 78362
rect 6146 78310 6198 78362
rect 6210 78310 6262 78362
rect 86546 78310 86598 78362
rect 86610 78310 86662 78362
rect 86674 78310 86726 78362
rect 86738 78310 86790 78362
rect 86802 78310 86854 78362
rect 88284 78049 88336 78058
rect 7140 77972 7192 78024
rect 88284 78015 88299 78049
rect 88299 78015 88336 78049
rect 88284 78006 88336 78015
rect 2908 77904 2960 77956
rect 87824 77904 87876 77956
rect 6690 77766 6742 77818
rect 6754 77766 6806 77818
rect 6818 77766 6870 77818
rect 6882 77766 6934 77818
rect 6946 77766 6998 77818
rect 87282 77766 87334 77818
rect 87346 77766 87398 77818
rect 87410 77766 87462 77818
rect 87474 77766 87526 77818
rect 87538 77766 87590 77818
rect 5954 77222 6006 77274
rect 6018 77222 6070 77274
rect 6082 77222 6134 77274
rect 6146 77222 6198 77274
rect 6210 77222 6262 77274
rect 86546 77222 86598 77274
rect 86610 77222 86662 77274
rect 86674 77222 86726 77274
rect 86738 77222 86790 77274
rect 86802 77222 86854 77274
rect 7140 76884 7192 76936
rect 2724 76816 2776 76868
rect 86628 76816 86680 76868
rect 88008 76859 88060 76868
rect 88008 76825 88017 76859
rect 88017 76825 88051 76859
rect 88051 76825 88060 76859
rect 88008 76816 88060 76825
rect 6690 76678 6742 76730
rect 6754 76678 6806 76730
rect 6818 76678 6870 76730
rect 6882 76678 6934 76730
rect 6946 76678 6998 76730
rect 87282 76678 87334 76730
rect 87346 76678 87398 76730
rect 87410 76678 87462 76730
rect 87474 76678 87526 76730
rect 87538 76678 87590 76730
rect 5954 76134 6006 76186
rect 6018 76134 6070 76186
rect 6082 76134 6134 76186
rect 6146 76134 6198 76186
rect 6210 76134 6262 76186
rect 86546 76134 86598 76186
rect 86610 76134 86662 76186
rect 86674 76134 86726 76186
rect 86738 76134 86790 76186
rect 86802 76134 86854 76186
rect 86904 75932 86956 75984
rect 7140 75796 7192 75848
rect 88468 75796 88520 75848
rect 2908 75728 2960 75780
rect 6690 75590 6742 75642
rect 6754 75590 6806 75642
rect 6818 75590 6870 75642
rect 6882 75590 6934 75642
rect 6946 75590 6998 75642
rect 87282 75590 87334 75642
rect 87346 75590 87398 75642
rect 87410 75590 87462 75642
rect 87474 75590 87526 75642
rect 87538 75590 87590 75642
rect 5954 75046 6006 75098
rect 6018 75046 6070 75098
rect 6082 75046 6134 75098
rect 6146 75046 6198 75098
rect 6210 75046 6262 75098
rect 86546 75046 86598 75098
rect 86610 75046 86662 75098
rect 86674 75046 86726 75098
rect 86738 75046 86790 75098
rect 86802 75046 86854 75098
rect 4380 74844 4432 74896
rect 84420 74844 84472 74896
rect 5668 74742 5720 74794
rect 88560 74776 88612 74828
rect 6690 74502 6742 74554
rect 6754 74502 6806 74554
rect 6818 74502 6870 74554
rect 6882 74502 6934 74554
rect 6946 74502 6998 74554
rect 87282 74502 87334 74554
rect 87346 74502 87398 74554
rect 87410 74502 87462 74554
rect 87474 74502 87526 74554
rect 87538 74502 87590 74554
rect 5954 73958 6006 74010
rect 6018 73958 6070 74010
rect 6082 73958 6134 74010
rect 6146 73958 6198 74010
rect 6210 73958 6262 74010
rect 86546 73958 86598 74010
rect 86610 73958 86662 74010
rect 86674 73958 86726 74010
rect 86738 73958 86790 74010
rect 86802 73958 86854 74010
rect 6690 73414 6742 73466
rect 6754 73414 6806 73466
rect 6818 73414 6870 73466
rect 6882 73414 6934 73466
rect 6946 73414 6998 73466
rect 87282 73414 87334 73466
rect 87346 73414 87398 73466
rect 87410 73414 87462 73466
rect 87474 73414 87526 73466
rect 87538 73414 87590 73466
rect 7140 73212 7192 73264
rect 88284 73221 88336 73230
rect 88008 73144 88060 73196
rect 88284 73187 88299 73221
rect 88299 73187 88336 73221
rect 88284 73178 88336 73187
rect 2908 73008 2960 73060
rect 5954 72870 6006 72922
rect 6018 72870 6070 72922
rect 6082 72870 6134 72922
rect 6146 72870 6198 72922
rect 6210 72870 6262 72922
rect 86546 72870 86598 72922
rect 86610 72870 86662 72922
rect 86674 72870 86726 72922
rect 86738 72870 86790 72922
rect 86802 72870 86854 72922
rect 88284 72603 88336 72612
rect 7140 72532 7192 72584
rect 87180 72532 87232 72584
rect 88284 72569 88299 72603
rect 88299 72569 88336 72603
rect 88284 72560 88336 72569
rect 2908 72464 2960 72516
rect 6690 72326 6742 72378
rect 6754 72326 6806 72378
rect 6818 72326 6870 72378
rect 6882 72326 6934 72378
rect 6946 72326 6998 72378
rect 87282 72326 87334 72378
rect 87346 72326 87398 72378
rect 87410 72326 87462 72378
rect 87474 72326 87526 72378
rect 87538 72326 87590 72378
rect 5954 71782 6006 71834
rect 6018 71782 6070 71834
rect 6082 71782 6134 71834
rect 6146 71782 6198 71834
rect 6210 71782 6262 71834
rect 86546 71782 86598 71834
rect 86610 71782 86662 71834
rect 86674 71782 86726 71834
rect 86738 71782 86790 71834
rect 86802 71782 86854 71834
rect 86904 71580 86956 71632
rect 88284 71521 88336 71530
rect 7140 71444 7192 71496
rect 88284 71487 88299 71521
rect 88299 71487 88336 71521
rect 88284 71478 88336 71487
rect 2724 71376 2776 71428
rect 6690 71238 6742 71290
rect 6754 71238 6806 71290
rect 6818 71238 6870 71290
rect 6882 71238 6934 71290
rect 6946 71238 6998 71290
rect 87282 71238 87334 71290
rect 87346 71238 87398 71290
rect 87410 71238 87462 71290
rect 87474 71238 87526 71290
rect 87538 71238 87590 71290
rect 5954 70694 6006 70746
rect 6018 70694 6070 70746
rect 6082 70694 6134 70746
rect 6146 70694 6198 70746
rect 6210 70694 6262 70746
rect 86546 70694 86598 70746
rect 86610 70694 86662 70746
rect 86674 70694 86726 70746
rect 86738 70694 86790 70746
rect 86802 70694 86854 70746
rect 86904 70492 86956 70544
rect 88192 70433 88244 70476
rect 88192 70424 88233 70433
rect 88233 70424 88244 70433
rect 7140 70356 7192 70408
rect 2908 70288 2960 70340
rect 6690 70150 6742 70202
rect 6754 70150 6806 70202
rect 6818 70150 6870 70202
rect 6882 70150 6934 70202
rect 6946 70150 6998 70202
rect 87282 70150 87334 70202
rect 87346 70150 87398 70202
rect 87410 70150 87462 70202
rect 87474 70150 87526 70202
rect 87538 70150 87590 70202
rect 5954 69606 6006 69658
rect 6018 69606 6070 69658
rect 6082 69606 6134 69658
rect 6146 69606 6198 69658
rect 6210 69606 6262 69658
rect 86546 69606 86598 69658
rect 86610 69606 86662 69658
rect 86674 69606 86726 69658
rect 86738 69606 86790 69658
rect 86802 69606 86854 69658
rect 5668 69302 5720 69354
rect 86904 69268 86956 69320
rect 4380 69200 4432 69252
rect 88560 69268 88612 69320
rect 6690 69062 6742 69114
rect 6754 69062 6806 69114
rect 6818 69062 6870 69114
rect 6882 69062 6934 69114
rect 6946 69062 6998 69114
rect 87282 69062 87334 69114
rect 87346 69062 87398 69114
rect 87410 69062 87462 69114
rect 87474 69062 87526 69114
rect 87538 69062 87590 69114
rect 5954 68518 6006 68570
rect 6018 68518 6070 68570
rect 6082 68518 6134 68570
rect 6146 68518 6198 68570
rect 6210 68518 6262 68570
rect 86546 68518 86598 68570
rect 86610 68518 86662 68570
rect 86674 68518 86726 68570
rect 86738 68518 86790 68570
rect 86802 68518 86854 68570
rect 6690 67974 6742 68026
rect 6754 67974 6806 68026
rect 6818 67974 6870 68026
rect 6882 67974 6934 68026
rect 6946 67974 6998 68026
rect 87282 67974 87334 68026
rect 87346 67974 87398 68026
rect 87410 67974 87462 68026
rect 87474 67974 87526 68026
rect 87538 67974 87590 68026
rect 5668 67738 5720 67790
rect 88284 67781 88336 67790
rect 88284 67747 88299 67781
rect 88299 67747 88336 67781
rect 88284 67738 88336 67747
rect 84420 67636 84472 67688
rect 2908 67568 2960 67620
rect 5954 67430 6006 67482
rect 6018 67430 6070 67482
rect 6082 67430 6134 67482
rect 6146 67430 6198 67482
rect 6210 67430 6262 67482
rect 86546 67430 86598 67482
rect 86610 67430 86662 67482
rect 86674 67430 86726 67482
rect 86738 67430 86790 67482
rect 86802 67430 86854 67482
rect 88284 67163 88336 67172
rect 7140 67092 7192 67144
rect 86904 67092 86956 67144
rect 88284 67129 88299 67163
rect 88299 67129 88336 67163
rect 88284 67120 88336 67129
rect 2908 67024 2960 67076
rect 6690 66886 6742 66938
rect 6754 66886 6806 66938
rect 6818 66886 6870 66938
rect 6882 66886 6934 66938
rect 6946 66886 6998 66938
rect 87282 66886 87334 66938
rect 87346 66886 87398 66938
rect 87410 66886 87462 66938
rect 87474 66886 87526 66938
rect 87538 66886 87590 66938
rect 5954 66342 6006 66394
rect 6018 66342 6070 66394
rect 6082 66342 6134 66394
rect 6146 66342 6198 66394
rect 6210 66342 6262 66394
rect 86546 66342 86598 66394
rect 86610 66342 86662 66394
rect 86674 66342 86726 66394
rect 86738 66342 86790 66394
rect 86802 66342 86854 66394
rect 2908 65936 2960 65988
rect 7232 66004 7284 66056
rect 87088 66004 87140 66056
rect 88192 65979 88244 65988
rect 88192 65945 88215 65979
rect 88215 65945 88244 65979
rect 88192 65936 88244 65945
rect 6690 65798 6742 65850
rect 6754 65798 6806 65850
rect 6818 65798 6870 65850
rect 6882 65798 6934 65850
rect 6946 65798 6998 65850
rect 87282 65798 87334 65850
rect 87346 65798 87398 65850
rect 87410 65798 87462 65850
rect 87474 65798 87526 65850
rect 87538 65798 87590 65850
rect 5954 65254 6006 65306
rect 6018 65254 6070 65306
rect 6082 65254 6134 65306
rect 6146 65254 6198 65306
rect 6210 65254 6262 65306
rect 86546 65254 86598 65306
rect 86610 65254 86662 65306
rect 86674 65254 86726 65306
rect 86738 65254 86790 65306
rect 86802 65254 86854 65306
rect 2908 64848 2960 64900
rect 7232 64916 7284 64968
rect 87088 64916 87140 64968
rect 88376 64848 88428 64900
rect 6690 64710 6742 64762
rect 6754 64710 6806 64762
rect 6818 64710 6870 64762
rect 6882 64710 6934 64762
rect 6946 64710 6998 64762
rect 87282 64710 87334 64762
rect 87346 64710 87398 64762
rect 87410 64710 87462 64762
rect 87474 64710 87526 64762
rect 87538 64710 87590 64762
rect 7416 64576 7468 64628
rect 5954 64166 6006 64218
rect 6018 64166 6070 64218
rect 6082 64166 6134 64218
rect 6146 64166 6198 64218
rect 6210 64166 6262 64218
rect 86546 64166 86598 64218
rect 86610 64166 86662 64218
rect 86674 64166 86726 64218
rect 86738 64166 86790 64218
rect 86802 64166 86854 64218
rect 5208 63905 5260 63914
rect 5208 63871 5217 63905
rect 5217 63871 5251 63905
rect 5251 63871 5260 63905
rect 5208 63862 5260 63871
rect 9624 63896 9676 63948
rect 7416 63871 7468 63880
rect 7416 63837 7435 63871
rect 7435 63837 7468 63871
rect 7416 63828 7468 63837
rect 84420 63828 84472 63880
rect 7232 63760 7284 63812
rect 7784 63760 7836 63812
rect 88560 63760 88612 63812
rect 6690 63622 6742 63674
rect 6754 63622 6806 63674
rect 6818 63622 6870 63674
rect 6882 63622 6934 63674
rect 6946 63622 6998 63674
rect 87282 63622 87334 63674
rect 87346 63622 87398 63674
rect 87410 63622 87462 63674
rect 87474 63622 87526 63674
rect 87538 63622 87590 63674
rect 7324 63216 7376 63268
rect 5954 63078 6006 63130
rect 6018 63078 6070 63130
rect 6082 63078 6134 63130
rect 6146 63078 6198 63130
rect 6210 63078 6262 63130
rect 86546 63078 86598 63130
rect 86610 63078 86662 63130
rect 86674 63078 86726 63130
rect 86738 63078 86790 63130
rect 86802 63078 86854 63130
rect 6690 62534 6742 62586
rect 6754 62534 6806 62586
rect 6818 62534 6870 62586
rect 6882 62534 6934 62586
rect 6946 62534 6998 62586
rect 87282 62534 87334 62586
rect 87346 62534 87398 62586
rect 87410 62534 87462 62586
rect 87474 62534 87526 62586
rect 87538 62534 87590 62586
rect 7232 62400 7284 62452
rect 4932 62298 4984 62350
rect 87088 62332 87140 62384
rect 88560 62332 88612 62384
rect 5954 61990 6006 62042
rect 6018 61990 6070 62042
rect 6082 61990 6134 62042
rect 6146 61990 6198 62042
rect 6210 61990 6262 62042
rect 86546 61990 86598 62042
rect 86610 61990 86662 62042
rect 86674 61990 86726 62042
rect 86738 61990 86790 62042
rect 86802 61990 86854 62042
rect 2908 61584 2960 61636
rect 7232 61652 7284 61704
rect 87088 61652 87140 61704
rect 88192 61627 88244 61636
rect 88192 61593 88215 61627
rect 88215 61593 88244 61627
rect 88192 61584 88244 61593
rect 6690 61446 6742 61498
rect 6754 61446 6806 61498
rect 6818 61446 6870 61498
rect 6882 61446 6934 61498
rect 6946 61446 6998 61498
rect 87282 61446 87334 61498
rect 87346 61446 87398 61498
rect 87410 61446 87462 61498
rect 87474 61446 87526 61498
rect 87538 61446 87590 61498
rect 5954 60902 6006 60954
rect 6018 60902 6070 60954
rect 6082 60902 6134 60954
rect 6146 60902 6198 60954
rect 6210 60902 6262 60954
rect 86546 60902 86598 60954
rect 86610 60902 86662 60954
rect 86674 60902 86726 60954
rect 86738 60902 86790 60954
rect 86802 60902 86854 60954
rect 2908 60496 2960 60548
rect 7232 60564 7284 60616
rect 87088 60564 87140 60616
rect 88192 60539 88244 60548
rect 88192 60505 88215 60539
rect 88215 60505 88244 60539
rect 88192 60496 88244 60505
rect 6690 60358 6742 60410
rect 6754 60358 6806 60410
rect 6818 60358 6870 60410
rect 6882 60358 6934 60410
rect 6946 60358 6998 60410
rect 87282 60358 87334 60410
rect 87346 60358 87398 60410
rect 87410 60358 87462 60410
rect 87474 60358 87526 60410
rect 87538 60358 87590 60410
rect 5954 59814 6006 59866
rect 6018 59814 6070 59866
rect 6082 59814 6134 59866
rect 6146 59814 6198 59866
rect 6210 59814 6262 59866
rect 86546 59814 86598 59866
rect 86610 59814 86662 59866
rect 86674 59814 86726 59866
rect 86738 59814 86790 59866
rect 86802 59814 86854 59866
rect 5208 59519 5217 59528
rect 5217 59519 5251 59528
rect 5251 59519 5260 59528
rect 5208 59476 5260 59519
rect 7232 59476 7284 59528
rect 87640 59476 87692 59528
rect 88376 59408 88428 59460
rect 6690 59270 6742 59322
rect 6754 59270 6806 59322
rect 6818 59270 6870 59322
rect 6882 59270 6934 59322
rect 6946 59270 6998 59322
rect 87282 59270 87334 59322
rect 87346 59270 87398 59322
rect 87410 59270 87462 59322
rect 87474 59270 87526 59322
rect 87538 59270 87590 59322
rect 5954 58726 6006 58778
rect 6018 58726 6070 58778
rect 6082 58726 6134 58778
rect 6146 58726 6198 58778
rect 6210 58726 6262 58778
rect 86546 58726 86598 58778
rect 86610 58726 86662 58778
rect 86674 58726 86726 58778
rect 86738 58726 86790 58778
rect 86802 58726 86854 58778
rect 5208 58465 5260 58474
rect 5208 58431 5217 58465
rect 5217 58431 5251 58465
rect 5251 58431 5260 58465
rect 5208 58422 5260 58431
rect 88008 58465 88060 58474
rect 88008 58431 88017 58465
rect 88017 58431 88051 58465
rect 88051 58431 88060 58465
rect 88008 58422 88060 58431
rect 5392 58363 5444 58372
rect 5392 58329 5410 58363
rect 5410 58329 5444 58363
rect 5392 58320 5444 58329
rect 88560 58320 88612 58372
rect 6690 58182 6742 58234
rect 6754 58182 6806 58234
rect 6818 58182 6870 58234
rect 6882 58182 6934 58234
rect 6946 58182 6998 58234
rect 87282 58182 87334 58234
rect 87346 58182 87398 58234
rect 87410 58182 87462 58234
rect 87474 58182 87526 58234
rect 87538 58182 87590 58234
rect 5954 57638 6006 57690
rect 6018 57638 6070 57690
rect 6082 57638 6134 57690
rect 6146 57638 6198 57690
rect 6210 57638 6262 57690
rect 86546 57638 86598 57690
rect 86610 57638 86662 57690
rect 86674 57638 86726 57690
rect 86738 57638 86790 57690
rect 86802 57638 86854 57690
rect 6690 57094 6742 57146
rect 6754 57094 6806 57146
rect 6818 57094 6870 57146
rect 6882 57094 6934 57146
rect 6946 57094 6998 57146
rect 87282 57094 87334 57146
rect 87346 57094 87398 57146
rect 87410 57094 87462 57146
rect 87474 57094 87526 57146
rect 87538 57094 87590 57146
rect 7232 56960 7284 57012
rect 4932 56858 4984 56910
rect 88008 56901 88060 56910
rect 88008 56867 88017 56901
rect 88017 56867 88051 56901
rect 88051 56867 88060 56901
rect 88008 56858 88060 56867
rect 88836 56824 88888 56876
rect 5954 56550 6006 56602
rect 6018 56550 6070 56602
rect 6082 56550 6134 56602
rect 6146 56550 6198 56602
rect 6210 56550 6262 56602
rect 86546 56550 86598 56602
rect 86610 56550 86662 56602
rect 86674 56550 86726 56602
rect 86738 56550 86790 56602
rect 86802 56550 86854 56602
rect 2908 56212 2960 56264
rect 7232 56212 7284 56264
rect 87088 56212 87140 56264
rect 88192 56187 88244 56196
rect 88192 56153 88215 56187
rect 88215 56153 88244 56187
rect 88192 56144 88244 56153
rect 6690 56006 6742 56058
rect 6754 56006 6806 56058
rect 6818 56006 6870 56058
rect 6882 56006 6934 56058
rect 6946 56006 6998 56058
rect 87282 56006 87334 56058
rect 87346 56006 87398 56058
rect 87410 56006 87462 56058
rect 87474 56006 87526 56058
rect 87538 56006 87590 56058
rect 5954 55462 6006 55514
rect 6018 55462 6070 55514
rect 6082 55462 6134 55514
rect 6146 55462 6198 55514
rect 6210 55462 6262 55514
rect 86546 55462 86598 55514
rect 86610 55462 86662 55514
rect 86674 55462 86726 55514
rect 86738 55462 86790 55514
rect 86802 55462 86854 55514
rect 2908 55124 2960 55176
rect 7232 55124 7284 55176
rect 87088 55124 87140 55176
rect 88192 55099 88244 55108
rect 88192 55065 88215 55099
rect 88215 55065 88244 55099
rect 88192 55056 88244 55065
rect 6690 54918 6742 54970
rect 6754 54918 6806 54970
rect 6818 54918 6870 54970
rect 6882 54918 6934 54970
rect 6946 54918 6998 54970
rect 87282 54918 87334 54970
rect 87346 54918 87398 54970
rect 87410 54918 87462 54970
rect 87474 54918 87526 54970
rect 87538 54918 87590 54970
rect 5954 54374 6006 54426
rect 6018 54374 6070 54426
rect 6082 54374 6134 54426
rect 6146 54374 6198 54426
rect 6210 54374 6262 54426
rect 86546 54374 86598 54426
rect 86610 54374 86662 54426
rect 86674 54374 86726 54426
rect 86738 54374 86790 54426
rect 86802 54374 86854 54426
rect 5116 54036 5168 54088
rect 5668 54036 5720 54088
rect 84420 54036 84472 54088
rect 88652 54036 88704 54088
rect 6690 53830 6742 53882
rect 6754 53830 6806 53882
rect 6818 53830 6870 53882
rect 6882 53830 6934 53882
rect 6946 53830 6998 53882
rect 87282 53830 87334 53882
rect 87346 53830 87398 53882
rect 87410 53830 87462 53882
rect 87474 53830 87526 53882
rect 87538 53830 87590 53882
rect 5954 53286 6006 53338
rect 6018 53286 6070 53338
rect 6082 53286 6134 53338
rect 6146 53286 6198 53338
rect 6210 53286 6262 53338
rect 86546 53286 86598 53338
rect 86610 53286 86662 53338
rect 86674 53286 86726 53338
rect 86738 53286 86790 53338
rect 86802 53286 86854 53338
rect 2908 52948 2960 53000
rect 7232 52948 7284 53000
rect 87088 52948 87140 53000
rect 88284 52880 88336 52932
rect 6690 52742 6742 52794
rect 6754 52742 6806 52794
rect 6818 52742 6870 52794
rect 6882 52742 6934 52794
rect 6946 52742 6998 52794
rect 87282 52742 87334 52794
rect 87346 52742 87398 52794
rect 87410 52742 87462 52794
rect 87474 52742 87526 52794
rect 87538 52742 87590 52794
rect 5954 52198 6006 52250
rect 6018 52198 6070 52250
rect 6082 52198 6134 52250
rect 6146 52198 6198 52250
rect 6210 52198 6262 52250
rect 86546 52198 86598 52250
rect 86610 52198 86662 52250
rect 86674 52198 86726 52250
rect 86738 52198 86790 52250
rect 86802 52198 86854 52250
rect 6690 51654 6742 51706
rect 6754 51654 6806 51706
rect 6818 51654 6870 51706
rect 6882 51654 6934 51706
rect 6946 51654 6998 51706
rect 87282 51654 87334 51706
rect 87346 51654 87398 51706
rect 87410 51654 87462 51706
rect 87474 51654 87526 51706
rect 87538 51654 87590 51706
rect 7232 51520 7284 51572
rect 2908 51384 2960 51436
rect 85800 51452 85852 51504
rect 88192 51359 88244 51368
rect 88192 51325 88215 51359
rect 88215 51325 88244 51359
rect 88192 51316 88244 51325
rect 5954 51110 6006 51162
rect 6018 51110 6070 51162
rect 6082 51110 6134 51162
rect 6146 51110 6198 51162
rect 6210 51110 6262 51162
rect 86546 51110 86598 51162
rect 86610 51110 86662 51162
rect 86674 51110 86726 51162
rect 86738 51110 86790 51162
rect 86802 51110 86854 51162
rect 85432 50704 85484 50756
rect 6690 50566 6742 50618
rect 6754 50566 6806 50618
rect 6818 50566 6870 50618
rect 6882 50566 6934 50618
rect 6946 50566 6998 50618
rect 87282 50566 87334 50618
rect 87346 50566 87398 50618
rect 87410 50566 87462 50618
rect 87474 50566 87526 50618
rect 87538 50566 87590 50618
rect 5954 50022 6006 50074
rect 6018 50022 6070 50074
rect 6082 50022 6134 50074
rect 6146 50022 6198 50074
rect 6210 50022 6262 50074
rect 86546 50022 86598 50074
rect 86610 50022 86662 50074
rect 86674 50022 86726 50074
rect 86738 50022 86790 50074
rect 86802 50022 86854 50074
rect 85524 49616 85576 49668
rect 6690 49478 6742 49530
rect 6754 49478 6806 49530
rect 6818 49478 6870 49530
rect 6882 49478 6934 49530
rect 6946 49478 6998 49530
rect 87282 49478 87334 49530
rect 87346 49478 87398 49530
rect 87410 49478 87462 49530
rect 87474 49478 87526 49530
rect 87538 49478 87590 49530
rect 5954 48934 6006 48986
rect 6018 48934 6070 48986
rect 6082 48934 6134 48986
rect 6146 48934 6198 48986
rect 6210 48934 6262 48986
rect 86546 48934 86598 48986
rect 86610 48934 86662 48986
rect 86674 48934 86726 48986
rect 86738 48934 86790 48986
rect 86802 48934 86854 48986
rect 88192 48639 88244 48648
rect 88192 48605 88201 48639
rect 88201 48605 88235 48639
rect 88235 48605 88244 48639
rect 88192 48596 88244 48605
rect 85340 48528 85392 48580
rect 6690 48390 6742 48442
rect 6754 48390 6806 48442
rect 6818 48390 6870 48442
rect 6882 48390 6934 48442
rect 6946 48390 6998 48442
rect 87282 48390 87334 48442
rect 87346 48390 87398 48442
rect 87410 48390 87462 48442
rect 87474 48390 87526 48442
rect 87538 48390 87590 48442
rect 88192 48027 88244 48036
rect 88192 47993 88201 48027
rect 88201 47993 88235 48027
rect 88235 47993 88244 48027
rect 88192 47984 88244 47993
rect 5954 47846 6006 47898
rect 6018 47846 6070 47898
rect 6082 47846 6134 47898
rect 6146 47846 6198 47898
rect 6210 47846 6262 47898
rect 86546 47846 86598 47898
rect 86610 47846 86662 47898
rect 86674 47846 86726 47898
rect 86738 47846 86790 47898
rect 86802 47846 86854 47898
rect 85800 47508 85852 47560
rect 88192 47483 88244 47492
rect 88192 47449 88215 47483
rect 88215 47449 88244 47483
rect 88192 47440 88244 47449
rect 6690 47302 6742 47354
rect 6754 47302 6806 47354
rect 6818 47302 6870 47354
rect 6882 47302 6934 47354
rect 6946 47302 6998 47354
rect 87282 47302 87334 47354
rect 87346 47302 87398 47354
rect 87410 47302 87462 47354
rect 87474 47302 87526 47354
rect 87538 47302 87590 47354
rect 88192 46939 88244 46948
rect 88192 46905 88201 46939
rect 88201 46905 88235 46939
rect 88235 46905 88244 46939
rect 88192 46896 88244 46905
rect 5954 46758 6006 46810
rect 6018 46758 6070 46810
rect 6082 46758 6134 46810
rect 6146 46758 6198 46810
rect 6210 46758 6262 46810
rect 86546 46758 86598 46810
rect 86610 46758 86662 46810
rect 86674 46758 86726 46810
rect 86738 46758 86790 46810
rect 86802 46758 86854 46810
rect 6690 46214 6742 46266
rect 6754 46214 6806 46266
rect 6818 46214 6870 46266
rect 6882 46214 6934 46266
rect 6946 46214 6998 46266
rect 87282 46214 87334 46266
rect 87346 46214 87398 46266
rect 87410 46214 87462 46266
rect 87474 46214 87526 46266
rect 87538 46214 87590 46266
rect 5392 45876 5444 45928
rect 13884 45876 13936 45928
rect 46424 45876 46476 45928
rect 51284 45876 51336 45928
rect 85800 45876 85852 45928
rect 88192 45851 88244 45860
rect 88192 45817 88201 45851
rect 88201 45817 88235 45851
rect 88235 45817 88244 45851
rect 88192 45808 88244 45817
rect 5954 45670 6006 45722
rect 6018 45670 6070 45722
rect 6082 45670 6134 45722
rect 6146 45670 6198 45722
rect 6210 45670 6262 45722
rect 86546 45670 86598 45722
rect 86610 45670 86662 45722
rect 86674 45670 86726 45722
rect 86738 45670 86790 45722
rect 86802 45670 86854 45722
rect 5392 45579 5444 45588
rect 5392 45545 5410 45579
rect 5410 45545 5444 45579
rect 5392 45536 5444 45545
rect 7324 45579 7376 45588
rect 7324 45545 7333 45579
rect 7333 45545 7367 45579
rect 7367 45545 7376 45579
rect 7324 45536 7376 45545
rect 9992 45536 10044 45588
rect 85800 45579 85852 45588
rect 85800 45545 85809 45579
rect 85809 45545 85843 45579
rect 85843 45545 85852 45579
rect 85800 45536 85852 45545
rect 7140 45511 7192 45520
rect 7140 45477 7149 45511
rect 7149 45477 7183 45511
rect 7183 45477 7192 45511
rect 7140 45468 7192 45477
rect 85984 45511 86036 45520
rect 85984 45477 85993 45511
rect 85993 45477 86027 45511
rect 86027 45477 86036 45511
rect 85984 45468 86036 45477
rect 2908 45332 2960 45384
rect 86168 45375 86220 45384
rect 86168 45341 86177 45375
rect 86177 45341 86211 45375
rect 86211 45341 86220 45375
rect 86168 45332 86220 45341
rect 88192 45375 88244 45384
rect 88192 45341 88201 45375
rect 88201 45341 88235 45375
rect 88235 45341 88244 45375
rect 88192 45332 88244 45341
rect 85616 45307 85668 45316
rect 85616 45273 85625 45307
rect 85625 45273 85659 45307
rect 85659 45273 85668 45307
rect 85616 45264 85668 45273
rect 6690 45126 6742 45178
rect 6754 45126 6806 45178
rect 6818 45126 6870 45178
rect 6882 45126 6934 45178
rect 6946 45126 6998 45178
rect 87282 45126 87334 45178
rect 87346 45126 87398 45178
rect 87410 45126 87462 45178
rect 87474 45126 87526 45178
rect 87538 45126 87590 45178
rect 7508 45035 7560 45044
rect 7508 45001 7517 45035
rect 7517 45001 7551 45035
rect 7551 45001 7560 45035
rect 7508 44992 7560 45001
rect 88284 44933 88336 44942
rect 7140 44856 7192 44908
rect 88284 44899 88299 44933
rect 88299 44899 88336 44933
rect 88284 44890 88336 44899
rect 87180 44788 87232 44840
rect 2908 44720 2960 44772
rect 5954 44582 6006 44634
rect 6018 44582 6070 44634
rect 6082 44582 6134 44634
rect 6146 44582 6198 44634
rect 6210 44582 6262 44634
rect 86546 44582 86598 44634
rect 86610 44582 86662 44634
rect 86674 44582 86726 44634
rect 86738 44582 86790 44634
rect 86802 44582 86854 44634
rect 88284 44315 88336 44324
rect 8152 44244 8204 44296
rect 85800 44244 85852 44296
rect 88284 44281 88299 44315
rect 88299 44281 88336 44315
rect 88284 44272 88336 44281
rect 2724 44176 2776 44228
rect 6690 44038 6742 44090
rect 6754 44038 6806 44090
rect 6818 44038 6870 44090
rect 6882 44038 6934 44090
rect 6946 44038 6998 44090
rect 87282 44038 87334 44090
rect 87346 44038 87398 44090
rect 87410 44038 87462 44090
rect 87474 44038 87526 44090
rect 87538 44038 87590 44090
rect 5954 43494 6006 43546
rect 6018 43494 6070 43546
rect 6082 43494 6134 43546
rect 6146 43494 6198 43546
rect 6210 43494 6262 43546
rect 86546 43494 86598 43546
rect 86610 43494 86662 43546
rect 86674 43494 86726 43546
rect 86738 43494 86790 43546
rect 86802 43494 86854 43546
rect 6690 42950 6742 43002
rect 6754 42950 6806 43002
rect 6818 42950 6870 43002
rect 6882 42950 6934 43002
rect 6946 42950 6998 43002
rect 87282 42950 87334 43002
rect 87346 42950 87398 43002
rect 87410 42950 87462 43002
rect 87474 42950 87526 43002
rect 87538 42950 87590 43002
rect 88284 42757 88336 42766
rect 7140 42680 7192 42732
rect 88284 42723 88299 42757
rect 88299 42723 88336 42757
rect 88284 42714 88336 42723
rect 86352 42612 86404 42664
rect 2908 42544 2960 42596
rect 5954 42406 6006 42458
rect 6018 42406 6070 42458
rect 6082 42406 6134 42458
rect 6146 42406 6198 42458
rect 6210 42406 6262 42458
rect 86546 42406 86598 42458
rect 86610 42406 86662 42458
rect 86674 42406 86726 42458
rect 86738 42406 86790 42458
rect 86802 42406 86854 42458
rect 6690 41862 6742 41914
rect 6754 41862 6806 41914
rect 6818 41862 6870 41914
rect 6882 41862 6934 41914
rect 6946 41862 6998 41914
rect 87282 41862 87334 41914
rect 87346 41862 87398 41914
rect 87410 41862 87462 41914
rect 87474 41862 87526 41914
rect 87538 41862 87590 41914
rect 4380 41728 4432 41780
rect 87180 41728 87232 41780
rect 5668 41626 5720 41678
rect 88284 41669 88336 41678
rect 88284 41635 88299 41669
rect 88299 41635 88336 41669
rect 88284 41626 88336 41635
rect 5954 41318 6006 41370
rect 6018 41318 6070 41370
rect 6082 41318 6134 41370
rect 6146 41318 6198 41370
rect 6210 41318 6262 41370
rect 86546 41318 86598 41370
rect 86610 41318 86662 41370
rect 86674 41318 86726 41370
rect 86738 41318 86790 41370
rect 86802 41318 86854 41370
rect 6690 40774 6742 40826
rect 6754 40774 6806 40826
rect 6818 40774 6870 40826
rect 6882 40774 6934 40826
rect 6946 40774 6998 40826
rect 87282 40774 87334 40826
rect 87346 40774 87398 40826
rect 87410 40774 87462 40826
rect 87474 40774 87526 40826
rect 87538 40774 87590 40826
rect 7140 40504 7192 40556
rect 87916 40547 87968 40556
rect 87916 40513 87925 40547
rect 87925 40513 87959 40547
rect 87959 40513 87968 40547
rect 87916 40504 87968 40513
rect 88284 40547 88336 40556
rect 88284 40513 88303 40547
rect 88303 40513 88336 40547
rect 88284 40504 88336 40513
rect 2908 40368 2960 40420
rect 5954 40230 6006 40282
rect 6018 40230 6070 40282
rect 6082 40230 6134 40282
rect 6146 40230 6198 40282
rect 6210 40230 6262 40282
rect 86546 40230 86598 40282
rect 86610 40230 86662 40282
rect 86674 40230 86726 40282
rect 86738 40230 86790 40282
rect 86802 40230 86854 40282
rect 88284 40096 88336 40148
rect 6690 39686 6742 39738
rect 6754 39686 6806 39738
rect 6818 39686 6870 39738
rect 6882 39686 6934 39738
rect 6946 39686 6998 39738
rect 87282 39686 87334 39738
rect 87346 39686 87398 39738
rect 87410 39686 87462 39738
rect 87474 39686 87526 39738
rect 87538 39686 87590 39738
rect 88284 39493 88336 39502
rect 7140 39416 7192 39468
rect 88284 39459 88303 39493
rect 88303 39459 88336 39493
rect 88284 39450 88336 39459
rect 87180 39348 87232 39400
rect 2908 39280 2960 39332
rect 5954 39142 6006 39194
rect 6018 39142 6070 39194
rect 6082 39142 6134 39194
rect 6146 39142 6198 39194
rect 6210 39142 6262 39194
rect 86546 39142 86598 39194
rect 86610 39142 86662 39194
rect 86674 39142 86726 39194
rect 86738 39142 86790 39194
rect 86802 39142 86854 39194
rect 4380 38940 4432 38992
rect 84420 38940 84472 38992
rect 88284 38881 88336 38890
rect 7784 38804 7836 38856
rect 88284 38847 88303 38881
rect 88303 38847 88336 38881
rect 88284 38838 88336 38847
rect 6690 38598 6742 38650
rect 6754 38598 6806 38650
rect 6818 38598 6870 38650
rect 6882 38598 6934 38650
rect 6946 38598 6998 38650
rect 87282 38598 87334 38650
rect 87346 38598 87398 38650
rect 87410 38598 87462 38650
rect 87474 38598 87526 38650
rect 87538 38598 87590 38650
rect 5954 38054 6006 38106
rect 6018 38054 6070 38106
rect 6082 38054 6134 38106
rect 6146 38054 6198 38106
rect 6210 38054 6262 38106
rect 86546 38054 86598 38106
rect 86610 38054 86662 38106
rect 86674 38054 86726 38106
rect 86738 38054 86790 38106
rect 86802 38054 86854 38106
rect 6690 37510 6742 37562
rect 6754 37510 6806 37562
rect 6818 37510 6870 37562
rect 6882 37510 6934 37562
rect 6946 37510 6998 37562
rect 87282 37510 87334 37562
rect 87346 37510 87398 37562
rect 87410 37510 87462 37562
rect 87474 37510 87526 37562
rect 87538 37510 87590 37562
rect 88284 37317 88336 37326
rect 7232 37240 7284 37292
rect 88284 37283 88299 37317
rect 88299 37283 88336 37317
rect 88284 37274 88336 37283
rect 86352 37172 86404 37224
rect 2908 37104 2960 37156
rect 5954 36966 6006 37018
rect 6018 36966 6070 37018
rect 6082 36966 6134 37018
rect 6146 36966 6198 37018
rect 6210 36966 6262 37018
rect 86546 36966 86598 37018
rect 86610 36966 86662 37018
rect 86674 36966 86726 37018
rect 86738 36966 86790 37018
rect 86802 36966 86854 37018
rect 6690 36422 6742 36474
rect 6754 36422 6806 36474
rect 6818 36422 6870 36474
rect 6882 36422 6934 36474
rect 6946 36422 6998 36474
rect 87282 36422 87334 36474
rect 87346 36422 87398 36474
rect 87410 36422 87462 36474
rect 87474 36422 87526 36474
rect 87538 36422 87590 36474
rect 5668 36186 5720 36238
rect 88560 36152 88612 36204
rect 4380 36084 4432 36136
rect 84420 36084 84472 36136
rect 5954 35878 6006 35930
rect 6018 35878 6070 35930
rect 6082 35878 6134 35930
rect 6146 35878 6198 35930
rect 6210 35878 6262 35930
rect 86546 35878 86598 35930
rect 86610 35878 86662 35930
rect 86674 35878 86726 35930
rect 86738 35878 86790 35930
rect 86802 35878 86854 35930
rect 6690 35334 6742 35386
rect 6754 35334 6806 35386
rect 6818 35334 6870 35386
rect 6882 35334 6934 35386
rect 6946 35334 6998 35386
rect 87282 35334 87334 35386
rect 87346 35334 87398 35386
rect 87410 35334 87462 35386
rect 87474 35334 87526 35386
rect 87538 35334 87590 35386
rect 88284 35141 88336 35150
rect 7232 35064 7284 35116
rect 88284 35107 88299 35141
rect 88299 35107 88336 35141
rect 88284 35098 88336 35107
rect 86352 34996 86404 35048
rect 2908 34928 2960 34980
rect 5954 34790 6006 34842
rect 6018 34790 6070 34842
rect 6082 34790 6134 34842
rect 6146 34790 6198 34842
rect 6210 34790 6262 34842
rect 86546 34790 86598 34842
rect 86610 34790 86662 34842
rect 86674 34790 86726 34842
rect 86738 34790 86790 34842
rect 86802 34790 86854 34842
rect 6690 34246 6742 34298
rect 6754 34246 6806 34298
rect 6818 34246 6870 34298
rect 6882 34246 6934 34298
rect 6946 34246 6998 34298
rect 87282 34246 87334 34298
rect 87346 34246 87398 34298
rect 87410 34246 87462 34298
rect 87474 34246 87526 34298
rect 87538 34246 87590 34298
rect 88284 34053 88336 34062
rect 7232 33976 7284 34028
rect 88284 34019 88299 34053
rect 88299 34019 88336 34053
rect 88284 34010 88336 34019
rect 86352 33908 86404 33960
rect 2908 33840 2960 33892
rect 5954 33702 6006 33754
rect 6018 33702 6070 33754
rect 6082 33702 6134 33754
rect 6146 33702 6198 33754
rect 6210 33702 6262 33754
rect 86546 33702 86598 33754
rect 86610 33702 86662 33754
rect 86674 33702 86726 33754
rect 86738 33702 86790 33754
rect 86802 33702 86854 33754
rect 4380 33500 4432 33552
rect 5668 33398 5720 33450
rect 84420 33364 84472 33416
rect 88560 33364 88612 33416
rect 6690 33158 6742 33210
rect 6754 33158 6806 33210
rect 6818 33158 6870 33210
rect 6882 33158 6934 33210
rect 6946 33158 6998 33210
rect 87282 33158 87334 33210
rect 87346 33158 87398 33210
rect 87410 33158 87462 33210
rect 87474 33158 87526 33210
rect 87538 33158 87590 33210
rect 5954 32614 6006 32666
rect 6018 32614 6070 32666
rect 6082 32614 6134 32666
rect 6146 32614 6198 32666
rect 6210 32614 6262 32666
rect 86546 32614 86598 32666
rect 86610 32614 86662 32666
rect 86674 32614 86726 32666
rect 86738 32614 86790 32666
rect 86802 32614 86854 32666
rect 6690 32070 6742 32122
rect 6754 32070 6806 32122
rect 6818 32070 6870 32122
rect 6882 32070 6934 32122
rect 6946 32070 6998 32122
rect 87282 32070 87334 32122
rect 87346 32070 87398 32122
rect 87410 32070 87462 32122
rect 87474 32070 87526 32122
rect 87538 32070 87590 32122
rect 88284 31877 88336 31886
rect 7232 31800 7284 31852
rect 88284 31843 88299 31877
rect 88299 31843 88336 31877
rect 88284 31834 88336 31843
rect 86352 31732 86404 31784
rect 2908 31664 2960 31716
rect 5954 31526 6006 31578
rect 6018 31526 6070 31578
rect 6082 31526 6134 31578
rect 6146 31526 6198 31578
rect 6210 31526 6262 31578
rect 86546 31526 86598 31578
rect 86610 31526 86662 31578
rect 86674 31526 86726 31578
rect 86738 31526 86790 31578
rect 86802 31526 86854 31578
rect 6690 30982 6742 31034
rect 6754 30982 6806 31034
rect 6818 30982 6870 31034
rect 6882 30982 6934 31034
rect 6946 30982 6998 31034
rect 87282 30982 87334 31034
rect 87346 30982 87398 31034
rect 87410 30982 87462 31034
rect 87474 30982 87526 31034
rect 87538 30982 87590 31034
rect 5668 30746 5720 30798
rect 88560 30712 88612 30764
rect 4380 30576 4432 30628
rect 84420 30576 84472 30628
rect 5954 30438 6006 30490
rect 6018 30438 6070 30490
rect 6082 30438 6134 30490
rect 6146 30438 6198 30490
rect 6210 30438 6262 30490
rect 86546 30438 86598 30490
rect 86610 30438 86662 30490
rect 86674 30438 86726 30490
rect 86738 30438 86790 30490
rect 86802 30438 86854 30490
rect 6690 29894 6742 29946
rect 6754 29894 6806 29946
rect 6818 29894 6870 29946
rect 6882 29894 6934 29946
rect 6946 29894 6998 29946
rect 87282 29894 87334 29946
rect 87346 29894 87398 29946
rect 87410 29894 87462 29946
rect 87474 29894 87526 29946
rect 87538 29894 87590 29946
rect 2908 29624 2960 29676
rect 86352 29624 86404 29676
rect 7232 29556 7284 29608
rect 88284 29488 88336 29540
rect 5954 29350 6006 29402
rect 6018 29350 6070 29402
rect 6082 29350 6134 29402
rect 6146 29350 6198 29402
rect 6210 29350 6262 29402
rect 86546 29350 86598 29402
rect 86610 29350 86662 29402
rect 86674 29350 86726 29402
rect 86738 29350 86790 29402
rect 86802 29350 86854 29402
rect 6690 28806 6742 28858
rect 6754 28806 6806 28858
rect 6818 28806 6870 28858
rect 6882 28806 6934 28858
rect 6946 28806 6998 28858
rect 87282 28806 87334 28858
rect 87346 28806 87398 28858
rect 87410 28806 87462 28858
rect 87474 28806 87526 28858
rect 87538 28806 87590 28858
rect 2908 28536 2960 28588
rect 86352 28536 86404 28588
rect 7232 28468 7284 28520
rect 88192 28443 88244 28452
rect 88192 28409 88215 28443
rect 88215 28409 88244 28443
rect 88192 28400 88244 28409
rect 5954 28262 6006 28314
rect 6018 28262 6070 28314
rect 6082 28262 6134 28314
rect 6146 28262 6198 28314
rect 6210 28262 6262 28314
rect 86546 28262 86598 28314
rect 86610 28262 86662 28314
rect 86674 28262 86726 28314
rect 86738 28262 86790 28314
rect 86802 28262 86854 28314
rect 5116 28060 5168 28112
rect 85248 27924 85300 27976
rect 5392 27899 5444 27908
rect 5392 27865 5411 27899
rect 5411 27865 5444 27899
rect 5392 27856 5444 27865
rect 88928 27856 88980 27908
rect 6690 27718 6742 27770
rect 6754 27718 6806 27770
rect 6818 27718 6870 27770
rect 6882 27718 6934 27770
rect 6946 27718 6998 27770
rect 87282 27718 87334 27770
rect 87346 27718 87398 27770
rect 87410 27718 87462 27770
rect 87474 27718 87526 27770
rect 87538 27718 87590 27770
rect 5954 27174 6006 27226
rect 6018 27174 6070 27226
rect 6082 27174 6134 27226
rect 6146 27174 6198 27226
rect 6210 27174 6262 27226
rect 86546 27174 86598 27226
rect 86610 27174 86662 27226
rect 86674 27174 86726 27226
rect 86738 27174 86790 27226
rect 86802 27174 86854 27226
rect 6690 26630 6742 26682
rect 6754 26630 6806 26682
rect 6818 26630 6870 26682
rect 6882 26630 6934 26682
rect 6946 26630 6998 26682
rect 87282 26630 87334 26682
rect 87346 26630 87398 26682
rect 87410 26630 87462 26682
rect 87474 26630 87526 26682
rect 87538 26630 87590 26682
rect 2908 26360 2960 26412
rect 87732 26394 87784 26446
rect 7140 26292 7192 26344
rect 88192 26267 88244 26276
rect 88192 26233 88215 26267
rect 88215 26233 88244 26267
rect 88192 26224 88244 26233
rect 5954 26086 6006 26138
rect 6018 26086 6070 26138
rect 6082 26086 6134 26138
rect 6146 26086 6198 26138
rect 6210 26086 6262 26138
rect 86546 26086 86598 26138
rect 86610 26086 86662 26138
rect 86674 26086 86726 26138
rect 86738 26086 86790 26138
rect 86802 26086 86854 26138
rect 6690 25542 6742 25594
rect 6754 25542 6806 25594
rect 6818 25542 6870 25594
rect 6882 25542 6934 25594
rect 6946 25542 6998 25594
rect 87282 25542 87334 25594
rect 87346 25542 87398 25594
rect 87410 25542 87462 25594
rect 87474 25542 87526 25594
rect 87538 25542 87590 25594
rect 4932 25306 4984 25358
rect 87732 25306 87784 25358
rect 7140 25204 7192 25256
rect 88560 25136 88612 25188
rect 5954 24998 6006 25050
rect 6018 24998 6070 25050
rect 6082 24998 6134 25050
rect 6146 24998 6198 25050
rect 6210 24998 6262 25050
rect 86546 24998 86598 25050
rect 86610 24998 86662 25050
rect 86674 24998 86726 25050
rect 86738 24998 86790 25050
rect 86802 24998 86854 25050
rect 6690 24454 6742 24506
rect 6754 24454 6806 24506
rect 6818 24454 6870 24506
rect 6882 24454 6934 24506
rect 6946 24454 6998 24506
rect 87282 24454 87334 24506
rect 87346 24454 87398 24506
rect 87410 24454 87462 24506
rect 87474 24454 87526 24506
rect 87538 24454 87590 24506
rect 2908 24184 2960 24236
rect 87732 24218 87784 24270
rect 7140 24116 7192 24168
rect 88284 24048 88336 24100
rect 5954 23910 6006 23962
rect 6018 23910 6070 23962
rect 6082 23910 6134 23962
rect 6146 23910 6198 23962
rect 6210 23910 6262 23962
rect 86546 23910 86598 23962
rect 86610 23910 86662 23962
rect 86674 23910 86726 23962
rect 86738 23910 86790 23962
rect 86802 23910 86854 23962
rect 6690 23366 6742 23418
rect 6754 23366 6806 23418
rect 6818 23366 6870 23418
rect 6882 23366 6934 23418
rect 6946 23366 6998 23418
rect 87282 23366 87334 23418
rect 87346 23366 87398 23418
rect 87410 23366 87462 23418
rect 87474 23366 87526 23418
rect 87538 23366 87590 23418
rect 2908 23096 2960 23148
rect 86352 23096 86404 23148
rect 7140 23028 7192 23080
rect 88284 22960 88336 23012
rect 5954 22822 6006 22874
rect 6018 22822 6070 22874
rect 6082 22822 6134 22874
rect 6146 22822 6198 22874
rect 6210 22822 6262 22874
rect 86546 22822 86598 22874
rect 86610 22822 86662 22874
rect 86674 22822 86726 22874
rect 86738 22822 86790 22874
rect 86802 22822 86854 22874
rect 4932 22518 4984 22570
rect 9164 22484 9216 22536
rect 84420 22484 84472 22536
rect 88560 22416 88612 22468
rect 6690 22278 6742 22330
rect 6754 22278 6806 22330
rect 6818 22278 6870 22330
rect 6882 22278 6934 22330
rect 6946 22278 6998 22330
rect 87282 22278 87334 22330
rect 87346 22278 87398 22330
rect 87410 22278 87462 22330
rect 87474 22278 87526 22330
rect 87538 22278 87590 22330
rect 5954 21734 6006 21786
rect 6018 21734 6070 21786
rect 6082 21734 6134 21786
rect 6146 21734 6198 21786
rect 6210 21734 6262 21786
rect 86546 21734 86598 21786
rect 86610 21734 86662 21786
rect 86674 21734 86726 21786
rect 86738 21734 86790 21786
rect 86802 21734 86854 21786
rect 6690 21190 6742 21242
rect 6754 21190 6806 21242
rect 6818 21190 6870 21242
rect 6882 21190 6934 21242
rect 6946 21190 6998 21242
rect 87282 21190 87334 21242
rect 87346 21190 87398 21242
rect 87410 21190 87462 21242
rect 87474 21190 87526 21242
rect 87538 21190 87590 21242
rect 9256 21056 9308 21108
rect 5208 20997 5260 21006
rect 5208 20963 5217 20997
rect 5217 20963 5251 20997
rect 5251 20963 5260 20997
rect 5208 20954 5260 20963
rect 84420 20920 84472 20972
rect 88560 20920 88612 20972
rect 5954 20646 6006 20698
rect 6018 20646 6070 20698
rect 6082 20646 6134 20698
rect 6146 20646 6198 20698
rect 6210 20646 6262 20698
rect 86546 20646 86598 20698
rect 86610 20646 86662 20698
rect 86674 20646 86726 20698
rect 86738 20646 86790 20698
rect 86802 20646 86854 20698
rect 6690 20102 6742 20154
rect 6754 20102 6806 20154
rect 6818 20102 6870 20154
rect 6882 20102 6934 20154
rect 6946 20102 6998 20154
rect 87282 20102 87334 20154
rect 87346 20102 87398 20154
rect 87410 20102 87462 20154
rect 87474 20102 87526 20154
rect 87538 20102 87590 20154
rect 4932 19866 4984 19918
rect 87732 19866 87784 19918
rect 7140 19764 7192 19816
rect 88560 19696 88612 19748
rect 5954 19558 6006 19610
rect 6018 19558 6070 19610
rect 6082 19558 6134 19610
rect 6146 19558 6198 19610
rect 6210 19558 6262 19610
rect 86546 19558 86598 19610
rect 86610 19558 86662 19610
rect 86674 19558 86726 19610
rect 86738 19558 86790 19610
rect 86802 19558 86854 19610
rect 6690 19014 6742 19066
rect 6754 19014 6806 19066
rect 6818 19014 6870 19066
rect 6882 19014 6934 19066
rect 6946 19014 6998 19066
rect 87282 19014 87334 19066
rect 87346 19014 87398 19066
rect 87410 19014 87462 19066
rect 87474 19014 87526 19066
rect 87538 19014 87590 19066
rect 2908 18744 2960 18796
rect 87732 18778 87784 18830
rect 7140 18676 7192 18728
rect 88284 18608 88336 18660
rect 5954 18470 6006 18522
rect 6018 18470 6070 18522
rect 6082 18470 6134 18522
rect 6146 18470 6198 18522
rect 6210 18470 6262 18522
rect 86546 18470 86598 18522
rect 86610 18470 86662 18522
rect 86674 18470 86726 18522
rect 86738 18470 86790 18522
rect 86802 18470 86854 18522
rect 6690 17926 6742 17978
rect 6754 17926 6806 17978
rect 6818 17926 6870 17978
rect 6882 17926 6934 17978
rect 6946 17926 6998 17978
rect 87282 17926 87334 17978
rect 87346 17926 87398 17978
rect 87410 17926 87462 17978
rect 87474 17926 87526 17978
rect 87538 17926 87590 17978
rect 2908 17656 2960 17708
rect 86352 17656 86404 17708
rect 7232 17588 7284 17640
rect 88192 17563 88244 17572
rect 88192 17529 88215 17563
rect 88215 17529 88244 17563
rect 88192 17520 88244 17529
rect 5954 17382 6006 17434
rect 6018 17382 6070 17434
rect 6082 17382 6134 17434
rect 6146 17382 6198 17434
rect 6210 17382 6262 17434
rect 86546 17382 86598 17434
rect 86610 17382 86662 17434
rect 86674 17382 86726 17434
rect 86738 17382 86790 17434
rect 86802 17382 86854 17434
rect 5208 17121 5260 17130
rect 5208 17087 5217 17121
rect 5217 17087 5251 17121
rect 5251 17087 5260 17121
rect 5208 17078 5260 17087
rect 88008 17121 88060 17130
rect 88008 17087 88017 17121
rect 88017 17087 88051 17121
rect 88051 17087 88060 17121
rect 88008 17078 88060 17087
rect 5392 17019 5444 17028
rect 5392 16985 5411 17019
rect 5411 16985 5444 17019
rect 5392 16976 5444 16985
rect 88560 16976 88612 17028
rect 6690 16838 6742 16890
rect 6754 16838 6806 16890
rect 6818 16838 6870 16890
rect 6882 16838 6934 16890
rect 6946 16838 6998 16890
rect 87282 16838 87334 16890
rect 87346 16838 87398 16890
rect 87410 16838 87462 16890
rect 87474 16838 87526 16890
rect 87538 16838 87590 16890
rect 5954 16294 6006 16346
rect 6018 16294 6070 16346
rect 6082 16294 6134 16346
rect 6146 16294 6198 16346
rect 6210 16294 6262 16346
rect 86546 16294 86598 16346
rect 86610 16294 86662 16346
rect 86674 16294 86726 16346
rect 86738 16294 86790 16346
rect 86802 16294 86854 16346
rect 6690 15750 6742 15802
rect 6754 15750 6806 15802
rect 6818 15750 6870 15802
rect 6882 15750 6934 15802
rect 6946 15750 6998 15802
rect 87282 15750 87334 15802
rect 87346 15750 87398 15802
rect 87410 15750 87462 15802
rect 87474 15750 87526 15802
rect 87538 15750 87590 15802
rect 5208 15557 5260 15566
rect 5208 15523 5217 15557
rect 5217 15523 5251 15557
rect 5251 15523 5260 15557
rect 5208 15514 5260 15523
rect 84420 15480 84472 15532
rect 5668 15412 5720 15464
rect 88560 15412 88612 15464
rect 5954 15206 6006 15258
rect 6018 15206 6070 15258
rect 6082 15206 6134 15258
rect 6146 15206 6198 15258
rect 6210 15206 6262 15258
rect 86546 15206 86598 15258
rect 86610 15206 86662 15258
rect 86674 15206 86726 15258
rect 86738 15206 86790 15258
rect 86802 15206 86854 15258
rect 85432 14936 85484 14988
rect 85616 14936 85668 14988
rect 88008 14843 88060 14852
rect 88008 14809 88017 14843
rect 88017 14809 88051 14843
rect 88051 14809 88060 14843
rect 88008 14800 88060 14809
rect 6690 14662 6742 14714
rect 6754 14662 6806 14714
rect 6818 14662 6870 14714
rect 6882 14662 6934 14714
rect 6946 14662 6998 14714
rect 87282 14662 87334 14714
rect 87346 14662 87398 14714
rect 87410 14662 87462 14714
rect 87474 14662 87526 14714
rect 87538 14662 87590 14714
rect 83684 14256 83736 14308
rect 85616 14299 85668 14308
rect 85616 14265 85625 14299
rect 85625 14265 85659 14299
rect 85659 14265 85668 14299
rect 85616 14256 85668 14265
rect 5954 14118 6006 14170
rect 6018 14118 6070 14170
rect 6082 14118 6134 14170
rect 6146 14118 6198 14170
rect 6210 14118 6262 14170
rect 86546 14118 86598 14170
rect 86610 14118 86662 14170
rect 86674 14118 86726 14170
rect 86738 14118 86790 14170
rect 86802 14118 86854 14170
rect 6690 13574 6742 13626
rect 6754 13574 6806 13626
rect 6818 13574 6870 13626
rect 6882 13574 6934 13626
rect 6946 13574 6998 13626
rect 87282 13574 87334 13626
rect 87346 13574 87398 13626
rect 87410 13574 87462 13626
rect 87474 13574 87526 13626
rect 87538 13574 87590 13626
rect 83500 13440 83552 13492
rect 85524 13440 85576 13492
rect 88192 13381 88244 13390
rect 87916 13347 87968 13356
rect 87916 13313 87925 13347
rect 87925 13313 87959 13347
rect 87959 13313 87968 13347
rect 87916 13304 87968 13313
rect 88192 13347 88226 13381
rect 88226 13347 88244 13381
rect 88192 13338 88244 13347
rect 5954 13030 6006 13082
rect 6018 13030 6070 13082
rect 6082 13030 6134 13082
rect 6146 13030 6198 13082
rect 6210 13030 6262 13082
rect 86546 13030 86598 13082
rect 86610 13030 86662 13082
rect 86674 13030 86726 13082
rect 86738 13030 86790 13082
rect 86802 13030 86854 13082
rect 87916 12896 87968 12948
rect 87180 12692 87232 12744
rect 88560 12692 88612 12744
rect 6690 12486 6742 12538
rect 6754 12486 6806 12538
rect 6818 12486 6870 12538
rect 6882 12486 6934 12538
rect 6946 12486 6998 12538
rect 87282 12486 87334 12538
rect 87346 12486 87398 12538
rect 87410 12486 87462 12538
rect 87474 12486 87526 12538
rect 87538 12486 87590 12538
rect 83500 12352 83552 12404
rect 85340 12352 85392 12404
rect 87180 12352 87232 12404
rect 5954 11942 6006 11994
rect 6018 11942 6070 11994
rect 6082 11942 6134 11994
rect 6146 11942 6198 11994
rect 6210 11942 6262 11994
rect 86546 11942 86598 11994
rect 86610 11942 86662 11994
rect 86674 11942 86726 11994
rect 86738 11942 86790 11994
rect 86802 11942 86854 11994
rect 83408 11740 83460 11792
rect 83684 11740 83736 11792
rect 6690 11398 6742 11450
rect 6754 11398 6806 11450
rect 6818 11398 6870 11450
rect 6882 11398 6934 11450
rect 6946 11398 6998 11450
rect 87282 11398 87334 11450
rect 87346 11398 87398 11450
rect 87410 11398 87462 11450
rect 87474 11398 87526 11450
rect 87538 11398 87590 11450
rect 83316 11196 83368 11248
rect 5954 10854 6006 10906
rect 6018 10854 6070 10906
rect 6082 10854 6134 10906
rect 6146 10854 6198 10906
rect 6210 10854 6262 10906
rect 86546 10854 86598 10906
rect 86610 10854 86662 10906
rect 86674 10854 86726 10906
rect 86738 10854 86790 10906
rect 86802 10854 86854 10906
rect 88376 10524 88428 10576
rect 6690 10310 6742 10362
rect 6754 10310 6806 10362
rect 6818 10310 6870 10362
rect 6882 10310 6934 10362
rect 6946 10310 6998 10362
rect 87282 10310 87334 10362
rect 87346 10310 87398 10362
rect 87410 10310 87462 10362
rect 87474 10310 87526 10362
rect 87538 10310 87590 10362
rect 45596 10176 45648 10228
rect 46056 10176 46108 10228
rect 82488 10176 82540 10228
rect 88560 10040 88612 10092
rect 81384 9972 81436 10024
rect 5954 9766 6006 9818
rect 6018 9766 6070 9818
rect 6082 9766 6134 9818
rect 6146 9766 6198 9818
rect 6210 9766 6262 9818
rect 86546 9766 86598 9818
rect 86610 9766 86662 9818
rect 86674 9766 86726 9818
rect 86738 9766 86790 9818
rect 86802 9766 86854 9818
rect 6690 9222 6742 9274
rect 6754 9222 6806 9274
rect 6818 9222 6870 9274
rect 6882 9222 6934 9274
rect 6946 9222 6998 9274
rect 87282 9222 87334 9274
rect 87346 9222 87398 9274
rect 87410 9222 87462 9274
rect 87474 9222 87526 9274
rect 87538 9222 87590 9274
rect 5954 8678 6006 8730
rect 6018 8678 6070 8730
rect 6082 8678 6134 8730
rect 6146 8678 6198 8730
rect 6210 8678 6262 8730
rect 86546 8678 86598 8730
rect 86610 8678 86662 8730
rect 86674 8678 86726 8730
rect 86738 8678 86790 8730
rect 86802 8678 86854 8730
rect 6690 8134 6742 8186
rect 6754 8134 6806 8186
rect 6818 8134 6870 8186
rect 6882 8134 6934 8186
rect 6946 8134 6998 8186
rect 87282 8134 87334 8186
rect 87346 8134 87398 8186
rect 87410 8134 87462 8186
rect 87474 8134 87526 8186
rect 87538 8134 87590 8186
rect 5954 7590 6006 7642
rect 6018 7590 6070 7642
rect 6082 7590 6134 7642
rect 6146 7590 6198 7642
rect 6210 7590 6262 7642
rect 17722 7590 17774 7642
rect 17786 7590 17838 7642
rect 17850 7590 17902 7642
rect 17914 7590 17966 7642
rect 17978 7590 18030 7642
rect 36122 7590 36174 7642
rect 36186 7590 36238 7642
rect 36250 7590 36302 7642
rect 36314 7590 36366 7642
rect 36378 7590 36430 7642
rect 54522 7590 54574 7642
rect 54586 7590 54638 7642
rect 54650 7590 54702 7642
rect 54714 7590 54766 7642
rect 54778 7590 54830 7642
rect 72922 7590 72974 7642
rect 72986 7590 73038 7642
rect 73050 7590 73102 7642
rect 73114 7590 73166 7642
rect 73178 7590 73230 7642
rect 86546 7590 86598 7642
rect 86610 7590 86662 7642
rect 86674 7590 86726 7642
rect 86738 7590 86790 7642
rect 86802 7590 86854 7642
rect 45688 7456 45740 7508
rect 45964 7499 46016 7508
rect 45964 7465 45973 7499
rect 45973 7465 46007 7499
rect 46007 7465 46016 7499
rect 45964 7456 46016 7465
rect 45596 7431 45648 7440
rect 45596 7397 45605 7431
rect 45605 7397 45639 7431
rect 45639 7397 45648 7431
rect 45596 7388 45648 7397
rect 46056 7388 46108 7440
rect 83500 7320 83552 7372
rect 45964 7252 46016 7304
rect 83408 7252 83460 7304
rect 45596 7184 45648 7236
rect 83592 7184 83644 7236
rect 6690 7046 6742 7098
rect 6754 7046 6806 7098
rect 6818 7046 6870 7098
rect 6882 7046 6934 7098
rect 6946 7046 6998 7098
rect 18382 7046 18434 7098
rect 18446 7046 18498 7098
rect 18510 7046 18562 7098
rect 18574 7046 18626 7098
rect 18638 7046 18690 7098
rect 36782 7046 36834 7098
rect 36846 7046 36898 7098
rect 36910 7046 36962 7098
rect 36974 7046 37026 7098
rect 37038 7046 37090 7098
rect 55182 7046 55234 7098
rect 55246 7046 55298 7098
rect 55310 7046 55362 7098
rect 55374 7046 55426 7098
rect 55438 7046 55490 7098
rect 73582 7046 73634 7098
rect 73646 7046 73698 7098
rect 73710 7046 73762 7098
rect 73774 7046 73826 7098
rect 73838 7046 73890 7098
rect 87282 7046 87334 7098
rect 87346 7046 87398 7098
rect 87410 7046 87462 7098
rect 87474 7046 87526 7098
rect 87538 7046 87590 7098
rect 17722 6502 17774 6554
rect 17786 6502 17838 6554
rect 17850 6502 17902 6554
rect 17914 6502 17966 6554
rect 17978 6502 18030 6554
rect 36122 6502 36174 6554
rect 36186 6502 36238 6554
rect 36250 6502 36302 6554
rect 36314 6502 36366 6554
rect 36378 6502 36430 6554
rect 54522 6502 54574 6554
rect 54586 6502 54638 6554
rect 54650 6502 54702 6554
rect 54714 6502 54766 6554
rect 54778 6502 54830 6554
rect 72922 6502 72974 6554
rect 72986 6502 73038 6554
rect 73050 6502 73102 6554
rect 73114 6502 73166 6554
rect 73178 6502 73230 6554
rect 18382 5958 18434 6010
rect 18446 5958 18498 6010
rect 18510 5958 18562 6010
rect 18574 5958 18626 6010
rect 18638 5958 18690 6010
rect 36782 5958 36834 6010
rect 36846 5958 36898 6010
rect 36910 5958 36962 6010
rect 36974 5958 37026 6010
rect 37038 5958 37090 6010
rect 55182 5958 55234 6010
rect 55246 5958 55298 6010
rect 55310 5958 55362 6010
rect 55374 5958 55426 6010
rect 55438 5958 55490 6010
rect 73582 5958 73634 6010
rect 73646 5958 73698 6010
rect 73710 5958 73762 6010
rect 73774 5958 73826 6010
rect 73838 5958 73890 6010
rect 17722 5414 17774 5466
rect 17786 5414 17838 5466
rect 17850 5414 17902 5466
rect 17914 5414 17966 5466
rect 17978 5414 18030 5466
rect 36122 5414 36174 5466
rect 36186 5414 36238 5466
rect 36250 5414 36302 5466
rect 36314 5414 36366 5466
rect 36378 5414 36430 5466
rect 54522 5414 54574 5466
rect 54586 5414 54638 5466
rect 54650 5414 54702 5466
rect 54714 5414 54766 5466
rect 54778 5414 54830 5466
rect 72922 5414 72974 5466
rect 72986 5414 73038 5466
rect 73050 5414 73102 5466
rect 73114 5414 73166 5466
rect 73178 5414 73230 5466
rect 30692 5280 30744 5332
rect 31520 5323 31572 5332
rect 31520 5289 31538 5323
rect 31538 5289 31572 5323
rect 31520 5280 31572 5289
rect 33820 5280 33872 5332
rect 35108 5280 35160 5332
rect 35936 5280 35988 5332
rect 37132 5280 37184 5332
rect 38420 5280 38472 5332
rect 39248 5323 39300 5332
rect 39248 5289 39266 5323
rect 39266 5289 39300 5323
rect 39248 5280 39300 5289
rect 41640 5280 41692 5332
rect 42836 5280 42888 5332
rect 43664 5280 43716 5332
rect 44768 5280 44820 5332
rect 67860 5280 67912 5332
rect 69332 5280 69384 5332
rect 71172 5280 71224 5332
rect 72276 5280 72328 5332
rect 73380 5323 73432 5332
rect 73380 5289 73399 5323
rect 73399 5289 73432 5323
rect 73380 5280 73432 5289
rect 74484 5280 74536 5332
rect 75588 5280 75640 5332
rect 76692 5280 76744 5332
rect 78900 5280 78952 5332
rect 80280 5280 80332 5332
rect 32716 5212 32768 5264
rect 40444 5212 40496 5264
rect 70068 5212 70120 5264
rect 77796 5212 77848 5264
rect 15236 5110 15288 5162
rect 16064 5153 16116 5162
rect 16064 5119 16104 5153
rect 16104 5119 16116 5153
rect 16064 5110 16116 5119
rect 17168 5153 17220 5162
rect 17168 5119 17177 5153
rect 17177 5119 17211 5153
rect 17211 5119 17220 5153
rect 17168 5110 17220 5119
rect 18272 5110 18324 5162
rect 19652 5110 19704 5162
rect 20480 5153 20532 5162
rect 20480 5119 20489 5153
rect 20489 5119 20523 5153
rect 20523 5119 20532 5153
rect 20480 5110 20532 5119
rect 21584 5110 21636 5162
rect 22964 5110 23016 5162
rect 23792 5153 23844 5162
rect 23792 5119 23832 5153
rect 23832 5119 23844 5153
rect 23792 5110 23844 5119
rect 24896 5153 24948 5162
rect 24896 5119 24905 5153
rect 24905 5119 24939 5153
rect 24939 5119 24948 5153
rect 24896 5110 24948 5119
rect 26092 5110 26144 5162
rect 27380 5110 27432 5162
rect 28208 5153 28260 5162
rect 28208 5119 28217 5153
rect 28217 5119 28251 5153
rect 28251 5119 28260 5153
rect 28208 5110 28260 5119
rect 29312 5110 29364 5162
rect 35752 5076 35804 5128
rect 43480 5076 43532 5128
rect 52404 5110 52456 5162
rect 53692 5110 53744 5162
rect 54888 5110 54940 5162
rect 55716 5110 55768 5162
rect 56820 5110 56872 5162
rect 57924 5153 57976 5162
rect 57924 5119 57964 5153
rect 57964 5119 57976 5153
rect 57924 5110 57976 5119
rect 59028 5110 59080 5162
rect 60132 5110 60184 5162
rect 61420 5110 61472 5162
rect 62340 5110 62392 5162
rect 63444 5110 63496 5162
rect 64548 5110 64600 5162
rect 65652 5153 65704 5162
rect 65652 5119 65692 5153
rect 65692 5119 65704 5153
rect 65652 5110 65704 5119
rect 66756 5110 66808 5162
rect 69240 5076 69292 5128
rect 69884 5110 69936 5162
rect 74392 5076 74444 5128
rect 76968 5076 77020 5128
rect 77612 5110 77664 5162
rect 15144 5008 15196 5060
rect 15788 5008 15840 5060
rect 17076 5008 17128 5060
rect 18272 5008 18324 5060
rect 19652 5008 19704 5060
rect 20296 5008 20348 5060
rect 21584 5008 21636 5060
rect 22872 5008 22924 5060
rect 23516 5008 23568 5060
rect 24804 5008 24856 5060
rect 26092 5008 26144 5060
rect 27380 5008 27432 5060
rect 28024 5008 28076 5060
rect 29312 5008 29364 5060
rect 30600 5008 30652 5060
rect 31244 5008 31296 5060
rect 32532 5008 32584 5060
rect 33820 5008 33872 5060
rect 35108 5008 35160 5060
rect 37132 5008 37184 5060
rect 38328 5008 38380 5060
rect 38972 5008 39024 5060
rect 40260 5008 40312 5060
rect 41548 5008 41600 5060
rect 42836 5008 42888 5060
rect 44768 5008 44820 5060
rect 52496 5008 52548 5060
rect 53784 5008 53836 5060
rect 54428 5008 54480 5060
rect 55716 5008 55768 5060
rect 57004 5008 57056 5060
rect 57648 5008 57700 5060
rect 58936 5008 58988 5060
rect 60224 5008 60276 5060
rect 61512 5008 61564 5060
rect 62156 5008 62208 5060
rect 63444 5008 63496 5060
rect 64732 5008 64784 5060
rect 65376 5008 65428 5060
rect 66664 5008 66716 5060
rect 67952 5008 68004 5060
rect 71172 5008 71224 5060
rect 72460 5008 72512 5060
rect 73104 5008 73156 5060
rect 75680 5008 75732 5060
rect 78900 5008 78952 5060
rect 80188 5008 80240 5060
rect 18382 4870 18434 4922
rect 18446 4870 18498 4922
rect 18510 4870 18562 4922
rect 18574 4870 18626 4922
rect 18638 4870 18690 4922
rect 36782 4870 36834 4922
rect 36846 4870 36898 4922
rect 36910 4870 36962 4922
rect 36974 4870 37026 4922
rect 37038 4870 37090 4922
rect 55182 4870 55234 4922
rect 55246 4870 55298 4922
rect 55310 4870 55362 4922
rect 55374 4870 55426 4922
rect 55438 4870 55490 4922
rect 73582 4870 73634 4922
rect 73646 4870 73698 4922
rect 73710 4870 73762 4922
rect 73774 4870 73826 4922
rect 73838 4870 73890 4922
<< metal2 >>
rect 10634 88000 10690 88800
rect 15142 88000 15198 88800
rect 15786 88000 15842 88800
rect 17074 88000 17130 88800
rect 18362 88000 18418 88800
rect 19650 88000 19706 88800
rect 20294 88000 20350 88800
rect 21582 88000 21638 88800
rect 22870 88000 22926 88800
rect 23514 88000 23570 88800
rect 24802 88000 24858 88800
rect 26090 88000 26146 88800
rect 27378 88000 27434 88800
rect 28022 88000 28078 88800
rect 29310 88000 29366 88800
rect 30598 88000 30654 88800
rect 31242 88000 31298 88800
rect 32530 88000 32586 88800
rect 33818 88000 33874 88800
rect 35106 88000 35162 88800
rect 35750 88000 35806 88800
rect 37038 88000 37094 88800
rect 37682 88000 37738 88800
rect 38326 88000 38382 88800
rect 38970 88000 39026 88800
rect 39614 88000 39670 88800
rect 40258 88000 40314 88800
rect 40902 88000 40958 88800
rect 41546 88000 41602 88800
rect 42190 88000 42246 88800
rect 42834 88000 42890 88800
rect 43478 88000 43534 88800
rect 44122 88000 44178 88800
rect 44766 88000 44822 88800
rect 45410 88000 45466 88800
rect 46054 88000 46110 88800
rect 46698 88000 46754 88800
rect 47342 88000 47398 88800
rect 47986 88000 48042 88800
rect 48630 88000 48686 88800
rect 49274 88000 49330 88800
rect 49918 88000 49974 88800
rect 50562 88000 50618 88800
rect 52494 88000 52550 88800
rect 53782 88000 53838 88800
rect 54426 88000 54482 88800
rect 55714 88000 55770 88800
rect 57002 88000 57058 88800
rect 57646 88000 57702 88800
rect 58934 88000 58990 88800
rect 60222 88000 60278 88800
rect 61510 88000 61566 88800
rect 62154 88000 62210 88800
rect 63442 88000 63498 88800
rect 64730 88000 64786 88800
rect 65374 88000 65430 88800
rect 66662 88000 66718 88800
rect 67950 88000 68006 88800
rect 69238 88000 69294 88800
rect 69882 88000 69938 88800
rect 71170 88000 71226 88800
rect 72458 88000 72514 88800
rect 73102 88000 73158 88800
rect 74390 88000 74446 88800
rect 75678 88000 75734 88800
rect 76966 88000 77022 88800
rect 77610 88000 77666 88800
rect 78898 88000 78954 88800
rect 80186 88000 80242 88800
rect 80830 88000 80886 88800
rect 82118 88000 82174 88800
rect 10648 87482 10676 88000
rect 15156 87482 15184 88000
rect 10636 87476 10688 87482
rect 10636 87418 10688 87424
rect 15144 87476 15196 87482
rect 15144 87418 15196 87424
rect 15800 87414 15828 88000
rect 17088 87482 17116 88000
rect 18376 87770 18404 88000
rect 18284 87742 18404 87770
rect 18284 87482 18312 87742
rect 18382 87612 18690 87621
rect 18382 87610 18388 87612
rect 18444 87610 18468 87612
rect 18524 87610 18548 87612
rect 18604 87610 18628 87612
rect 18684 87610 18690 87612
rect 18444 87558 18446 87610
rect 18626 87558 18628 87610
rect 18382 87556 18388 87558
rect 18444 87556 18468 87558
rect 18524 87556 18548 87558
rect 18604 87556 18628 87558
rect 18684 87556 18690 87558
rect 18382 87547 18690 87556
rect 19664 87482 19692 88000
rect 17076 87476 17128 87482
rect 17076 87418 17128 87424
rect 18272 87476 18324 87482
rect 18272 87418 18324 87424
rect 19652 87476 19704 87482
rect 19652 87418 19704 87424
rect 20308 87414 20336 88000
rect 21596 87482 21624 88000
rect 22884 87482 22912 88000
rect 23528 87482 23556 88000
rect 24816 87482 24844 88000
rect 26104 87482 26132 88000
rect 27392 87482 27420 88000
rect 21584 87476 21636 87482
rect 21584 87418 21636 87424
rect 22872 87476 22924 87482
rect 22872 87418 22924 87424
rect 23516 87476 23568 87482
rect 23516 87418 23568 87424
rect 24804 87476 24856 87482
rect 24804 87418 24856 87424
rect 26092 87476 26144 87482
rect 26092 87418 26144 87424
rect 27380 87476 27432 87482
rect 27380 87418 27432 87424
rect 28036 87414 28064 88000
rect 29324 87482 29352 88000
rect 30612 87482 30640 88000
rect 31256 87482 31284 88000
rect 32544 87482 32572 88000
rect 33832 87482 33860 88000
rect 35120 87482 35148 88000
rect 35764 87482 35792 88000
rect 37052 87770 37080 88000
rect 37052 87742 37172 87770
rect 36782 87612 37090 87621
rect 36782 87610 36788 87612
rect 36844 87610 36868 87612
rect 36924 87610 36948 87612
rect 37004 87610 37028 87612
rect 37084 87610 37090 87612
rect 36844 87558 36846 87610
rect 37026 87558 37028 87610
rect 36782 87556 36788 87558
rect 36844 87556 36868 87558
rect 36924 87556 36948 87558
rect 37004 87556 37028 87558
rect 37084 87556 37090 87558
rect 36782 87547 37090 87556
rect 37144 87482 37172 87742
rect 37696 87482 37724 88000
rect 38340 87482 38368 88000
rect 38984 87482 39012 88000
rect 29312 87476 29364 87482
rect 29312 87418 29364 87424
rect 30600 87476 30652 87482
rect 30600 87418 30652 87424
rect 31244 87476 31296 87482
rect 31244 87418 31296 87424
rect 32532 87476 32584 87482
rect 32532 87418 32584 87424
rect 33820 87476 33872 87482
rect 33820 87418 33872 87424
rect 35108 87476 35160 87482
rect 35108 87418 35160 87424
rect 35752 87476 35804 87482
rect 35752 87418 35804 87424
rect 37132 87476 37184 87482
rect 37132 87418 37184 87424
rect 37684 87476 37736 87482
rect 37684 87418 37736 87424
rect 38328 87476 38380 87482
rect 38328 87418 38380 87424
rect 38972 87476 39024 87482
rect 38972 87418 39024 87424
rect 15788 87408 15840 87414
rect 10726 87376 10782 87385
rect 15788 87350 15840 87356
rect 20296 87408 20348 87414
rect 20296 87350 20348 87356
rect 28024 87408 28076 87414
rect 28024 87350 28076 87356
rect 30600 87374 30652 87380
rect 10726 87311 10782 87320
rect 18272 87340 18324 87346
rect 18272 87282 18324 87288
rect 19560 87340 19612 87346
rect 30600 87316 30652 87322
rect 31520 87374 31572 87380
rect 31520 87316 31572 87322
rect 32624 87374 32676 87380
rect 32624 87316 32676 87322
rect 33728 87374 33780 87380
rect 33728 87316 33780 87322
rect 34924 87374 34976 87380
rect 34924 87316 34976 87322
rect 35936 87374 35988 87380
rect 35936 87316 35988 87322
rect 37132 87374 37184 87380
rect 37132 87316 37184 87322
rect 38144 87374 38196 87380
rect 38144 87316 38196 87322
rect 39248 87374 39300 87380
rect 39248 87316 39300 87322
rect 19560 87282 19612 87288
rect 15512 87204 15564 87210
rect 15512 87146 15564 87152
rect 16064 87204 16116 87210
rect 16064 87146 16116 87152
rect 17168 87204 17220 87210
rect 17168 87146 17220 87152
rect 5954 84892 6262 84901
rect 5954 84890 5960 84892
rect 6016 84890 6040 84892
rect 6096 84890 6120 84892
rect 6176 84890 6200 84892
rect 6256 84890 6262 84892
rect 6016 84838 6018 84890
rect 6198 84838 6200 84890
rect 5954 84836 5960 84838
rect 6016 84836 6040 84838
rect 6096 84836 6120 84838
rect 6176 84836 6200 84838
rect 6256 84836 6262 84838
rect 5954 84827 6262 84836
rect 12752 84688 12804 84694
rect 12752 84630 12804 84636
rect 11648 84620 11700 84626
rect 11648 84562 11700 84568
rect 7416 84552 7468 84558
rect 7416 84494 7468 84500
rect 6690 84348 6998 84357
rect 6690 84346 6696 84348
rect 6752 84346 6776 84348
rect 6832 84346 6856 84348
rect 6912 84346 6936 84348
rect 6992 84346 6998 84348
rect 6752 84294 6754 84346
rect 6934 84294 6936 84346
rect 6690 84292 6696 84294
rect 6752 84292 6776 84294
rect 6832 84292 6856 84294
rect 6912 84292 6936 84294
rect 6992 84292 6998 84294
rect 6690 84283 6998 84292
rect 5954 83804 6262 83813
rect 5954 83802 5960 83804
rect 6016 83802 6040 83804
rect 6096 83802 6120 83804
rect 6176 83802 6200 83804
rect 6256 83802 6262 83804
rect 6016 83750 6018 83802
rect 6198 83750 6200 83802
rect 5954 83748 5960 83750
rect 6016 83748 6040 83750
rect 6096 83748 6120 83750
rect 6176 83748 6200 83750
rect 6256 83748 6262 83750
rect 5954 83739 6262 83748
rect 6690 83260 6998 83269
rect 6690 83258 6696 83260
rect 6752 83258 6776 83260
rect 6832 83258 6856 83260
rect 6912 83258 6936 83260
rect 6992 83258 6998 83260
rect 6752 83206 6754 83258
rect 6934 83206 6936 83258
rect 6690 83204 6696 83206
rect 6752 83204 6776 83206
rect 6832 83204 6856 83206
rect 6912 83204 6936 83206
rect 6992 83204 6998 83206
rect 6690 83195 6998 83204
rect 5954 82716 6262 82725
rect 5954 82714 5960 82716
rect 6016 82714 6040 82716
rect 6096 82714 6120 82716
rect 6176 82714 6200 82716
rect 6256 82714 6262 82716
rect 6016 82662 6018 82714
rect 6198 82662 6200 82714
rect 5954 82660 5960 82662
rect 6016 82660 6040 82662
rect 6096 82660 6120 82662
rect 6176 82660 6200 82662
rect 6256 82660 6262 82662
rect 5954 82651 6262 82660
rect 7232 82308 7284 82314
rect 7232 82250 7284 82256
rect 6690 82172 6998 82181
rect 6690 82170 6696 82172
rect 6752 82170 6776 82172
rect 6832 82170 6856 82172
rect 6912 82170 6936 82172
rect 6992 82170 6998 82172
rect 6752 82118 6754 82170
rect 6934 82118 6936 82170
rect 6690 82116 6696 82118
rect 6752 82116 6776 82118
rect 6832 82116 6856 82118
rect 6912 82116 6936 82118
rect 6992 82116 6998 82118
rect 6690 82107 6998 82116
rect 5954 81628 6262 81637
rect 5954 81626 5960 81628
rect 6016 81626 6040 81628
rect 6096 81626 6120 81628
rect 6176 81626 6200 81628
rect 6256 81626 6262 81628
rect 6016 81574 6018 81626
rect 6198 81574 6200 81626
rect 5954 81572 5960 81574
rect 6016 81572 6040 81574
rect 6096 81572 6120 81574
rect 6176 81572 6200 81574
rect 6256 81572 6262 81574
rect 5954 81563 6262 81572
rect 6690 81084 6998 81093
rect 6690 81082 6696 81084
rect 6752 81082 6776 81084
rect 6832 81082 6856 81084
rect 6912 81082 6936 81084
rect 6992 81082 6998 81084
rect 6752 81030 6754 81082
rect 6934 81030 6936 81082
rect 6690 81028 6696 81030
rect 6752 81028 6776 81030
rect 6832 81028 6856 81030
rect 6912 81028 6936 81030
rect 6992 81028 6998 81030
rect 6690 81019 6998 81028
rect 5954 80540 6262 80549
rect 5954 80538 5960 80540
rect 6016 80538 6040 80540
rect 6096 80538 6120 80540
rect 6176 80538 6200 80540
rect 6256 80538 6262 80540
rect 6016 80486 6018 80538
rect 6198 80486 6200 80538
rect 5954 80484 5960 80486
rect 6016 80484 6040 80486
rect 6096 80484 6120 80486
rect 6176 80484 6200 80486
rect 6256 80484 6262 80486
rect 5954 80475 6262 80484
rect 7140 80200 7192 80206
rect 7138 80168 7140 80177
rect 7192 80168 7194 80177
rect 2908 80132 2960 80138
rect 7138 80103 7194 80112
rect 2908 80074 2960 80080
rect 2920 79905 2948 80074
rect 6690 79996 6998 80005
rect 6690 79994 6696 79996
rect 6752 79994 6776 79996
rect 6832 79994 6856 79996
rect 6912 79994 6936 79996
rect 6992 79994 6998 79996
rect 6752 79942 6754 79994
rect 6934 79942 6936 79994
rect 6690 79940 6696 79942
rect 6752 79940 6776 79942
rect 6832 79940 6856 79942
rect 6912 79940 6936 79942
rect 6992 79940 6998 79942
rect 6690 79931 6998 79940
rect 2906 79896 2962 79905
rect 2906 79831 2962 79840
rect 5954 79452 6262 79461
rect 5954 79450 5960 79452
rect 6016 79450 6040 79452
rect 6096 79450 6120 79452
rect 6176 79450 6200 79452
rect 6256 79450 6262 79452
rect 6016 79398 6018 79450
rect 6198 79398 6200 79450
rect 5954 79396 5960 79398
rect 6016 79396 6040 79398
rect 6096 79396 6120 79398
rect 6176 79396 6200 79398
rect 6256 79396 6262 79398
rect 5954 79387 6262 79396
rect 6690 78908 6998 78917
rect 6690 78906 6696 78908
rect 6752 78906 6776 78908
rect 6832 78906 6856 78908
rect 6912 78906 6936 78908
rect 6992 78906 6998 78908
rect 6752 78854 6754 78906
rect 6934 78854 6936 78906
rect 6690 78852 6696 78854
rect 6752 78852 6776 78854
rect 6832 78852 6856 78854
rect 6912 78852 6936 78854
rect 6992 78852 6998 78854
rect 6690 78843 6998 78852
rect 7138 78808 7194 78817
rect 7138 78743 7194 78752
rect 7152 78710 7180 78743
rect 7140 78704 7192 78710
rect 7140 78646 7192 78652
rect 2906 78536 2962 78545
rect 2906 78471 2908 78480
rect 2960 78471 2962 78480
rect 2908 78442 2960 78448
rect 5954 78364 6262 78373
rect 5954 78362 5960 78364
rect 6016 78362 6040 78364
rect 6096 78362 6120 78364
rect 6176 78362 6200 78364
rect 6256 78362 6262 78364
rect 6016 78310 6018 78362
rect 6198 78310 6200 78362
rect 5954 78308 5960 78310
rect 6016 78308 6040 78310
rect 6096 78308 6120 78310
rect 6176 78308 6200 78310
rect 6256 78308 6262 78310
rect 5954 78299 6262 78308
rect 7140 78024 7192 78030
rect 7138 77992 7140 78001
rect 7192 77992 7194 78001
rect 2908 77956 2960 77962
rect 7138 77927 7194 77936
rect 2908 77898 2960 77904
rect 2920 77865 2948 77898
rect 2906 77856 2962 77865
rect 2906 77791 2962 77800
rect 6690 77820 6998 77829
rect 6690 77818 6696 77820
rect 6752 77818 6776 77820
rect 6832 77818 6856 77820
rect 6912 77818 6936 77820
rect 6992 77818 6998 77820
rect 6752 77766 6754 77818
rect 6934 77766 6936 77818
rect 6690 77764 6696 77766
rect 6752 77764 6776 77766
rect 6832 77764 6856 77766
rect 6912 77764 6936 77766
rect 6992 77764 6998 77766
rect 6690 77755 6998 77764
rect 5954 77276 6262 77285
rect 5954 77274 5960 77276
rect 6016 77274 6040 77276
rect 6096 77274 6120 77276
rect 6176 77274 6200 77276
rect 6256 77274 6262 77276
rect 6016 77222 6018 77274
rect 6198 77222 6200 77274
rect 5954 77220 5960 77222
rect 6016 77220 6040 77222
rect 6096 77220 6120 77222
rect 6176 77220 6200 77222
rect 6256 77220 6262 77222
rect 5954 77211 6262 77220
rect 7140 76936 7192 76942
rect 7138 76904 7140 76913
rect 7192 76904 7194 76913
rect 2724 76868 2776 76874
rect 7138 76839 7194 76848
rect 2724 76810 2776 76816
rect 2736 76505 2764 76810
rect 6690 76732 6998 76741
rect 6690 76730 6696 76732
rect 6752 76730 6776 76732
rect 6832 76730 6856 76732
rect 6912 76730 6936 76732
rect 6992 76730 6998 76732
rect 6752 76678 6754 76730
rect 6934 76678 6936 76730
rect 6690 76676 6696 76678
rect 6752 76676 6776 76678
rect 6832 76676 6856 76678
rect 6912 76676 6936 76678
rect 6992 76676 6998 76678
rect 6690 76667 6998 76676
rect 2722 76496 2778 76505
rect 2722 76431 2778 76440
rect 5954 76188 6262 76197
rect 5954 76186 5960 76188
rect 6016 76186 6040 76188
rect 6096 76186 6120 76188
rect 6176 76186 6200 76188
rect 6256 76186 6262 76188
rect 6016 76134 6018 76186
rect 6198 76134 6200 76186
rect 5954 76132 5960 76134
rect 6016 76132 6040 76134
rect 6096 76132 6120 76134
rect 6176 76132 6200 76134
rect 6256 76132 6262 76134
rect 5954 76123 6262 76132
rect 7140 75848 7192 75854
rect 2906 75816 2962 75825
rect 2906 75751 2908 75760
rect 2960 75751 2962 75760
rect 7138 75816 7140 75825
rect 7192 75816 7194 75825
rect 7138 75751 7194 75760
rect 2908 75722 2960 75728
rect 6690 75644 6998 75653
rect 6690 75642 6696 75644
rect 6752 75642 6776 75644
rect 6832 75642 6856 75644
rect 6912 75642 6936 75644
rect 6992 75642 6998 75644
rect 6752 75590 6754 75642
rect 6934 75590 6936 75642
rect 6690 75588 6696 75590
rect 6752 75588 6776 75590
rect 6832 75588 6856 75590
rect 6912 75588 6936 75590
rect 6992 75588 6998 75590
rect 6690 75579 6998 75588
rect 5954 75100 6262 75109
rect 5954 75098 5960 75100
rect 6016 75098 6040 75100
rect 6096 75098 6120 75100
rect 6176 75098 6200 75100
rect 6256 75098 6262 75100
rect 6016 75046 6018 75098
rect 6198 75046 6200 75098
rect 5954 75044 5960 75046
rect 6016 75044 6040 75046
rect 6096 75044 6120 75046
rect 6176 75044 6200 75046
rect 6256 75044 6262 75046
rect 5954 75035 6262 75044
rect 4380 74896 4432 74902
rect 4380 74838 4432 74844
rect 4392 74465 4420 74838
rect 5668 74794 5720 74800
rect 5668 74736 5720 74742
rect 5680 74601 5708 74736
rect 5666 74592 5722 74601
rect 5666 74527 5722 74536
rect 6690 74556 6998 74565
rect 6690 74554 6696 74556
rect 6752 74554 6776 74556
rect 6832 74554 6856 74556
rect 6912 74554 6936 74556
rect 6992 74554 6998 74556
rect 6752 74502 6754 74554
rect 6934 74502 6936 74554
rect 6690 74500 6696 74502
rect 6752 74500 6776 74502
rect 6832 74500 6856 74502
rect 6912 74500 6936 74502
rect 6992 74500 6998 74502
rect 6690 74491 6998 74500
rect 4378 74456 4434 74465
rect 4378 74391 4434 74400
rect 5954 74012 6262 74021
rect 5954 74010 5960 74012
rect 6016 74010 6040 74012
rect 6096 74010 6120 74012
rect 6176 74010 6200 74012
rect 6256 74010 6262 74012
rect 6016 73958 6018 74010
rect 6198 73958 6200 74010
rect 5954 73956 5960 73958
rect 6016 73956 6040 73958
rect 6096 73956 6120 73958
rect 6176 73956 6200 73958
rect 6256 73956 6262 73958
rect 5954 73947 6262 73956
rect 6690 73468 6998 73477
rect 6690 73466 6696 73468
rect 6752 73466 6776 73468
rect 6832 73466 6856 73468
rect 6912 73466 6936 73468
rect 6992 73466 6998 73468
rect 6752 73414 6754 73466
rect 6934 73414 6936 73466
rect 6690 73412 6696 73414
rect 6752 73412 6776 73414
rect 6832 73412 6856 73414
rect 6912 73412 6936 73414
rect 6992 73412 6998 73414
rect 6690 73403 6998 73412
rect 7138 73368 7194 73377
rect 7138 73303 7194 73312
rect 7152 73270 7180 73303
rect 7140 73264 7192 73270
rect 7140 73206 7192 73212
rect 2906 73096 2962 73105
rect 2906 73031 2908 73040
rect 2960 73031 2962 73040
rect 2908 73002 2960 73008
rect 5954 72924 6262 72933
rect 5954 72922 5960 72924
rect 6016 72922 6040 72924
rect 6096 72922 6120 72924
rect 6176 72922 6200 72924
rect 6256 72922 6262 72924
rect 6016 72870 6018 72922
rect 6198 72870 6200 72922
rect 5954 72868 5960 72870
rect 6016 72868 6040 72870
rect 6096 72868 6120 72870
rect 6176 72868 6200 72870
rect 6256 72868 6262 72870
rect 5954 72859 6262 72868
rect 7140 72584 7192 72590
rect 7138 72552 7140 72561
rect 7192 72552 7194 72561
rect 2908 72516 2960 72522
rect 7138 72487 7194 72496
rect 2908 72458 2960 72464
rect 2920 72425 2948 72458
rect 2906 72416 2962 72425
rect 2906 72351 2962 72360
rect 6690 72380 6998 72389
rect 6690 72378 6696 72380
rect 6752 72378 6776 72380
rect 6832 72378 6856 72380
rect 6912 72378 6936 72380
rect 6992 72378 6998 72380
rect 6752 72326 6754 72378
rect 6934 72326 6936 72378
rect 6690 72324 6696 72326
rect 6752 72324 6776 72326
rect 6832 72324 6856 72326
rect 6912 72324 6936 72326
rect 6992 72324 6998 72326
rect 6690 72315 6998 72324
rect 5954 71836 6262 71845
rect 5954 71834 5960 71836
rect 6016 71834 6040 71836
rect 6096 71834 6120 71836
rect 6176 71834 6200 71836
rect 6256 71834 6262 71836
rect 6016 71782 6018 71834
rect 6198 71782 6200 71834
rect 5954 71780 5960 71782
rect 6016 71780 6040 71782
rect 6096 71780 6120 71782
rect 6176 71780 6200 71782
rect 6256 71780 6262 71782
rect 5954 71771 6262 71780
rect 7140 71496 7192 71502
rect 7138 71464 7140 71473
rect 7192 71464 7194 71473
rect 2724 71428 2776 71434
rect 7138 71399 7194 71408
rect 2724 71370 2776 71376
rect 2736 71065 2764 71370
rect 6690 71292 6998 71301
rect 6690 71290 6696 71292
rect 6752 71290 6776 71292
rect 6832 71290 6856 71292
rect 6912 71290 6936 71292
rect 6992 71290 6998 71292
rect 6752 71238 6754 71290
rect 6934 71238 6936 71290
rect 6690 71236 6696 71238
rect 6752 71236 6776 71238
rect 6832 71236 6856 71238
rect 6912 71236 6936 71238
rect 6992 71236 6998 71238
rect 6690 71227 6998 71236
rect 2722 71056 2778 71065
rect 2722 70991 2778 71000
rect 5954 70748 6262 70757
rect 5954 70746 5960 70748
rect 6016 70746 6040 70748
rect 6096 70746 6120 70748
rect 6176 70746 6200 70748
rect 6256 70746 6262 70748
rect 6016 70694 6018 70746
rect 6198 70694 6200 70746
rect 5954 70692 5960 70694
rect 6016 70692 6040 70694
rect 6096 70692 6120 70694
rect 6176 70692 6200 70694
rect 6256 70692 6262 70694
rect 5954 70683 6262 70692
rect 7140 70408 7192 70414
rect 2906 70376 2962 70385
rect 2906 70311 2908 70320
rect 2960 70311 2962 70320
rect 7138 70376 7140 70385
rect 7192 70376 7194 70385
rect 7138 70311 7194 70320
rect 2908 70282 2960 70288
rect 6690 70204 6998 70213
rect 6690 70202 6696 70204
rect 6752 70202 6776 70204
rect 6832 70202 6856 70204
rect 6912 70202 6936 70204
rect 6992 70202 6998 70204
rect 6752 70150 6754 70202
rect 6934 70150 6936 70202
rect 6690 70148 6696 70150
rect 6752 70148 6776 70150
rect 6832 70148 6856 70150
rect 6912 70148 6936 70150
rect 6992 70148 6998 70150
rect 6690 70139 6998 70148
rect 5954 69660 6262 69669
rect 5954 69658 5960 69660
rect 6016 69658 6040 69660
rect 6096 69658 6120 69660
rect 6176 69658 6200 69660
rect 6256 69658 6262 69660
rect 6016 69606 6018 69658
rect 6198 69606 6200 69658
rect 5954 69604 5960 69606
rect 6016 69604 6040 69606
rect 6096 69604 6120 69606
rect 6176 69604 6200 69606
rect 6256 69604 6262 69606
rect 5954 69595 6262 69604
rect 5668 69354 5720 69360
rect 5668 69296 5720 69302
rect 4380 69252 4432 69258
rect 4380 69194 4432 69200
rect 4392 69025 4420 69194
rect 4378 69016 4434 69025
rect 4378 68951 4434 68960
rect 5680 68889 5708 69296
rect 6690 69116 6998 69125
rect 6690 69114 6696 69116
rect 6752 69114 6776 69116
rect 6832 69114 6856 69116
rect 6912 69114 6936 69116
rect 6992 69114 6998 69116
rect 6752 69062 6754 69114
rect 6934 69062 6936 69114
rect 6690 69060 6696 69062
rect 6752 69060 6776 69062
rect 6832 69060 6856 69062
rect 6912 69060 6936 69062
rect 6992 69060 6998 69062
rect 6690 69051 6998 69060
rect 5666 68880 5722 68889
rect 5666 68815 5722 68824
rect 5954 68572 6262 68581
rect 5954 68570 5960 68572
rect 6016 68570 6040 68572
rect 6096 68570 6120 68572
rect 6176 68570 6200 68572
rect 6256 68570 6262 68572
rect 6016 68518 6018 68570
rect 6198 68518 6200 68570
rect 5954 68516 5960 68518
rect 6016 68516 6040 68518
rect 6096 68516 6120 68518
rect 6176 68516 6200 68518
rect 6256 68516 6262 68518
rect 5954 68507 6262 68516
rect 5666 68200 5722 68209
rect 5666 68135 5722 68144
rect 5680 67796 5708 68135
rect 6690 68028 6998 68037
rect 6690 68026 6696 68028
rect 6752 68026 6776 68028
rect 6832 68026 6856 68028
rect 6912 68026 6936 68028
rect 6992 68026 6998 68028
rect 6752 67974 6754 68026
rect 6934 67974 6936 68026
rect 6690 67972 6696 67974
rect 6752 67972 6776 67974
rect 6832 67972 6856 67974
rect 6912 67972 6936 67974
rect 6992 67972 6998 67974
rect 6690 67963 6998 67972
rect 5668 67790 5720 67796
rect 5668 67732 5720 67738
rect 2906 67656 2962 67665
rect 2906 67591 2908 67600
rect 2960 67591 2962 67600
rect 2908 67562 2960 67568
rect 5954 67484 6262 67493
rect 5954 67482 5960 67484
rect 6016 67482 6040 67484
rect 6096 67482 6120 67484
rect 6176 67482 6200 67484
rect 6256 67482 6262 67484
rect 6016 67430 6018 67482
rect 6198 67430 6200 67482
rect 5954 67428 5960 67430
rect 6016 67428 6040 67430
rect 6096 67428 6120 67430
rect 6176 67428 6200 67430
rect 6256 67428 6262 67430
rect 5954 67419 6262 67428
rect 7140 67144 7192 67150
rect 7138 67112 7140 67121
rect 7192 67112 7194 67121
rect 2908 67076 2960 67082
rect 7138 67047 7194 67056
rect 2908 67018 2960 67024
rect 2920 66985 2948 67018
rect 2906 66976 2962 66985
rect 2906 66911 2962 66920
rect 6690 66940 6998 66949
rect 6690 66938 6696 66940
rect 6752 66938 6776 66940
rect 6832 66938 6856 66940
rect 6912 66938 6936 66940
rect 6992 66938 6998 66940
rect 6752 66886 6754 66938
rect 6934 66886 6936 66938
rect 6690 66884 6696 66886
rect 6752 66884 6776 66886
rect 6832 66884 6856 66886
rect 6912 66884 6936 66886
rect 6992 66884 6998 66886
rect 6690 66875 6998 66884
rect 7244 66474 7272 82250
rect 7152 66446 7272 66474
rect 5954 66396 6262 66405
rect 5954 66394 5960 66396
rect 6016 66394 6040 66396
rect 6096 66394 6120 66396
rect 6176 66394 6200 66396
rect 6256 66394 6262 66396
rect 6016 66342 6018 66394
rect 6198 66342 6200 66394
rect 5954 66340 5960 66342
rect 6016 66340 6040 66342
rect 6096 66340 6120 66342
rect 6176 66340 6200 66342
rect 6256 66340 6262 66342
rect 5954 66331 6262 66340
rect 2908 65988 2960 65994
rect 2908 65930 2960 65936
rect 2920 65625 2948 65930
rect 6690 65852 6998 65861
rect 6690 65850 6696 65852
rect 6752 65850 6776 65852
rect 6832 65850 6856 65852
rect 6912 65850 6936 65852
rect 6992 65850 6998 65852
rect 6752 65798 6754 65850
rect 6934 65798 6936 65850
rect 6690 65796 6696 65798
rect 6752 65796 6776 65798
rect 6832 65796 6856 65798
rect 6912 65796 6936 65798
rect 6992 65796 6998 65798
rect 6690 65787 6998 65796
rect 2906 65616 2962 65625
rect 2906 65551 2962 65560
rect 5954 65308 6262 65317
rect 5954 65306 5960 65308
rect 6016 65306 6040 65308
rect 6096 65306 6120 65308
rect 6176 65306 6200 65308
rect 6256 65306 6262 65308
rect 6016 65254 6018 65306
rect 6198 65254 6200 65306
rect 5954 65252 5960 65254
rect 6016 65252 6040 65254
rect 6096 65252 6120 65254
rect 6176 65252 6200 65254
rect 6256 65252 6262 65254
rect 5954 65243 6262 65252
rect 2906 64936 2962 64945
rect 2906 64871 2908 64880
rect 2960 64871 2962 64880
rect 2908 64842 2960 64848
rect 6690 64764 6998 64773
rect 6690 64762 6696 64764
rect 6752 64762 6776 64764
rect 6832 64762 6856 64764
rect 6912 64762 6936 64764
rect 6992 64762 6998 64764
rect 6752 64710 6754 64762
rect 6934 64710 6936 64762
rect 6690 64708 6696 64710
rect 6752 64708 6776 64710
rect 6832 64708 6856 64710
rect 6912 64708 6936 64710
rect 6992 64708 6998 64710
rect 6690 64699 6998 64708
rect 5954 64220 6262 64229
rect 5954 64218 5960 64220
rect 6016 64218 6040 64220
rect 6096 64218 6120 64220
rect 6176 64218 6200 64220
rect 6256 64218 6262 64220
rect 6016 64166 6018 64218
rect 6198 64166 6200 64218
rect 5954 64164 5960 64166
rect 6016 64164 6040 64166
rect 6096 64164 6120 64166
rect 6176 64164 6200 64166
rect 6256 64164 6262 64166
rect 5954 64155 6262 64164
rect 5208 63914 5260 63920
rect 5208 63856 5260 63862
rect 5220 63585 5248 63856
rect 6690 63676 6998 63685
rect 6690 63674 6696 63676
rect 6752 63674 6776 63676
rect 6832 63674 6856 63676
rect 6912 63674 6936 63676
rect 6992 63674 6998 63676
rect 6752 63622 6754 63674
rect 6934 63622 6936 63674
rect 6690 63620 6696 63622
rect 6752 63620 6776 63622
rect 6832 63620 6856 63622
rect 6912 63620 6936 63622
rect 6992 63620 6998 63622
rect 6690 63611 6998 63620
rect 5206 63576 5262 63585
rect 5206 63511 5262 63520
rect 5954 63132 6262 63141
rect 5954 63130 5960 63132
rect 6016 63130 6040 63132
rect 6096 63130 6120 63132
rect 6176 63130 6200 63132
rect 6256 63130 6262 63132
rect 6016 63078 6018 63130
rect 6198 63078 6200 63130
rect 5954 63076 5960 63078
rect 6016 63076 6040 63078
rect 6096 63076 6120 63078
rect 6176 63076 6200 63078
rect 6256 63076 6262 63078
rect 5954 63067 6262 63076
rect 6690 62588 6998 62597
rect 6690 62586 6696 62588
rect 6752 62586 6776 62588
rect 6832 62586 6856 62588
rect 6912 62586 6936 62588
rect 6992 62586 6998 62588
rect 6752 62534 6754 62586
rect 6934 62534 6936 62586
rect 6690 62532 6696 62534
rect 6752 62532 6776 62534
rect 6832 62532 6856 62534
rect 6912 62532 6936 62534
rect 6992 62532 6998 62534
rect 6690 62523 6998 62532
rect 4932 62350 4984 62356
rect 4932 62292 4984 62298
rect 4944 62225 4972 62292
rect 4930 62216 4986 62225
rect 4930 62151 4986 62160
rect 5954 62044 6262 62053
rect 5954 62042 5960 62044
rect 6016 62042 6040 62044
rect 6096 62042 6120 62044
rect 6176 62042 6200 62044
rect 6256 62042 6262 62044
rect 6016 61990 6018 62042
rect 6198 61990 6200 62042
rect 5954 61988 5960 61990
rect 6016 61988 6040 61990
rect 6096 61988 6120 61990
rect 6176 61988 6200 61990
rect 6256 61988 6262 61990
rect 5954 61979 6262 61988
rect 2908 61636 2960 61642
rect 2908 61578 2960 61584
rect 2920 61545 2948 61578
rect 2906 61536 2962 61545
rect 2906 61471 2962 61480
rect 6690 61500 6998 61509
rect 6690 61498 6696 61500
rect 6752 61498 6776 61500
rect 6832 61498 6856 61500
rect 6912 61498 6936 61500
rect 6992 61498 6998 61500
rect 6752 61446 6754 61498
rect 6934 61446 6936 61498
rect 6690 61444 6696 61446
rect 6752 61444 6776 61446
rect 6832 61444 6856 61446
rect 6912 61444 6936 61446
rect 6992 61444 6998 61446
rect 6690 61435 6998 61444
rect 5954 60956 6262 60965
rect 5954 60954 5960 60956
rect 6016 60954 6040 60956
rect 6096 60954 6120 60956
rect 6176 60954 6200 60956
rect 6256 60954 6262 60956
rect 6016 60902 6018 60954
rect 6198 60902 6200 60954
rect 5954 60900 5960 60902
rect 6016 60900 6040 60902
rect 6096 60900 6120 60902
rect 6176 60900 6200 60902
rect 6256 60900 6262 60902
rect 5954 60891 6262 60900
rect 2908 60548 2960 60554
rect 2908 60490 2960 60496
rect 2920 60185 2948 60490
rect 6690 60412 6998 60421
rect 6690 60410 6696 60412
rect 6752 60410 6776 60412
rect 6832 60410 6856 60412
rect 6912 60410 6936 60412
rect 6992 60410 6998 60412
rect 6752 60358 6754 60410
rect 6934 60358 6936 60410
rect 6690 60356 6696 60358
rect 6752 60356 6776 60358
rect 6832 60356 6856 60358
rect 6912 60356 6936 60358
rect 6992 60356 6998 60358
rect 6690 60347 6998 60356
rect 2906 60176 2962 60185
rect 2906 60111 2962 60120
rect 5954 59868 6262 59877
rect 5954 59866 5960 59868
rect 6016 59866 6040 59868
rect 6096 59866 6120 59868
rect 6176 59866 6200 59868
rect 6256 59866 6262 59868
rect 6016 59814 6018 59866
rect 6198 59814 6200 59866
rect 5954 59812 5960 59814
rect 6016 59812 6040 59814
rect 6096 59812 6120 59814
rect 6176 59812 6200 59814
rect 6256 59812 6262 59814
rect 5954 59803 6262 59812
rect 5208 59528 5260 59534
rect 5206 59496 5208 59505
rect 5260 59496 5262 59505
rect 5206 59431 5262 59440
rect 6690 59324 6998 59333
rect 6690 59322 6696 59324
rect 6752 59322 6776 59324
rect 6832 59322 6856 59324
rect 6912 59322 6936 59324
rect 6992 59322 6998 59324
rect 6752 59270 6754 59322
rect 6934 59270 6936 59322
rect 6690 59268 6696 59270
rect 6752 59268 6776 59270
rect 6832 59268 6856 59270
rect 6912 59268 6936 59270
rect 6992 59268 6998 59270
rect 6690 59259 6998 59268
rect 5954 58780 6262 58789
rect 5954 58778 5960 58780
rect 6016 58778 6040 58780
rect 6096 58778 6120 58780
rect 6176 58778 6200 58780
rect 6256 58778 6262 58780
rect 6016 58726 6018 58778
rect 6198 58726 6200 58778
rect 5954 58724 5960 58726
rect 6016 58724 6040 58726
rect 6096 58724 6120 58726
rect 6176 58724 6200 58726
rect 6256 58724 6262 58726
rect 5954 58715 6262 58724
rect 5208 58474 5260 58480
rect 5208 58416 5260 58422
rect 5220 58145 5248 58416
rect 5392 58372 5444 58378
rect 5392 58314 5444 58320
rect 5206 58136 5262 58145
rect 5206 58071 5262 58080
rect 5404 58009 5432 58314
rect 6690 58236 6998 58245
rect 6690 58234 6696 58236
rect 6752 58234 6776 58236
rect 6832 58234 6856 58236
rect 6912 58234 6936 58236
rect 6992 58234 6998 58236
rect 6752 58182 6754 58234
rect 6934 58182 6936 58234
rect 6690 58180 6696 58182
rect 6752 58180 6776 58182
rect 6832 58180 6856 58182
rect 6912 58180 6936 58182
rect 6992 58180 6998 58182
rect 6690 58171 6998 58180
rect 5390 58000 5446 58009
rect 5390 57935 5446 57944
rect 5954 57692 6262 57701
rect 5954 57690 5960 57692
rect 6016 57690 6040 57692
rect 6096 57690 6120 57692
rect 6176 57690 6200 57692
rect 6256 57690 6262 57692
rect 6016 57638 6018 57690
rect 6198 57638 6200 57690
rect 5954 57636 5960 57638
rect 6016 57636 6040 57638
rect 6096 57636 6120 57638
rect 6176 57636 6200 57638
rect 6256 57636 6262 57638
rect 5954 57627 6262 57636
rect 6690 57148 6998 57157
rect 6690 57146 6696 57148
rect 6752 57146 6776 57148
rect 6832 57146 6856 57148
rect 6912 57146 6936 57148
rect 6992 57146 6998 57148
rect 6752 57094 6754 57146
rect 6934 57094 6936 57146
rect 6690 57092 6696 57094
rect 6752 57092 6776 57094
rect 6832 57092 6856 57094
rect 6912 57092 6936 57094
rect 6992 57092 6998 57094
rect 6690 57083 6998 57092
rect 4932 56910 4984 56916
rect 4932 56852 4984 56858
rect 4944 56785 4972 56852
rect 4930 56776 4986 56785
rect 4930 56711 4986 56720
rect 5954 56604 6262 56613
rect 5954 56602 5960 56604
rect 6016 56602 6040 56604
rect 6096 56602 6120 56604
rect 6176 56602 6200 56604
rect 6256 56602 6262 56604
rect 6016 56550 6018 56602
rect 6198 56550 6200 56602
rect 5954 56548 5960 56550
rect 6016 56548 6040 56550
rect 6096 56548 6120 56550
rect 6176 56548 6200 56550
rect 6256 56548 6262 56550
rect 5954 56539 6262 56548
rect 2908 56264 2960 56270
rect 2908 56206 2960 56212
rect 2920 56105 2948 56206
rect 2906 56096 2962 56105
rect 2906 56031 2962 56040
rect 6690 56060 6998 56069
rect 6690 56058 6696 56060
rect 6752 56058 6776 56060
rect 6832 56058 6856 56060
rect 6912 56058 6936 56060
rect 6992 56058 6998 56060
rect 6752 56006 6754 56058
rect 6934 56006 6936 56058
rect 6690 56004 6696 56006
rect 6752 56004 6776 56006
rect 6832 56004 6856 56006
rect 6912 56004 6936 56006
rect 6992 56004 6998 56006
rect 6690 55995 6998 56004
rect 5954 55516 6262 55525
rect 5954 55514 5960 55516
rect 6016 55514 6040 55516
rect 6096 55514 6120 55516
rect 6176 55514 6200 55516
rect 6256 55514 6262 55516
rect 6016 55462 6018 55514
rect 6198 55462 6200 55514
rect 5954 55460 5960 55462
rect 6016 55460 6040 55462
rect 6096 55460 6120 55462
rect 6176 55460 6200 55462
rect 6256 55460 6262 55462
rect 5954 55451 6262 55460
rect 2908 55176 2960 55182
rect 2908 55118 2960 55124
rect 2920 54745 2948 55118
rect 6690 54972 6998 54981
rect 6690 54970 6696 54972
rect 6752 54970 6776 54972
rect 6832 54970 6856 54972
rect 6912 54970 6936 54972
rect 6992 54970 6998 54972
rect 6752 54918 6754 54970
rect 6934 54918 6936 54970
rect 6690 54916 6696 54918
rect 6752 54916 6776 54918
rect 6832 54916 6856 54918
rect 6912 54916 6936 54918
rect 6992 54916 6998 54918
rect 6690 54907 6998 54916
rect 2906 54736 2962 54745
rect 2906 54671 2962 54680
rect 5954 54428 6262 54437
rect 5954 54426 5960 54428
rect 6016 54426 6040 54428
rect 6096 54426 6120 54428
rect 6176 54426 6200 54428
rect 6256 54426 6262 54428
rect 6016 54374 6018 54426
rect 6198 54374 6200 54426
rect 5954 54372 5960 54374
rect 6016 54372 6040 54374
rect 6096 54372 6120 54374
rect 6176 54372 6200 54374
rect 6256 54372 6262 54374
rect 5954 54363 6262 54372
rect 5116 54088 5168 54094
rect 5114 54056 5116 54065
rect 5668 54088 5720 54094
rect 5168 54056 5170 54065
rect 5114 53991 5170 54000
rect 5666 54056 5668 54065
rect 5720 54056 5722 54065
rect 5666 53991 5722 54000
rect 6690 53884 6998 53893
rect 6690 53882 6696 53884
rect 6752 53882 6776 53884
rect 6832 53882 6856 53884
rect 6912 53882 6936 53884
rect 6992 53882 6998 53884
rect 6752 53830 6754 53882
rect 6934 53830 6936 53882
rect 6690 53828 6696 53830
rect 6752 53828 6776 53830
rect 6832 53828 6856 53830
rect 6912 53828 6936 53830
rect 6992 53828 6998 53830
rect 6690 53819 6998 53828
rect 5954 53340 6262 53349
rect 5954 53338 5960 53340
rect 6016 53338 6040 53340
rect 6096 53338 6120 53340
rect 6176 53338 6200 53340
rect 6256 53338 6262 53340
rect 6016 53286 6018 53338
rect 6198 53286 6200 53338
rect 5954 53284 5960 53286
rect 6016 53284 6040 53286
rect 6096 53284 6120 53286
rect 6176 53284 6200 53286
rect 6256 53284 6262 53286
rect 5954 53275 6262 53284
rect 2908 53000 2960 53006
rect 2908 52942 2960 52948
rect 2920 52705 2948 52942
rect 6690 52796 6998 52805
rect 6690 52794 6696 52796
rect 6752 52794 6776 52796
rect 6832 52794 6856 52796
rect 6912 52794 6936 52796
rect 6992 52794 6998 52796
rect 6752 52742 6754 52794
rect 6934 52742 6936 52794
rect 6690 52740 6696 52742
rect 6752 52740 6776 52742
rect 6832 52740 6856 52742
rect 6912 52740 6936 52742
rect 6992 52740 6998 52742
rect 6690 52731 6998 52740
rect 2906 52696 2962 52705
rect 2906 52631 2962 52640
rect 5954 52252 6262 52261
rect 5954 52250 5960 52252
rect 6016 52250 6040 52252
rect 6096 52250 6120 52252
rect 6176 52250 6200 52252
rect 6256 52250 6262 52252
rect 6016 52198 6018 52250
rect 6198 52198 6200 52250
rect 5954 52196 5960 52198
rect 6016 52196 6040 52198
rect 6096 52196 6120 52198
rect 6176 52196 6200 52198
rect 6256 52196 6262 52198
rect 5954 52187 6262 52196
rect 6690 51708 6998 51717
rect 6690 51706 6696 51708
rect 6752 51706 6776 51708
rect 6832 51706 6856 51708
rect 6912 51706 6936 51708
rect 6992 51706 6998 51708
rect 6752 51654 6754 51706
rect 6934 51654 6936 51706
rect 6690 51652 6696 51654
rect 6752 51652 6776 51654
rect 6832 51652 6856 51654
rect 6912 51652 6936 51654
rect 6992 51652 6998 51654
rect 6690 51643 6998 51652
rect 2908 51436 2960 51442
rect 2908 51378 2960 51384
rect 2920 51345 2948 51378
rect 2906 51336 2962 51345
rect 2906 51271 2962 51280
rect 5954 51164 6262 51173
rect 5954 51162 5960 51164
rect 6016 51162 6040 51164
rect 6096 51162 6120 51164
rect 6176 51162 6200 51164
rect 6256 51162 6262 51164
rect 6016 51110 6018 51162
rect 6198 51110 6200 51162
rect 5954 51108 5960 51110
rect 6016 51108 6040 51110
rect 6096 51108 6120 51110
rect 6176 51108 6200 51110
rect 6256 51108 6262 51110
rect 5954 51099 6262 51108
rect 6690 50620 6998 50629
rect 6690 50618 6696 50620
rect 6752 50618 6776 50620
rect 6832 50618 6856 50620
rect 6912 50618 6936 50620
rect 6992 50618 6998 50620
rect 6752 50566 6754 50618
rect 6934 50566 6936 50618
rect 6690 50564 6696 50566
rect 6752 50564 6776 50566
rect 6832 50564 6856 50566
rect 6912 50564 6936 50566
rect 6992 50564 6998 50566
rect 6690 50555 6998 50564
rect 5954 50076 6262 50085
rect 5954 50074 5960 50076
rect 6016 50074 6040 50076
rect 6096 50074 6120 50076
rect 6176 50074 6200 50076
rect 6256 50074 6262 50076
rect 6016 50022 6018 50074
rect 6198 50022 6200 50074
rect 5954 50020 5960 50022
rect 6016 50020 6040 50022
rect 6096 50020 6120 50022
rect 6176 50020 6200 50022
rect 6256 50020 6262 50022
rect 5954 50011 6262 50020
rect 6690 49532 6998 49541
rect 6690 49530 6696 49532
rect 6752 49530 6776 49532
rect 6832 49530 6856 49532
rect 6912 49530 6936 49532
rect 6992 49530 6998 49532
rect 6752 49478 6754 49530
rect 6934 49478 6936 49530
rect 6690 49476 6696 49478
rect 6752 49476 6776 49478
rect 6832 49476 6856 49478
rect 6912 49476 6936 49478
rect 6992 49476 6998 49478
rect 6690 49467 6998 49476
rect 5954 48988 6262 48997
rect 5954 48986 5960 48988
rect 6016 48986 6040 48988
rect 6096 48986 6120 48988
rect 6176 48986 6200 48988
rect 6256 48986 6262 48988
rect 6016 48934 6018 48986
rect 6198 48934 6200 48986
rect 5954 48932 5960 48934
rect 6016 48932 6040 48934
rect 6096 48932 6120 48934
rect 6176 48932 6200 48934
rect 6256 48932 6262 48934
rect 5954 48923 6262 48932
rect 6690 48444 6998 48453
rect 6690 48442 6696 48444
rect 6752 48442 6776 48444
rect 6832 48442 6856 48444
rect 6912 48442 6936 48444
rect 6992 48442 6998 48444
rect 6752 48390 6754 48442
rect 6934 48390 6936 48442
rect 6690 48388 6696 48390
rect 6752 48388 6776 48390
rect 6832 48388 6856 48390
rect 6912 48388 6936 48390
rect 6992 48388 6998 48390
rect 6690 48379 6998 48388
rect 5954 47900 6262 47909
rect 5954 47898 5960 47900
rect 6016 47898 6040 47900
rect 6096 47898 6120 47900
rect 6176 47898 6200 47900
rect 6256 47898 6262 47900
rect 6016 47846 6018 47898
rect 6198 47846 6200 47898
rect 5954 47844 5960 47846
rect 6016 47844 6040 47846
rect 6096 47844 6120 47846
rect 6176 47844 6200 47846
rect 6256 47844 6262 47846
rect 5954 47835 6262 47844
rect 6690 47356 6998 47365
rect 6690 47354 6696 47356
rect 6752 47354 6776 47356
rect 6832 47354 6856 47356
rect 6912 47354 6936 47356
rect 6992 47354 6998 47356
rect 6752 47302 6754 47354
rect 6934 47302 6936 47354
rect 6690 47300 6696 47302
rect 6752 47300 6776 47302
rect 6832 47300 6856 47302
rect 6912 47300 6936 47302
rect 6992 47300 6998 47302
rect 6690 47291 6998 47300
rect 5954 46812 6262 46821
rect 5954 46810 5960 46812
rect 6016 46810 6040 46812
rect 6096 46810 6120 46812
rect 6176 46810 6200 46812
rect 6256 46810 6262 46812
rect 6016 46758 6018 46810
rect 6198 46758 6200 46810
rect 5954 46756 5960 46758
rect 6016 46756 6040 46758
rect 6096 46756 6120 46758
rect 6176 46756 6200 46758
rect 6256 46756 6262 46758
rect 5954 46747 6262 46756
rect 6690 46268 6998 46277
rect 6690 46266 6696 46268
rect 6752 46266 6776 46268
rect 6832 46266 6856 46268
rect 6912 46266 6936 46268
rect 6992 46266 6998 46268
rect 6752 46214 6754 46266
rect 6934 46214 6936 46266
rect 6690 46212 6696 46214
rect 6752 46212 6776 46214
rect 6832 46212 6856 46214
rect 6912 46212 6936 46214
rect 6992 46212 6998 46214
rect 6690 46203 6998 46212
rect 5392 45928 5444 45934
rect 5392 45870 5444 45876
rect 5404 45594 5432 45870
rect 5954 45724 6262 45733
rect 5954 45722 5960 45724
rect 6016 45722 6040 45724
rect 6096 45722 6120 45724
rect 6176 45722 6200 45724
rect 6256 45722 6262 45724
rect 6016 45670 6018 45722
rect 6198 45670 6200 45722
rect 5954 45668 5960 45670
rect 6016 45668 6040 45670
rect 6096 45668 6120 45670
rect 6176 45668 6200 45670
rect 6256 45668 6262 45670
rect 5954 45659 6262 45668
rect 5392 45588 5444 45594
rect 5392 45530 5444 45536
rect 7152 45526 7180 66446
rect 7232 66056 7284 66062
rect 7232 65998 7284 66004
rect 7244 65897 7272 65998
rect 7230 65888 7286 65897
rect 7230 65823 7286 65832
rect 7232 64968 7284 64974
rect 7232 64910 7284 64916
rect 7244 64809 7272 64910
rect 7230 64800 7286 64809
rect 7230 64735 7286 64744
rect 7428 64634 7456 84494
rect 10544 84484 10596 84490
rect 10544 84426 10596 84432
rect 7600 82376 7652 82382
rect 10556 82353 10584 84426
rect 11660 82466 11688 84562
rect 12764 82466 12792 84630
rect 13856 84484 13908 84490
rect 13856 84426 13908 84432
rect 13868 83130 13896 84426
rect 13856 83124 13908 83130
rect 13856 83066 13908 83072
rect 13868 82466 13896 83066
rect 11660 82438 11716 82466
rect 12764 82438 12820 82466
rect 13868 82438 13924 82466
rect 15524 82450 15552 87146
rect 16076 82466 16104 87146
rect 17180 82466 17208 87146
rect 17722 87068 18030 87077
rect 17722 87066 17728 87068
rect 17784 87066 17808 87068
rect 17864 87066 17888 87068
rect 17944 87066 17968 87068
rect 18024 87066 18030 87068
rect 17784 87014 17786 87066
rect 17966 87014 17968 87066
rect 17722 87012 17728 87014
rect 17784 87012 17808 87014
rect 17864 87012 17888 87014
rect 17944 87012 17968 87014
rect 18024 87012 18030 87014
rect 17722 87003 18030 87012
rect 17722 85980 18030 85989
rect 17722 85978 17728 85980
rect 17784 85978 17808 85980
rect 17864 85978 17888 85980
rect 17944 85978 17968 85980
rect 18024 85978 18030 85980
rect 17784 85926 17786 85978
rect 17966 85926 17968 85978
rect 17722 85924 17728 85926
rect 17784 85924 17808 85926
rect 17864 85924 17888 85926
rect 17944 85924 17968 85926
rect 18024 85924 18030 85926
rect 17722 85915 18030 85924
rect 17722 84892 18030 84901
rect 17722 84890 17728 84892
rect 17784 84890 17808 84892
rect 17864 84890 17888 84892
rect 17944 84890 17968 84892
rect 18024 84890 18030 84892
rect 17784 84838 17786 84890
rect 17966 84838 17968 84890
rect 17722 84836 17728 84838
rect 17784 84836 17808 84838
rect 17864 84836 17888 84838
rect 17944 84836 17968 84838
rect 18024 84836 18030 84838
rect 17722 84827 18030 84836
rect 18284 82466 18312 87282
rect 18382 86524 18690 86533
rect 18382 86522 18388 86524
rect 18444 86522 18468 86524
rect 18524 86522 18548 86524
rect 18604 86522 18628 86524
rect 18684 86522 18690 86524
rect 18444 86470 18446 86522
rect 18626 86470 18628 86522
rect 18382 86468 18388 86470
rect 18444 86468 18468 86470
rect 18524 86468 18548 86470
rect 18604 86468 18628 86470
rect 18684 86468 18690 86470
rect 18382 86459 18690 86468
rect 18382 85436 18690 85445
rect 18382 85434 18388 85436
rect 18444 85434 18468 85436
rect 18524 85434 18548 85436
rect 18604 85434 18628 85436
rect 18684 85434 18690 85436
rect 18444 85382 18446 85434
rect 18626 85382 18628 85434
rect 18382 85380 18388 85382
rect 18444 85380 18468 85382
rect 18524 85380 18548 85382
rect 18604 85380 18628 85382
rect 18684 85380 18690 85382
rect 18382 85371 18690 85380
rect 18382 84348 18690 84357
rect 18382 84346 18388 84348
rect 18444 84346 18468 84348
rect 18524 84346 18548 84348
rect 18604 84346 18628 84348
rect 18684 84346 18690 84348
rect 18444 84294 18446 84346
rect 18626 84294 18628 84346
rect 18382 84292 18388 84294
rect 18444 84292 18468 84294
rect 18524 84292 18548 84294
rect 18604 84292 18628 84294
rect 18684 84292 18690 84294
rect 18382 84283 18690 84292
rect 19572 82466 19600 87282
rect 22688 87272 22740 87278
rect 22688 87214 22740 87220
rect 27104 87272 27156 87278
rect 27104 87214 27156 87220
rect 20480 87204 20532 87210
rect 20480 87146 20532 87152
rect 21584 87204 21636 87210
rect 21584 87146 21636 87152
rect 11688 82382 11716 82438
rect 11676 82376 11728 82382
rect 7600 82318 7652 82324
rect 10542 82344 10598 82353
rect 7416 64628 7468 64634
rect 7416 64570 7468 64576
rect 7428 63886 7456 64570
rect 7416 63880 7468 63886
rect 7416 63822 7468 63828
rect 7232 63812 7284 63818
rect 7232 63754 7284 63760
rect 7244 63698 7272 63754
rect 7244 63670 7364 63698
rect 7336 63274 7364 63670
rect 7324 63268 7376 63274
rect 7324 63210 7376 63216
rect 7230 62488 7286 62497
rect 7230 62423 7232 62432
rect 7284 62423 7286 62432
rect 7232 62394 7284 62400
rect 7232 61704 7284 61710
rect 7232 61646 7284 61652
rect 7244 61545 7272 61646
rect 7230 61536 7286 61545
rect 7230 61471 7286 61480
rect 7232 60616 7284 60622
rect 7232 60558 7284 60564
rect 7244 60457 7272 60558
rect 7230 60448 7286 60457
rect 7230 60383 7286 60392
rect 7232 59528 7284 59534
rect 7232 59470 7284 59476
rect 7244 59369 7272 59470
rect 7230 59360 7286 59369
rect 7230 59295 7286 59304
rect 7230 57048 7286 57057
rect 7230 56983 7232 56992
rect 7284 56983 7286 56992
rect 7232 56954 7284 56960
rect 7232 56264 7284 56270
rect 7232 56206 7284 56212
rect 7244 56105 7272 56206
rect 7230 56096 7286 56105
rect 7230 56031 7286 56040
rect 7232 55176 7284 55182
rect 7232 55118 7284 55124
rect 7244 55017 7272 55118
rect 7230 55008 7286 55017
rect 7230 54943 7286 54952
rect 7232 53000 7284 53006
rect 7232 52942 7284 52948
rect 7244 52841 7272 52942
rect 7230 52832 7286 52841
rect 7230 52767 7286 52776
rect 7230 51608 7286 51617
rect 7230 51543 7232 51552
rect 7284 51543 7286 51552
rect 7232 51514 7284 51520
rect 7336 45594 7364 63210
rect 7612 47154 7640 82318
rect 11676 82318 11728 82324
rect 10542 82279 10598 82288
rect 11688 82180 11716 82318
rect 12792 82314 12820 82438
rect 12780 82308 12832 82314
rect 12780 82250 12832 82256
rect 12792 82180 12820 82250
rect 13896 82180 13924 82438
rect 14988 82444 15040 82450
rect 14988 82386 15040 82392
rect 15512 82444 15564 82450
rect 16076 82438 16132 82466
rect 17180 82438 17236 82466
rect 18284 82438 18340 82466
rect 15512 82386 15564 82392
rect 15000 82180 15028 82386
rect 16104 82180 16132 82438
rect 17208 82180 17236 82438
rect 18312 82180 18340 82438
rect 19416 82438 19600 82466
rect 20492 82466 20520 87146
rect 21596 82466 21624 87146
rect 22700 82466 22728 87214
rect 23792 87204 23844 87210
rect 23792 87146 23844 87152
rect 25080 87204 25132 87210
rect 25080 87146 25132 87152
rect 26092 87204 26144 87210
rect 26092 87146 26144 87152
rect 23804 82466 23832 87146
rect 25092 82466 25120 87146
rect 26104 82466 26132 87146
rect 20492 82438 20548 82466
rect 21596 82438 21652 82466
rect 22700 82438 22756 82466
rect 23804 82438 23860 82466
rect 19416 82180 19444 82438
rect 20520 82180 20548 82438
rect 21624 82180 21652 82438
rect 22728 82180 22756 82438
rect 23832 82180 23860 82438
rect 24936 82438 25120 82466
rect 26040 82438 26132 82466
rect 27116 82466 27144 87214
rect 28208 87204 28260 87210
rect 28208 87146 28260 87152
rect 29312 87204 29364 87210
rect 29312 87146 29364 87152
rect 28220 82466 28248 87146
rect 29324 82466 29352 87146
rect 30612 82466 30640 87316
rect 30704 84762 31284 84778
rect 30692 84756 31284 84762
rect 30744 84750 31284 84756
rect 30692 84698 30744 84704
rect 31256 84694 31284 84750
rect 31244 84688 31296 84694
rect 30704 84626 31192 84642
rect 31244 84630 31296 84636
rect 30692 84620 31204 84626
rect 30744 84614 31152 84620
rect 30692 84562 30744 84568
rect 31152 84562 31204 84568
rect 27116 82438 27172 82466
rect 28220 82438 28276 82466
rect 29324 82438 29380 82466
rect 24936 82180 24964 82438
rect 26040 82180 26068 82438
rect 27144 82180 27172 82438
rect 28248 82180 28276 82438
rect 29352 82180 29380 82438
rect 30456 82438 30640 82466
rect 31532 82466 31560 87316
rect 32636 82466 32664 87316
rect 33740 82466 33768 87316
rect 34936 82466 34964 87316
rect 31532 82438 31588 82466
rect 32636 82438 32692 82466
rect 33740 82438 33796 82466
rect 30456 82180 30484 82438
rect 31560 82180 31588 82438
rect 32664 82180 32692 82438
rect 33768 82180 33796 82438
rect 34872 82438 34964 82466
rect 35948 82466 35976 87316
rect 36122 87068 36430 87077
rect 36122 87066 36128 87068
rect 36184 87066 36208 87068
rect 36264 87066 36288 87068
rect 36344 87066 36368 87068
rect 36424 87066 36430 87068
rect 36184 87014 36186 87066
rect 36366 87014 36368 87066
rect 36122 87012 36128 87014
rect 36184 87012 36208 87014
rect 36264 87012 36288 87014
rect 36344 87012 36368 87014
rect 36424 87012 36430 87014
rect 36122 87003 36430 87012
rect 36782 86524 37090 86533
rect 36782 86522 36788 86524
rect 36844 86522 36868 86524
rect 36924 86522 36948 86524
rect 37004 86522 37028 86524
rect 37084 86522 37090 86524
rect 36844 86470 36846 86522
rect 37026 86470 37028 86522
rect 36782 86468 36788 86470
rect 36844 86468 36868 86470
rect 36924 86468 36948 86470
rect 37004 86468 37028 86470
rect 37084 86468 37090 86470
rect 36782 86459 37090 86468
rect 36122 85980 36430 85989
rect 36122 85978 36128 85980
rect 36184 85978 36208 85980
rect 36264 85978 36288 85980
rect 36344 85978 36368 85980
rect 36424 85978 36430 85980
rect 36184 85926 36186 85978
rect 36366 85926 36368 85978
rect 36122 85924 36128 85926
rect 36184 85924 36208 85926
rect 36264 85924 36288 85926
rect 36344 85924 36368 85926
rect 36424 85924 36430 85926
rect 36122 85915 36430 85924
rect 36782 85436 37090 85445
rect 36782 85434 36788 85436
rect 36844 85434 36868 85436
rect 36924 85434 36948 85436
rect 37004 85434 37028 85436
rect 37084 85434 37090 85436
rect 36844 85382 36846 85434
rect 37026 85382 37028 85434
rect 36782 85380 36788 85382
rect 36844 85380 36868 85382
rect 36924 85380 36948 85382
rect 37004 85380 37028 85382
rect 37084 85380 37090 85382
rect 36782 85371 37090 85380
rect 36122 84892 36430 84901
rect 36122 84890 36128 84892
rect 36184 84890 36208 84892
rect 36264 84890 36288 84892
rect 36344 84890 36368 84892
rect 36424 84890 36430 84892
rect 36184 84838 36186 84890
rect 36366 84838 36368 84890
rect 36122 84836 36128 84838
rect 36184 84836 36208 84838
rect 36264 84836 36288 84838
rect 36344 84836 36368 84838
rect 36424 84836 36430 84838
rect 36122 84827 36430 84836
rect 36782 84348 37090 84357
rect 36782 84346 36788 84348
rect 36844 84346 36868 84348
rect 36924 84346 36948 84348
rect 37004 84346 37028 84348
rect 37084 84346 37090 84348
rect 36844 84294 36846 84346
rect 37026 84294 37028 84346
rect 36782 84292 36788 84294
rect 36844 84292 36868 84294
rect 36924 84292 36948 84294
rect 37004 84292 37028 84294
rect 37084 84292 37090 84294
rect 36782 84283 37090 84292
rect 37144 82466 37172 87316
rect 35948 82438 36004 82466
rect 34872 82180 34900 82438
rect 35976 82180 36004 82438
rect 37080 82438 37172 82466
rect 38156 82466 38184 87316
rect 39064 87272 39116 87278
rect 39064 87214 39116 87220
rect 39076 84694 39104 87214
rect 39064 84688 39116 84694
rect 39064 84630 39116 84636
rect 39260 82466 39288 87316
rect 39628 84762 39656 88000
rect 40272 87482 40300 88000
rect 40916 87482 40944 88000
rect 40260 87476 40312 87482
rect 40260 87418 40312 87424
rect 40904 87476 40956 87482
rect 40904 87418 40956 87424
rect 40352 87374 40404 87380
rect 40352 87316 40404 87322
rect 39616 84756 39668 84762
rect 39616 84698 39668 84704
rect 40364 82466 40392 87316
rect 41560 86938 41588 88000
rect 42204 87482 42232 88000
rect 42192 87476 42244 87482
rect 42192 87418 42244 87424
rect 42848 87414 42876 88000
rect 43492 87482 43520 88000
rect 44136 87482 44164 88000
rect 43480 87476 43532 87482
rect 43480 87418 43532 87424
rect 44124 87476 44176 87482
rect 44124 87418 44176 87424
rect 44780 87414 44808 88000
rect 45424 87414 45452 88000
rect 46068 87414 46096 88000
rect 46712 87414 46740 88000
rect 47356 87414 47384 88000
rect 48000 87414 48028 88000
rect 48644 87414 48672 88000
rect 49288 87414 49316 88000
rect 49932 87414 49960 88000
rect 50576 87414 50604 88000
rect 52508 87482 52536 88000
rect 52496 87476 52548 87482
rect 52496 87418 52548 87424
rect 53796 87414 53824 88000
rect 42836 87408 42888 87414
rect 42560 87374 42612 87380
rect 44768 87408 44820 87414
rect 42836 87350 42888 87356
rect 43664 87374 43716 87380
rect 42560 87316 42612 87322
rect 43664 87316 43716 87322
rect 44676 87374 44728 87380
rect 44768 87350 44820 87356
rect 45412 87408 45464 87414
rect 45412 87350 45464 87356
rect 46056 87408 46108 87414
rect 46056 87350 46108 87356
rect 46700 87408 46752 87414
rect 46700 87350 46752 87356
rect 47344 87408 47396 87414
rect 47344 87350 47396 87356
rect 47988 87408 48040 87414
rect 47988 87350 48040 87356
rect 48632 87408 48684 87414
rect 48632 87350 48684 87356
rect 49276 87408 49328 87414
rect 49276 87350 49328 87356
rect 49920 87408 49972 87414
rect 49920 87350 49972 87356
rect 50564 87408 50616 87414
rect 50564 87350 50616 87356
rect 53784 87408 53836 87414
rect 54440 87380 54468 88000
rect 55182 87612 55490 87621
rect 55182 87610 55188 87612
rect 55244 87610 55268 87612
rect 55324 87610 55348 87612
rect 55404 87610 55428 87612
rect 55484 87610 55490 87612
rect 55244 87558 55246 87610
rect 55426 87558 55428 87610
rect 55182 87556 55188 87558
rect 55244 87556 55268 87558
rect 55324 87556 55348 87558
rect 55404 87556 55428 87558
rect 55484 87556 55490 87558
rect 55182 87547 55490 87556
rect 55728 87482 55756 88000
rect 57016 87482 57044 88000
rect 57660 87482 57688 88000
rect 55716 87476 55768 87482
rect 55716 87418 55768 87424
rect 57004 87476 57056 87482
rect 57004 87418 57056 87424
rect 57648 87476 57700 87482
rect 57648 87418 57700 87424
rect 58948 87414 58976 88000
rect 60236 87482 60264 88000
rect 60224 87476 60276 87482
rect 60224 87418 60276 87424
rect 61524 87414 61552 88000
rect 58936 87408 58988 87414
rect 53784 87350 53836 87356
rect 54428 87374 54480 87380
rect 44676 87316 44728 87322
rect 58936 87350 58988 87356
rect 61512 87408 61564 87414
rect 62168 87380 62196 88000
rect 63456 87482 63484 88000
rect 64744 87482 64772 88000
rect 65388 87482 65416 88000
rect 63444 87476 63496 87482
rect 63444 87418 63496 87424
rect 64732 87476 64784 87482
rect 64732 87418 64784 87424
rect 65376 87476 65428 87482
rect 65376 87418 65428 87424
rect 66676 87414 66704 88000
rect 67964 87482 67992 88000
rect 69252 87482 69280 88000
rect 69896 87482 69924 88000
rect 71184 87482 71212 88000
rect 72472 87482 72500 88000
rect 73116 87482 73144 88000
rect 73582 87612 73890 87621
rect 73582 87610 73588 87612
rect 73644 87610 73668 87612
rect 73724 87610 73748 87612
rect 73804 87610 73828 87612
rect 73884 87610 73890 87612
rect 73644 87558 73646 87610
rect 73826 87558 73828 87610
rect 73582 87556 73588 87558
rect 73644 87556 73668 87558
rect 73724 87556 73748 87558
rect 73804 87556 73828 87558
rect 73884 87556 73890 87558
rect 73582 87547 73890 87556
rect 74404 87482 74432 88000
rect 75692 87482 75720 88000
rect 76980 87482 77008 88000
rect 77624 87482 77652 88000
rect 78912 87482 78940 88000
rect 80200 87482 80228 88000
rect 80844 87482 80872 88000
rect 82132 87482 82160 88000
rect 67952 87476 68004 87482
rect 67952 87418 68004 87424
rect 69240 87476 69292 87482
rect 69240 87418 69292 87424
rect 69884 87476 69936 87482
rect 69884 87418 69936 87424
rect 71172 87476 71224 87482
rect 71172 87418 71224 87424
rect 72460 87476 72512 87482
rect 72460 87418 72512 87424
rect 73104 87476 73156 87482
rect 73104 87418 73156 87424
rect 74392 87476 74444 87482
rect 74392 87418 74444 87424
rect 75680 87476 75732 87482
rect 75680 87418 75732 87424
rect 76968 87476 77020 87482
rect 76968 87418 77020 87424
rect 77612 87476 77664 87482
rect 77612 87418 77664 87424
rect 78900 87476 78952 87482
rect 78900 87418 78952 87424
rect 80188 87476 80240 87482
rect 80188 87418 80240 87424
rect 80832 87476 80884 87482
rect 80832 87418 80884 87424
rect 82120 87476 82172 87482
rect 82120 87418 82172 87424
rect 66664 87408 66716 87414
rect 61512 87350 61564 87356
rect 62156 87374 62208 87380
rect 54428 87316 54480 87322
rect 60132 87340 60184 87346
rect 41824 87204 41876 87210
rect 41824 87146 41876 87152
rect 41548 86932 41600 86938
rect 41548 86874 41600 86880
rect 41456 86762 41508 86768
rect 41456 86704 41508 86710
rect 41468 82466 41496 86704
rect 41836 85034 41864 87146
rect 41824 85028 41876 85034
rect 41824 84970 41876 84976
rect 41836 84626 41864 84970
rect 41824 84620 41876 84626
rect 41824 84562 41876 84568
rect 42572 82466 42600 87316
rect 43676 82466 43704 87316
rect 44688 85794 44716 87316
rect 66664 87350 66716 87356
rect 67860 87374 67912 87380
rect 62156 87316 62208 87322
rect 67860 87316 67912 87322
rect 69332 87374 69384 87380
rect 69332 87316 69384 87322
rect 70068 87374 70120 87380
rect 70068 87316 70120 87322
rect 71172 87374 71224 87380
rect 71172 87316 71224 87322
rect 72276 87374 72328 87380
rect 72276 87316 72328 87322
rect 73380 87374 73432 87380
rect 73380 87316 73432 87322
rect 74484 87374 74536 87380
rect 74484 87316 74536 87322
rect 75588 87374 75640 87380
rect 77796 87374 77848 87380
rect 75588 87316 75640 87322
rect 76692 87340 76744 87346
rect 60132 87282 60184 87288
rect 56820 87272 56872 87278
rect 56820 87214 56872 87220
rect 52680 87204 52732 87210
rect 52680 87146 52732 87152
rect 53508 87204 53560 87210
rect 53508 87146 53560 87152
rect 54428 87204 54480 87210
rect 54428 87146 54480 87152
rect 55716 87204 55768 87210
rect 55716 87146 55768 87152
rect 44688 85766 44808 85794
rect 44780 82466 44808 85766
rect 49092 85028 49144 85034
rect 49092 84970 49144 84976
rect 46148 84756 46200 84762
rect 46148 84698 46200 84704
rect 46160 84626 46188 84698
rect 46056 84620 46108 84626
rect 46056 84562 46108 84568
rect 46148 84620 46200 84626
rect 46148 84562 46200 84568
rect 45872 84484 45924 84490
rect 45872 84426 45924 84432
rect 45964 84484 46016 84490
rect 45964 84426 46016 84432
rect 38156 82438 38212 82466
rect 39260 82438 39316 82466
rect 40364 82438 40420 82466
rect 41468 82438 41524 82466
rect 42572 82438 42628 82466
rect 43676 82438 43732 82466
rect 44780 82438 44836 82466
rect 37080 82180 37108 82438
rect 38184 82180 38212 82438
rect 39288 82180 39316 82438
rect 40392 82180 40420 82438
rect 41496 82180 41524 82438
rect 42600 82180 42628 82438
rect 43704 82180 43732 82438
rect 44808 82180 44836 82438
rect 9990 82072 10046 82081
rect 9990 82007 10046 82016
rect 10542 82072 10598 82081
rect 10542 82007 10598 82016
rect 10004 81770 10032 82007
rect 7784 81764 7836 81770
rect 7784 81706 7836 81712
rect 9992 81764 10044 81770
rect 9992 81706 10044 81712
rect 7796 63818 7824 81706
rect 9624 63948 9676 63954
rect 9624 63890 9676 63896
rect 7784 63812 7836 63818
rect 7784 63754 7836 63760
rect 9636 63653 9664 63890
rect 9622 63644 9678 63653
rect 9622 63579 9678 63588
rect 45884 49509 45912 84426
rect 45976 50597 46004 84426
rect 45962 50588 46018 50597
rect 45962 50523 46018 50532
rect 45870 49500 45926 49509
rect 45870 49435 45926 49444
rect 7520 47126 7640 47154
rect 7324 45588 7376 45594
rect 7324 45530 7376 45536
rect 7140 45520 7192 45526
rect 7138 45488 7140 45497
rect 7192 45488 7194 45497
rect 7138 45423 7194 45432
rect 2908 45384 2960 45390
rect 7520 45361 7548 47126
rect 13884 45928 13936 45934
rect 13884 45870 13936 45876
rect 14972 45882 15000 46548
rect 16076 45882 16104 46548
rect 17180 45882 17208 46548
rect 18284 45882 18312 46548
rect 19388 45882 19416 46548
rect 20492 45882 20520 46548
rect 21596 45882 21624 46548
rect 22700 45882 22728 46548
rect 23804 45882 23832 46548
rect 24908 45882 24936 46548
rect 26012 45882 26040 46548
rect 27116 45882 27144 46548
rect 28220 45882 28248 46548
rect 29324 45882 29352 46548
rect 30428 45882 30456 46548
rect 31532 45882 31560 46548
rect 32636 45882 32664 46548
rect 33740 45882 33768 46548
rect 34844 45882 34872 46548
rect 35948 45882 35976 46548
rect 37052 45882 37080 46548
rect 38156 45882 38184 46548
rect 39260 45882 39288 46548
rect 40364 45882 40392 46548
rect 41468 45882 41496 46548
rect 42572 45882 42600 46548
rect 43676 45882 43704 46548
rect 44780 45882 44808 46548
rect 13896 45732 13924 45870
rect 14972 45854 15028 45882
rect 16076 45854 16132 45882
rect 17180 45854 17236 45882
rect 18284 45854 18340 45882
rect 19388 45854 19444 45882
rect 20492 45854 20548 45882
rect 21596 45854 21652 45882
rect 22700 45854 22756 45882
rect 23804 45854 23860 45882
rect 24908 45854 24964 45882
rect 26012 45854 26068 45882
rect 27116 45854 27172 45882
rect 28220 45854 28276 45882
rect 29324 45854 29380 45882
rect 30428 45854 30484 45882
rect 31532 45854 31588 45882
rect 32636 45854 32692 45882
rect 33740 45854 33796 45882
rect 34844 45854 34900 45882
rect 35948 45854 36004 45882
rect 37052 45854 37108 45882
rect 38156 45854 38212 45882
rect 39260 45854 39316 45882
rect 40364 45854 40420 45882
rect 41468 45854 41524 45882
rect 42572 45854 42628 45882
rect 43676 45854 43732 45882
rect 44780 45854 44836 45882
rect 15000 45732 15028 45854
rect 16104 45732 16132 45854
rect 17208 45732 17236 45854
rect 18312 45732 18340 45854
rect 19416 45732 19444 45854
rect 20520 45732 20548 45854
rect 21624 45732 21652 45854
rect 22728 45732 22756 45854
rect 23832 45732 23860 45854
rect 24936 45732 24964 45854
rect 26040 45732 26068 45854
rect 27144 45732 27172 45854
rect 28248 45732 28276 45854
rect 29352 45732 29380 45854
rect 30456 45732 30484 45854
rect 31560 45732 31588 45854
rect 32664 45732 32692 45854
rect 33768 45732 33796 45854
rect 34872 45732 34900 45854
rect 35976 45732 36004 45854
rect 37080 45732 37108 45854
rect 38184 45732 38212 45854
rect 39288 45732 39316 45854
rect 40392 45732 40420 45854
rect 41496 45732 41524 45854
rect 42600 45732 42628 45854
rect 43704 45732 43732 45854
rect 44808 45732 44836 45854
rect 9990 45624 10046 45633
rect 9990 45559 9992 45568
rect 10044 45559 10046 45568
rect 10542 45624 10598 45633
rect 10542 45559 10598 45568
rect 9992 45530 10044 45536
rect 12778 45488 12834 45497
rect 12778 45423 12834 45432
rect 2908 45326 2960 45332
rect 7506 45352 7562 45361
rect 2920 45225 2948 45326
rect 7506 45287 7562 45296
rect 11674 45352 11730 45361
rect 11674 45287 11730 45296
rect 2906 45216 2962 45225
rect 2906 45151 2962 45160
rect 6690 45180 6998 45189
rect 6690 45178 6696 45180
rect 6752 45178 6776 45180
rect 6832 45178 6856 45180
rect 6912 45178 6936 45180
rect 6992 45178 6998 45180
rect 6752 45126 6754 45178
rect 6934 45126 6936 45178
rect 6690 45124 6696 45126
rect 6752 45124 6776 45126
rect 6832 45124 6856 45126
rect 6912 45124 6936 45126
rect 6992 45124 6998 45126
rect 6690 45115 6998 45124
rect 7520 45050 7548 45287
rect 7508 45044 7560 45050
rect 7508 44986 7560 44992
rect 7140 44908 7192 44914
rect 7140 44850 7192 44856
rect 2908 44772 2960 44778
rect 2908 44714 2960 44720
rect 2920 44545 2948 44714
rect 7152 44681 7180 44850
rect 7138 44672 7194 44681
rect 5954 44636 6262 44645
rect 5954 44634 5960 44636
rect 6016 44634 6040 44636
rect 6096 44634 6120 44636
rect 6176 44634 6200 44636
rect 6256 44634 6262 44636
rect 6016 44582 6018 44634
rect 6198 44582 6200 44634
rect 7138 44607 7194 44616
rect 5954 44580 5960 44582
rect 6016 44580 6040 44582
rect 6096 44580 6120 44582
rect 6176 44580 6200 44582
rect 6256 44580 6262 44582
rect 5954 44571 6262 44580
rect 2906 44536 2962 44545
rect 2906 44471 2962 44480
rect 8152 44296 8204 44302
rect 8152 44238 8204 44244
rect 2724 44228 2776 44234
rect 2724 44170 2776 44176
rect 2736 43865 2764 44170
rect 6690 44092 6998 44101
rect 6690 44090 6696 44092
rect 6752 44090 6776 44092
rect 6832 44090 6856 44092
rect 6912 44090 6936 44092
rect 6992 44090 6998 44092
rect 6752 44038 6754 44090
rect 6934 44038 6936 44090
rect 6690 44036 6696 44038
rect 6752 44036 6776 44038
rect 6832 44036 6856 44038
rect 6912 44036 6936 44038
rect 6992 44036 6998 44038
rect 6690 44027 6998 44036
rect 2722 43856 2778 43865
rect 2722 43791 2778 43800
rect 8164 43593 8192 44238
rect 8150 43584 8206 43593
rect 5954 43548 6262 43557
rect 5954 43546 5960 43548
rect 6016 43546 6040 43548
rect 6096 43546 6120 43548
rect 6176 43546 6200 43548
rect 6256 43546 6262 43548
rect 6016 43494 6018 43546
rect 6198 43494 6200 43546
rect 8150 43519 8206 43528
rect 5954 43492 5960 43494
rect 6016 43492 6040 43494
rect 6096 43492 6120 43494
rect 6176 43492 6200 43494
rect 6256 43492 6262 43494
rect 5954 43483 6262 43492
rect 6690 43004 6998 43013
rect 6690 43002 6696 43004
rect 6752 43002 6776 43004
rect 6832 43002 6856 43004
rect 6912 43002 6936 43004
rect 6992 43002 6998 43004
rect 6752 42950 6754 43002
rect 6934 42950 6936 43002
rect 6690 42948 6696 42950
rect 6752 42948 6776 42950
rect 6832 42948 6856 42950
rect 6912 42948 6936 42950
rect 6992 42948 6998 42950
rect 6690 42939 6998 42948
rect 7140 42732 7192 42738
rect 7140 42674 7192 42680
rect 2908 42596 2960 42602
rect 2908 42538 2960 42544
rect 2920 42505 2948 42538
rect 7152 42505 7180 42674
rect 2906 42496 2962 42505
rect 7138 42496 7194 42505
rect 2906 42431 2962 42440
rect 5954 42460 6262 42469
rect 5954 42458 5960 42460
rect 6016 42458 6040 42460
rect 6096 42458 6120 42460
rect 6176 42458 6200 42460
rect 6256 42458 6262 42460
rect 6016 42406 6018 42458
rect 6198 42406 6200 42458
rect 7138 42431 7194 42440
rect 5954 42404 5960 42406
rect 6016 42404 6040 42406
rect 6096 42404 6120 42406
rect 6176 42404 6200 42406
rect 6256 42404 6262 42406
rect 5954 42395 6262 42404
rect 6690 41916 6998 41925
rect 6690 41914 6696 41916
rect 6752 41914 6776 41916
rect 6832 41914 6856 41916
rect 6912 41914 6936 41916
rect 6992 41914 6998 41916
rect 6752 41862 6754 41914
rect 6934 41862 6936 41914
rect 6690 41860 6696 41862
rect 6752 41860 6776 41862
rect 6832 41860 6856 41862
rect 6912 41860 6936 41862
rect 6992 41860 6998 41862
rect 6690 41851 6998 41860
rect 4380 41780 4432 41786
rect 4380 41722 4432 41728
rect 4392 41145 4420 41722
rect 5668 41678 5720 41684
rect 5668 41620 5720 41626
rect 5680 41553 5708 41620
rect 5666 41544 5722 41553
rect 5666 41479 5722 41488
rect 5954 41372 6262 41381
rect 5954 41370 5960 41372
rect 6016 41370 6040 41372
rect 6096 41370 6120 41372
rect 6176 41370 6200 41372
rect 6256 41370 6262 41372
rect 6016 41318 6018 41370
rect 6198 41318 6200 41370
rect 5954 41316 5960 41318
rect 6016 41316 6040 41318
rect 6096 41316 6120 41318
rect 6176 41316 6200 41318
rect 6256 41316 6262 41318
rect 5954 41307 6262 41316
rect 4378 41136 4434 41145
rect 4378 41071 4434 41080
rect 6690 40828 6998 40837
rect 6690 40826 6696 40828
rect 6752 40826 6776 40828
rect 6832 40826 6856 40828
rect 6912 40826 6936 40828
rect 6992 40826 6998 40828
rect 6752 40774 6754 40826
rect 6934 40774 6936 40826
rect 6690 40772 6696 40774
rect 6752 40772 6776 40774
rect 6832 40772 6856 40774
rect 6912 40772 6936 40774
rect 6992 40772 6998 40774
rect 6690 40763 6998 40772
rect 7140 40556 7192 40562
rect 7140 40498 7192 40504
rect 2906 40456 2962 40465
rect 2906 40391 2908 40400
rect 2960 40391 2962 40400
rect 2908 40362 2960 40368
rect 7152 40329 7180 40498
rect 7138 40320 7194 40329
rect 5954 40284 6262 40293
rect 5954 40282 5960 40284
rect 6016 40282 6040 40284
rect 6096 40282 6120 40284
rect 6176 40282 6200 40284
rect 6256 40282 6262 40284
rect 6016 40230 6018 40282
rect 6198 40230 6200 40282
rect 7138 40255 7194 40264
rect 5954 40228 5960 40230
rect 6016 40228 6040 40230
rect 6096 40228 6120 40230
rect 6176 40228 6200 40230
rect 6256 40228 6262 40230
rect 5954 40219 6262 40228
rect 6690 39740 6998 39749
rect 6690 39738 6696 39740
rect 6752 39738 6776 39740
rect 6832 39738 6856 39740
rect 6912 39738 6936 39740
rect 6992 39738 6998 39740
rect 6752 39686 6754 39738
rect 6934 39686 6936 39738
rect 6690 39684 6696 39686
rect 6752 39684 6776 39686
rect 6832 39684 6856 39686
rect 6912 39684 6936 39686
rect 6992 39684 6998 39686
rect 6690 39675 6998 39684
rect 7140 39468 7192 39474
rect 7140 39410 7192 39416
rect 2908 39332 2960 39338
rect 2908 39274 2960 39280
rect 2920 39105 2948 39274
rect 7152 39241 7180 39410
rect 7138 39232 7194 39241
rect 5954 39196 6262 39205
rect 5954 39194 5960 39196
rect 6016 39194 6040 39196
rect 6096 39194 6120 39196
rect 6176 39194 6200 39196
rect 6256 39194 6262 39196
rect 6016 39142 6018 39194
rect 6198 39142 6200 39194
rect 7138 39167 7194 39176
rect 5954 39140 5960 39142
rect 6016 39140 6040 39142
rect 6096 39140 6120 39142
rect 6176 39140 6200 39142
rect 6256 39140 6262 39142
rect 5954 39131 6262 39140
rect 2906 39096 2962 39105
rect 2906 39031 2962 39040
rect 4380 38992 4432 38998
rect 4380 38934 4432 38940
rect 4392 38425 4420 38934
rect 7784 38856 7836 38862
rect 7784 38798 7836 38804
rect 6690 38652 6998 38661
rect 6690 38650 6696 38652
rect 6752 38650 6776 38652
rect 6832 38650 6856 38652
rect 6912 38650 6936 38652
rect 6992 38650 6998 38652
rect 6752 38598 6754 38650
rect 6934 38598 6936 38650
rect 6690 38596 6696 38598
rect 6752 38596 6776 38598
rect 6832 38596 6856 38598
rect 6912 38596 6936 38598
rect 6992 38596 6998 38598
rect 6690 38587 6998 38596
rect 4378 38416 4434 38425
rect 4378 38351 4434 38360
rect 7796 38153 7824 38798
rect 7782 38144 7838 38153
rect 5954 38108 6262 38117
rect 5954 38106 5960 38108
rect 6016 38106 6040 38108
rect 6096 38106 6120 38108
rect 6176 38106 6200 38108
rect 6256 38106 6262 38108
rect 6016 38054 6018 38106
rect 6198 38054 6200 38106
rect 7782 38079 7838 38088
rect 5954 38052 5960 38054
rect 6016 38052 6040 38054
rect 6096 38052 6120 38054
rect 6176 38052 6200 38054
rect 6256 38052 6262 38054
rect 5954 38043 6262 38052
rect 6690 37564 6998 37573
rect 6690 37562 6696 37564
rect 6752 37562 6776 37564
rect 6832 37562 6856 37564
rect 6912 37562 6936 37564
rect 6992 37562 6998 37564
rect 6752 37510 6754 37562
rect 6934 37510 6936 37562
rect 6690 37508 6696 37510
rect 6752 37508 6776 37510
rect 6832 37508 6856 37510
rect 6912 37508 6936 37510
rect 6992 37508 6998 37510
rect 6690 37499 6998 37508
rect 7232 37292 7284 37298
rect 7232 37234 7284 37240
rect 2908 37156 2960 37162
rect 2908 37098 2960 37104
rect 2920 37065 2948 37098
rect 7244 37065 7272 37234
rect 2906 37056 2962 37065
rect 7230 37056 7286 37065
rect 2906 36991 2962 37000
rect 5954 37020 6262 37029
rect 5954 37018 5960 37020
rect 6016 37018 6040 37020
rect 6096 37018 6120 37020
rect 6176 37018 6200 37020
rect 6256 37018 6262 37020
rect 6016 36966 6018 37018
rect 6198 36966 6200 37018
rect 7230 36991 7286 37000
rect 5954 36964 5960 36966
rect 6016 36964 6040 36966
rect 6096 36964 6120 36966
rect 6176 36964 6200 36966
rect 6256 36964 6262 36966
rect 5954 36955 6262 36964
rect 6690 36476 6998 36485
rect 6690 36474 6696 36476
rect 6752 36474 6776 36476
rect 6832 36474 6856 36476
rect 6912 36474 6936 36476
rect 6992 36474 6998 36476
rect 6752 36422 6754 36474
rect 6934 36422 6936 36474
rect 6690 36420 6696 36422
rect 6752 36420 6776 36422
rect 6832 36420 6856 36422
rect 6912 36420 6936 36422
rect 6992 36420 6998 36422
rect 6690 36411 6998 36420
rect 5668 36238 5720 36244
rect 5668 36180 5720 36186
rect 4380 36136 4432 36142
rect 5680 36113 5708 36180
rect 4380 36078 4432 36084
rect 5666 36104 5722 36113
rect 4392 35705 4420 36078
rect 5666 36039 5722 36048
rect 5954 35932 6262 35941
rect 5954 35930 5960 35932
rect 6016 35930 6040 35932
rect 6096 35930 6120 35932
rect 6176 35930 6200 35932
rect 6256 35930 6262 35932
rect 6016 35878 6018 35930
rect 6198 35878 6200 35930
rect 5954 35876 5960 35878
rect 6016 35876 6040 35878
rect 6096 35876 6120 35878
rect 6176 35876 6200 35878
rect 6256 35876 6262 35878
rect 5954 35867 6262 35876
rect 4378 35696 4434 35705
rect 4378 35631 4434 35640
rect 6690 35388 6998 35397
rect 6690 35386 6696 35388
rect 6752 35386 6776 35388
rect 6832 35386 6856 35388
rect 6912 35386 6936 35388
rect 6992 35386 6998 35388
rect 6752 35334 6754 35386
rect 6934 35334 6936 35386
rect 6690 35332 6696 35334
rect 6752 35332 6776 35334
rect 6832 35332 6856 35334
rect 6912 35332 6936 35334
rect 6992 35332 6998 35334
rect 6690 35323 6998 35332
rect 7232 35116 7284 35122
rect 7232 35058 7284 35064
rect 2906 35016 2962 35025
rect 2906 34951 2908 34960
rect 2960 34951 2962 34960
rect 2908 34922 2960 34928
rect 7244 34889 7272 35058
rect 7230 34880 7286 34889
rect 5954 34844 6262 34853
rect 5954 34842 5960 34844
rect 6016 34842 6040 34844
rect 6096 34842 6120 34844
rect 6176 34842 6200 34844
rect 6256 34842 6262 34844
rect 6016 34790 6018 34842
rect 6198 34790 6200 34842
rect 7230 34815 7286 34824
rect 5954 34788 5960 34790
rect 6016 34788 6040 34790
rect 6096 34788 6120 34790
rect 6176 34788 6200 34790
rect 6256 34788 6262 34790
rect 5954 34779 6262 34788
rect 6690 34300 6998 34309
rect 6690 34298 6696 34300
rect 6752 34298 6776 34300
rect 6832 34298 6856 34300
rect 6912 34298 6936 34300
rect 6992 34298 6998 34300
rect 6752 34246 6754 34298
rect 6934 34246 6936 34298
rect 6690 34244 6696 34246
rect 6752 34244 6776 34246
rect 6832 34244 6856 34246
rect 6912 34244 6936 34246
rect 6992 34244 6998 34246
rect 6690 34235 6998 34244
rect 7232 34028 7284 34034
rect 7232 33970 7284 33976
rect 2908 33892 2960 33898
rect 2908 33834 2960 33840
rect 2920 33665 2948 33834
rect 7244 33801 7272 33970
rect 7230 33792 7286 33801
rect 5954 33756 6262 33765
rect 5954 33754 5960 33756
rect 6016 33754 6040 33756
rect 6096 33754 6120 33756
rect 6176 33754 6200 33756
rect 6256 33754 6262 33756
rect 6016 33702 6018 33754
rect 6198 33702 6200 33754
rect 7230 33727 7286 33736
rect 5954 33700 5960 33702
rect 6016 33700 6040 33702
rect 6096 33700 6120 33702
rect 6176 33700 6200 33702
rect 6256 33700 6262 33702
rect 5954 33691 6262 33700
rect 2906 33656 2962 33665
rect 2906 33591 2962 33600
rect 4380 33552 4432 33558
rect 4380 33494 4432 33500
rect 4392 32985 4420 33494
rect 5668 33450 5720 33456
rect 5668 33392 5720 33398
rect 5680 32985 5708 33392
rect 6690 33212 6998 33221
rect 6690 33210 6696 33212
rect 6752 33210 6776 33212
rect 6832 33210 6856 33212
rect 6912 33210 6936 33212
rect 6992 33210 6998 33212
rect 6752 33158 6754 33210
rect 6934 33158 6936 33210
rect 6690 33156 6696 33158
rect 6752 33156 6776 33158
rect 6832 33156 6856 33158
rect 6912 33156 6936 33158
rect 6992 33156 6998 33158
rect 6690 33147 6998 33156
rect 4378 32976 4434 32985
rect 4378 32911 4434 32920
rect 5666 32976 5722 32985
rect 5666 32911 5722 32920
rect 5954 32668 6262 32677
rect 5954 32666 5960 32668
rect 6016 32666 6040 32668
rect 6096 32666 6120 32668
rect 6176 32666 6200 32668
rect 6256 32666 6262 32668
rect 6016 32614 6018 32666
rect 6198 32614 6200 32666
rect 5954 32612 5960 32614
rect 6016 32612 6040 32614
rect 6096 32612 6120 32614
rect 6176 32612 6200 32614
rect 6256 32612 6262 32614
rect 5954 32603 6262 32612
rect 6690 32124 6998 32133
rect 6690 32122 6696 32124
rect 6752 32122 6776 32124
rect 6832 32122 6856 32124
rect 6912 32122 6936 32124
rect 6992 32122 6998 32124
rect 6752 32070 6754 32122
rect 6934 32070 6936 32122
rect 6690 32068 6696 32070
rect 6752 32068 6776 32070
rect 6832 32068 6856 32070
rect 6912 32068 6936 32070
rect 6992 32068 6998 32070
rect 6690 32059 6998 32068
rect 7232 31852 7284 31858
rect 7232 31794 7284 31800
rect 2908 31716 2960 31722
rect 2908 31658 2960 31664
rect 2920 31625 2948 31658
rect 7244 31625 7272 31794
rect 2906 31616 2962 31625
rect 7230 31616 7286 31625
rect 2906 31551 2962 31560
rect 5954 31580 6262 31589
rect 5954 31578 5960 31580
rect 6016 31578 6040 31580
rect 6096 31578 6120 31580
rect 6176 31578 6200 31580
rect 6256 31578 6262 31580
rect 6016 31526 6018 31578
rect 6198 31526 6200 31578
rect 7230 31551 7286 31560
rect 5954 31524 5960 31526
rect 6016 31524 6040 31526
rect 6096 31524 6120 31526
rect 6176 31524 6200 31526
rect 6256 31524 6262 31526
rect 5954 31515 6262 31524
rect 6690 31036 6998 31045
rect 6690 31034 6696 31036
rect 6752 31034 6776 31036
rect 6832 31034 6856 31036
rect 6912 31034 6936 31036
rect 6992 31034 6998 31036
rect 6752 30982 6754 31034
rect 6934 30982 6936 31034
rect 6690 30980 6696 30982
rect 6752 30980 6776 30982
rect 6832 30980 6856 30982
rect 6912 30980 6936 30982
rect 6992 30980 6998 30982
rect 6690 30971 6998 30980
rect 5668 30798 5720 30804
rect 5668 30740 5720 30746
rect 4380 30628 4432 30634
rect 4380 30570 4432 30576
rect 4392 30265 4420 30570
rect 5680 30265 5708 30740
rect 5954 30492 6262 30501
rect 5954 30490 5960 30492
rect 6016 30490 6040 30492
rect 6096 30490 6120 30492
rect 6176 30490 6200 30492
rect 6256 30490 6262 30492
rect 6016 30438 6018 30490
rect 6198 30438 6200 30490
rect 5954 30436 5960 30438
rect 6016 30436 6040 30438
rect 6096 30436 6120 30438
rect 6176 30436 6200 30438
rect 6256 30436 6262 30438
rect 5954 30427 6262 30436
rect 4378 30256 4434 30265
rect 4378 30191 4434 30200
rect 5666 30256 5722 30265
rect 5666 30191 5722 30200
rect 6690 29948 6998 29957
rect 6690 29946 6696 29948
rect 6752 29946 6776 29948
rect 6832 29946 6856 29948
rect 6912 29946 6936 29948
rect 6992 29946 6998 29948
rect 6752 29894 6754 29946
rect 6934 29894 6936 29946
rect 6690 29892 6696 29894
rect 6752 29892 6776 29894
rect 6832 29892 6856 29894
rect 6912 29892 6936 29894
rect 6992 29892 6998 29894
rect 6690 29883 6998 29892
rect 2908 29676 2960 29682
rect 2908 29618 2960 29624
rect 2920 29585 2948 29618
rect 7232 29608 7284 29614
rect 2906 29576 2962 29585
rect 7232 29550 7284 29556
rect 2906 29511 2962 29520
rect 7244 29449 7272 29550
rect 7230 29440 7286 29449
rect 5954 29404 6262 29413
rect 5954 29402 5960 29404
rect 6016 29402 6040 29404
rect 6096 29402 6120 29404
rect 6176 29402 6200 29404
rect 6256 29402 6262 29404
rect 6016 29350 6018 29402
rect 6198 29350 6200 29402
rect 7230 29375 7286 29384
rect 5954 29348 5960 29350
rect 6016 29348 6040 29350
rect 6096 29348 6120 29350
rect 6176 29348 6200 29350
rect 6256 29348 6262 29350
rect 5954 29339 6262 29348
rect 6690 28860 6998 28869
rect 6690 28858 6696 28860
rect 6752 28858 6776 28860
rect 6832 28858 6856 28860
rect 6912 28858 6936 28860
rect 6992 28858 6998 28860
rect 6752 28806 6754 28858
rect 6934 28806 6936 28858
rect 6690 28804 6696 28806
rect 6752 28804 6776 28806
rect 6832 28804 6856 28806
rect 6912 28804 6936 28806
rect 6992 28804 6998 28806
rect 6690 28795 6998 28804
rect 2908 28588 2960 28594
rect 2908 28530 2960 28536
rect 2920 28225 2948 28530
rect 7232 28520 7284 28526
rect 7232 28462 7284 28468
rect 7244 28361 7272 28462
rect 7230 28352 7286 28361
rect 5954 28316 6262 28325
rect 5954 28314 5960 28316
rect 6016 28314 6040 28316
rect 6096 28314 6120 28316
rect 6176 28314 6200 28316
rect 6256 28314 6262 28316
rect 6016 28262 6018 28314
rect 6198 28262 6200 28314
rect 7230 28287 7286 28296
rect 5954 28260 5960 28262
rect 6016 28260 6040 28262
rect 6096 28260 6120 28262
rect 6176 28260 6200 28262
rect 6256 28260 6262 28262
rect 5954 28251 6262 28260
rect 2906 28216 2962 28225
rect 2906 28151 2962 28160
rect 5116 28112 5168 28118
rect 5116 28054 5168 28060
rect 5128 27545 5156 28054
rect 5392 27908 5444 27914
rect 5392 27850 5444 27856
rect 5404 27545 5432 27850
rect 6690 27772 6998 27781
rect 6690 27770 6696 27772
rect 6752 27770 6776 27772
rect 6832 27770 6856 27772
rect 6912 27770 6936 27772
rect 6992 27770 6998 27772
rect 6752 27718 6754 27770
rect 6934 27718 6936 27770
rect 6690 27716 6696 27718
rect 6752 27716 6776 27718
rect 6832 27716 6856 27718
rect 6912 27716 6936 27718
rect 6992 27716 6998 27718
rect 6690 27707 6998 27716
rect 5114 27536 5170 27545
rect 5114 27471 5170 27480
rect 5390 27536 5446 27545
rect 5390 27471 5446 27480
rect 5954 27228 6262 27237
rect 5954 27226 5960 27228
rect 6016 27226 6040 27228
rect 6096 27226 6120 27228
rect 6176 27226 6200 27228
rect 6256 27226 6262 27228
rect 6016 27174 6018 27226
rect 6198 27174 6200 27226
rect 5954 27172 5960 27174
rect 6016 27172 6040 27174
rect 6096 27172 6120 27174
rect 6176 27172 6200 27174
rect 6256 27172 6262 27174
rect 5954 27163 6262 27172
rect 6690 26684 6998 26693
rect 6690 26682 6696 26684
rect 6752 26682 6776 26684
rect 6832 26682 6856 26684
rect 6912 26682 6936 26684
rect 6992 26682 6998 26684
rect 6752 26630 6754 26682
rect 6934 26630 6936 26682
rect 6690 26628 6696 26630
rect 6752 26628 6776 26630
rect 6832 26628 6856 26630
rect 6912 26628 6936 26630
rect 6992 26628 6998 26630
rect 6690 26619 6998 26628
rect 2908 26412 2960 26418
rect 2908 26354 2960 26360
rect 2920 26185 2948 26354
rect 7140 26344 7192 26350
rect 7140 26286 7192 26292
rect 7152 26185 7180 26286
rect 2906 26176 2962 26185
rect 7138 26176 7194 26185
rect 2906 26111 2962 26120
rect 5954 26140 6262 26149
rect 5954 26138 5960 26140
rect 6016 26138 6040 26140
rect 6096 26138 6120 26140
rect 6176 26138 6200 26140
rect 6256 26138 6262 26140
rect 6016 26086 6018 26138
rect 6198 26086 6200 26138
rect 7138 26111 7194 26120
rect 5954 26084 5960 26086
rect 6016 26084 6040 26086
rect 6096 26084 6120 26086
rect 6176 26084 6200 26086
rect 6256 26084 6262 26086
rect 5954 26075 6262 26084
rect 6690 25596 6998 25605
rect 6690 25594 6696 25596
rect 6752 25594 6776 25596
rect 6832 25594 6856 25596
rect 6912 25594 6936 25596
rect 6992 25594 6998 25596
rect 6752 25542 6754 25594
rect 6934 25542 6936 25594
rect 6690 25540 6696 25542
rect 6752 25540 6776 25542
rect 6832 25540 6856 25542
rect 6912 25540 6936 25542
rect 6992 25540 6998 25542
rect 6690 25531 6998 25540
rect 4932 25358 4984 25364
rect 4932 25300 4984 25306
rect 4944 24825 4972 25300
rect 7140 25256 7192 25262
rect 7140 25198 7192 25204
rect 7152 25097 7180 25198
rect 7138 25088 7194 25097
rect 5954 25052 6262 25061
rect 5954 25050 5960 25052
rect 6016 25050 6040 25052
rect 6096 25050 6120 25052
rect 6176 25050 6200 25052
rect 6256 25050 6262 25052
rect 6016 24998 6018 25050
rect 6198 24998 6200 25050
rect 7138 25023 7194 25032
rect 5954 24996 5960 24998
rect 6016 24996 6040 24998
rect 6096 24996 6120 24998
rect 6176 24996 6200 24998
rect 6256 24996 6262 24998
rect 5954 24987 6262 24996
rect 4930 24816 4986 24825
rect 4930 24751 4986 24760
rect 6690 24508 6998 24517
rect 6690 24506 6696 24508
rect 6752 24506 6776 24508
rect 6832 24506 6856 24508
rect 6912 24506 6936 24508
rect 6992 24506 6998 24508
rect 6752 24454 6754 24506
rect 6934 24454 6936 24506
rect 6690 24452 6696 24454
rect 6752 24452 6776 24454
rect 6832 24452 6856 24454
rect 6912 24452 6936 24454
rect 6992 24452 6998 24454
rect 6690 24443 6998 24452
rect 2908 24236 2960 24242
rect 2908 24178 2960 24184
rect 2920 24145 2948 24178
rect 7140 24168 7192 24174
rect 2906 24136 2962 24145
rect 7140 24110 7192 24116
rect 2906 24071 2962 24080
rect 7152 24009 7180 24110
rect 7138 24000 7194 24009
rect 5954 23964 6262 23973
rect 5954 23962 5960 23964
rect 6016 23962 6040 23964
rect 6096 23962 6120 23964
rect 6176 23962 6200 23964
rect 6256 23962 6262 23964
rect 6016 23910 6018 23962
rect 6198 23910 6200 23962
rect 7138 23935 7194 23944
rect 5954 23908 5960 23910
rect 6016 23908 6040 23910
rect 6096 23908 6120 23910
rect 6176 23908 6200 23910
rect 6256 23908 6262 23910
rect 5954 23899 6262 23908
rect 6690 23420 6998 23429
rect 6690 23418 6696 23420
rect 6752 23418 6776 23420
rect 6832 23418 6856 23420
rect 6912 23418 6936 23420
rect 6992 23418 6998 23420
rect 6752 23366 6754 23418
rect 6934 23366 6936 23418
rect 6690 23364 6696 23366
rect 6752 23364 6776 23366
rect 6832 23364 6856 23366
rect 6912 23364 6936 23366
rect 6992 23364 6998 23366
rect 6690 23355 6998 23364
rect 2908 23148 2960 23154
rect 2908 23090 2960 23096
rect 2920 22785 2948 23090
rect 7140 23080 7192 23086
rect 7140 23022 7192 23028
rect 7152 22921 7180 23022
rect 7138 22912 7194 22921
rect 5954 22876 6262 22885
rect 5954 22874 5960 22876
rect 6016 22874 6040 22876
rect 6096 22874 6120 22876
rect 6176 22874 6200 22876
rect 6256 22874 6262 22876
rect 6016 22822 6018 22874
rect 6198 22822 6200 22874
rect 7138 22847 7194 22856
rect 5954 22820 5960 22822
rect 6016 22820 6040 22822
rect 6096 22820 6120 22822
rect 6176 22820 6200 22822
rect 6256 22820 6262 22822
rect 5954 22811 6262 22820
rect 2906 22776 2962 22785
rect 2906 22711 2962 22720
rect 4932 22570 4984 22576
rect 4932 22512 4984 22518
rect 9164 22536 9216 22542
rect 4944 22105 4972 22512
rect 9164 22478 9216 22484
rect 6690 22332 6998 22341
rect 6690 22330 6696 22332
rect 6752 22330 6776 22332
rect 6832 22330 6856 22332
rect 6912 22330 6936 22332
rect 6992 22330 6998 22332
rect 6752 22278 6754 22330
rect 6934 22278 6936 22330
rect 6690 22276 6696 22278
rect 6752 22276 6776 22278
rect 6832 22276 6856 22278
rect 6912 22276 6936 22278
rect 6992 22276 6998 22278
rect 6690 22267 6998 22276
rect 4930 22096 4986 22105
rect 4930 22031 4986 22040
rect 9176 21833 9204 22478
rect 9162 21824 9218 21833
rect 5954 21788 6262 21797
rect 5954 21786 5960 21788
rect 6016 21786 6040 21788
rect 6096 21786 6120 21788
rect 6176 21786 6200 21788
rect 6256 21786 6262 21788
rect 6016 21734 6018 21786
rect 6198 21734 6200 21786
rect 9162 21759 9218 21768
rect 5954 21732 5960 21734
rect 6016 21732 6040 21734
rect 6096 21732 6120 21734
rect 6176 21732 6200 21734
rect 6256 21732 6262 21734
rect 5954 21723 6262 21732
rect 6690 21244 6998 21253
rect 6690 21242 6696 21244
rect 6752 21242 6776 21244
rect 6832 21242 6856 21244
rect 6912 21242 6936 21244
rect 6992 21242 6998 21244
rect 6752 21190 6754 21242
rect 6934 21190 6936 21242
rect 6690 21188 6696 21190
rect 6752 21188 6776 21190
rect 6832 21188 6856 21190
rect 6912 21188 6936 21190
rect 6992 21188 6998 21190
rect 6690 21179 6998 21188
rect 9256 21108 9308 21114
rect 9256 21050 9308 21056
rect 5208 21006 5260 21012
rect 5208 20948 5260 20954
rect 5220 20745 5248 20948
rect 9268 20745 9296 21050
rect 5206 20736 5262 20745
rect 9254 20736 9310 20745
rect 5206 20671 5262 20680
rect 5954 20700 6262 20709
rect 5954 20698 5960 20700
rect 6016 20698 6040 20700
rect 6096 20698 6120 20700
rect 6176 20698 6200 20700
rect 6256 20698 6262 20700
rect 6016 20646 6018 20698
rect 6198 20646 6200 20698
rect 9254 20671 9310 20680
rect 5954 20644 5960 20646
rect 6016 20644 6040 20646
rect 6096 20644 6120 20646
rect 6176 20644 6200 20646
rect 6256 20644 6262 20646
rect 5954 20635 6262 20644
rect 6690 20156 6998 20165
rect 6690 20154 6696 20156
rect 6752 20154 6776 20156
rect 6832 20154 6856 20156
rect 6912 20154 6936 20156
rect 6992 20154 6998 20156
rect 6752 20102 6754 20154
rect 6934 20102 6936 20154
rect 6690 20100 6696 20102
rect 6752 20100 6776 20102
rect 6832 20100 6856 20102
rect 6912 20100 6936 20102
rect 6992 20100 6998 20102
rect 6690 20091 6998 20100
rect 4932 19918 4984 19924
rect 4932 19860 4984 19866
rect 4944 19385 4972 19860
rect 7140 19816 7192 19822
rect 7140 19758 7192 19764
rect 7152 19657 7180 19758
rect 7138 19648 7194 19657
rect 5954 19612 6262 19621
rect 5954 19610 5960 19612
rect 6016 19610 6040 19612
rect 6096 19610 6120 19612
rect 6176 19610 6200 19612
rect 6256 19610 6262 19612
rect 6016 19558 6018 19610
rect 6198 19558 6200 19610
rect 7138 19583 7194 19592
rect 5954 19556 5960 19558
rect 6016 19556 6040 19558
rect 6096 19556 6120 19558
rect 6176 19556 6200 19558
rect 6256 19556 6262 19558
rect 5954 19547 6262 19556
rect 4930 19376 4986 19385
rect 4930 19311 4986 19320
rect 6690 19068 6998 19077
rect 6690 19066 6696 19068
rect 6752 19066 6776 19068
rect 6832 19066 6856 19068
rect 6912 19066 6936 19068
rect 6992 19066 6998 19068
rect 6752 19014 6754 19066
rect 6934 19014 6936 19066
rect 6690 19012 6696 19014
rect 6752 19012 6776 19014
rect 6832 19012 6856 19014
rect 6912 19012 6936 19014
rect 6992 19012 6998 19014
rect 6690 19003 6998 19012
rect 2908 18796 2960 18802
rect 2908 18738 2960 18744
rect 2920 18705 2948 18738
rect 7140 18728 7192 18734
rect 2906 18696 2962 18705
rect 7140 18670 7192 18676
rect 2906 18631 2962 18640
rect 7152 18569 7180 18670
rect 7138 18560 7194 18569
rect 5954 18524 6262 18533
rect 5954 18522 5960 18524
rect 6016 18522 6040 18524
rect 6096 18522 6120 18524
rect 6176 18522 6200 18524
rect 6256 18522 6262 18524
rect 6016 18470 6018 18522
rect 6198 18470 6200 18522
rect 7138 18495 7194 18504
rect 5954 18468 5960 18470
rect 6016 18468 6040 18470
rect 6096 18468 6120 18470
rect 6176 18468 6200 18470
rect 6256 18468 6262 18470
rect 5954 18459 6262 18468
rect 6690 17980 6998 17989
rect 6690 17978 6696 17980
rect 6752 17978 6776 17980
rect 6832 17978 6856 17980
rect 6912 17978 6936 17980
rect 6992 17978 6998 17980
rect 6752 17926 6754 17978
rect 6934 17926 6936 17978
rect 6690 17924 6696 17926
rect 6752 17924 6776 17926
rect 6832 17924 6856 17926
rect 6912 17924 6936 17926
rect 6992 17924 6998 17926
rect 6690 17915 6998 17924
rect 2908 17708 2960 17714
rect 2908 17650 2960 17656
rect 2920 17345 2948 17650
rect 7232 17640 7284 17646
rect 7232 17582 7284 17588
rect 7244 17481 7272 17582
rect 7230 17472 7286 17481
rect 5954 17436 6262 17445
rect 5954 17434 5960 17436
rect 6016 17434 6040 17436
rect 6096 17434 6120 17436
rect 6176 17434 6200 17436
rect 6256 17434 6262 17436
rect 6016 17382 6018 17434
rect 6198 17382 6200 17434
rect 7230 17407 7286 17416
rect 5954 17380 5960 17382
rect 6016 17380 6040 17382
rect 6096 17380 6120 17382
rect 6176 17380 6200 17382
rect 6256 17380 6262 17382
rect 5954 17371 6262 17380
rect 2906 17336 2962 17345
rect 2906 17271 2962 17280
rect 5208 17130 5260 17136
rect 5208 17072 5260 17078
rect 5220 16665 5248 17072
rect 5392 17028 5444 17034
rect 5392 16970 5444 16976
rect 5404 16665 5432 16970
rect 6690 16892 6998 16901
rect 6690 16890 6696 16892
rect 6752 16890 6776 16892
rect 6832 16890 6856 16892
rect 6912 16890 6936 16892
rect 6992 16890 6998 16892
rect 6752 16838 6754 16890
rect 6934 16838 6936 16890
rect 6690 16836 6696 16838
rect 6752 16836 6776 16838
rect 6832 16836 6856 16838
rect 6912 16836 6936 16838
rect 6992 16836 6998 16838
rect 6690 16827 6998 16836
rect 5206 16656 5262 16665
rect 5206 16591 5262 16600
rect 5390 16656 5446 16665
rect 5390 16591 5446 16600
rect 5954 16348 6262 16357
rect 5954 16346 5960 16348
rect 6016 16346 6040 16348
rect 6096 16346 6120 16348
rect 6176 16346 6200 16348
rect 6256 16346 6262 16348
rect 6016 16294 6018 16346
rect 6198 16294 6200 16346
rect 5954 16292 5960 16294
rect 6016 16292 6040 16294
rect 6096 16292 6120 16294
rect 6176 16292 6200 16294
rect 6256 16292 6262 16294
rect 5954 16283 6262 16292
rect 6690 15804 6998 15813
rect 6690 15802 6696 15804
rect 6752 15802 6776 15804
rect 6832 15802 6856 15804
rect 6912 15802 6936 15804
rect 6992 15802 6998 15804
rect 6752 15750 6754 15802
rect 6934 15750 6936 15802
rect 6690 15748 6696 15750
rect 6752 15748 6776 15750
rect 6832 15748 6856 15750
rect 6912 15748 6936 15750
rect 6992 15748 6998 15750
rect 6690 15739 6998 15748
rect 5208 15566 5260 15572
rect 5208 15508 5260 15514
rect 5220 15305 5248 15508
rect 5668 15464 5720 15470
rect 5668 15406 5720 15412
rect 5206 15296 5262 15305
rect 5206 15231 5262 15240
rect 5680 15033 5708 15406
rect 5954 15260 6262 15269
rect 5954 15258 5960 15260
rect 6016 15258 6040 15260
rect 6096 15258 6120 15260
rect 6176 15258 6200 15260
rect 6256 15258 6262 15260
rect 6016 15206 6018 15258
rect 6198 15206 6200 15258
rect 5954 15204 5960 15206
rect 6016 15204 6040 15206
rect 6096 15204 6120 15206
rect 6176 15204 6200 15206
rect 6256 15204 6262 15206
rect 5954 15195 6262 15204
rect 5666 15024 5722 15033
rect 5666 14959 5722 14968
rect 6690 14716 6998 14725
rect 6690 14714 6696 14716
rect 6752 14714 6776 14716
rect 6832 14714 6856 14716
rect 6912 14714 6936 14716
rect 6992 14714 6998 14716
rect 6752 14662 6754 14714
rect 6934 14662 6936 14714
rect 6690 14660 6696 14662
rect 6752 14660 6776 14662
rect 6832 14660 6856 14662
rect 6912 14660 6936 14662
rect 6992 14660 6998 14662
rect 6690 14651 6998 14660
rect 5954 14172 6262 14181
rect 5954 14170 5960 14172
rect 6016 14170 6040 14172
rect 6096 14170 6120 14172
rect 6176 14170 6200 14172
rect 6256 14170 6262 14172
rect 6016 14118 6018 14170
rect 6198 14118 6200 14170
rect 5954 14116 5960 14118
rect 6016 14116 6040 14118
rect 6096 14116 6120 14118
rect 6176 14116 6200 14118
rect 6256 14116 6262 14118
rect 5954 14107 6262 14116
rect 6690 13628 6998 13637
rect 6690 13626 6696 13628
rect 6752 13626 6776 13628
rect 6832 13626 6856 13628
rect 6912 13626 6936 13628
rect 6992 13626 6998 13628
rect 6752 13574 6754 13626
rect 6934 13574 6936 13626
rect 6690 13572 6696 13574
rect 6752 13572 6776 13574
rect 6832 13572 6856 13574
rect 6912 13572 6936 13574
rect 6992 13572 6998 13574
rect 6690 13563 6998 13572
rect 45884 13097 45912 49435
rect 45976 14185 46004 50523
rect 46068 48421 46096 84562
rect 46054 48412 46110 48421
rect 46054 48347 46110 48356
rect 45962 14176 46018 14185
rect 45962 14111 46018 14120
rect 5954 13084 6262 13093
rect 5954 13082 5960 13084
rect 6016 13082 6040 13084
rect 6096 13082 6120 13084
rect 6176 13082 6200 13084
rect 6256 13082 6262 13084
rect 6016 13030 6018 13082
rect 6198 13030 6200 13082
rect 5954 13028 5960 13030
rect 6016 13028 6040 13030
rect 6096 13028 6120 13030
rect 6176 13028 6200 13030
rect 6256 13028 6262 13030
rect 5954 13019 6262 13028
rect 45870 13088 45926 13097
rect 45870 13023 45926 13032
rect 6690 12540 6998 12549
rect 6690 12538 6696 12540
rect 6752 12538 6776 12540
rect 6832 12538 6856 12540
rect 6912 12538 6936 12540
rect 6992 12538 6998 12540
rect 6752 12486 6754 12538
rect 6934 12486 6936 12538
rect 6690 12484 6696 12486
rect 6752 12484 6776 12486
rect 6832 12484 6856 12486
rect 6912 12484 6936 12486
rect 6992 12484 6998 12486
rect 6690 12475 6998 12484
rect 5954 11996 6262 12005
rect 5954 11994 5960 11996
rect 6016 11994 6040 11996
rect 6096 11994 6120 11996
rect 6176 11994 6200 11996
rect 6256 11994 6262 11996
rect 6016 11942 6018 11994
rect 6198 11942 6200 11994
rect 5954 11940 5960 11942
rect 6016 11940 6040 11942
rect 6096 11940 6120 11942
rect 6176 11940 6200 11942
rect 6256 11940 6262 11942
rect 5954 11931 6262 11940
rect 6690 11452 6998 11461
rect 6690 11450 6696 11452
rect 6752 11450 6776 11452
rect 6832 11450 6856 11452
rect 6912 11450 6936 11452
rect 6992 11450 6998 11452
rect 6752 11398 6754 11450
rect 6934 11398 6936 11450
rect 6690 11396 6696 11398
rect 6752 11396 6776 11398
rect 6832 11396 6856 11398
rect 6912 11396 6936 11398
rect 6992 11396 6998 11398
rect 6690 11387 6998 11396
rect 5954 10908 6262 10917
rect 5954 10906 5960 10908
rect 6016 10906 6040 10908
rect 6096 10906 6120 10908
rect 6176 10906 6200 10908
rect 6256 10906 6262 10908
rect 6016 10854 6018 10906
rect 6198 10854 6200 10906
rect 5954 10852 5960 10854
rect 6016 10852 6040 10854
rect 6096 10852 6120 10854
rect 6176 10852 6200 10854
rect 6256 10852 6262 10854
rect 5954 10843 6262 10852
rect 45870 10876 45926 10885
rect 45870 10811 45926 10820
rect 6690 10364 6998 10373
rect 6690 10362 6696 10364
rect 6752 10362 6776 10364
rect 6832 10362 6856 10364
rect 6912 10362 6936 10364
rect 6992 10362 6998 10364
rect 6752 10310 6754 10362
rect 6934 10310 6936 10362
rect 6690 10308 6696 10310
rect 6752 10308 6776 10310
rect 6832 10308 6856 10310
rect 6912 10308 6936 10310
rect 6992 10308 6998 10310
rect 6690 10299 6998 10308
rect 45596 10228 45648 10234
rect 45596 10170 45648 10176
rect 15032 10086 15276 10114
rect 5954 9820 6262 9829
rect 5954 9818 5960 9820
rect 6016 9818 6040 9820
rect 6096 9818 6120 9820
rect 6176 9818 6200 9820
rect 6256 9818 6262 9820
rect 6016 9766 6018 9818
rect 6198 9766 6200 9818
rect 5954 9764 5960 9766
rect 6016 9764 6040 9766
rect 6096 9764 6120 9766
rect 6176 9764 6200 9766
rect 6256 9764 6262 9766
rect 5954 9755 6262 9764
rect 6690 9276 6998 9285
rect 6690 9274 6696 9276
rect 6752 9274 6776 9276
rect 6832 9274 6856 9276
rect 6912 9274 6936 9276
rect 6992 9274 6998 9276
rect 6752 9222 6754 9274
rect 6934 9222 6936 9274
rect 6690 9220 6696 9222
rect 6752 9220 6776 9222
rect 6832 9220 6856 9222
rect 6912 9220 6936 9222
rect 6992 9220 6998 9222
rect 6690 9211 6998 9220
rect 5954 8732 6262 8741
rect 5954 8730 5960 8732
rect 6016 8730 6040 8732
rect 6096 8730 6120 8732
rect 6176 8730 6200 8732
rect 6256 8730 6262 8732
rect 6016 8678 6018 8730
rect 6198 8678 6200 8730
rect 5954 8676 5960 8678
rect 6016 8676 6040 8678
rect 6096 8676 6120 8678
rect 6176 8676 6200 8678
rect 6256 8676 6262 8678
rect 5954 8667 6262 8676
rect 6690 8188 6998 8197
rect 6690 8186 6696 8188
rect 6752 8186 6776 8188
rect 6832 8186 6856 8188
rect 6912 8186 6936 8188
rect 6992 8186 6998 8188
rect 6752 8134 6754 8186
rect 6934 8134 6936 8186
rect 6690 8132 6696 8134
rect 6752 8132 6776 8134
rect 6832 8132 6856 8134
rect 6912 8132 6936 8134
rect 6992 8132 6998 8134
rect 6690 8123 6998 8132
rect 5954 7644 6262 7653
rect 5954 7642 5960 7644
rect 6016 7642 6040 7644
rect 6096 7642 6120 7644
rect 6176 7642 6200 7644
rect 6256 7642 6262 7644
rect 6016 7590 6018 7642
rect 6198 7590 6200 7642
rect 5954 7588 5960 7590
rect 6016 7588 6040 7590
rect 6096 7588 6120 7590
rect 6176 7588 6200 7590
rect 6256 7588 6262 7590
rect 5954 7579 6262 7588
rect 6690 7100 6998 7109
rect 6690 7098 6696 7100
rect 6752 7098 6776 7100
rect 6832 7098 6856 7100
rect 6912 7098 6936 7100
rect 6992 7098 6998 7100
rect 6752 7046 6754 7098
rect 6934 7046 6936 7098
rect 6690 7044 6696 7046
rect 6752 7044 6776 7046
rect 6832 7044 6856 7046
rect 6912 7044 6936 7046
rect 6992 7044 6998 7046
rect 6690 7035 6998 7044
rect 15248 5168 15276 10086
rect 16076 5168 16104 10100
rect 17180 5168 17208 10100
rect 17722 7644 18030 7653
rect 17722 7642 17728 7644
rect 17784 7642 17808 7644
rect 17864 7642 17888 7644
rect 17944 7642 17968 7644
rect 18024 7642 18030 7644
rect 17784 7590 17786 7642
rect 17966 7590 17968 7642
rect 17722 7588 17728 7590
rect 17784 7588 17808 7590
rect 17864 7588 17888 7590
rect 17944 7588 17968 7590
rect 18024 7588 18030 7590
rect 17722 7579 18030 7588
rect 17722 6556 18030 6565
rect 17722 6554 17728 6556
rect 17784 6554 17808 6556
rect 17864 6554 17888 6556
rect 17944 6554 17968 6556
rect 18024 6554 18030 6556
rect 17784 6502 17786 6554
rect 17966 6502 17968 6554
rect 17722 6500 17728 6502
rect 17784 6500 17808 6502
rect 17864 6500 17888 6502
rect 17944 6500 17968 6502
rect 18024 6500 18030 6502
rect 17722 6491 18030 6500
rect 17722 5468 18030 5477
rect 17722 5466 17728 5468
rect 17784 5466 17808 5468
rect 17864 5466 17888 5468
rect 17944 5466 17968 5468
rect 18024 5466 18030 5468
rect 17784 5414 17786 5466
rect 17966 5414 17968 5466
rect 17722 5412 17728 5414
rect 17784 5412 17808 5414
rect 17864 5412 17888 5414
rect 17944 5412 17968 5414
rect 18024 5412 18030 5414
rect 17722 5403 18030 5412
rect 18284 5168 18312 10100
rect 19448 10086 19692 10114
rect 18382 7100 18690 7109
rect 18382 7098 18388 7100
rect 18444 7098 18468 7100
rect 18524 7098 18548 7100
rect 18604 7098 18628 7100
rect 18684 7098 18690 7100
rect 18444 7046 18446 7098
rect 18626 7046 18628 7098
rect 18382 7044 18388 7046
rect 18444 7044 18468 7046
rect 18524 7044 18548 7046
rect 18604 7044 18628 7046
rect 18684 7044 18690 7046
rect 18382 7035 18690 7044
rect 18382 6012 18690 6021
rect 18382 6010 18388 6012
rect 18444 6010 18468 6012
rect 18524 6010 18548 6012
rect 18604 6010 18628 6012
rect 18684 6010 18690 6012
rect 18444 5958 18446 6010
rect 18626 5958 18628 6010
rect 18382 5956 18388 5958
rect 18444 5956 18468 5958
rect 18524 5956 18548 5958
rect 18604 5956 18628 5958
rect 18684 5956 18690 5958
rect 18382 5947 18690 5956
rect 19664 5168 19692 10086
rect 20492 5168 20520 10100
rect 21596 5168 21624 10100
rect 22760 10086 23004 10114
rect 22976 5168 23004 10086
rect 23804 5168 23832 10100
rect 24908 5168 24936 10100
rect 26058 9842 26086 10100
rect 27176 10086 27420 10114
rect 26058 9814 26132 9842
rect 26104 5168 26132 9814
rect 27392 5168 27420 10086
rect 28220 5168 28248 10100
rect 29324 5168 29352 10100
rect 30488 10086 30732 10114
rect 30704 5338 30732 10086
rect 31532 5338 31560 10100
rect 32682 9842 32710 10100
rect 33786 9842 33814 10100
rect 34904 10086 35148 10114
rect 32682 9814 32756 9842
rect 33786 9814 33860 9842
rect 30692 5332 30744 5338
rect 30692 5274 30744 5280
rect 31520 5332 31572 5338
rect 31520 5274 31572 5280
rect 32728 5270 32756 9814
rect 33832 5338 33860 9814
rect 35120 5338 35148 10086
rect 35948 5338 35976 10100
rect 37098 9842 37126 10100
rect 38216 10086 38460 10114
rect 37098 9814 37172 9842
rect 36122 7644 36430 7653
rect 36122 7642 36128 7644
rect 36184 7642 36208 7644
rect 36264 7642 36288 7644
rect 36344 7642 36368 7644
rect 36424 7642 36430 7644
rect 36184 7590 36186 7642
rect 36366 7590 36368 7642
rect 36122 7588 36128 7590
rect 36184 7588 36208 7590
rect 36264 7588 36288 7590
rect 36344 7588 36368 7590
rect 36424 7588 36430 7590
rect 36122 7579 36430 7588
rect 36782 7100 37090 7109
rect 36782 7098 36788 7100
rect 36844 7098 36868 7100
rect 36924 7098 36948 7100
rect 37004 7098 37028 7100
rect 37084 7098 37090 7100
rect 36844 7046 36846 7098
rect 37026 7046 37028 7098
rect 36782 7044 36788 7046
rect 36844 7044 36868 7046
rect 36924 7044 36948 7046
rect 37004 7044 37028 7046
rect 37084 7044 37090 7046
rect 36782 7035 37090 7044
rect 36122 6556 36430 6565
rect 36122 6554 36128 6556
rect 36184 6554 36208 6556
rect 36264 6554 36288 6556
rect 36344 6554 36368 6556
rect 36424 6554 36430 6556
rect 36184 6502 36186 6554
rect 36366 6502 36368 6554
rect 36122 6500 36128 6502
rect 36184 6500 36208 6502
rect 36264 6500 36288 6502
rect 36344 6500 36368 6502
rect 36424 6500 36430 6502
rect 36122 6491 36430 6500
rect 36782 6012 37090 6021
rect 36782 6010 36788 6012
rect 36844 6010 36868 6012
rect 36924 6010 36948 6012
rect 37004 6010 37028 6012
rect 37084 6010 37090 6012
rect 36844 5958 36846 6010
rect 37026 5958 37028 6010
rect 36782 5956 36788 5958
rect 36844 5956 36868 5958
rect 36924 5956 36948 5958
rect 37004 5956 37028 5958
rect 37084 5956 37090 5958
rect 36782 5947 37090 5956
rect 36122 5468 36430 5477
rect 36122 5466 36128 5468
rect 36184 5466 36208 5468
rect 36264 5466 36288 5468
rect 36344 5466 36368 5468
rect 36424 5466 36430 5468
rect 36184 5414 36186 5466
rect 36366 5414 36368 5466
rect 36122 5412 36128 5414
rect 36184 5412 36208 5414
rect 36264 5412 36288 5414
rect 36344 5412 36368 5414
rect 36424 5412 36430 5414
rect 36122 5403 36430 5412
rect 37144 5338 37172 9814
rect 38432 5338 38460 10086
rect 39260 5338 39288 10100
rect 40410 9842 40438 10100
rect 41528 10086 41680 10114
rect 42632 10086 42876 10114
rect 40410 9814 40484 9842
rect 33820 5332 33872 5338
rect 33820 5274 33872 5280
rect 35108 5332 35160 5338
rect 35108 5274 35160 5280
rect 35936 5332 35988 5338
rect 35936 5274 35988 5280
rect 37132 5332 37184 5338
rect 37132 5274 37184 5280
rect 38420 5332 38472 5338
rect 38420 5274 38472 5280
rect 39248 5332 39300 5338
rect 39248 5274 39300 5280
rect 40456 5270 40484 9814
rect 41652 5338 41680 10086
rect 42848 5338 42876 10086
rect 43676 5338 43704 10100
rect 44780 5338 44808 10100
rect 45608 7446 45636 10170
rect 45884 8514 45912 10811
rect 45700 8486 45912 8514
rect 45700 7514 45728 8486
rect 45976 7514 46004 14111
rect 46068 12009 46096 48347
rect 46160 47333 46188 84562
rect 47160 84552 47212 84558
rect 47160 84494 47212 84500
rect 47172 83062 47200 84494
rect 49104 84490 49132 84970
rect 50196 84688 50248 84694
rect 50196 84630 50248 84636
rect 50208 84490 50236 84630
rect 51300 84620 51352 84626
rect 51300 84562 51352 84568
rect 49092 84484 49144 84490
rect 49092 84426 49144 84432
rect 50196 84484 50248 84490
rect 50196 84426 50248 84432
rect 47068 83056 47120 83062
rect 47068 82998 47120 83004
rect 47160 83056 47212 83062
rect 47160 82998 47212 83004
rect 47988 83056 48040 83062
rect 47988 82998 48040 83004
rect 46146 47324 46202 47333
rect 46146 47259 46202 47268
rect 46424 45928 46476 45934
rect 46424 45870 46476 45876
rect 46146 13088 46202 13097
rect 46146 13023 46202 13032
rect 46054 12000 46110 12009
rect 46054 11935 46110 11944
rect 46068 10234 46096 11935
rect 46056 10228 46108 10234
rect 46056 10170 46108 10176
rect 46160 8514 46188 13023
rect 46436 10953 46464 45870
rect 47080 45769 47108 82998
rect 48000 82466 48028 82998
rect 49104 82466 49132 84426
rect 50208 82466 50236 84426
rect 51312 82466 51340 84562
rect 52692 82466 52720 87146
rect 53520 82466 53548 87146
rect 47984 82438 48028 82466
rect 49088 82438 49132 82466
rect 50192 82438 50236 82466
rect 51296 82438 51340 82466
rect 52400 82438 52720 82466
rect 53504 82438 53548 82466
rect 54440 82466 54468 87146
rect 54522 87068 54830 87077
rect 54522 87066 54528 87068
rect 54584 87066 54608 87068
rect 54664 87066 54688 87068
rect 54744 87066 54768 87068
rect 54824 87066 54830 87068
rect 54584 87014 54586 87066
rect 54766 87014 54768 87066
rect 54522 87012 54528 87014
rect 54584 87012 54608 87014
rect 54664 87012 54688 87014
rect 54744 87012 54768 87014
rect 54824 87012 54830 87014
rect 54522 87003 54830 87012
rect 55182 86524 55490 86533
rect 55182 86522 55188 86524
rect 55244 86522 55268 86524
rect 55324 86522 55348 86524
rect 55404 86522 55428 86524
rect 55484 86522 55490 86524
rect 55244 86470 55246 86522
rect 55426 86470 55428 86522
rect 55182 86468 55188 86470
rect 55244 86468 55268 86470
rect 55324 86468 55348 86470
rect 55404 86468 55428 86470
rect 55484 86468 55490 86470
rect 55182 86459 55490 86468
rect 54522 85980 54830 85989
rect 54522 85978 54528 85980
rect 54584 85978 54608 85980
rect 54664 85978 54688 85980
rect 54744 85978 54768 85980
rect 54824 85978 54830 85980
rect 54584 85926 54586 85978
rect 54766 85926 54768 85978
rect 54522 85924 54528 85926
rect 54584 85924 54608 85926
rect 54664 85924 54688 85926
rect 54744 85924 54768 85926
rect 54824 85924 54830 85926
rect 54522 85915 54830 85924
rect 55182 85436 55490 85445
rect 55182 85434 55188 85436
rect 55244 85434 55268 85436
rect 55324 85434 55348 85436
rect 55404 85434 55428 85436
rect 55484 85434 55490 85436
rect 55244 85382 55246 85434
rect 55426 85382 55428 85434
rect 55182 85380 55188 85382
rect 55244 85380 55268 85382
rect 55324 85380 55348 85382
rect 55404 85380 55428 85382
rect 55484 85380 55490 85382
rect 55182 85371 55490 85380
rect 54522 84892 54830 84901
rect 54522 84890 54528 84892
rect 54584 84890 54608 84892
rect 54664 84890 54688 84892
rect 54744 84890 54768 84892
rect 54824 84890 54830 84892
rect 54584 84838 54586 84890
rect 54766 84838 54768 84890
rect 54522 84836 54528 84838
rect 54584 84836 54608 84838
rect 54664 84836 54688 84838
rect 54744 84836 54768 84838
rect 54824 84836 54830 84838
rect 54522 84827 54830 84836
rect 55182 84348 55490 84357
rect 55182 84346 55188 84348
rect 55244 84346 55268 84348
rect 55324 84346 55348 84348
rect 55404 84346 55428 84348
rect 55484 84346 55490 84348
rect 55244 84294 55246 84346
rect 55426 84294 55428 84346
rect 55182 84292 55188 84294
rect 55244 84292 55268 84294
rect 55324 84292 55348 84294
rect 55404 84292 55428 84294
rect 55484 84292 55490 84294
rect 55182 84283 55490 84292
rect 55728 82466 55756 87146
rect 56832 82466 56860 87214
rect 57924 87204 57976 87210
rect 57924 87146 57976 87152
rect 59028 87204 59080 87210
rect 59028 87146 59080 87152
rect 57936 82466 57964 87146
rect 59040 82466 59068 87146
rect 60144 82466 60172 87282
rect 62340 87272 62392 87278
rect 62340 87214 62392 87220
rect 64548 87272 64600 87278
rect 64548 87214 64600 87220
rect 61236 87204 61288 87210
rect 61236 87146 61288 87152
rect 61248 82466 61276 87146
rect 62352 82466 62380 87214
rect 63444 87204 63496 87210
rect 63444 87146 63496 87152
rect 63456 82466 63484 87146
rect 64560 82466 64588 87214
rect 65652 87204 65704 87210
rect 65652 87146 65704 87152
rect 66756 87204 66808 87210
rect 66756 87146 66808 87152
rect 65664 82466 65692 87146
rect 66768 82466 66796 87146
rect 67872 82466 67900 87316
rect 54440 82438 54636 82466
rect 47984 82180 48012 82438
rect 49088 82180 49116 82438
rect 50192 82180 50220 82438
rect 51296 82180 51324 82438
rect 52400 82180 52428 82438
rect 53504 82180 53532 82438
rect 54608 82180 54636 82438
rect 55712 82438 55756 82466
rect 56816 82438 56860 82466
rect 57920 82438 57964 82466
rect 59024 82438 59068 82466
rect 60128 82438 60172 82466
rect 61232 82438 61276 82466
rect 62336 82438 62380 82466
rect 63440 82438 63484 82466
rect 64544 82438 64588 82466
rect 65648 82438 65692 82466
rect 66752 82438 66796 82466
rect 67856 82438 67900 82466
rect 69344 82450 69372 87316
rect 70080 82466 70108 87316
rect 71184 82466 71212 87316
rect 72288 82466 72316 87316
rect 72922 87068 73230 87077
rect 72922 87066 72928 87068
rect 72984 87066 73008 87068
rect 73064 87066 73088 87068
rect 73144 87066 73168 87068
rect 73224 87066 73230 87068
rect 72984 87014 72986 87066
rect 73166 87014 73168 87066
rect 72922 87012 72928 87014
rect 72984 87012 73008 87014
rect 73064 87012 73088 87014
rect 73144 87012 73168 87014
rect 73224 87012 73230 87014
rect 72922 87003 73230 87012
rect 72922 85980 73230 85989
rect 72922 85978 72928 85980
rect 72984 85978 73008 85980
rect 73064 85978 73088 85980
rect 73144 85978 73168 85980
rect 73224 85978 73230 85980
rect 72984 85926 72986 85978
rect 73166 85926 73168 85978
rect 72922 85924 72928 85926
rect 72984 85924 73008 85926
rect 73064 85924 73088 85926
rect 73144 85924 73168 85926
rect 73224 85924 73230 85926
rect 72922 85915 73230 85924
rect 72922 84892 73230 84901
rect 72922 84890 72928 84892
rect 72984 84890 73008 84892
rect 73064 84890 73088 84892
rect 73144 84890 73168 84892
rect 73224 84890 73230 84892
rect 72984 84838 72986 84890
rect 73166 84838 73168 84890
rect 72922 84836 72928 84838
rect 72984 84836 73008 84838
rect 73064 84836 73088 84838
rect 73144 84836 73168 84838
rect 73224 84836 73230 84838
rect 72922 84827 73230 84836
rect 73392 82466 73420 87316
rect 73582 86524 73890 86533
rect 73582 86522 73588 86524
rect 73644 86522 73668 86524
rect 73724 86522 73748 86524
rect 73804 86522 73828 86524
rect 73884 86522 73890 86524
rect 73644 86470 73646 86522
rect 73826 86470 73828 86522
rect 73582 86468 73588 86470
rect 73644 86468 73668 86470
rect 73724 86468 73748 86470
rect 73804 86468 73828 86470
rect 73884 86468 73890 86470
rect 73582 86459 73890 86468
rect 73582 85436 73890 85445
rect 73582 85434 73588 85436
rect 73644 85434 73668 85436
rect 73724 85434 73748 85436
rect 73804 85434 73828 85436
rect 73884 85434 73890 85436
rect 73644 85382 73646 85434
rect 73826 85382 73828 85434
rect 73582 85380 73588 85382
rect 73644 85380 73668 85382
rect 73724 85380 73748 85382
rect 73804 85380 73828 85382
rect 73884 85380 73890 85382
rect 73582 85371 73890 85380
rect 73582 84348 73890 84357
rect 73582 84346 73588 84348
rect 73644 84346 73668 84348
rect 73724 84346 73748 84348
rect 73804 84346 73828 84348
rect 73884 84346 73890 84348
rect 73644 84294 73646 84346
rect 73826 84294 73828 84346
rect 73582 84292 73588 84294
rect 73644 84292 73668 84294
rect 73724 84292 73748 84294
rect 73804 84292 73828 84294
rect 73884 84292 73890 84294
rect 73582 84283 73890 84292
rect 74496 82466 74524 87316
rect 75600 82466 75628 87316
rect 77796 87316 77848 87322
rect 78900 87374 78952 87380
rect 78900 87316 78952 87322
rect 80280 87374 80332 87380
rect 80280 87316 80332 87322
rect 81108 87374 81160 87380
rect 81108 87316 81160 87322
rect 82212 87374 82264 87380
rect 82212 87316 82264 87322
rect 76692 87282 76744 87288
rect 76704 82466 76732 87282
rect 77808 82466 77836 87316
rect 78912 82466 78940 87316
rect 80292 82466 80320 87316
rect 81120 82466 81148 87316
rect 82224 82466 82252 87316
rect 86546 84892 86854 84901
rect 86546 84890 86552 84892
rect 86608 84890 86632 84892
rect 86688 84890 86712 84892
rect 86768 84890 86792 84892
rect 86848 84890 86854 84892
rect 86608 84838 86610 84890
rect 86790 84838 86792 84890
rect 86546 84836 86552 84838
rect 86608 84836 86632 84838
rect 86688 84836 86712 84838
rect 86768 84836 86792 84838
rect 86848 84836 86854 84838
rect 86546 84827 86854 84836
rect 87282 84348 87590 84357
rect 87282 84346 87288 84348
rect 87344 84346 87368 84348
rect 87424 84346 87448 84348
rect 87504 84346 87528 84348
rect 87584 84346 87590 84348
rect 87344 84294 87346 84346
rect 87526 84294 87528 84346
rect 87282 84292 87288 84294
rect 87344 84292 87368 84294
rect 87424 84292 87448 84294
rect 87504 84292 87528 84294
rect 87584 84292 87590 84294
rect 87282 84283 87590 84292
rect 86546 83804 86854 83813
rect 86546 83802 86552 83804
rect 86608 83802 86632 83804
rect 86688 83802 86712 83804
rect 86768 83802 86792 83804
rect 86848 83802 86854 83804
rect 86608 83750 86610 83802
rect 86790 83750 86792 83802
rect 86546 83748 86552 83750
rect 86608 83748 86632 83750
rect 86688 83748 86712 83750
rect 86768 83748 86792 83750
rect 86848 83748 86854 83750
rect 86546 83739 86854 83748
rect 87282 83260 87590 83269
rect 87282 83258 87288 83260
rect 87344 83258 87368 83260
rect 87424 83258 87448 83260
rect 87504 83258 87528 83260
rect 87584 83258 87590 83260
rect 87344 83206 87346 83258
rect 87526 83206 87528 83258
rect 87282 83204 87288 83206
rect 87344 83204 87368 83206
rect 87424 83204 87448 83206
rect 87504 83204 87528 83206
rect 87584 83204 87590 83206
rect 87282 83195 87590 83204
rect 83316 83124 83368 83130
rect 83316 83066 83368 83072
rect 68948 82444 69000 82450
rect 55712 82180 55740 82438
rect 56816 82180 56844 82438
rect 57920 82180 57948 82438
rect 59024 82180 59052 82438
rect 60128 82180 60156 82438
rect 61232 82180 61260 82438
rect 62336 82180 62364 82438
rect 63440 82180 63468 82438
rect 64544 82180 64572 82438
rect 65648 82180 65676 82438
rect 66752 82180 66780 82438
rect 67856 82180 67884 82438
rect 68948 82386 69000 82392
rect 69332 82444 69384 82450
rect 69332 82386 69384 82392
rect 70064 82438 70108 82466
rect 71168 82438 71212 82466
rect 72272 82438 72316 82466
rect 73376 82438 73420 82466
rect 74480 82438 74524 82466
rect 75584 82438 75628 82466
rect 76688 82438 76732 82466
rect 77792 82438 77836 82466
rect 78896 82438 78940 82466
rect 80000 82438 80320 82466
rect 81104 82438 81148 82466
rect 82208 82438 82252 82466
rect 68960 82180 68988 82386
rect 70064 82180 70092 82438
rect 71168 82180 71196 82438
rect 72272 82180 72300 82438
rect 73376 82180 73404 82438
rect 74480 82180 74508 82438
rect 75584 82180 75612 82438
rect 76688 82180 76716 82438
rect 77792 82180 77820 82438
rect 78896 82180 78924 82438
rect 80000 82180 80028 82438
rect 81104 82180 81132 82438
rect 82208 82180 82236 82438
rect 51284 45928 51336 45934
rect 52416 45882 52444 46548
rect 53520 45882 53548 46548
rect 54624 45882 54652 46548
rect 55728 45882 55756 46548
rect 56832 45882 56860 46548
rect 57936 45882 57964 46548
rect 59040 45882 59068 46548
rect 60144 45882 60172 46548
rect 61248 45882 61276 46548
rect 62352 45882 62380 46548
rect 63456 45882 63484 46548
rect 64560 45882 64588 46548
rect 65664 45882 65692 46548
rect 66768 45882 66796 46548
rect 67872 45882 67900 46548
rect 68976 45882 69004 46548
rect 70080 45882 70108 46548
rect 71184 45882 71212 46548
rect 72288 45882 72316 46548
rect 73392 45882 73420 46548
rect 74496 45882 74524 46548
rect 75600 45882 75628 46548
rect 76704 45882 76732 46548
rect 77808 45882 77836 46548
rect 78912 45882 78940 46548
rect 80016 45882 80044 46548
rect 81120 45882 81148 46548
rect 82224 45882 82252 46548
rect 51284 45870 51336 45876
rect 47066 45760 47122 45769
rect 47066 45695 47122 45704
rect 47342 45760 47398 45769
rect 51296 45732 51324 45870
rect 52400 45854 52444 45882
rect 53504 45854 53548 45882
rect 54608 45854 54652 45882
rect 55712 45854 55756 45882
rect 56816 45854 56860 45882
rect 57920 45854 57964 45882
rect 59024 45854 59068 45882
rect 60128 45854 60172 45882
rect 61232 45854 61276 45882
rect 62336 45854 62380 45882
rect 63440 45854 63484 45882
rect 64544 45854 64588 45882
rect 65648 45854 65692 45882
rect 66752 45854 66796 45882
rect 67856 45854 67900 45882
rect 68960 45854 69004 45882
rect 70064 45854 70108 45882
rect 71168 45854 71212 45882
rect 72272 45854 72316 45882
rect 73376 45854 73420 45882
rect 74480 45854 74524 45882
rect 75584 45854 75628 45882
rect 76688 45854 76732 45882
rect 77792 45854 77836 45882
rect 78896 45854 78940 45882
rect 80000 45854 80044 45882
rect 81104 45854 81148 45882
rect 82208 45854 82252 45882
rect 52400 45732 52428 45854
rect 53504 45732 53532 45854
rect 54608 45732 54636 45854
rect 55712 45732 55740 45854
rect 56816 45732 56844 45854
rect 57920 45732 57948 45854
rect 59024 45732 59052 45854
rect 60128 45732 60156 45854
rect 61232 45732 61260 45854
rect 62336 45732 62364 45854
rect 63440 45732 63468 45854
rect 64544 45732 64572 45854
rect 65648 45732 65676 45854
rect 66752 45732 66780 45854
rect 67856 45732 67884 45854
rect 68960 45732 68988 45854
rect 70064 45732 70092 45854
rect 71168 45732 71196 45854
rect 72272 45732 72300 45854
rect 73376 45732 73404 45854
rect 74480 45732 74508 45854
rect 75584 45732 75612 45854
rect 76688 45732 76716 45854
rect 77792 45732 77820 45854
rect 78896 45732 78924 45854
rect 80000 45732 80028 45854
rect 81104 45732 81132 45854
rect 82208 45732 82236 45854
rect 47342 45695 47398 45704
rect 47356 45225 47384 45695
rect 50178 45488 50234 45497
rect 50178 45423 50234 45432
rect 49074 45352 49130 45361
rect 49074 45287 49130 45296
rect 47342 45216 47398 45225
rect 47342 45151 47398 45160
rect 47970 45216 48026 45225
rect 47970 45151 48026 45160
rect 83328 11254 83356 83066
rect 86546 82716 86854 82725
rect 86546 82714 86552 82716
rect 86608 82714 86632 82716
rect 86688 82714 86712 82716
rect 86768 82714 86792 82716
rect 86848 82714 86854 82716
rect 86608 82662 86610 82714
rect 86790 82662 86792 82714
rect 86546 82660 86552 82662
rect 86608 82660 86632 82662
rect 86688 82660 86712 82662
rect 86768 82660 86792 82662
rect 86848 82660 86854 82662
rect 86546 82651 86854 82660
rect 87282 82172 87590 82181
rect 87282 82170 87288 82172
rect 87344 82170 87368 82172
rect 87424 82170 87448 82172
rect 87504 82170 87528 82172
rect 87584 82170 87590 82172
rect 87344 82118 87346 82170
rect 87526 82118 87528 82170
rect 87282 82116 87288 82118
rect 87344 82116 87368 82118
rect 87424 82116 87448 82118
rect 87504 82116 87528 82118
rect 87584 82116 87590 82118
rect 87282 82107 87590 82116
rect 86546 81628 86854 81637
rect 86546 81626 86552 81628
rect 86608 81626 86632 81628
rect 86688 81626 86712 81628
rect 86768 81626 86792 81628
rect 86848 81626 86854 81628
rect 86608 81574 86610 81626
rect 86790 81574 86792 81626
rect 86546 81572 86552 81574
rect 86608 81572 86632 81574
rect 86688 81572 86712 81574
rect 86768 81572 86792 81574
rect 86848 81572 86854 81574
rect 86546 81563 86854 81572
rect 83500 81424 83552 81430
rect 83500 81366 83552 81372
rect 83512 81061 83540 81366
rect 88376 81296 88428 81302
rect 88374 81256 88376 81265
rect 88428 81256 88430 81265
rect 88374 81191 88430 81200
rect 87282 81084 87590 81093
rect 87282 81082 87288 81084
rect 87344 81082 87368 81084
rect 87424 81082 87448 81084
rect 87504 81082 87528 81084
rect 87584 81082 87590 81084
rect 83498 81052 83554 81061
rect 87344 81030 87346 81082
rect 87526 81030 87528 81082
rect 87282 81028 87288 81030
rect 87344 81028 87368 81030
rect 87424 81028 87448 81030
rect 87504 81028 87528 81030
rect 87584 81028 87590 81030
rect 87282 81019 87590 81028
rect 83498 80987 83554 80996
rect 86546 80540 86854 80549
rect 86546 80538 86552 80540
rect 86608 80538 86632 80540
rect 86688 80538 86712 80540
rect 86768 80538 86792 80540
rect 86848 80538 86854 80540
rect 86608 80486 86610 80538
rect 86790 80486 86792 80538
rect 86546 80484 86552 80486
rect 86608 80484 86632 80486
rect 86688 80484 86712 80486
rect 86768 80484 86792 80486
rect 86848 80484 86854 80486
rect 86546 80475 86854 80484
rect 88284 80234 88336 80240
rect 83500 80200 83552 80206
rect 88284 80176 88336 80182
rect 83500 80142 83552 80148
rect 83512 79973 83540 80142
rect 87282 79996 87590 80005
rect 87282 79994 87288 79996
rect 87344 79994 87368 79996
rect 87424 79994 87448 79996
rect 87504 79994 87528 79996
rect 87584 79994 87590 79996
rect 83498 79964 83554 79973
rect 87344 79942 87346 79994
rect 87526 79942 87528 79994
rect 87282 79940 87288 79942
rect 87344 79940 87368 79942
rect 87424 79940 87448 79942
rect 87504 79940 87528 79942
rect 87584 79940 87590 79942
rect 87282 79931 87590 79940
rect 83498 79899 83554 79908
rect 88296 79905 88324 80176
rect 88282 79896 88338 79905
rect 88282 79831 88338 79840
rect 86546 79452 86854 79461
rect 86546 79450 86552 79452
rect 86608 79450 86632 79452
rect 86688 79450 86712 79452
rect 86768 79450 86792 79452
rect 86848 79450 86854 79452
rect 86608 79398 86610 79450
rect 86790 79398 86792 79450
rect 86546 79396 86552 79398
rect 86608 79396 86632 79398
rect 86688 79396 86712 79398
rect 86768 79396 86792 79398
rect 86848 79396 86854 79398
rect 86546 79387 86854 79396
rect 87282 78908 87590 78917
rect 87282 78906 87288 78908
rect 87344 78906 87368 78908
rect 87424 78906 87448 78908
rect 87504 78906 87528 78908
rect 87584 78906 87590 78908
rect 87344 78854 87346 78906
rect 87526 78854 87528 78906
rect 87282 78852 87288 78854
rect 87344 78852 87368 78854
rect 87424 78852 87448 78854
rect 87504 78852 87528 78854
rect 87584 78852 87590 78854
rect 87282 78843 87590 78852
rect 88006 78672 88062 78681
rect 88006 78607 88062 78616
rect 88284 78670 88336 78676
rect 88284 78612 88336 78618
rect 88020 78574 88048 78607
rect 88008 78568 88060 78574
rect 88296 78545 88324 78612
rect 88008 78510 88060 78516
rect 88282 78536 88338 78545
rect 88282 78471 88338 78480
rect 86546 78364 86854 78373
rect 86546 78362 86552 78364
rect 86608 78362 86632 78364
rect 86688 78362 86712 78364
rect 86768 78362 86792 78364
rect 86848 78362 86854 78364
rect 86608 78310 86610 78362
rect 86790 78310 86792 78362
rect 86546 78308 86552 78310
rect 86608 78308 86632 78310
rect 86688 78308 86712 78310
rect 86768 78308 86792 78310
rect 86848 78308 86854 78310
rect 86546 78299 86854 78308
rect 88284 78058 88336 78064
rect 87822 77992 87878 78001
rect 88284 78000 88336 78006
rect 87822 77927 87824 77936
rect 87876 77927 87878 77936
rect 87824 77898 87876 77904
rect 88296 77865 88324 78000
rect 88282 77856 88338 77865
rect 87282 77820 87590 77829
rect 87282 77818 87288 77820
rect 87344 77818 87368 77820
rect 87424 77818 87448 77820
rect 87504 77818 87528 77820
rect 87584 77818 87590 77820
rect 87344 77766 87346 77818
rect 87526 77766 87528 77818
rect 88282 77791 88338 77800
rect 87282 77764 87288 77766
rect 87344 77764 87368 77766
rect 87424 77764 87448 77766
rect 87504 77764 87528 77766
rect 87584 77764 87590 77766
rect 87282 77755 87590 77764
rect 86546 77276 86854 77285
rect 86546 77274 86552 77276
rect 86608 77274 86632 77276
rect 86688 77274 86712 77276
rect 86768 77274 86792 77276
rect 86848 77274 86854 77276
rect 86608 77222 86610 77274
rect 86790 77222 86792 77274
rect 86546 77220 86552 77222
rect 86608 77220 86632 77222
rect 86688 77220 86712 77222
rect 86768 77220 86792 77222
rect 86848 77220 86854 77222
rect 86546 77211 86854 77220
rect 86628 76868 86680 76874
rect 86628 76810 86680 76816
rect 88008 76868 88060 76874
rect 88008 76810 88060 76816
rect 86640 76777 86668 76810
rect 86626 76768 86682 76777
rect 86626 76703 86682 76712
rect 87282 76732 87590 76741
rect 87282 76730 87288 76732
rect 87344 76730 87368 76732
rect 87424 76730 87448 76732
rect 87504 76730 87528 76732
rect 87584 76730 87590 76732
rect 87344 76678 87346 76730
rect 87526 76678 87528 76730
rect 87282 76676 87288 76678
rect 87344 76676 87368 76678
rect 87424 76676 87448 76678
rect 87504 76676 87528 76678
rect 87584 76676 87590 76678
rect 87282 76667 87590 76676
rect 88020 76505 88048 76810
rect 88006 76496 88062 76505
rect 88006 76431 88062 76440
rect 86546 76188 86854 76197
rect 86546 76186 86552 76188
rect 86608 76186 86632 76188
rect 86688 76186 86712 76188
rect 86768 76186 86792 76188
rect 86848 76186 86854 76188
rect 86608 76134 86610 76186
rect 86790 76134 86792 76186
rect 86546 76132 86552 76134
rect 86608 76132 86632 76134
rect 86688 76132 86712 76134
rect 86768 76132 86792 76134
rect 86848 76132 86854 76134
rect 86546 76123 86854 76132
rect 86904 75984 86956 75990
rect 86904 75926 86956 75932
rect 86916 75689 86944 75926
rect 88468 75848 88520 75854
rect 88466 75816 88468 75825
rect 88520 75816 88522 75825
rect 88466 75751 88522 75760
rect 86902 75680 86958 75689
rect 86902 75615 86958 75624
rect 87282 75644 87590 75653
rect 87282 75642 87288 75644
rect 87344 75642 87368 75644
rect 87424 75642 87448 75644
rect 87504 75642 87528 75644
rect 87584 75642 87590 75644
rect 87344 75590 87346 75642
rect 87526 75590 87528 75642
rect 87282 75588 87288 75590
rect 87344 75588 87368 75590
rect 87424 75588 87448 75590
rect 87504 75588 87528 75590
rect 87584 75588 87590 75590
rect 87282 75579 87590 75588
rect 86546 75100 86854 75109
rect 86546 75098 86552 75100
rect 86608 75098 86632 75100
rect 86688 75098 86712 75100
rect 86768 75098 86792 75100
rect 86848 75098 86854 75100
rect 86608 75046 86610 75098
rect 86790 75046 86792 75098
rect 86546 75044 86552 75046
rect 86608 75044 86632 75046
rect 86688 75044 86712 75046
rect 86768 75044 86792 75046
rect 86848 75044 86854 75046
rect 86546 75035 86854 75044
rect 84420 74896 84472 74902
rect 84420 74838 84472 74844
rect 84432 74601 84460 74838
rect 88560 74828 88612 74834
rect 88560 74770 88612 74776
rect 84418 74592 84474 74601
rect 84418 74527 84474 74536
rect 87282 74556 87590 74565
rect 87282 74554 87288 74556
rect 87344 74554 87368 74556
rect 87424 74554 87448 74556
rect 87504 74554 87528 74556
rect 87584 74554 87590 74556
rect 87344 74502 87346 74554
rect 87526 74502 87528 74554
rect 87282 74500 87288 74502
rect 87344 74500 87368 74502
rect 87424 74500 87448 74502
rect 87504 74500 87528 74502
rect 87584 74500 87590 74502
rect 87282 74491 87590 74500
rect 88572 74465 88600 74770
rect 88558 74456 88614 74465
rect 88558 74391 88614 74400
rect 86546 74012 86854 74021
rect 86546 74010 86552 74012
rect 86608 74010 86632 74012
rect 86688 74010 86712 74012
rect 86768 74010 86792 74012
rect 86848 74010 86854 74012
rect 86608 73958 86610 74010
rect 86790 73958 86792 74010
rect 86546 73956 86552 73958
rect 86608 73956 86632 73958
rect 86688 73956 86712 73958
rect 86768 73956 86792 73958
rect 86848 73956 86854 73958
rect 86546 73947 86854 73956
rect 87282 73468 87590 73477
rect 87282 73466 87288 73468
rect 87344 73466 87368 73468
rect 87424 73466 87448 73468
rect 87504 73466 87528 73468
rect 87584 73466 87590 73468
rect 87344 73414 87346 73466
rect 87526 73414 87528 73466
rect 87282 73412 87288 73414
rect 87344 73412 87368 73414
rect 87424 73412 87448 73414
rect 87504 73412 87528 73414
rect 87584 73412 87590 73414
rect 87282 73403 87590 73412
rect 88006 73232 88062 73241
rect 88006 73167 88008 73176
rect 88060 73167 88062 73176
rect 88284 73230 88336 73236
rect 88284 73172 88336 73178
rect 88008 73138 88060 73144
rect 88296 73105 88324 73172
rect 88282 73096 88338 73105
rect 88282 73031 88338 73040
rect 86546 72924 86854 72933
rect 86546 72922 86552 72924
rect 86608 72922 86632 72924
rect 86688 72922 86712 72924
rect 86768 72922 86792 72924
rect 86848 72922 86854 72924
rect 86608 72870 86610 72922
rect 86790 72870 86792 72922
rect 86546 72868 86552 72870
rect 86608 72868 86632 72870
rect 86688 72868 86712 72870
rect 86768 72868 86792 72870
rect 86848 72868 86854 72870
rect 86546 72859 86854 72868
rect 88284 72612 88336 72618
rect 87180 72584 87232 72590
rect 87178 72552 87180 72561
rect 87232 72552 87234 72561
rect 88284 72554 88336 72560
rect 87178 72487 87234 72496
rect 88296 72425 88324 72554
rect 88282 72416 88338 72425
rect 87282 72380 87590 72389
rect 87282 72378 87288 72380
rect 87344 72378 87368 72380
rect 87424 72378 87448 72380
rect 87504 72378 87528 72380
rect 87584 72378 87590 72380
rect 87344 72326 87346 72378
rect 87526 72326 87528 72378
rect 88282 72351 88338 72360
rect 87282 72324 87288 72326
rect 87344 72324 87368 72326
rect 87424 72324 87448 72326
rect 87504 72324 87528 72326
rect 87584 72324 87590 72326
rect 87282 72315 87590 72324
rect 86546 71836 86854 71845
rect 86546 71834 86552 71836
rect 86608 71834 86632 71836
rect 86688 71834 86712 71836
rect 86768 71834 86792 71836
rect 86848 71834 86854 71836
rect 86608 71782 86610 71834
rect 86790 71782 86792 71834
rect 86546 71780 86552 71782
rect 86608 71780 86632 71782
rect 86688 71780 86712 71782
rect 86768 71780 86792 71782
rect 86848 71780 86854 71782
rect 86546 71771 86854 71780
rect 86904 71632 86956 71638
rect 86904 71574 86956 71580
rect 86916 71337 86944 71574
rect 88284 71530 88336 71536
rect 88284 71472 88336 71478
rect 86902 71328 86958 71337
rect 86902 71263 86958 71272
rect 87282 71292 87590 71301
rect 87282 71290 87288 71292
rect 87344 71290 87368 71292
rect 87424 71290 87448 71292
rect 87504 71290 87528 71292
rect 87584 71290 87590 71292
rect 87344 71238 87346 71290
rect 87526 71238 87528 71290
rect 87282 71236 87288 71238
rect 87344 71236 87368 71238
rect 87424 71236 87448 71238
rect 87504 71236 87528 71238
rect 87584 71236 87590 71238
rect 87282 71227 87590 71236
rect 88296 71065 88324 71472
rect 88282 71056 88338 71065
rect 88282 70991 88338 71000
rect 86546 70748 86854 70757
rect 86546 70746 86552 70748
rect 86608 70746 86632 70748
rect 86688 70746 86712 70748
rect 86768 70746 86792 70748
rect 86848 70746 86854 70748
rect 86608 70694 86610 70746
rect 86790 70694 86792 70746
rect 86546 70692 86552 70694
rect 86608 70692 86632 70694
rect 86688 70692 86712 70694
rect 86768 70692 86792 70694
rect 86848 70692 86854 70694
rect 86546 70683 86854 70692
rect 86904 70544 86956 70550
rect 86904 70486 86956 70492
rect 86916 70249 86944 70486
rect 88192 70476 88244 70482
rect 88192 70418 88244 70424
rect 88204 70385 88232 70418
rect 88190 70376 88246 70385
rect 88190 70311 88246 70320
rect 86902 70240 86958 70249
rect 86902 70175 86958 70184
rect 87282 70204 87590 70213
rect 87282 70202 87288 70204
rect 87344 70202 87368 70204
rect 87424 70202 87448 70204
rect 87504 70202 87528 70204
rect 87584 70202 87590 70204
rect 87344 70150 87346 70202
rect 87526 70150 87528 70202
rect 87282 70148 87288 70150
rect 87344 70148 87368 70150
rect 87424 70148 87448 70150
rect 87504 70148 87528 70150
rect 87584 70148 87590 70150
rect 87282 70139 87590 70148
rect 86546 69660 86854 69669
rect 86546 69658 86552 69660
rect 86608 69658 86632 69660
rect 86688 69658 86712 69660
rect 86768 69658 86792 69660
rect 86848 69658 86854 69660
rect 86608 69606 86610 69658
rect 86790 69606 86792 69658
rect 86546 69604 86552 69606
rect 86608 69604 86632 69606
rect 86688 69604 86712 69606
rect 86768 69604 86792 69606
rect 86848 69604 86854 69606
rect 86546 69595 86854 69604
rect 86904 69320 86956 69326
rect 86904 69262 86956 69268
rect 88560 69320 88612 69326
rect 88560 69262 88612 69268
rect 86916 69161 86944 69262
rect 86902 69152 86958 69161
rect 86902 69087 86958 69096
rect 87282 69116 87590 69125
rect 87282 69114 87288 69116
rect 87344 69114 87368 69116
rect 87424 69114 87448 69116
rect 87504 69114 87528 69116
rect 87584 69114 87590 69116
rect 87344 69062 87346 69114
rect 87526 69062 87528 69114
rect 87282 69060 87288 69062
rect 87344 69060 87368 69062
rect 87424 69060 87448 69062
rect 87504 69060 87528 69062
rect 87584 69060 87590 69062
rect 87282 69051 87590 69060
rect 88572 69025 88600 69262
rect 88558 69016 88614 69025
rect 88558 68951 88614 68960
rect 86546 68572 86854 68581
rect 86546 68570 86552 68572
rect 86608 68570 86632 68572
rect 86688 68570 86712 68572
rect 86768 68570 86792 68572
rect 86848 68570 86854 68572
rect 86608 68518 86610 68570
rect 86790 68518 86792 68570
rect 86546 68516 86552 68518
rect 86608 68516 86632 68518
rect 86688 68516 86712 68518
rect 86768 68516 86792 68518
rect 86848 68516 86854 68518
rect 86546 68507 86854 68516
rect 87282 68028 87590 68037
rect 87282 68026 87288 68028
rect 87344 68026 87368 68028
rect 87424 68026 87448 68028
rect 87504 68026 87528 68028
rect 87584 68026 87590 68028
rect 87344 67974 87346 68026
rect 87526 67974 87528 68026
rect 87282 67972 87288 67974
rect 87344 67972 87368 67974
rect 87424 67972 87448 67974
rect 87504 67972 87528 67974
rect 87584 67972 87590 67974
rect 87282 67963 87590 67972
rect 84418 67928 84474 67937
rect 84418 67863 84474 67872
rect 84432 67694 84460 67863
rect 88284 67790 88336 67796
rect 88284 67732 88336 67738
rect 84420 67688 84472 67694
rect 88296 67665 88324 67732
rect 84420 67630 84472 67636
rect 88282 67656 88338 67665
rect 88282 67591 88338 67600
rect 86546 67484 86854 67493
rect 86546 67482 86552 67484
rect 86608 67482 86632 67484
rect 86688 67482 86712 67484
rect 86768 67482 86792 67484
rect 86848 67482 86854 67484
rect 86608 67430 86610 67482
rect 86790 67430 86792 67482
rect 86546 67428 86552 67430
rect 86608 67428 86632 67430
rect 86688 67428 86712 67430
rect 86768 67428 86792 67430
rect 86848 67428 86854 67430
rect 86546 67419 86854 67428
rect 88284 67172 88336 67178
rect 86904 67144 86956 67150
rect 88284 67114 88336 67120
rect 86904 67086 86956 67092
rect 86916 66985 86944 67086
rect 88296 66985 88324 67114
rect 86902 66976 86958 66985
rect 88282 66976 88338 66985
rect 86902 66911 86958 66920
rect 87282 66940 87590 66949
rect 87282 66938 87288 66940
rect 87344 66938 87368 66940
rect 87424 66938 87448 66940
rect 87504 66938 87528 66940
rect 87584 66938 87590 66940
rect 87344 66886 87346 66938
rect 87526 66886 87528 66938
rect 88282 66911 88338 66920
rect 87282 66884 87288 66886
rect 87344 66884 87368 66886
rect 87424 66884 87448 66886
rect 87504 66884 87528 66886
rect 87584 66884 87590 66886
rect 87282 66875 87590 66884
rect 86546 66396 86854 66405
rect 86546 66394 86552 66396
rect 86608 66394 86632 66396
rect 86688 66394 86712 66396
rect 86768 66394 86792 66396
rect 86848 66394 86854 66396
rect 86608 66342 86610 66394
rect 86790 66342 86792 66394
rect 86546 66340 86552 66342
rect 86608 66340 86632 66342
rect 86688 66340 86712 66342
rect 86768 66340 86792 66342
rect 86848 66340 86854 66342
rect 86546 66331 86854 66340
rect 87088 66056 87140 66062
rect 87088 65998 87140 66004
rect 87100 65897 87128 65998
rect 88192 65988 88244 65994
rect 88192 65930 88244 65936
rect 87086 65888 87142 65897
rect 87086 65823 87142 65832
rect 87282 65852 87590 65861
rect 87282 65850 87288 65852
rect 87344 65850 87368 65852
rect 87424 65850 87448 65852
rect 87504 65850 87528 65852
rect 87584 65850 87590 65852
rect 87344 65798 87346 65850
rect 87526 65798 87528 65850
rect 87282 65796 87288 65798
rect 87344 65796 87368 65798
rect 87424 65796 87448 65798
rect 87504 65796 87528 65798
rect 87584 65796 87590 65798
rect 87282 65787 87590 65796
rect 88204 65625 88232 65930
rect 88190 65616 88246 65625
rect 88190 65551 88246 65560
rect 86546 65308 86854 65317
rect 86546 65306 86552 65308
rect 86608 65306 86632 65308
rect 86688 65306 86712 65308
rect 86768 65306 86792 65308
rect 86848 65306 86854 65308
rect 86608 65254 86610 65306
rect 86790 65254 86792 65306
rect 86546 65252 86552 65254
rect 86608 65252 86632 65254
rect 86688 65252 86712 65254
rect 86768 65252 86792 65254
rect 86848 65252 86854 65254
rect 86546 65243 86854 65252
rect 87088 64968 87140 64974
rect 87088 64910 87140 64916
rect 88374 64936 88430 64945
rect 87100 64809 87128 64910
rect 88374 64871 88376 64880
rect 88428 64871 88430 64880
rect 88376 64842 88428 64848
rect 87086 64800 87142 64809
rect 87086 64735 87142 64744
rect 87282 64764 87590 64773
rect 87282 64762 87288 64764
rect 87344 64762 87368 64764
rect 87424 64762 87448 64764
rect 87504 64762 87528 64764
rect 87584 64762 87590 64764
rect 87344 64710 87346 64762
rect 87526 64710 87528 64762
rect 87282 64708 87288 64710
rect 87344 64708 87368 64710
rect 87424 64708 87448 64710
rect 87504 64708 87528 64710
rect 87584 64708 87590 64710
rect 87282 64699 87590 64708
rect 86546 64220 86854 64229
rect 86546 64218 86552 64220
rect 86608 64218 86632 64220
rect 86688 64218 86712 64220
rect 86768 64218 86792 64220
rect 86848 64218 86854 64220
rect 86608 64166 86610 64218
rect 86790 64166 86792 64218
rect 86546 64164 86552 64166
rect 86608 64164 86632 64166
rect 86688 64164 86712 64166
rect 86768 64164 86792 64166
rect 86848 64164 86854 64166
rect 86546 64155 86854 64164
rect 84420 63880 84472 63886
rect 84420 63822 84472 63828
rect 84432 63721 84460 63822
rect 88560 63812 88612 63818
rect 88560 63754 88612 63760
rect 84418 63712 84474 63721
rect 84418 63647 84474 63656
rect 87282 63676 87590 63685
rect 87282 63674 87288 63676
rect 87344 63674 87368 63676
rect 87424 63674 87448 63676
rect 87504 63674 87528 63676
rect 87584 63674 87590 63676
rect 87344 63622 87346 63674
rect 87526 63622 87528 63674
rect 87282 63620 87288 63622
rect 87344 63620 87368 63622
rect 87424 63620 87448 63622
rect 87504 63620 87528 63622
rect 87584 63620 87590 63622
rect 87282 63611 87590 63620
rect 88572 63585 88600 63754
rect 88558 63576 88614 63585
rect 88558 63511 88614 63520
rect 86546 63132 86854 63141
rect 86546 63130 86552 63132
rect 86608 63130 86632 63132
rect 86688 63130 86712 63132
rect 86768 63130 86792 63132
rect 86848 63130 86854 63132
rect 86608 63078 86610 63130
rect 86790 63078 86792 63130
rect 86546 63076 86552 63078
rect 86608 63076 86632 63078
rect 86688 63076 86712 63078
rect 86768 63076 86792 63078
rect 86848 63076 86854 63078
rect 86546 63067 86854 63076
rect 87282 62588 87590 62597
rect 87282 62586 87288 62588
rect 87344 62586 87368 62588
rect 87424 62586 87448 62588
rect 87504 62586 87528 62588
rect 87584 62586 87590 62588
rect 87344 62534 87346 62586
rect 87526 62534 87528 62586
rect 87282 62532 87288 62534
rect 87344 62532 87368 62534
rect 87424 62532 87448 62534
rect 87504 62532 87528 62534
rect 87584 62532 87590 62534
rect 87282 62523 87590 62532
rect 87086 62488 87142 62497
rect 87086 62423 87142 62432
rect 87100 62390 87128 62423
rect 87088 62384 87140 62390
rect 87088 62326 87140 62332
rect 88560 62384 88612 62390
rect 88560 62326 88612 62332
rect 88572 62225 88600 62326
rect 88558 62216 88614 62225
rect 88558 62151 88614 62160
rect 86546 62044 86854 62053
rect 86546 62042 86552 62044
rect 86608 62042 86632 62044
rect 86688 62042 86712 62044
rect 86768 62042 86792 62044
rect 86848 62042 86854 62044
rect 86608 61990 86610 62042
rect 86790 61990 86792 62042
rect 86546 61988 86552 61990
rect 86608 61988 86632 61990
rect 86688 61988 86712 61990
rect 86768 61988 86792 61990
rect 86848 61988 86854 61990
rect 86546 61979 86854 61988
rect 87088 61704 87140 61710
rect 87088 61646 87140 61652
rect 87100 61545 87128 61646
rect 88192 61636 88244 61642
rect 88192 61578 88244 61584
rect 88204 61545 88232 61578
rect 87086 61536 87142 61545
rect 88190 61536 88246 61545
rect 87086 61471 87142 61480
rect 87282 61500 87590 61509
rect 87282 61498 87288 61500
rect 87344 61498 87368 61500
rect 87424 61498 87448 61500
rect 87504 61498 87528 61500
rect 87584 61498 87590 61500
rect 87344 61446 87346 61498
rect 87526 61446 87528 61498
rect 88190 61471 88246 61480
rect 87282 61444 87288 61446
rect 87344 61444 87368 61446
rect 87424 61444 87448 61446
rect 87504 61444 87528 61446
rect 87584 61444 87590 61446
rect 87282 61435 87590 61444
rect 86546 60956 86854 60965
rect 86546 60954 86552 60956
rect 86608 60954 86632 60956
rect 86688 60954 86712 60956
rect 86768 60954 86792 60956
rect 86848 60954 86854 60956
rect 86608 60902 86610 60954
rect 86790 60902 86792 60954
rect 86546 60900 86552 60902
rect 86608 60900 86632 60902
rect 86688 60900 86712 60902
rect 86768 60900 86792 60902
rect 86848 60900 86854 60902
rect 86546 60891 86854 60900
rect 87088 60616 87140 60622
rect 87088 60558 87140 60564
rect 87100 60457 87128 60558
rect 88192 60548 88244 60554
rect 88192 60490 88244 60496
rect 87086 60448 87142 60457
rect 87086 60383 87142 60392
rect 87282 60412 87590 60421
rect 87282 60410 87288 60412
rect 87344 60410 87368 60412
rect 87424 60410 87448 60412
rect 87504 60410 87528 60412
rect 87584 60410 87590 60412
rect 87344 60358 87346 60410
rect 87526 60358 87528 60410
rect 87282 60356 87288 60358
rect 87344 60356 87368 60358
rect 87424 60356 87448 60358
rect 87504 60356 87528 60358
rect 87584 60356 87590 60358
rect 87282 60347 87590 60356
rect 88204 60185 88232 60490
rect 88190 60176 88246 60185
rect 88190 60111 88246 60120
rect 86546 59868 86854 59877
rect 86546 59866 86552 59868
rect 86608 59866 86632 59868
rect 86688 59866 86712 59868
rect 86768 59866 86792 59868
rect 86848 59866 86854 59868
rect 86608 59814 86610 59866
rect 86790 59814 86792 59866
rect 86546 59812 86552 59814
rect 86608 59812 86632 59814
rect 86688 59812 86712 59814
rect 86768 59812 86792 59814
rect 86848 59812 86854 59814
rect 86546 59803 86854 59812
rect 87640 59528 87692 59534
rect 87638 59496 87640 59505
rect 87692 59496 87694 59505
rect 87638 59431 87694 59440
rect 88374 59496 88430 59505
rect 88374 59431 88376 59440
rect 88428 59431 88430 59440
rect 88376 59402 88428 59408
rect 87282 59324 87590 59333
rect 87282 59322 87288 59324
rect 87344 59322 87368 59324
rect 87424 59322 87448 59324
rect 87504 59322 87528 59324
rect 87584 59322 87590 59324
rect 87344 59270 87346 59322
rect 87526 59270 87528 59322
rect 87282 59268 87288 59270
rect 87344 59268 87368 59270
rect 87424 59268 87448 59270
rect 87504 59268 87528 59270
rect 87584 59268 87590 59270
rect 87282 59259 87590 59268
rect 86546 58780 86854 58789
rect 86546 58778 86552 58780
rect 86608 58778 86632 58780
rect 86688 58778 86712 58780
rect 86768 58778 86792 58780
rect 86848 58778 86854 58780
rect 86608 58726 86610 58778
rect 86790 58726 86792 58778
rect 86546 58724 86552 58726
rect 86608 58724 86632 58726
rect 86688 58724 86712 58726
rect 86768 58724 86792 58726
rect 86848 58724 86854 58726
rect 86546 58715 86854 58724
rect 88008 58474 88060 58480
rect 88008 58416 88060 58422
rect 87282 58236 87590 58245
rect 87282 58234 87288 58236
rect 87344 58234 87368 58236
rect 87424 58234 87448 58236
rect 87504 58234 87528 58236
rect 87584 58234 87590 58236
rect 87344 58182 87346 58234
rect 87526 58182 87528 58234
rect 87282 58180 87288 58182
rect 87344 58180 87368 58182
rect 87424 58180 87448 58182
rect 87504 58180 87528 58182
rect 87584 58180 87590 58182
rect 87282 58171 87590 58180
rect 88020 58009 88048 58416
rect 88560 58372 88612 58378
rect 88560 58314 88612 58320
rect 88572 58145 88600 58314
rect 88558 58136 88614 58145
rect 88558 58071 88614 58080
rect 88006 58000 88062 58009
rect 88006 57935 88062 57944
rect 86546 57692 86854 57701
rect 86546 57690 86552 57692
rect 86608 57690 86632 57692
rect 86688 57690 86712 57692
rect 86768 57690 86792 57692
rect 86848 57690 86854 57692
rect 86608 57638 86610 57690
rect 86790 57638 86792 57690
rect 86546 57636 86552 57638
rect 86608 57636 86632 57638
rect 86688 57636 86712 57638
rect 86768 57636 86792 57638
rect 86848 57636 86854 57638
rect 86546 57627 86854 57636
rect 87282 57148 87590 57157
rect 87282 57146 87288 57148
rect 87344 57146 87368 57148
rect 87424 57146 87448 57148
rect 87504 57146 87528 57148
rect 87584 57146 87590 57148
rect 87344 57094 87346 57146
rect 87526 57094 87528 57146
rect 87282 57092 87288 57094
rect 87344 57092 87368 57094
rect 87424 57092 87448 57094
rect 87504 57092 87528 57094
rect 87584 57092 87590 57094
rect 87282 57083 87590 57092
rect 88006 56912 88062 56921
rect 88006 56847 88062 56856
rect 88836 56876 88888 56882
rect 88836 56818 88888 56824
rect 88848 56785 88876 56818
rect 88834 56776 88890 56785
rect 88834 56711 88890 56720
rect 86546 56604 86854 56613
rect 86546 56602 86552 56604
rect 86608 56602 86632 56604
rect 86688 56602 86712 56604
rect 86768 56602 86792 56604
rect 86848 56602 86854 56604
rect 86608 56550 86610 56602
rect 86790 56550 86792 56602
rect 86546 56548 86552 56550
rect 86608 56548 86632 56550
rect 86688 56548 86712 56550
rect 86768 56548 86792 56550
rect 86848 56548 86854 56550
rect 86546 56539 86854 56548
rect 87088 56264 87140 56270
rect 87088 56206 87140 56212
rect 87100 56105 87128 56206
rect 88192 56196 88244 56202
rect 88192 56138 88244 56144
rect 88204 56105 88232 56138
rect 87086 56096 87142 56105
rect 88190 56096 88246 56105
rect 87086 56031 87142 56040
rect 87282 56060 87590 56069
rect 87282 56058 87288 56060
rect 87344 56058 87368 56060
rect 87424 56058 87448 56060
rect 87504 56058 87528 56060
rect 87584 56058 87590 56060
rect 87344 56006 87346 56058
rect 87526 56006 87528 56058
rect 88190 56031 88246 56040
rect 87282 56004 87288 56006
rect 87344 56004 87368 56006
rect 87424 56004 87448 56006
rect 87504 56004 87528 56006
rect 87584 56004 87590 56006
rect 87282 55995 87590 56004
rect 86546 55516 86854 55525
rect 86546 55514 86552 55516
rect 86608 55514 86632 55516
rect 86688 55514 86712 55516
rect 86768 55514 86792 55516
rect 86848 55514 86854 55516
rect 86608 55462 86610 55514
rect 86790 55462 86792 55514
rect 86546 55460 86552 55462
rect 86608 55460 86632 55462
rect 86688 55460 86712 55462
rect 86768 55460 86792 55462
rect 86848 55460 86854 55462
rect 86546 55451 86854 55460
rect 87088 55176 87140 55182
rect 87088 55118 87140 55124
rect 87100 55017 87128 55118
rect 88192 55108 88244 55114
rect 88192 55050 88244 55056
rect 87086 55008 87142 55017
rect 87086 54943 87142 54952
rect 87282 54972 87590 54981
rect 87282 54970 87288 54972
rect 87344 54970 87368 54972
rect 87424 54970 87448 54972
rect 87504 54970 87528 54972
rect 87584 54970 87590 54972
rect 87344 54918 87346 54970
rect 87526 54918 87528 54970
rect 87282 54916 87288 54918
rect 87344 54916 87368 54918
rect 87424 54916 87448 54918
rect 87504 54916 87528 54918
rect 87584 54916 87590 54918
rect 87282 54907 87590 54916
rect 88204 54745 88232 55050
rect 88190 54736 88246 54745
rect 88190 54671 88246 54680
rect 86546 54428 86854 54437
rect 86546 54426 86552 54428
rect 86608 54426 86632 54428
rect 86688 54426 86712 54428
rect 86768 54426 86792 54428
rect 86848 54426 86854 54428
rect 86608 54374 86610 54426
rect 86790 54374 86792 54426
rect 86546 54372 86552 54374
rect 86608 54372 86632 54374
rect 86688 54372 86712 54374
rect 86768 54372 86792 54374
rect 86848 54372 86854 54374
rect 86546 54363 86854 54372
rect 84420 54088 84472 54094
rect 88652 54088 88704 54094
rect 84420 54030 84472 54036
rect 88650 54056 88652 54065
rect 88704 54056 88706 54065
rect 84432 53929 84460 54030
rect 88650 53991 88706 54000
rect 84418 53920 84474 53929
rect 84418 53855 84474 53864
rect 87282 53884 87590 53893
rect 87282 53882 87288 53884
rect 87344 53882 87368 53884
rect 87424 53882 87448 53884
rect 87504 53882 87528 53884
rect 87584 53882 87590 53884
rect 87344 53830 87346 53882
rect 87526 53830 87528 53882
rect 87282 53828 87288 53830
rect 87344 53828 87368 53830
rect 87424 53828 87448 53830
rect 87504 53828 87528 53830
rect 87584 53828 87590 53830
rect 87282 53819 87590 53828
rect 86546 53340 86854 53349
rect 86546 53338 86552 53340
rect 86608 53338 86632 53340
rect 86688 53338 86712 53340
rect 86768 53338 86792 53340
rect 86848 53338 86854 53340
rect 86608 53286 86610 53338
rect 86790 53286 86792 53338
rect 86546 53284 86552 53286
rect 86608 53284 86632 53286
rect 86688 53284 86712 53286
rect 86768 53284 86792 53286
rect 86848 53284 86854 53286
rect 86546 53275 86854 53284
rect 87088 53000 87140 53006
rect 87088 52942 87140 52948
rect 87100 52841 87128 52942
rect 88284 52932 88336 52938
rect 88284 52874 88336 52880
rect 87086 52832 87142 52841
rect 87086 52767 87142 52776
rect 87282 52796 87590 52805
rect 87282 52794 87288 52796
rect 87344 52794 87368 52796
rect 87424 52794 87448 52796
rect 87504 52794 87528 52796
rect 87584 52794 87590 52796
rect 87344 52742 87346 52794
rect 87526 52742 87528 52794
rect 87282 52740 87288 52742
rect 87344 52740 87368 52742
rect 87424 52740 87448 52742
rect 87504 52740 87528 52742
rect 87584 52740 87590 52742
rect 87282 52731 87590 52740
rect 88296 52705 88324 52874
rect 88282 52696 88338 52705
rect 88282 52631 88338 52640
rect 86546 52252 86854 52261
rect 86546 52250 86552 52252
rect 86608 52250 86632 52252
rect 86688 52250 86712 52252
rect 86768 52250 86792 52252
rect 86848 52250 86854 52252
rect 86608 52198 86610 52250
rect 86790 52198 86792 52250
rect 86546 52196 86552 52198
rect 86608 52196 86632 52198
rect 86688 52196 86712 52198
rect 86768 52196 86792 52198
rect 86848 52196 86854 52198
rect 86546 52187 86854 52196
rect 87282 51708 87590 51717
rect 87282 51706 87288 51708
rect 87344 51706 87368 51708
rect 87424 51706 87448 51708
rect 87504 51706 87528 51708
rect 87584 51706 87590 51708
rect 87344 51654 87346 51706
rect 87526 51654 87528 51706
rect 87282 51652 87288 51654
rect 87344 51652 87368 51654
rect 87424 51652 87448 51654
rect 87504 51652 87528 51654
rect 87584 51652 87590 51654
rect 87282 51643 87590 51652
rect 85798 51608 85854 51617
rect 85798 51543 85854 51552
rect 85812 51510 85840 51543
rect 85800 51504 85852 51510
rect 85800 51446 85852 51452
rect 88192 51368 88244 51374
rect 88190 51336 88192 51345
rect 88244 51336 88246 51345
rect 88190 51271 88246 51280
rect 86546 51164 86854 51173
rect 86546 51162 86552 51164
rect 86608 51162 86632 51164
rect 86688 51162 86712 51164
rect 86768 51162 86792 51164
rect 86848 51162 86854 51164
rect 86608 51110 86610 51162
rect 86790 51110 86792 51162
rect 86546 51108 86552 51110
rect 86608 51108 86632 51110
rect 86688 51108 86712 51110
rect 86768 51108 86792 51110
rect 86848 51108 86854 51110
rect 86546 51099 86854 51108
rect 85432 50756 85484 50762
rect 85432 50698 85484 50704
rect 85444 50529 85472 50698
rect 87282 50620 87590 50629
rect 87282 50618 87288 50620
rect 87344 50618 87368 50620
rect 87424 50618 87448 50620
rect 87504 50618 87528 50620
rect 87584 50618 87590 50620
rect 87344 50566 87346 50618
rect 87526 50566 87528 50618
rect 87282 50564 87288 50566
rect 87344 50564 87368 50566
rect 87424 50564 87448 50566
rect 87504 50564 87528 50566
rect 87584 50564 87590 50566
rect 87282 50555 87590 50564
rect 85430 50520 85486 50529
rect 85430 50455 85486 50464
rect 85340 48580 85392 48586
rect 85340 48522 85392 48528
rect 85352 48353 85380 48522
rect 85338 48344 85394 48353
rect 85338 48279 85394 48288
rect 84420 38992 84472 38998
rect 84420 38934 84472 38940
rect 84432 38153 84460 38934
rect 84418 38144 84474 38153
rect 84418 38079 84474 38088
rect 84420 36136 84472 36142
rect 84420 36078 84472 36084
rect 84432 35977 84460 36078
rect 84418 35968 84474 35977
rect 84418 35903 84474 35912
rect 84420 33416 84472 33422
rect 84420 33358 84472 33364
rect 84432 32713 84460 33358
rect 84418 32704 84474 32713
rect 84418 32639 84474 32648
rect 84420 30628 84472 30634
rect 84420 30570 84472 30576
rect 84432 30537 84460 30570
rect 84418 30528 84474 30537
rect 84418 30463 84474 30472
rect 85248 27976 85300 27982
rect 85248 27918 85300 27924
rect 85260 27273 85288 27918
rect 85246 27264 85302 27273
rect 85246 27199 85302 27208
rect 84420 22536 84472 22542
rect 84420 22478 84472 22484
rect 84432 21833 84460 22478
rect 84418 21824 84474 21833
rect 84418 21759 84474 21768
rect 84420 20972 84472 20978
rect 84420 20914 84472 20920
rect 84432 20745 84460 20914
rect 84418 20736 84474 20745
rect 84418 20671 84474 20680
rect 84420 15532 84472 15538
rect 84420 15474 84472 15480
rect 84432 15305 84460 15474
rect 84418 15296 84474 15305
rect 84418 15231 84474 15240
rect 83684 14308 83736 14314
rect 83684 14250 83736 14256
rect 83696 14217 83724 14250
rect 83682 14208 83738 14217
rect 83682 14143 83738 14152
rect 83500 13492 83552 13498
rect 83500 13434 83552 13440
rect 83512 13097 83540 13434
rect 83498 13088 83554 13097
rect 83420 13046 83498 13074
rect 83420 11882 83448 13046
rect 83498 13023 83554 13032
rect 83500 12404 83552 12410
rect 83500 12346 83552 12352
rect 83512 12009 83540 12346
rect 83498 12000 83554 12009
rect 83554 11958 83632 11986
rect 83498 11935 83554 11944
rect 83420 11854 83540 11882
rect 83408 11792 83460 11798
rect 83408 11734 83460 11740
rect 83316 11248 83368 11254
rect 83316 11190 83368 11196
rect 46422 10944 46478 10953
rect 46422 10879 46478 10888
rect 83328 10885 83356 11190
rect 83314 10876 83370 10885
rect 83314 10811 83370 10820
rect 82488 10228 82540 10234
rect 82488 10170 82540 10176
rect 82500 10114 82528 10170
rect 46068 8486 46188 8514
rect 45688 7508 45740 7514
rect 45688 7450 45740 7456
rect 45964 7508 46016 7514
rect 45964 7450 46016 7456
rect 45596 7440 45648 7446
rect 45596 7382 45648 7388
rect 45608 7242 45636 7382
rect 45976 7310 46004 7450
rect 46068 7446 46096 8486
rect 46056 7440 46108 7446
rect 46056 7382 46108 7388
rect 45964 7304 46016 7310
rect 45964 7246 46016 7252
rect 45596 7236 45648 7242
rect 45596 7178 45648 7184
rect 41640 5332 41692 5338
rect 41640 5274 41692 5280
rect 42836 5332 42888 5338
rect 42836 5274 42888 5280
rect 43664 5332 43716 5338
rect 43664 5274 43716 5280
rect 44768 5332 44820 5338
rect 44768 5274 44820 5280
rect 32716 5264 32768 5270
rect 32716 5206 32768 5212
rect 40444 5264 40496 5270
rect 40444 5206 40496 5212
rect 52416 5168 52444 10100
rect 53534 10086 53732 10114
rect 54638 10086 54928 10114
rect 53704 5168 53732 10086
rect 54522 7644 54830 7653
rect 54522 7642 54528 7644
rect 54584 7642 54608 7644
rect 54664 7642 54688 7644
rect 54744 7642 54768 7644
rect 54824 7642 54830 7644
rect 54584 7590 54586 7642
rect 54766 7590 54768 7642
rect 54522 7588 54528 7590
rect 54584 7588 54608 7590
rect 54664 7588 54688 7590
rect 54744 7588 54768 7590
rect 54824 7588 54830 7590
rect 54522 7579 54830 7588
rect 54522 6556 54830 6565
rect 54522 6554 54528 6556
rect 54584 6554 54608 6556
rect 54664 6554 54688 6556
rect 54744 6554 54768 6556
rect 54824 6554 54830 6556
rect 54584 6502 54586 6554
rect 54766 6502 54768 6554
rect 54522 6500 54528 6502
rect 54584 6500 54608 6502
rect 54664 6500 54688 6502
rect 54744 6500 54768 6502
rect 54824 6500 54830 6502
rect 54522 6491 54830 6500
rect 54522 5468 54830 5477
rect 54522 5466 54528 5468
rect 54584 5466 54608 5468
rect 54664 5466 54688 5468
rect 54744 5466 54768 5468
rect 54824 5466 54830 5468
rect 54584 5414 54586 5466
rect 54766 5414 54768 5466
rect 54522 5412 54528 5414
rect 54584 5412 54608 5414
rect 54664 5412 54688 5414
rect 54744 5412 54768 5414
rect 54824 5412 54830 5414
rect 54522 5403 54830 5412
rect 54900 5168 54928 10086
rect 55182 7100 55490 7109
rect 55182 7098 55188 7100
rect 55244 7098 55268 7100
rect 55324 7098 55348 7100
rect 55404 7098 55428 7100
rect 55484 7098 55490 7100
rect 55244 7046 55246 7098
rect 55426 7046 55428 7098
rect 55182 7044 55188 7046
rect 55244 7044 55268 7046
rect 55324 7044 55348 7046
rect 55404 7044 55428 7046
rect 55484 7044 55490 7046
rect 55182 7035 55490 7044
rect 55182 6012 55490 6021
rect 55182 6010 55188 6012
rect 55244 6010 55268 6012
rect 55324 6010 55348 6012
rect 55404 6010 55428 6012
rect 55484 6010 55490 6012
rect 55244 5958 55246 6010
rect 55426 5958 55428 6010
rect 55182 5956 55188 5958
rect 55244 5956 55268 5958
rect 55324 5956 55348 5958
rect 55404 5956 55428 5958
rect 55484 5956 55490 5958
rect 55182 5947 55490 5956
rect 55728 5168 55756 10100
rect 56832 5168 56860 10100
rect 57936 5168 57964 10100
rect 59040 5168 59068 10100
rect 60144 5168 60172 10100
rect 61262 10086 61460 10114
rect 61432 5168 61460 10086
rect 62352 5168 62380 10100
rect 63456 5168 63484 10100
rect 64560 5168 64588 10100
rect 65664 5168 65692 10100
rect 66768 5168 66796 10100
rect 67872 5338 67900 10100
rect 68990 10086 69372 10114
rect 69344 5338 69372 10086
rect 67860 5332 67912 5338
rect 67860 5274 67912 5280
rect 69332 5332 69384 5338
rect 69332 5274 69384 5280
rect 70080 5270 70108 10100
rect 71184 5338 71212 10100
rect 72288 5338 72316 10100
rect 72922 7644 73230 7653
rect 72922 7642 72928 7644
rect 72984 7642 73008 7644
rect 73064 7642 73088 7644
rect 73144 7642 73168 7644
rect 73224 7642 73230 7644
rect 72984 7590 72986 7642
rect 73166 7590 73168 7642
rect 72922 7588 72928 7590
rect 72984 7588 73008 7590
rect 73064 7588 73088 7590
rect 73144 7588 73168 7590
rect 73224 7588 73230 7590
rect 72922 7579 73230 7588
rect 72922 6556 73230 6565
rect 72922 6554 72928 6556
rect 72984 6554 73008 6556
rect 73064 6554 73088 6556
rect 73144 6554 73168 6556
rect 73224 6554 73230 6556
rect 72984 6502 72986 6554
rect 73166 6502 73168 6554
rect 72922 6500 72928 6502
rect 72984 6500 73008 6502
rect 73064 6500 73088 6502
rect 73144 6500 73168 6502
rect 73224 6500 73230 6502
rect 72922 6491 73230 6500
rect 72922 5468 73230 5477
rect 72922 5466 72928 5468
rect 72984 5466 73008 5468
rect 73064 5466 73088 5468
rect 73144 5466 73168 5468
rect 73224 5466 73230 5468
rect 72984 5414 72986 5466
rect 73166 5414 73168 5466
rect 72922 5412 72928 5414
rect 72984 5412 73008 5414
rect 73064 5412 73088 5414
rect 73144 5412 73168 5414
rect 73224 5412 73230 5414
rect 72922 5403 73230 5412
rect 73392 5338 73420 10100
rect 73582 7100 73890 7109
rect 73582 7098 73588 7100
rect 73644 7098 73668 7100
rect 73724 7098 73748 7100
rect 73804 7098 73828 7100
rect 73884 7098 73890 7100
rect 73644 7046 73646 7098
rect 73826 7046 73828 7098
rect 73582 7044 73588 7046
rect 73644 7044 73668 7046
rect 73724 7044 73748 7046
rect 73804 7044 73828 7046
rect 73884 7044 73890 7046
rect 73582 7035 73890 7044
rect 73582 6012 73890 6021
rect 73582 6010 73588 6012
rect 73644 6010 73668 6012
rect 73724 6010 73748 6012
rect 73804 6010 73828 6012
rect 73884 6010 73890 6012
rect 73644 5958 73646 6010
rect 73826 5958 73828 6010
rect 73582 5956 73588 5958
rect 73644 5956 73668 5958
rect 73724 5956 73748 5958
rect 73804 5956 73828 5958
rect 73884 5956 73890 5958
rect 73582 5947 73890 5956
rect 74496 5338 74524 10100
rect 75600 5338 75628 10100
rect 76704 5338 76732 10100
rect 71172 5332 71224 5338
rect 71172 5274 71224 5280
rect 72276 5332 72328 5338
rect 72276 5274 72328 5280
rect 73380 5332 73432 5338
rect 73380 5274 73432 5280
rect 74484 5332 74536 5338
rect 74484 5274 74536 5280
rect 75588 5332 75640 5338
rect 75588 5274 75640 5280
rect 76692 5332 76744 5338
rect 76692 5274 76744 5280
rect 77808 5270 77836 10100
rect 78912 5338 78940 10100
rect 80030 10086 80320 10114
rect 81134 10086 81424 10114
rect 82238 10086 82528 10114
rect 80292 5338 80320 10086
rect 81396 10030 81424 10086
rect 81384 10024 81436 10030
rect 81384 9966 81436 9972
rect 83420 7310 83448 11734
rect 83512 7378 83540 11854
rect 83500 7372 83552 7378
rect 83500 7314 83552 7320
rect 83408 7304 83460 7310
rect 83408 7246 83460 7252
rect 83604 7242 83632 11958
rect 83696 11798 83724 14143
rect 85352 12410 85380 48279
rect 85444 14994 85472 50455
rect 86546 50076 86854 50085
rect 86546 50074 86552 50076
rect 86608 50074 86632 50076
rect 86688 50074 86712 50076
rect 86768 50074 86792 50076
rect 86848 50074 86854 50076
rect 86608 50022 86610 50074
rect 86790 50022 86792 50074
rect 86546 50020 86552 50022
rect 86608 50020 86632 50022
rect 86688 50020 86712 50022
rect 86768 50020 86792 50022
rect 86848 50020 86854 50022
rect 86546 50011 86854 50020
rect 85524 49668 85576 49674
rect 85524 49610 85576 49616
rect 85536 49441 85564 49610
rect 87282 49532 87590 49541
rect 87282 49530 87288 49532
rect 87344 49530 87368 49532
rect 87424 49530 87448 49532
rect 87504 49530 87528 49532
rect 87584 49530 87590 49532
rect 87344 49478 87346 49530
rect 87526 49478 87528 49530
rect 87282 49476 87288 49478
rect 87344 49476 87368 49478
rect 87424 49476 87448 49478
rect 87504 49476 87528 49478
rect 87584 49476 87590 49478
rect 87282 49467 87590 49476
rect 85522 49432 85578 49441
rect 85522 49367 85578 49376
rect 85432 14988 85484 14994
rect 85432 14930 85484 14936
rect 85536 13498 85564 49367
rect 86546 48988 86854 48997
rect 86546 48986 86552 48988
rect 86608 48986 86632 48988
rect 86688 48986 86712 48988
rect 86768 48986 86792 48988
rect 86848 48986 86854 48988
rect 86608 48934 86610 48986
rect 86790 48934 86792 48986
rect 86546 48932 86552 48934
rect 86608 48932 86632 48934
rect 86688 48932 86712 48934
rect 86768 48932 86792 48934
rect 86848 48932 86854 48934
rect 86546 48923 86854 48932
rect 88192 48648 88244 48654
rect 88190 48616 88192 48625
rect 88244 48616 88246 48625
rect 88190 48551 88246 48560
rect 87282 48444 87590 48453
rect 87282 48442 87288 48444
rect 87344 48442 87368 48444
rect 87424 48442 87448 48444
rect 87504 48442 87528 48444
rect 87584 48442 87590 48444
rect 87344 48390 87346 48442
rect 87526 48390 87528 48442
rect 87282 48388 87288 48390
rect 87344 48388 87368 48390
rect 87424 48388 87448 48390
rect 87504 48388 87528 48390
rect 87584 48388 87590 48390
rect 87282 48379 87590 48388
rect 88192 48036 88244 48042
rect 88192 47978 88244 47984
rect 88204 47945 88232 47978
rect 88190 47936 88246 47945
rect 86546 47900 86854 47909
rect 86546 47898 86552 47900
rect 86608 47898 86632 47900
rect 86688 47898 86712 47900
rect 86768 47898 86792 47900
rect 86848 47898 86854 47900
rect 86608 47846 86610 47898
rect 86790 47846 86792 47898
rect 88190 47871 88246 47880
rect 86546 47844 86552 47846
rect 86608 47844 86632 47846
rect 86688 47844 86712 47846
rect 86768 47844 86792 47846
rect 86848 47844 86854 47846
rect 86546 47835 86854 47844
rect 85800 47560 85852 47566
rect 85800 47502 85852 47508
rect 85812 47401 85840 47502
rect 88192 47492 88244 47498
rect 88192 47434 88244 47440
rect 85798 47392 85854 47401
rect 85798 47327 85854 47336
rect 87282 47356 87590 47365
rect 87282 47354 87288 47356
rect 87344 47354 87368 47356
rect 87424 47354 87448 47356
rect 87504 47354 87528 47356
rect 87584 47354 87590 47356
rect 87344 47302 87346 47354
rect 87526 47302 87528 47354
rect 87282 47300 87288 47302
rect 87344 47300 87368 47302
rect 87424 47300 87448 47302
rect 87504 47300 87528 47302
rect 87584 47300 87590 47302
rect 87282 47291 87590 47300
rect 88204 47265 88232 47434
rect 88190 47256 88246 47265
rect 88190 47191 88246 47200
rect 88192 46948 88244 46954
rect 88192 46890 88244 46896
rect 86546 46812 86854 46821
rect 86546 46810 86552 46812
rect 86608 46810 86632 46812
rect 86688 46810 86712 46812
rect 86768 46810 86792 46812
rect 86848 46810 86854 46812
rect 86608 46758 86610 46810
rect 86790 46758 86792 46810
rect 86546 46756 86552 46758
rect 86608 46756 86632 46758
rect 86688 46756 86712 46758
rect 86768 46756 86792 46758
rect 86848 46756 86854 46758
rect 86546 46747 86854 46756
rect 88204 46585 88232 46890
rect 88190 46576 88246 46585
rect 88190 46511 88246 46520
rect 87282 46268 87590 46277
rect 87282 46266 87288 46268
rect 87344 46266 87368 46268
rect 87424 46266 87448 46268
rect 87504 46266 87528 46268
rect 87584 46266 87590 46268
rect 87344 46214 87346 46266
rect 87526 46214 87528 46266
rect 87282 46212 87288 46214
rect 87344 46212 87368 46214
rect 87424 46212 87448 46214
rect 87504 46212 87528 46214
rect 87584 46212 87590 46214
rect 87282 46203 87590 46212
rect 85800 45928 85852 45934
rect 85800 45870 85852 45876
rect 88190 45896 88246 45905
rect 85812 45594 85840 45870
rect 88190 45831 88192 45840
rect 88244 45831 88246 45840
rect 88192 45802 88244 45808
rect 86546 45724 86854 45733
rect 86546 45722 86552 45724
rect 86608 45722 86632 45724
rect 86688 45722 86712 45724
rect 86768 45722 86792 45724
rect 86848 45722 86854 45724
rect 86608 45670 86610 45722
rect 86790 45670 86792 45722
rect 86546 45668 86552 45670
rect 86608 45668 86632 45670
rect 86688 45668 86712 45670
rect 86768 45668 86792 45670
rect 86848 45668 86854 45670
rect 86546 45659 86854 45668
rect 85800 45588 85852 45594
rect 85800 45530 85852 45536
rect 85984 45520 86036 45526
rect 85982 45488 85984 45497
rect 86036 45488 86038 45497
rect 85982 45423 86038 45432
rect 86168 45384 86220 45390
rect 86166 45352 86168 45361
rect 88192 45384 88244 45390
rect 86220 45352 86222 45361
rect 85616 45316 85668 45322
rect 88192 45326 88244 45332
rect 86166 45287 86222 45296
rect 85616 45258 85668 45264
rect 85628 45225 85656 45258
rect 88204 45225 88232 45326
rect 85614 45216 85670 45225
rect 88190 45216 88246 45225
rect 85614 45151 85670 45160
rect 87282 45180 87590 45189
rect 87282 45178 87288 45180
rect 87344 45178 87368 45180
rect 87424 45178 87448 45180
rect 87504 45178 87528 45180
rect 87584 45178 87590 45180
rect 87344 45126 87346 45178
rect 87526 45126 87528 45178
rect 88190 45151 88246 45160
rect 87282 45124 87288 45126
rect 87344 45124 87368 45126
rect 87424 45124 87448 45126
rect 87504 45124 87528 45126
rect 87584 45124 87590 45126
rect 87282 45115 87590 45124
rect 88284 44942 88336 44948
rect 88284 44884 88336 44890
rect 87180 44840 87232 44846
rect 87178 44808 87180 44817
rect 87232 44808 87234 44817
rect 87178 44743 87234 44752
rect 86546 44636 86854 44645
rect 86546 44634 86552 44636
rect 86608 44634 86632 44636
rect 86688 44634 86712 44636
rect 86768 44634 86792 44636
rect 86848 44634 86854 44636
rect 86608 44582 86610 44634
rect 86790 44582 86792 44634
rect 86546 44580 86552 44582
rect 86608 44580 86632 44582
rect 86688 44580 86712 44582
rect 86768 44580 86792 44582
rect 86848 44580 86854 44582
rect 86546 44571 86854 44580
rect 88296 44545 88324 44884
rect 88282 44536 88338 44545
rect 88282 44471 88338 44480
rect 88284 44324 88336 44330
rect 85800 44296 85852 44302
rect 88284 44266 88336 44272
rect 85800 44238 85852 44244
rect 85812 43593 85840 44238
rect 87282 44092 87590 44101
rect 87282 44090 87288 44092
rect 87344 44090 87368 44092
rect 87424 44090 87448 44092
rect 87504 44090 87528 44092
rect 87584 44090 87590 44092
rect 87344 44038 87346 44090
rect 87526 44038 87528 44090
rect 87282 44036 87288 44038
rect 87344 44036 87368 44038
rect 87424 44036 87448 44038
rect 87504 44036 87528 44038
rect 87584 44036 87590 44038
rect 87282 44027 87590 44036
rect 88296 43865 88324 44266
rect 88282 43856 88338 43865
rect 88282 43791 88338 43800
rect 85798 43584 85854 43593
rect 85798 43519 85854 43528
rect 86546 43548 86854 43557
rect 86546 43546 86552 43548
rect 86608 43546 86632 43548
rect 86688 43546 86712 43548
rect 86768 43546 86792 43548
rect 86848 43546 86854 43548
rect 86608 43494 86610 43546
rect 86790 43494 86792 43546
rect 86546 43492 86552 43494
rect 86608 43492 86632 43494
rect 86688 43492 86712 43494
rect 86768 43492 86792 43494
rect 86848 43492 86854 43494
rect 86546 43483 86854 43492
rect 87282 43004 87590 43013
rect 87282 43002 87288 43004
rect 87344 43002 87368 43004
rect 87424 43002 87448 43004
rect 87504 43002 87528 43004
rect 87584 43002 87590 43004
rect 87344 42950 87346 43002
rect 87526 42950 87528 43002
rect 87282 42948 87288 42950
rect 87344 42948 87368 42950
rect 87424 42948 87448 42950
rect 87504 42948 87528 42950
rect 87584 42948 87590 42950
rect 87282 42939 87590 42948
rect 88284 42766 88336 42772
rect 88284 42708 88336 42714
rect 86352 42664 86404 42670
rect 86352 42606 86404 42612
rect 86364 42505 86392 42606
rect 88296 42505 88324 42708
rect 86350 42496 86406 42505
rect 88282 42496 88338 42505
rect 86350 42431 86406 42440
rect 86546 42460 86854 42469
rect 86546 42458 86552 42460
rect 86608 42458 86632 42460
rect 86688 42458 86712 42460
rect 86768 42458 86792 42460
rect 86848 42458 86854 42460
rect 86608 42406 86610 42458
rect 86790 42406 86792 42458
rect 88282 42431 88338 42440
rect 86546 42404 86552 42406
rect 86608 42404 86632 42406
rect 86688 42404 86712 42406
rect 86768 42404 86792 42406
rect 86848 42404 86854 42406
rect 86546 42395 86854 42404
rect 87282 41916 87590 41925
rect 87282 41914 87288 41916
rect 87344 41914 87368 41916
rect 87424 41914 87448 41916
rect 87504 41914 87528 41916
rect 87584 41914 87590 41916
rect 87344 41862 87346 41914
rect 87526 41862 87528 41914
rect 87282 41860 87288 41862
rect 87344 41860 87368 41862
rect 87424 41860 87448 41862
rect 87504 41860 87528 41862
rect 87584 41860 87590 41862
rect 87282 41851 87590 41860
rect 87180 41780 87232 41786
rect 87180 41722 87232 41728
rect 87192 41553 87220 41722
rect 88284 41678 88336 41684
rect 88284 41620 88336 41626
rect 87178 41544 87234 41553
rect 87178 41479 87234 41488
rect 86546 41372 86854 41381
rect 86546 41370 86552 41372
rect 86608 41370 86632 41372
rect 86688 41370 86712 41372
rect 86768 41370 86792 41372
rect 86848 41370 86854 41372
rect 86608 41318 86610 41370
rect 86790 41318 86792 41370
rect 86546 41316 86552 41318
rect 86608 41316 86632 41318
rect 86688 41316 86712 41318
rect 86768 41316 86792 41318
rect 86848 41316 86854 41318
rect 86546 41307 86854 41316
rect 88296 41145 88324 41620
rect 88282 41136 88338 41145
rect 88282 41071 88338 41080
rect 87282 40828 87590 40837
rect 87282 40826 87288 40828
rect 87344 40826 87368 40828
rect 87424 40826 87448 40828
rect 87504 40826 87528 40828
rect 87584 40826 87590 40828
rect 87344 40774 87346 40826
rect 87526 40774 87528 40826
rect 87282 40772 87288 40774
rect 87344 40772 87368 40774
rect 87424 40772 87448 40774
rect 87504 40772 87528 40774
rect 87584 40772 87590 40774
rect 87282 40763 87590 40772
rect 87916 40556 87968 40562
rect 87916 40498 87968 40504
rect 88284 40556 88336 40562
rect 88284 40498 88336 40504
rect 87928 40465 87956 40498
rect 88296 40465 88324 40498
rect 87914 40456 87970 40465
rect 87914 40391 87970 40400
rect 88282 40456 88338 40465
rect 88282 40391 88338 40400
rect 86546 40284 86854 40293
rect 86546 40282 86552 40284
rect 86608 40282 86632 40284
rect 86688 40282 86712 40284
rect 86768 40282 86792 40284
rect 86848 40282 86854 40284
rect 86608 40230 86610 40282
rect 86790 40230 86792 40282
rect 86546 40228 86552 40230
rect 86608 40228 86632 40230
rect 86688 40228 86712 40230
rect 86768 40228 86792 40230
rect 86848 40228 86854 40230
rect 86546 40219 86854 40228
rect 88296 40154 88324 40391
rect 88284 40148 88336 40154
rect 88284 40090 88336 40096
rect 87282 39740 87590 39749
rect 87282 39738 87288 39740
rect 87344 39738 87368 39740
rect 87424 39738 87448 39740
rect 87504 39738 87528 39740
rect 87584 39738 87590 39740
rect 87344 39686 87346 39738
rect 87526 39686 87528 39738
rect 87282 39684 87288 39686
rect 87344 39684 87368 39686
rect 87424 39684 87448 39686
rect 87504 39684 87528 39686
rect 87584 39684 87590 39686
rect 87282 39675 87590 39684
rect 88284 39502 88336 39508
rect 88284 39444 88336 39450
rect 87180 39400 87232 39406
rect 87178 39368 87180 39377
rect 87232 39368 87234 39377
rect 87178 39303 87234 39312
rect 86546 39196 86854 39205
rect 86546 39194 86552 39196
rect 86608 39194 86632 39196
rect 86688 39194 86712 39196
rect 86768 39194 86792 39196
rect 86848 39194 86854 39196
rect 86608 39142 86610 39194
rect 86790 39142 86792 39194
rect 86546 39140 86552 39142
rect 86608 39140 86632 39142
rect 86688 39140 86712 39142
rect 86768 39140 86792 39142
rect 86848 39140 86854 39142
rect 86546 39131 86854 39140
rect 88296 39105 88324 39444
rect 88282 39096 88338 39105
rect 88282 39031 88338 39040
rect 88284 38890 88336 38896
rect 88284 38832 88336 38838
rect 87282 38652 87590 38661
rect 87282 38650 87288 38652
rect 87344 38650 87368 38652
rect 87424 38650 87448 38652
rect 87504 38650 87528 38652
rect 87584 38650 87590 38652
rect 87344 38598 87346 38650
rect 87526 38598 87528 38650
rect 87282 38596 87288 38598
rect 87344 38596 87368 38598
rect 87424 38596 87448 38598
rect 87504 38596 87528 38598
rect 87584 38596 87590 38598
rect 87282 38587 87590 38596
rect 88296 38425 88324 38832
rect 88282 38416 88338 38425
rect 88282 38351 88338 38360
rect 86546 38108 86854 38117
rect 86546 38106 86552 38108
rect 86608 38106 86632 38108
rect 86688 38106 86712 38108
rect 86768 38106 86792 38108
rect 86848 38106 86854 38108
rect 86608 38054 86610 38106
rect 86790 38054 86792 38106
rect 86546 38052 86552 38054
rect 86608 38052 86632 38054
rect 86688 38052 86712 38054
rect 86768 38052 86792 38054
rect 86848 38052 86854 38054
rect 86546 38043 86854 38052
rect 87282 37564 87590 37573
rect 87282 37562 87288 37564
rect 87344 37562 87368 37564
rect 87424 37562 87448 37564
rect 87504 37562 87528 37564
rect 87584 37562 87590 37564
rect 87344 37510 87346 37562
rect 87526 37510 87528 37562
rect 87282 37508 87288 37510
rect 87344 37508 87368 37510
rect 87424 37508 87448 37510
rect 87504 37508 87528 37510
rect 87584 37508 87590 37510
rect 87282 37499 87590 37508
rect 88284 37326 88336 37332
rect 88284 37268 88336 37274
rect 86352 37224 86404 37230
rect 86352 37166 86404 37172
rect 86364 37065 86392 37166
rect 88296 37065 88324 37268
rect 86350 37056 86406 37065
rect 88282 37056 88338 37065
rect 86350 36991 86406 37000
rect 86546 37020 86854 37029
rect 86546 37018 86552 37020
rect 86608 37018 86632 37020
rect 86688 37018 86712 37020
rect 86768 37018 86792 37020
rect 86848 37018 86854 37020
rect 86608 36966 86610 37018
rect 86790 36966 86792 37018
rect 88282 36991 88338 37000
rect 86546 36964 86552 36966
rect 86608 36964 86632 36966
rect 86688 36964 86712 36966
rect 86768 36964 86792 36966
rect 86848 36964 86854 36966
rect 86546 36955 86854 36964
rect 87282 36476 87590 36485
rect 87282 36474 87288 36476
rect 87344 36474 87368 36476
rect 87424 36474 87448 36476
rect 87504 36474 87528 36476
rect 87584 36474 87590 36476
rect 87344 36422 87346 36474
rect 87526 36422 87528 36474
rect 87282 36420 87288 36422
rect 87344 36420 87368 36422
rect 87424 36420 87448 36422
rect 87504 36420 87528 36422
rect 87584 36420 87590 36422
rect 87282 36411 87590 36420
rect 88560 36204 88612 36210
rect 88560 36146 88612 36152
rect 86546 35932 86854 35941
rect 86546 35930 86552 35932
rect 86608 35930 86632 35932
rect 86688 35930 86712 35932
rect 86768 35930 86792 35932
rect 86848 35930 86854 35932
rect 86608 35878 86610 35930
rect 86790 35878 86792 35930
rect 86546 35876 86552 35878
rect 86608 35876 86632 35878
rect 86688 35876 86712 35878
rect 86768 35876 86792 35878
rect 86848 35876 86854 35878
rect 86546 35867 86854 35876
rect 88572 35705 88600 36146
rect 88558 35696 88614 35705
rect 88558 35631 88614 35640
rect 87282 35388 87590 35397
rect 87282 35386 87288 35388
rect 87344 35386 87368 35388
rect 87424 35386 87448 35388
rect 87504 35386 87528 35388
rect 87584 35386 87590 35388
rect 87344 35334 87346 35386
rect 87526 35334 87528 35386
rect 87282 35332 87288 35334
rect 87344 35332 87368 35334
rect 87424 35332 87448 35334
rect 87504 35332 87528 35334
rect 87584 35332 87590 35334
rect 87282 35323 87590 35332
rect 88284 35150 88336 35156
rect 88284 35092 88336 35098
rect 86352 35048 86404 35054
rect 88296 35025 88324 35092
rect 86352 34990 86404 34996
rect 88282 35016 88338 35025
rect 86364 34889 86392 34990
rect 88282 34951 88338 34960
rect 86350 34880 86406 34889
rect 86350 34815 86406 34824
rect 86546 34844 86854 34853
rect 86546 34842 86552 34844
rect 86608 34842 86632 34844
rect 86688 34842 86712 34844
rect 86768 34842 86792 34844
rect 86848 34842 86854 34844
rect 86608 34790 86610 34842
rect 86790 34790 86792 34842
rect 86546 34788 86552 34790
rect 86608 34788 86632 34790
rect 86688 34788 86712 34790
rect 86768 34788 86792 34790
rect 86848 34788 86854 34790
rect 86546 34779 86854 34788
rect 87282 34300 87590 34309
rect 87282 34298 87288 34300
rect 87344 34298 87368 34300
rect 87424 34298 87448 34300
rect 87504 34298 87528 34300
rect 87584 34298 87590 34300
rect 87344 34246 87346 34298
rect 87526 34246 87528 34298
rect 87282 34244 87288 34246
rect 87344 34244 87368 34246
rect 87424 34244 87448 34246
rect 87504 34244 87528 34246
rect 87584 34244 87590 34246
rect 87282 34235 87590 34244
rect 88284 34062 88336 34068
rect 88284 34004 88336 34010
rect 86352 33960 86404 33966
rect 86352 33902 86404 33908
rect 86364 33801 86392 33902
rect 86350 33792 86406 33801
rect 86350 33727 86406 33736
rect 86546 33756 86854 33765
rect 86546 33754 86552 33756
rect 86608 33754 86632 33756
rect 86688 33754 86712 33756
rect 86768 33754 86792 33756
rect 86848 33754 86854 33756
rect 86608 33702 86610 33754
rect 86790 33702 86792 33754
rect 86546 33700 86552 33702
rect 86608 33700 86632 33702
rect 86688 33700 86712 33702
rect 86768 33700 86792 33702
rect 86848 33700 86854 33702
rect 86546 33691 86854 33700
rect 88296 33665 88324 34004
rect 88282 33656 88338 33665
rect 88282 33591 88338 33600
rect 88560 33416 88612 33422
rect 88560 33358 88612 33364
rect 87282 33212 87590 33221
rect 87282 33210 87288 33212
rect 87344 33210 87368 33212
rect 87424 33210 87448 33212
rect 87504 33210 87528 33212
rect 87584 33210 87590 33212
rect 87344 33158 87346 33210
rect 87526 33158 87528 33210
rect 87282 33156 87288 33158
rect 87344 33156 87368 33158
rect 87424 33156 87448 33158
rect 87504 33156 87528 33158
rect 87584 33156 87590 33158
rect 87282 33147 87590 33156
rect 88572 32985 88600 33358
rect 88558 32976 88614 32985
rect 88558 32911 88614 32920
rect 86546 32668 86854 32677
rect 86546 32666 86552 32668
rect 86608 32666 86632 32668
rect 86688 32666 86712 32668
rect 86768 32666 86792 32668
rect 86848 32666 86854 32668
rect 86608 32614 86610 32666
rect 86790 32614 86792 32666
rect 86546 32612 86552 32614
rect 86608 32612 86632 32614
rect 86688 32612 86712 32614
rect 86768 32612 86792 32614
rect 86848 32612 86854 32614
rect 86546 32603 86854 32612
rect 87282 32124 87590 32133
rect 87282 32122 87288 32124
rect 87344 32122 87368 32124
rect 87424 32122 87448 32124
rect 87504 32122 87528 32124
rect 87584 32122 87590 32124
rect 87344 32070 87346 32122
rect 87526 32070 87528 32122
rect 87282 32068 87288 32070
rect 87344 32068 87368 32070
rect 87424 32068 87448 32070
rect 87504 32068 87528 32070
rect 87584 32068 87590 32070
rect 87282 32059 87590 32068
rect 88284 31886 88336 31892
rect 88284 31828 88336 31834
rect 86352 31784 86404 31790
rect 86352 31726 86404 31732
rect 86364 31625 86392 31726
rect 88296 31625 88324 31828
rect 86350 31616 86406 31625
rect 88282 31616 88338 31625
rect 86350 31551 86406 31560
rect 86546 31580 86854 31589
rect 86546 31578 86552 31580
rect 86608 31578 86632 31580
rect 86688 31578 86712 31580
rect 86768 31578 86792 31580
rect 86848 31578 86854 31580
rect 86608 31526 86610 31578
rect 86790 31526 86792 31578
rect 88282 31551 88338 31560
rect 86546 31524 86552 31526
rect 86608 31524 86632 31526
rect 86688 31524 86712 31526
rect 86768 31524 86792 31526
rect 86848 31524 86854 31526
rect 86546 31515 86854 31524
rect 87282 31036 87590 31045
rect 87282 31034 87288 31036
rect 87344 31034 87368 31036
rect 87424 31034 87448 31036
rect 87504 31034 87528 31036
rect 87584 31034 87590 31036
rect 87344 30982 87346 31034
rect 87526 30982 87528 31034
rect 87282 30980 87288 30982
rect 87344 30980 87368 30982
rect 87424 30980 87448 30982
rect 87504 30980 87528 30982
rect 87584 30980 87590 30982
rect 87282 30971 87590 30980
rect 88560 30764 88612 30770
rect 88560 30706 88612 30712
rect 86546 30492 86854 30501
rect 86546 30490 86552 30492
rect 86608 30490 86632 30492
rect 86688 30490 86712 30492
rect 86768 30490 86792 30492
rect 86848 30490 86854 30492
rect 86608 30438 86610 30490
rect 86790 30438 86792 30490
rect 86546 30436 86552 30438
rect 86608 30436 86632 30438
rect 86688 30436 86712 30438
rect 86768 30436 86792 30438
rect 86848 30436 86854 30438
rect 86546 30427 86854 30436
rect 88572 30265 88600 30706
rect 88558 30256 88614 30265
rect 88558 30191 88614 30200
rect 87282 29948 87590 29957
rect 87282 29946 87288 29948
rect 87344 29946 87368 29948
rect 87424 29946 87448 29948
rect 87504 29946 87528 29948
rect 87584 29946 87590 29948
rect 87344 29894 87346 29946
rect 87526 29894 87528 29946
rect 87282 29892 87288 29894
rect 87344 29892 87368 29894
rect 87424 29892 87448 29894
rect 87504 29892 87528 29894
rect 87584 29892 87590 29894
rect 87282 29883 87590 29892
rect 86352 29676 86404 29682
rect 86352 29618 86404 29624
rect 86364 29449 86392 29618
rect 88282 29576 88338 29585
rect 88282 29511 88284 29520
rect 88336 29511 88338 29520
rect 88284 29482 88336 29488
rect 86350 29440 86406 29449
rect 86350 29375 86406 29384
rect 86546 29404 86854 29413
rect 86546 29402 86552 29404
rect 86608 29402 86632 29404
rect 86688 29402 86712 29404
rect 86768 29402 86792 29404
rect 86848 29402 86854 29404
rect 86608 29350 86610 29402
rect 86790 29350 86792 29402
rect 86546 29348 86552 29350
rect 86608 29348 86632 29350
rect 86688 29348 86712 29350
rect 86768 29348 86792 29350
rect 86848 29348 86854 29350
rect 86546 29339 86854 29348
rect 87282 28860 87590 28869
rect 87282 28858 87288 28860
rect 87344 28858 87368 28860
rect 87424 28858 87448 28860
rect 87504 28858 87528 28860
rect 87584 28858 87590 28860
rect 87344 28806 87346 28858
rect 87526 28806 87528 28858
rect 87282 28804 87288 28806
rect 87344 28804 87368 28806
rect 87424 28804 87448 28806
rect 87504 28804 87528 28806
rect 87584 28804 87590 28806
rect 87282 28795 87590 28804
rect 86352 28588 86404 28594
rect 86352 28530 86404 28536
rect 86364 28361 86392 28530
rect 88192 28452 88244 28458
rect 88192 28394 88244 28400
rect 86350 28352 86406 28361
rect 86350 28287 86406 28296
rect 86546 28316 86854 28325
rect 86546 28314 86552 28316
rect 86608 28314 86632 28316
rect 86688 28314 86712 28316
rect 86768 28314 86792 28316
rect 86848 28314 86854 28316
rect 86608 28262 86610 28314
rect 86790 28262 86792 28314
rect 86546 28260 86552 28262
rect 86608 28260 86632 28262
rect 86688 28260 86712 28262
rect 86768 28260 86792 28262
rect 86848 28260 86854 28262
rect 86546 28251 86854 28260
rect 88204 28225 88232 28394
rect 88190 28216 88246 28225
rect 88190 28151 88246 28160
rect 88928 27908 88980 27914
rect 88928 27850 88980 27856
rect 87282 27772 87590 27781
rect 87282 27770 87288 27772
rect 87344 27770 87368 27772
rect 87424 27770 87448 27772
rect 87504 27770 87528 27772
rect 87584 27770 87590 27772
rect 87344 27718 87346 27770
rect 87526 27718 87528 27770
rect 87282 27716 87288 27718
rect 87344 27716 87368 27718
rect 87424 27716 87448 27718
rect 87504 27716 87528 27718
rect 87584 27716 87590 27718
rect 87282 27707 87590 27716
rect 88940 27545 88968 27850
rect 88926 27536 88982 27545
rect 88926 27471 88982 27480
rect 86546 27228 86854 27237
rect 86546 27226 86552 27228
rect 86608 27226 86632 27228
rect 86688 27226 86712 27228
rect 86768 27226 86792 27228
rect 86848 27226 86854 27228
rect 86608 27174 86610 27226
rect 86790 27174 86792 27226
rect 86546 27172 86552 27174
rect 86608 27172 86632 27174
rect 86688 27172 86712 27174
rect 86768 27172 86792 27174
rect 86848 27172 86854 27174
rect 86546 27163 86854 27172
rect 87282 26684 87590 26693
rect 87282 26682 87288 26684
rect 87344 26682 87368 26684
rect 87424 26682 87448 26684
rect 87504 26682 87528 26684
rect 87584 26682 87590 26684
rect 87344 26630 87346 26682
rect 87526 26630 87528 26682
rect 87282 26628 87288 26630
rect 87344 26628 87368 26630
rect 87424 26628 87448 26630
rect 87504 26628 87528 26630
rect 87584 26628 87590 26630
rect 87282 26619 87590 26628
rect 87732 26446 87784 26452
rect 87732 26388 87784 26394
rect 87744 26321 87772 26388
rect 87730 26312 87786 26321
rect 87730 26247 87786 26256
rect 88192 26276 88244 26282
rect 88192 26218 88244 26224
rect 88204 26185 88232 26218
rect 88190 26176 88246 26185
rect 86546 26140 86854 26149
rect 86546 26138 86552 26140
rect 86608 26138 86632 26140
rect 86688 26138 86712 26140
rect 86768 26138 86792 26140
rect 86848 26138 86854 26140
rect 86608 26086 86610 26138
rect 86790 26086 86792 26138
rect 88190 26111 88246 26120
rect 86546 26084 86552 26086
rect 86608 26084 86632 26086
rect 86688 26084 86712 26086
rect 86768 26084 86792 26086
rect 86848 26084 86854 26086
rect 86546 26075 86854 26084
rect 87282 25596 87590 25605
rect 87282 25594 87288 25596
rect 87344 25594 87368 25596
rect 87424 25594 87448 25596
rect 87504 25594 87528 25596
rect 87584 25594 87590 25596
rect 87344 25542 87346 25594
rect 87526 25542 87528 25594
rect 87282 25540 87288 25542
rect 87344 25540 87368 25542
rect 87424 25540 87448 25542
rect 87504 25540 87528 25542
rect 87584 25540 87590 25542
rect 87282 25531 87590 25540
rect 87732 25358 87784 25364
rect 87732 25300 87784 25306
rect 87744 25233 87772 25300
rect 87730 25224 87786 25233
rect 87730 25159 87786 25168
rect 88560 25188 88612 25194
rect 88560 25130 88612 25136
rect 86546 25052 86854 25061
rect 86546 25050 86552 25052
rect 86608 25050 86632 25052
rect 86688 25050 86712 25052
rect 86768 25050 86792 25052
rect 86848 25050 86854 25052
rect 86608 24998 86610 25050
rect 86790 24998 86792 25050
rect 86546 24996 86552 24998
rect 86608 24996 86632 24998
rect 86688 24996 86712 24998
rect 86768 24996 86792 24998
rect 86848 24996 86854 24998
rect 86546 24987 86854 24996
rect 88572 24825 88600 25130
rect 88558 24816 88614 24825
rect 88558 24751 88614 24760
rect 87282 24508 87590 24517
rect 87282 24506 87288 24508
rect 87344 24506 87368 24508
rect 87424 24506 87448 24508
rect 87504 24506 87528 24508
rect 87584 24506 87590 24508
rect 87344 24454 87346 24506
rect 87526 24454 87528 24506
rect 87282 24452 87288 24454
rect 87344 24452 87368 24454
rect 87424 24452 87448 24454
rect 87504 24452 87528 24454
rect 87584 24452 87590 24454
rect 87282 24443 87590 24452
rect 87732 24270 87784 24276
rect 87732 24212 87784 24218
rect 87744 24145 87772 24212
rect 87730 24136 87786 24145
rect 87730 24071 87786 24080
rect 88282 24136 88338 24145
rect 88282 24071 88284 24080
rect 88336 24071 88338 24080
rect 88284 24042 88336 24048
rect 86546 23964 86854 23973
rect 86546 23962 86552 23964
rect 86608 23962 86632 23964
rect 86688 23962 86712 23964
rect 86768 23962 86792 23964
rect 86848 23962 86854 23964
rect 86608 23910 86610 23962
rect 86790 23910 86792 23962
rect 86546 23908 86552 23910
rect 86608 23908 86632 23910
rect 86688 23908 86712 23910
rect 86768 23908 86792 23910
rect 86848 23908 86854 23910
rect 86546 23899 86854 23908
rect 87282 23420 87590 23429
rect 87282 23418 87288 23420
rect 87344 23418 87368 23420
rect 87424 23418 87448 23420
rect 87504 23418 87528 23420
rect 87584 23418 87590 23420
rect 87344 23366 87346 23418
rect 87526 23366 87528 23418
rect 87282 23364 87288 23366
rect 87344 23364 87368 23366
rect 87424 23364 87448 23366
rect 87504 23364 87528 23366
rect 87584 23364 87590 23366
rect 87282 23355 87590 23364
rect 86352 23148 86404 23154
rect 86352 23090 86404 23096
rect 86364 22921 86392 23090
rect 88284 23012 88336 23018
rect 88284 22954 88336 22960
rect 86350 22912 86406 22921
rect 86350 22847 86406 22856
rect 86546 22876 86854 22885
rect 86546 22874 86552 22876
rect 86608 22874 86632 22876
rect 86688 22874 86712 22876
rect 86768 22874 86792 22876
rect 86848 22874 86854 22876
rect 86608 22822 86610 22874
rect 86790 22822 86792 22874
rect 86546 22820 86552 22822
rect 86608 22820 86632 22822
rect 86688 22820 86712 22822
rect 86768 22820 86792 22822
rect 86848 22820 86854 22822
rect 86546 22811 86854 22820
rect 88296 22785 88324 22954
rect 88282 22776 88338 22785
rect 88282 22711 88338 22720
rect 88560 22468 88612 22474
rect 88560 22410 88612 22416
rect 87282 22332 87590 22341
rect 87282 22330 87288 22332
rect 87344 22330 87368 22332
rect 87424 22330 87448 22332
rect 87504 22330 87528 22332
rect 87584 22330 87590 22332
rect 87344 22278 87346 22330
rect 87526 22278 87528 22330
rect 87282 22276 87288 22278
rect 87344 22276 87368 22278
rect 87424 22276 87448 22278
rect 87504 22276 87528 22278
rect 87584 22276 87590 22278
rect 87282 22267 87590 22276
rect 88572 22105 88600 22410
rect 88558 22096 88614 22105
rect 88558 22031 88614 22040
rect 86546 21788 86854 21797
rect 86546 21786 86552 21788
rect 86608 21786 86632 21788
rect 86688 21786 86712 21788
rect 86768 21786 86792 21788
rect 86848 21786 86854 21788
rect 86608 21734 86610 21786
rect 86790 21734 86792 21786
rect 86546 21732 86552 21734
rect 86608 21732 86632 21734
rect 86688 21732 86712 21734
rect 86768 21732 86792 21734
rect 86848 21732 86854 21734
rect 86546 21723 86854 21732
rect 87282 21244 87590 21253
rect 87282 21242 87288 21244
rect 87344 21242 87368 21244
rect 87424 21242 87448 21244
rect 87504 21242 87528 21244
rect 87584 21242 87590 21244
rect 87344 21190 87346 21242
rect 87526 21190 87528 21242
rect 87282 21188 87288 21190
rect 87344 21188 87368 21190
rect 87424 21188 87448 21190
rect 87504 21188 87528 21190
rect 87584 21188 87590 21190
rect 87282 21179 87590 21188
rect 88560 20972 88612 20978
rect 88560 20914 88612 20920
rect 88572 20745 88600 20914
rect 88558 20736 88614 20745
rect 86546 20700 86854 20709
rect 86546 20698 86552 20700
rect 86608 20698 86632 20700
rect 86688 20698 86712 20700
rect 86768 20698 86792 20700
rect 86848 20698 86854 20700
rect 86608 20646 86610 20698
rect 86790 20646 86792 20698
rect 88558 20671 88614 20680
rect 86546 20644 86552 20646
rect 86608 20644 86632 20646
rect 86688 20644 86712 20646
rect 86768 20644 86792 20646
rect 86848 20644 86854 20646
rect 86546 20635 86854 20644
rect 87282 20156 87590 20165
rect 87282 20154 87288 20156
rect 87344 20154 87368 20156
rect 87424 20154 87448 20156
rect 87504 20154 87528 20156
rect 87584 20154 87590 20156
rect 87344 20102 87346 20154
rect 87526 20102 87528 20154
rect 87282 20100 87288 20102
rect 87344 20100 87368 20102
rect 87424 20100 87448 20102
rect 87504 20100 87528 20102
rect 87584 20100 87590 20102
rect 87282 20091 87590 20100
rect 87732 19918 87784 19924
rect 87732 19860 87784 19866
rect 87744 19793 87772 19860
rect 87730 19784 87786 19793
rect 87730 19719 87786 19728
rect 88560 19748 88612 19754
rect 88560 19690 88612 19696
rect 86546 19612 86854 19621
rect 86546 19610 86552 19612
rect 86608 19610 86632 19612
rect 86688 19610 86712 19612
rect 86768 19610 86792 19612
rect 86848 19610 86854 19612
rect 86608 19558 86610 19610
rect 86790 19558 86792 19610
rect 86546 19556 86552 19558
rect 86608 19556 86632 19558
rect 86688 19556 86712 19558
rect 86768 19556 86792 19558
rect 86848 19556 86854 19558
rect 86546 19547 86854 19556
rect 88572 19385 88600 19690
rect 88558 19376 88614 19385
rect 88558 19311 88614 19320
rect 87282 19068 87590 19077
rect 87282 19066 87288 19068
rect 87344 19066 87368 19068
rect 87424 19066 87448 19068
rect 87504 19066 87528 19068
rect 87584 19066 87590 19068
rect 87344 19014 87346 19066
rect 87526 19014 87528 19066
rect 87282 19012 87288 19014
rect 87344 19012 87368 19014
rect 87424 19012 87448 19014
rect 87504 19012 87528 19014
rect 87584 19012 87590 19014
rect 87282 19003 87590 19012
rect 87732 18830 87784 18836
rect 87732 18772 87784 18778
rect 87744 18705 87772 18772
rect 87730 18696 87786 18705
rect 87730 18631 87786 18640
rect 88282 18696 88338 18705
rect 88282 18631 88284 18640
rect 88336 18631 88338 18640
rect 88284 18602 88336 18608
rect 86546 18524 86854 18533
rect 86546 18522 86552 18524
rect 86608 18522 86632 18524
rect 86688 18522 86712 18524
rect 86768 18522 86792 18524
rect 86848 18522 86854 18524
rect 86608 18470 86610 18522
rect 86790 18470 86792 18522
rect 86546 18468 86552 18470
rect 86608 18468 86632 18470
rect 86688 18468 86712 18470
rect 86768 18468 86792 18470
rect 86848 18468 86854 18470
rect 86546 18459 86854 18468
rect 87282 17980 87590 17989
rect 87282 17978 87288 17980
rect 87344 17978 87368 17980
rect 87424 17978 87448 17980
rect 87504 17978 87528 17980
rect 87584 17978 87590 17980
rect 87344 17926 87346 17978
rect 87526 17926 87528 17978
rect 87282 17924 87288 17926
rect 87344 17924 87368 17926
rect 87424 17924 87448 17926
rect 87504 17924 87528 17926
rect 87584 17924 87590 17926
rect 87282 17915 87590 17924
rect 86352 17708 86404 17714
rect 86352 17650 86404 17656
rect 86364 17481 86392 17650
rect 88192 17572 88244 17578
rect 88192 17514 88244 17520
rect 86350 17472 86406 17481
rect 86350 17407 86406 17416
rect 86546 17436 86854 17445
rect 86546 17434 86552 17436
rect 86608 17434 86632 17436
rect 86688 17434 86712 17436
rect 86768 17434 86792 17436
rect 86848 17434 86854 17436
rect 86608 17382 86610 17434
rect 86790 17382 86792 17434
rect 86546 17380 86552 17382
rect 86608 17380 86632 17382
rect 86688 17380 86712 17382
rect 86768 17380 86792 17382
rect 86848 17380 86854 17382
rect 86546 17371 86854 17380
rect 88204 17345 88232 17514
rect 88190 17336 88246 17345
rect 88190 17271 88246 17280
rect 88008 17130 88060 17136
rect 88008 17072 88060 17078
rect 87282 16892 87590 16901
rect 87282 16890 87288 16892
rect 87344 16890 87368 16892
rect 87424 16890 87448 16892
rect 87504 16890 87528 16892
rect 87584 16890 87590 16892
rect 87344 16838 87346 16890
rect 87526 16838 87528 16890
rect 87282 16836 87288 16838
rect 87344 16836 87368 16838
rect 87424 16836 87448 16838
rect 87504 16836 87528 16838
rect 87584 16836 87590 16838
rect 87282 16827 87590 16836
rect 88020 16529 88048 17072
rect 88560 17028 88612 17034
rect 88560 16970 88612 16976
rect 88572 16665 88600 16970
rect 88558 16656 88614 16665
rect 88558 16591 88614 16600
rect 88006 16520 88062 16529
rect 88006 16455 88062 16464
rect 86546 16348 86854 16357
rect 86546 16346 86552 16348
rect 86608 16346 86632 16348
rect 86688 16346 86712 16348
rect 86768 16346 86792 16348
rect 86848 16346 86854 16348
rect 86608 16294 86610 16346
rect 86790 16294 86792 16346
rect 86546 16292 86552 16294
rect 86608 16292 86632 16294
rect 86688 16292 86712 16294
rect 86768 16292 86792 16294
rect 86848 16292 86854 16294
rect 86546 16283 86854 16292
rect 87282 15804 87590 15813
rect 87282 15802 87288 15804
rect 87344 15802 87368 15804
rect 87424 15802 87448 15804
rect 87504 15802 87528 15804
rect 87584 15802 87590 15804
rect 87344 15750 87346 15802
rect 87526 15750 87528 15802
rect 87282 15748 87288 15750
rect 87344 15748 87368 15750
rect 87424 15748 87448 15750
rect 87504 15748 87528 15750
rect 87584 15748 87590 15750
rect 87282 15739 87590 15748
rect 88560 15464 88612 15470
rect 88560 15406 88612 15412
rect 88572 15305 88600 15406
rect 88558 15296 88614 15305
rect 86546 15260 86854 15269
rect 86546 15258 86552 15260
rect 86608 15258 86632 15260
rect 86688 15258 86712 15260
rect 86768 15258 86792 15260
rect 86848 15258 86854 15260
rect 86608 15206 86610 15258
rect 86790 15206 86792 15258
rect 88558 15231 88614 15240
rect 86546 15204 86552 15206
rect 86608 15204 86632 15206
rect 86688 15204 86712 15206
rect 86768 15204 86792 15206
rect 86848 15204 86854 15206
rect 86546 15195 86854 15204
rect 85616 14988 85668 14994
rect 85616 14930 85668 14936
rect 85628 14314 85656 14930
rect 88008 14852 88060 14858
rect 88008 14794 88060 14800
rect 87282 14716 87590 14725
rect 87282 14714 87288 14716
rect 87344 14714 87368 14716
rect 87424 14714 87448 14716
rect 87504 14714 87528 14716
rect 87584 14714 87590 14716
rect 87344 14662 87346 14714
rect 87526 14662 87528 14714
rect 87282 14660 87288 14662
rect 87344 14660 87368 14662
rect 87424 14660 87448 14662
rect 87504 14660 87528 14662
rect 87584 14660 87590 14662
rect 87282 14651 87590 14660
rect 88020 14625 88048 14794
rect 88006 14616 88062 14625
rect 88006 14551 88062 14560
rect 85616 14308 85668 14314
rect 85616 14250 85668 14256
rect 86546 14172 86854 14181
rect 86546 14170 86552 14172
rect 86608 14170 86632 14172
rect 86688 14170 86712 14172
rect 86768 14170 86792 14172
rect 86848 14170 86854 14172
rect 86608 14118 86610 14170
rect 86790 14118 86792 14170
rect 86546 14116 86552 14118
rect 86608 14116 86632 14118
rect 86688 14116 86712 14118
rect 86768 14116 86792 14118
rect 86848 14116 86854 14118
rect 86546 14107 86854 14116
rect 87282 13628 87590 13637
rect 87282 13626 87288 13628
rect 87344 13626 87368 13628
rect 87424 13626 87448 13628
rect 87504 13626 87528 13628
rect 87584 13626 87590 13628
rect 87344 13574 87346 13626
rect 87526 13574 87528 13626
rect 87282 13572 87288 13574
rect 87344 13572 87368 13574
rect 87424 13572 87448 13574
rect 87504 13572 87528 13574
rect 87584 13572 87590 13574
rect 87282 13563 87590 13572
rect 85524 13492 85576 13498
rect 85524 13434 85576 13440
rect 88192 13390 88244 13396
rect 87916 13356 87968 13362
rect 88192 13332 88244 13338
rect 87916 13298 87968 13304
rect 86546 13084 86854 13093
rect 86546 13082 86552 13084
rect 86608 13082 86632 13084
rect 86688 13082 86712 13084
rect 86768 13082 86792 13084
rect 86848 13082 86854 13084
rect 86608 13030 86610 13082
rect 86790 13030 86792 13082
rect 86546 13028 86552 13030
rect 86608 13028 86632 13030
rect 86688 13028 86712 13030
rect 86768 13028 86792 13030
rect 86848 13028 86854 13030
rect 86546 13019 86854 13028
rect 87928 12954 87956 13298
rect 88204 13265 88232 13332
rect 88190 13256 88246 13265
rect 88190 13191 88246 13200
rect 87916 12948 87968 12954
rect 87916 12890 87968 12896
rect 87180 12744 87232 12750
rect 87180 12686 87232 12692
rect 88560 12744 88612 12750
rect 88560 12686 88612 12692
rect 87192 12410 87220 12686
rect 88572 12585 88600 12686
rect 88558 12576 88614 12585
rect 87282 12540 87590 12549
rect 87282 12538 87288 12540
rect 87344 12538 87368 12540
rect 87424 12538 87448 12540
rect 87504 12538 87528 12540
rect 87584 12538 87590 12540
rect 87344 12486 87346 12538
rect 87526 12486 87528 12538
rect 88558 12511 88614 12520
rect 87282 12484 87288 12486
rect 87344 12484 87368 12486
rect 87424 12484 87448 12486
rect 87504 12484 87528 12486
rect 87584 12484 87590 12486
rect 87282 12475 87590 12484
rect 85340 12404 85392 12410
rect 85340 12346 85392 12352
rect 87180 12404 87232 12410
rect 87180 12346 87232 12352
rect 86546 11996 86854 12005
rect 86546 11994 86552 11996
rect 86608 11994 86632 11996
rect 86688 11994 86712 11996
rect 86768 11994 86792 11996
rect 86848 11994 86854 11996
rect 86608 11942 86610 11994
rect 86790 11942 86792 11994
rect 86546 11940 86552 11942
rect 86608 11940 86632 11942
rect 86688 11940 86712 11942
rect 86768 11940 86792 11942
rect 86848 11940 86854 11942
rect 86546 11931 86854 11940
rect 83684 11792 83736 11798
rect 83684 11734 83736 11740
rect 87282 11452 87590 11461
rect 87282 11450 87288 11452
rect 87344 11450 87368 11452
rect 87424 11450 87448 11452
rect 87504 11450 87528 11452
rect 87584 11450 87590 11452
rect 87344 11398 87346 11450
rect 87526 11398 87528 11450
rect 87282 11396 87288 11398
rect 87344 11396 87368 11398
rect 87424 11396 87448 11398
rect 87504 11396 87528 11398
rect 87584 11396 87590 11398
rect 87282 11387 87590 11396
rect 86546 10908 86854 10917
rect 86546 10906 86552 10908
rect 86608 10906 86632 10908
rect 86688 10906 86712 10908
rect 86768 10906 86792 10908
rect 86848 10906 86854 10908
rect 86608 10854 86610 10906
rect 86790 10854 86792 10906
rect 86546 10852 86552 10854
rect 86608 10852 86632 10854
rect 86688 10852 86712 10854
rect 86768 10852 86792 10854
rect 86848 10852 86854 10854
rect 86546 10843 86854 10852
rect 88376 10576 88428 10582
rect 88374 10536 88376 10545
rect 88428 10536 88430 10545
rect 88374 10471 88430 10480
rect 87282 10364 87590 10373
rect 87282 10362 87288 10364
rect 87344 10362 87368 10364
rect 87424 10362 87448 10364
rect 87504 10362 87528 10364
rect 87584 10362 87590 10364
rect 87344 10310 87346 10362
rect 87526 10310 87528 10362
rect 87282 10308 87288 10310
rect 87344 10308 87368 10310
rect 87424 10308 87448 10310
rect 87504 10308 87528 10310
rect 87584 10308 87590 10310
rect 87282 10299 87590 10308
rect 88560 10092 88612 10098
rect 88560 10034 88612 10040
rect 88572 9865 88600 10034
rect 88558 9856 88614 9865
rect 86546 9820 86854 9829
rect 86546 9818 86552 9820
rect 86608 9818 86632 9820
rect 86688 9818 86712 9820
rect 86768 9818 86792 9820
rect 86848 9818 86854 9820
rect 86608 9766 86610 9818
rect 86790 9766 86792 9818
rect 88558 9791 88614 9800
rect 86546 9764 86552 9766
rect 86608 9764 86632 9766
rect 86688 9764 86712 9766
rect 86768 9764 86792 9766
rect 86848 9764 86854 9766
rect 86546 9755 86854 9764
rect 87282 9276 87590 9285
rect 87282 9274 87288 9276
rect 87344 9274 87368 9276
rect 87424 9274 87448 9276
rect 87504 9274 87528 9276
rect 87584 9274 87590 9276
rect 87344 9222 87346 9274
rect 87526 9222 87528 9274
rect 87282 9220 87288 9222
rect 87344 9220 87368 9222
rect 87424 9220 87448 9222
rect 87504 9220 87528 9222
rect 87584 9220 87590 9222
rect 87282 9211 87590 9220
rect 86546 8732 86854 8741
rect 86546 8730 86552 8732
rect 86608 8730 86632 8732
rect 86688 8730 86712 8732
rect 86768 8730 86792 8732
rect 86848 8730 86854 8732
rect 86608 8678 86610 8730
rect 86790 8678 86792 8730
rect 86546 8676 86552 8678
rect 86608 8676 86632 8678
rect 86688 8676 86712 8678
rect 86768 8676 86792 8678
rect 86848 8676 86854 8678
rect 86546 8667 86854 8676
rect 87282 8188 87590 8197
rect 87282 8186 87288 8188
rect 87344 8186 87368 8188
rect 87424 8186 87448 8188
rect 87504 8186 87528 8188
rect 87584 8186 87590 8188
rect 87344 8134 87346 8186
rect 87526 8134 87528 8186
rect 87282 8132 87288 8134
rect 87344 8132 87368 8134
rect 87424 8132 87448 8134
rect 87504 8132 87528 8134
rect 87584 8132 87590 8134
rect 87282 8123 87590 8132
rect 86546 7644 86854 7653
rect 86546 7642 86552 7644
rect 86608 7642 86632 7644
rect 86688 7642 86712 7644
rect 86768 7642 86792 7644
rect 86848 7642 86854 7644
rect 86608 7590 86610 7642
rect 86790 7590 86792 7642
rect 86546 7588 86552 7590
rect 86608 7588 86632 7590
rect 86688 7588 86712 7590
rect 86768 7588 86792 7590
rect 86848 7588 86854 7590
rect 86546 7579 86854 7588
rect 83592 7236 83644 7242
rect 83592 7178 83644 7184
rect 87282 7100 87590 7109
rect 87282 7098 87288 7100
rect 87344 7098 87368 7100
rect 87424 7098 87448 7100
rect 87504 7098 87528 7100
rect 87584 7098 87590 7100
rect 87344 7046 87346 7098
rect 87526 7046 87528 7098
rect 87282 7044 87288 7046
rect 87344 7044 87368 7046
rect 87424 7044 87448 7046
rect 87504 7044 87528 7046
rect 87584 7044 87590 7046
rect 87282 7035 87590 7044
rect 78900 5332 78952 5338
rect 78900 5274 78952 5280
rect 80280 5332 80332 5338
rect 80280 5274 80332 5280
rect 70068 5264 70120 5270
rect 70068 5206 70120 5212
rect 77796 5264 77848 5270
rect 77796 5206 77848 5212
rect 15236 5162 15288 5168
rect 15236 5104 15288 5110
rect 16064 5162 16116 5168
rect 16064 5104 16116 5110
rect 17168 5162 17220 5168
rect 17168 5104 17220 5110
rect 18272 5162 18324 5168
rect 18272 5104 18324 5110
rect 19652 5162 19704 5168
rect 19652 5104 19704 5110
rect 20480 5162 20532 5168
rect 20480 5104 20532 5110
rect 21584 5162 21636 5168
rect 21584 5104 21636 5110
rect 22964 5162 23016 5168
rect 22964 5104 23016 5110
rect 23792 5162 23844 5168
rect 23792 5104 23844 5110
rect 24896 5162 24948 5168
rect 24896 5104 24948 5110
rect 26092 5162 26144 5168
rect 26092 5104 26144 5110
rect 27380 5162 27432 5168
rect 27380 5104 27432 5110
rect 28208 5162 28260 5168
rect 28208 5104 28260 5110
rect 29312 5162 29364 5168
rect 52404 5162 52456 5168
rect 29312 5104 29364 5110
rect 35752 5128 35804 5134
rect 35752 5070 35804 5076
rect 43480 5128 43532 5134
rect 52404 5104 52456 5110
rect 53692 5162 53744 5168
rect 53692 5104 53744 5110
rect 54888 5162 54940 5168
rect 54888 5104 54940 5110
rect 55716 5162 55768 5168
rect 55716 5104 55768 5110
rect 56820 5162 56872 5168
rect 56820 5104 56872 5110
rect 57924 5162 57976 5168
rect 57924 5104 57976 5110
rect 59028 5162 59080 5168
rect 59028 5104 59080 5110
rect 60132 5162 60184 5168
rect 60132 5104 60184 5110
rect 61420 5162 61472 5168
rect 61420 5104 61472 5110
rect 62340 5162 62392 5168
rect 62340 5104 62392 5110
rect 63444 5162 63496 5168
rect 63444 5104 63496 5110
rect 64548 5162 64600 5168
rect 64548 5104 64600 5110
rect 65652 5162 65704 5168
rect 65652 5104 65704 5110
rect 66756 5162 66808 5168
rect 69884 5162 69936 5168
rect 66756 5104 66808 5110
rect 69240 5128 69292 5134
rect 43480 5070 43532 5076
rect 77612 5162 77664 5168
rect 69884 5104 69936 5110
rect 74392 5128 74444 5134
rect 69240 5070 69292 5076
rect 15144 5060 15196 5066
rect 15144 5002 15196 5008
rect 15788 5060 15840 5066
rect 15788 5002 15840 5008
rect 17076 5060 17128 5066
rect 17076 5002 17128 5008
rect 18272 5060 18324 5066
rect 18272 5002 18324 5008
rect 19652 5060 19704 5066
rect 19652 5002 19704 5008
rect 20296 5060 20348 5066
rect 20296 5002 20348 5008
rect 21584 5060 21636 5066
rect 21584 5002 21636 5008
rect 22872 5060 22924 5066
rect 22872 5002 22924 5008
rect 23516 5060 23568 5066
rect 23516 5002 23568 5008
rect 24804 5060 24856 5066
rect 24804 5002 24856 5008
rect 26092 5060 26144 5066
rect 26092 5002 26144 5008
rect 27380 5060 27432 5066
rect 27380 5002 27432 5008
rect 28024 5060 28076 5066
rect 28024 5002 28076 5008
rect 29312 5060 29364 5066
rect 29312 5002 29364 5008
rect 30600 5060 30652 5066
rect 30600 5002 30652 5008
rect 31244 5060 31296 5066
rect 31244 5002 31296 5008
rect 32532 5060 32584 5066
rect 32532 5002 32584 5008
rect 33820 5060 33872 5066
rect 33820 5002 33872 5008
rect 35108 5060 35160 5066
rect 35108 5002 35160 5008
rect 15156 2400 15184 5002
rect 15800 2400 15828 5002
rect 17088 2400 17116 5002
rect 18284 3314 18312 5002
rect 18382 4924 18690 4933
rect 18382 4922 18388 4924
rect 18444 4922 18468 4924
rect 18524 4922 18548 4924
rect 18604 4922 18628 4924
rect 18684 4922 18690 4924
rect 18444 4870 18446 4922
rect 18626 4870 18628 4922
rect 18382 4868 18388 4870
rect 18444 4868 18468 4870
rect 18524 4868 18548 4870
rect 18604 4868 18628 4870
rect 18684 4868 18690 4870
rect 18382 4859 18690 4868
rect 18284 3286 18404 3314
rect 18376 2400 18404 3286
rect 19664 2400 19692 5002
rect 20308 2400 20336 5002
rect 21596 2400 21624 5002
rect 22884 2400 22912 5002
rect 23528 2400 23556 5002
rect 24816 2400 24844 5002
rect 26104 2400 26132 5002
rect 27392 2400 27420 5002
rect 28036 2400 28064 5002
rect 29324 2400 29352 5002
rect 30612 2400 30640 5002
rect 31256 2400 31284 5002
rect 32544 2400 32572 5002
rect 33832 2400 33860 5002
rect 35120 2400 35148 5002
rect 35764 2400 35792 5070
rect 37132 5060 37184 5066
rect 37132 5002 37184 5008
rect 38328 5060 38380 5066
rect 38328 5002 38380 5008
rect 38972 5060 39024 5066
rect 38972 5002 39024 5008
rect 40260 5060 40312 5066
rect 40260 5002 40312 5008
rect 41548 5060 41600 5066
rect 41548 5002 41600 5008
rect 42836 5060 42888 5066
rect 42836 5002 42888 5008
rect 36782 4924 37090 4933
rect 36782 4922 36788 4924
rect 36844 4922 36868 4924
rect 36924 4922 36948 4924
rect 37004 4922 37028 4924
rect 37084 4922 37090 4924
rect 36844 4870 36846 4922
rect 37026 4870 37028 4922
rect 36782 4868 36788 4870
rect 36844 4868 36868 4870
rect 36924 4868 36948 4870
rect 37004 4868 37028 4870
rect 37084 4868 37090 4870
rect 36782 4859 37090 4868
rect 37144 4810 37172 5002
rect 37052 4782 37172 4810
rect 37052 2400 37080 4782
rect 38340 2400 38368 5002
rect 38984 2400 39012 5002
rect 40272 2400 40300 5002
rect 41560 2400 41588 5002
rect 42848 2400 42876 5002
rect 43492 2400 43520 5070
rect 44768 5060 44820 5066
rect 44768 5002 44820 5008
rect 52496 5060 52548 5066
rect 52496 5002 52548 5008
rect 53784 5060 53836 5066
rect 53784 5002 53836 5008
rect 54428 5060 54480 5066
rect 54428 5002 54480 5008
rect 55716 5060 55768 5066
rect 55716 5002 55768 5008
rect 57004 5060 57056 5066
rect 57004 5002 57056 5008
rect 57648 5060 57700 5066
rect 57648 5002 57700 5008
rect 58936 5060 58988 5066
rect 58936 5002 58988 5008
rect 60224 5060 60276 5066
rect 60224 5002 60276 5008
rect 61512 5060 61564 5066
rect 61512 5002 61564 5008
rect 62156 5060 62208 5066
rect 62156 5002 62208 5008
rect 63444 5060 63496 5066
rect 63444 5002 63496 5008
rect 64732 5060 64784 5066
rect 64732 5002 64784 5008
rect 65376 5060 65428 5066
rect 65376 5002 65428 5008
rect 66664 5060 66716 5066
rect 66664 5002 66716 5008
rect 67952 5060 68004 5066
rect 67952 5002 68004 5008
rect 44780 2400 44808 5002
rect 52508 2400 52536 5002
rect 53796 2400 53824 5002
rect 54440 2400 54468 5002
rect 55182 4924 55490 4933
rect 55182 4922 55188 4924
rect 55244 4922 55268 4924
rect 55324 4922 55348 4924
rect 55404 4922 55428 4924
rect 55484 4922 55490 4924
rect 55244 4870 55246 4922
rect 55426 4870 55428 4922
rect 55182 4868 55188 4870
rect 55244 4868 55268 4870
rect 55324 4868 55348 4870
rect 55404 4868 55428 4870
rect 55484 4868 55490 4870
rect 55182 4859 55490 4868
rect 55728 2400 55756 5002
rect 57016 2400 57044 5002
rect 57660 2400 57688 5002
rect 58948 2400 58976 5002
rect 60236 2400 60264 5002
rect 61524 2400 61552 5002
rect 62168 2400 62196 5002
rect 63456 2400 63484 5002
rect 64744 2400 64772 5002
rect 65388 2400 65416 5002
rect 66676 2400 66704 5002
rect 67964 2400 67992 5002
rect 69252 2400 69280 5070
rect 69896 2400 69924 5104
rect 74392 5070 74444 5076
rect 76968 5128 77020 5134
rect 77612 5104 77664 5110
rect 76968 5070 77020 5076
rect 71172 5060 71224 5066
rect 71172 5002 71224 5008
rect 72460 5060 72512 5066
rect 72460 5002 72512 5008
rect 73104 5060 73156 5066
rect 73104 5002 73156 5008
rect 71184 2400 71212 5002
rect 72472 2400 72500 5002
rect 73116 2400 73144 5002
rect 73582 4924 73890 4933
rect 73582 4922 73588 4924
rect 73644 4922 73668 4924
rect 73724 4922 73748 4924
rect 73804 4922 73828 4924
rect 73884 4922 73890 4924
rect 73644 4870 73646 4922
rect 73826 4870 73828 4922
rect 73582 4868 73588 4870
rect 73644 4868 73668 4870
rect 73724 4868 73748 4870
rect 73804 4868 73828 4870
rect 73884 4868 73890 4870
rect 73582 4859 73890 4868
rect 74404 2400 74432 5070
rect 75680 5060 75732 5066
rect 75680 5002 75732 5008
rect 75692 2400 75720 5002
rect 76980 2400 77008 5070
rect 77624 2400 77652 5104
rect 78900 5060 78952 5066
rect 78900 5002 78952 5008
rect 80188 5060 80240 5066
rect 80188 5002 80240 5008
rect 78912 2400 78940 5002
rect 80200 2400 80228 5002
rect 1618 1600 1674 2400
rect 2262 1600 2318 2400
rect 2906 1600 2962 2400
rect 3550 1600 3606 2400
rect 4194 1600 4250 2400
rect 4838 1600 4894 2400
rect 5482 1600 5538 2400
rect 6126 1600 6182 2400
rect 6770 1600 6826 2400
rect 7414 1600 7470 2400
rect 8058 1600 8114 2400
rect 8702 1600 8758 2400
rect 9346 1600 9402 2400
rect 9990 1600 10046 2400
rect 10634 1600 10690 2400
rect 11278 1600 11334 2400
rect 15142 1600 15198 2400
rect 15786 1600 15842 2400
rect 17074 1600 17130 2400
rect 18362 1600 18418 2400
rect 19650 1600 19706 2400
rect 20294 1600 20350 2400
rect 21582 1600 21638 2400
rect 22870 1600 22926 2400
rect 23514 1600 23570 2400
rect 24802 1600 24858 2400
rect 26090 1600 26146 2400
rect 27378 1600 27434 2400
rect 28022 1600 28078 2400
rect 29310 1600 29366 2400
rect 30598 1600 30654 2400
rect 31242 1600 31298 2400
rect 32530 1600 32586 2400
rect 33818 1600 33874 2400
rect 35106 1600 35162 2400
rect 35750 1600 35806 2400
rect 37038 1600 37094 2400
rect 38326 1600 38382 2400
rect 38970 1600 39026 2400
rect 40258 1600 40314 2400
rect 41546 1600 41602 2400
rect 42834 1600 42890 2400
rect 43478 1600 43534 2400
rect 44766 1600 44822 2400
rect 52494 1600 52550 2400
rect 53782 1600 53838 2400
rect 54426 1600 54482 2400
rect 55714 1600 55770 2400
rect 57002 1600 57058 2400
rect 57646 1600 57702 2400
rect 58934 1600 58990 2400
rect 60222 1600 60278 2400
rect 61510 1600 61566 2400
rect 62154 1600 62210 2400
rect 63442 1600 63498 2400
rect 64730 1600 64786 2400
rect 65374 1600 65430 2400
rect 66662 1600 66718 2400
rect 67950 1600 68006 2400
rect 69238 1600 69294 2400
rect 69882 1600 69938 2400
rect 71170 1600 71226 2400
rect 72458 1600 72514 2400
rect 73102 1600 73158 2400
rect 74390 1600 74446 2400
rect 75678 1600 75734 2400
rect 76966 1600 77022 2400
rect 77610 1600 77666 2400
rect 78898 1600 78954 2400
rect 80186 1600 80242 2400
<< via2 >>
rect 18388 87610 18444 87612
rect 18468 87610 18524 87612
rect 18548 87610 18604 87612
rect 18628 87610 18684 87612
rect 18388 87558 18434 87610
rect 18434 87558 18444 87610
rect 18468 87558 18498 87610
rect 18498 87558 18510 87610
rect 18510 87558 18524 87610
rect 18548 87558 18562 87610
rect 18562 87558 18574 87610
rect 18574 87558 18604 87610
rect 18628 87558 18638 87610
rect 18638 87558 18684 87610
rect 18388 87556 18444 87558
rect 18468 87556 18524 87558
rect 18548 87556 18604 87558
rect 18628 87556 18684 87558
rect 36788 87610 36844 87612
rect 36868 87610 36924 87612
rect 36948 87610 37004 87612
rect 37028 87610 37084 87612
rect 36788 87558 36834 87610
rect 36834 87558 36844 87610
rect 36868 87558 36898 87610
rect 36898 87558 36910 87610
rect 36910 87558 36924 87610
rect 36948 87558 36962 87610
rect 36962 87558 36974 87610
rect 36974 87558 37004 87610
rect 37028 87558 37038 87610
rect 37038 87558 37084 87610
rect 36788 87556 36844 87558
rect 36868 87556 36924 87558
rect 36948 87556 37004 87558
rect 37028 87556 37084 87558
rect 10726 87374 10782 87376
rect 10726 87322 10728 87374
rect 10728 87322 10780 87374
rect 10780 87322 10782 87374
rect 10726 87320 10782 87322
rect 5960 84890 6016 84892
rect 6040 84890 6096 84892
rect 6120 84890 6176 84892
rect 6200 84890 6256 84892
rect 5960 84838 6006 84890
rect 6006 84838 6016 84890
rect 6040 84838 6070 84890
rect 6070 84838 6082 84890
rect 6082 84838 6096 84890
rect 6120 84838 6134 84890
rect 6134 84838 6146 84890
rect 6146 84838 6176 84890
rect 6200 84838 6210 84890
rect 6210 84838 6256 84890
rect 5960 84836 6016 84838
rect 6040 84836 6096 84838
rect 6120 84836 6176 84838
rect 6200 84836 6256 84838
rect 6696 84346 6752 84348
rect 6776 84346 6832 84348
rect 6856 84346 6912 84348
rect 6936 84346 6992 84348
rect 6696 84294 6742 84346
rect 6742 84294 6752 84346
rect 6776 84294 6806 84346
rect 6806 84294 6818 84346
rect 6818 84294 6832 84346
rect 6856 84294 6870 84346
rect 6870 84294 6882 84346
rect 6882 84294 6912 84346
rect 6936 84294 6946 84346
rect 6946 84294 6992 84346
rect 6696 84292 6752 84294
rect 6776 84292 6832 84294
rect 6856 84292 6912 84294
rect 6936 84292 6992 84294
rect 5960 83802 6016 83804
rect 6040 83802 6096 83804
rect 6120 83802 6176 83804
rect 6200 83802 6256 83804
rect 5960 83750 6006 83802
rect 6006 83750 6016 83802
rect 6040 83750 6070 83802
rect 6070 83750 6082 83802
rect 6082 83750 6096 83802
rect 6120 83750 6134 83802
rect 6134 83750 6146 83802
rect 6146 83750 6176 83802
rect 6200 83750 6210 83802
rect 6210 83750 6256 83802
rect 5960 83748 6016 83750
rect 6040 83748 6096 83750
rect 6120 83748 6176 83750
rect 6200 83748 6256 83750
rect 6696 83258 6752 83260
rect 6776 83258 6832 83260
rect 6856 83258 6912 83260
rect 6936 83258 6992 83260
rect 6696 83206 6742 83258
rect 6742 83206 6752 83258
rect 6776 83206 6806 83258
rect 6806 83206 6818 83258
rect 6818 83206 6832 83258
rect 6856 83206 6870 83258
rect 6870 83206 6882 83258
rect 6882 83206 6912 83258
rect 6936 83206 6946 83258
rect 6946 83206 6992 83258
rect 6696 83204 6752 83206
rect 6776 83204 6832 83206
rect 6856 83204 6912 83206
rect 6936 83204 6992 83206
rect 5960 82714 6016 82716
rect 6040 82714 6096 82716
rect 6120 82714 6176 82716
rect 6200 82714 6256 82716
rect 5960 82662 6006 82714
rect 6006 82662 6016 82714
rect 6040 82662 6070 82714
rect 6070 82662 6082 82714
rect 6082 82662 6096 82714
rect 6120 82662 6134 82714
rect 6134 82662 6146 82714
rect 6146 82662 6176 82714
rect 6200 82662 6210 82714
rect 6210 82662 6256 82714
rect 5960 82660 6016 82662
rect 6040 82660 6096 82662
rect 6120 82660 6176 82662
rect 6200 82660 6256 82662
rect 6696 82170 6752 82172
rect 6776 82170 6832 82172
rect 6856 82170 6912 82172
rect 6936 82170 6992 82172
rect 6696 82118 6742 82170
rect 6742 82118 6752 82170
rect 6776 82118 6806 82170
rect 6806 82118 6818 82170
rect 6818 82118 6832 82170
rect 6856 82118 6870 82170
rect 6870 82118 6882 82170
rect 6882 82118 6912 82170
rect 6936 82118 6946 82170
rect 6946 82118 6992 82170
rect 6696 82116 6752 82118
rect 6776 82116 6832 82118
rect 6856 82116 6912 82118
rect 6936 82116 6992 82118
rect 5960 81626 6016 81628
rect 6040 81626 6096 81628
rect 6120 81626 6176 81628
rect 6200 81626 6256 81628
rect 5960 81574 6006 81626
rect 6006 81574 6016 81626
rect 6040 81574 6070 81626
rect 6070 81574 6082 81626
rect 6082 81574 6096 81626
rect 6120 81574 6134 81626
rect 6134 81574 6146 81626
rect 6146 81574 6176 81626
rect 6200 81574 6210 81626
rect 6210 81574 6256 81626
rect 5960 81572 6016 81574
rect 6040 81572 6096 81574
rect 6120 81572 6176 81574
rect 6200 81572 6256 81574
rect 6696 81082 6752 81084
rect 6776 81082 6832 81084
rect 6856 81082 6912 81084
rect 6936 81082 6992 81084
rect 6696 81030 6742 81082
rect 6742 81030 6752 81082
rect 6776 81030 6806 81082
rect 6806 81030 6818 81082
rect 6818 81030 6832 81082
rect 6856 81030 6870 81082
rect 6870 81030 6882 81082
rect 6882 81030 6912 81082
rect 6936 81030 6946 81082
rect 6946 81030 6992 81082
rect 6696 81028 6752 81030
rect 6776 81028 6832 81030
rect 6856 81028 6912 81030
rect 6936 81028 6992 81030
rect 5960 80538 6016 80540
rect 6040 80538 6096 80540
rect 6120 80538 6176 80540
rect 6200 80538 6256 80540
rect 5960 80486 6006 80538
rect 6006 80486 6016 80538
rect 6040 80486 6070 80538
rect 6070 80486 6082 80538
rect 6082 80486 6096 80538
rect 6120 80486 6134 80538
rect 6134 80486 6146 80538
rect 6146 80486 6176 80538
rect 6200 80486 6210 80538
rect 6210 80486 6256 80538
rect 5960 80484 6016 80486
rect 6040 80484 6096 80486
rect 6120 80484 6176 80486
rect 6200 80484 6256 80486
rect 7138 80148 7140 80168
rect 7140 80148 7192 80168
rect 7192 80148 7194 80168
rect 7138 80112 7194 80148
rect 6696 79994 6752 79996
rect 6776 79994 6832 79996
rect 6856 79994 6912 79996
rect 6936 79994 6992 79996
rect 6696 79942 6742 79994
rect 6742 79942 6752 79994
rect 6776 79942 6806 79994
rect 6806 79942 6818 79994
rect 6818 79942 6832 79994
rect 6856 79942 6870 79994
rect 6870 79942 6882 79994
rect 6882 79942 6912 79994
rect 6936 79942 6946 79994
rect 6946 79942 6992 79994
rect 6696 79940 6752 79942
rect 6776 79940 6832 79942
rect 6856 79940 6912 79942
rect 6936 79940 6992 79942
rect 2906 79840 2962 79896
rect 5960 79450 6016 79452
rect 6040 79450 6096 79452
rect 6120 79450 6176 79452
rect 6200 79450 6256 79452
rect 5960 79398 6006 79450
rect 6006 79398 6016 79450
rect 6040 79398 6070 79450
rect 6070 79398 6082 79450
rect 6082 79398 6096 79450
rect 6120 79398 6134 79450
rect 6134 79398 6146 79450
rect 6146 79398 6176 79450
rect 6200 79398 6210 79450
rect 6210 79398 6256 79450
rect 5960 79396 6016 79398
rect 6040 79396 6096 79398
rect 6120 79396 6176 79398
rect 6200 79396 6256 79398
rect 6696 78906 6752 78908
rect 6776 78906 6832 78908
rect 6856 78906 6912 78908
rect 6936 78906 6992 78908
rect 6696 78854 6742 78906
rect 6742 78854 6752 78906
rect 6776 78854 6806 78906
rect 6806 78854 6818 78906
rect 6818 78854 6832 78906
rect 6856 78854 6870 78906
rect 6870 78854 6882 78906
rect 6882 78854 6912 78906
rect 6936 78854 6946 78906
rect 6946 78854 6992 78906
rect 6696 78852 6752 78854
rect 6776 78852 6832 78854
rect 6856 78852 6912 78854
rect 6936 78852 6992 78854
rect 7138 78752 7194 78808
rect 2906 78500 2962 78536
rect 2906 78480 2908 78500
rect 2908 78480 2960 78500
rect 2960 78480 2962 78500
rect 5960 78362 6016 78364
rect 6040 78362 6096 78364
rect 6120 78362 6176 78364
rect 6200 78362 6256 78364
rect 5960 78310 6006 78362
rect 6006 78310 6016 78362
rect 6040 78310 6070 78362
rect 6070 78310 6082 78362
rect 6082 78310 6096 78362
rect 6120 78310 6134 78362
rect 6134 78310 6146 78362
rect 6146 78310 6176 78362
rect 6200 78310 6210 78362
rect 6210 78310 6256 78362
rect 5960 78308 6016 78310
rect 6040 78308 6096 78310
rect 6120 78308 6176 78310
rect 6200 78308 6256 78310
rect 7138 77972 7140 77992
rect 7140 77972 7192 77992
rect 7192 77972 7194 77992
rect 7138 77936 7194 77972
rect 2906 77800 2962 77856
rect 6696 77818 6752 77820
rect 6776 77818 6832 77820
rect 6856 77818 6912 77820
rect 6936 77818 6992 77820
rect 6696 77766 6742 77818
rect 6742 77766 6752 77818
rect 6776 77766 6806 77818
rect 6806 77766 6818 77818
rect 6818 77766 6832 77818
rect 6856 77766 6870 77818
rect 6870 77766 6882 77818
rect 6882 77766 6912 77818
rect 6936 77766 6946 77818
rect 6946 77766 6992 77818
rect 6696 77764 6752 77766
rect 6776 77764 6832 77766
rect 6856 77764 6912 77766
rect 6936 77764 6992 77766
rect 5960 77274 6016 77276
rect 6040 77274 6096 77276
rect 6120 77274 6176 77276
rect 6200 77274 6256 77276
rect 5960 77222 6006 77274
rect 6006 77222 6016 77274
rect 6040 77222 6070 77274
rect 6070 77222 6082 77274
rect 6082 77222 6096 77274
rect 6120 77222 6134 77274
rect 6134 77222 6146 77274
rect 6146 77222 6176 77274
rect 6200 77222 6210 77274
rect 6210 77222 6256 77274
rect 5960 77220 6016 77222
rect 6040 77220 6096 77222
rect 6120 77220 6176 77222
rect 6200 77220 6256 77222
rect 7138 76884 7140 76904
rect 7140 76884 7192 76904
rect 7192 76884 7194 76904
rect 7138 76848 7194 76884
rect 6696 76730 6752 76732
rect 6776 76730 6832 76732
rect 6856 76730 6912 76732
rect 6936 76730 6992 76732
rect 6696 76678 6742 76730
rect 6742 76678 6752 76730
rect 6776 76678 6806 76730
rect 6806 76678 6818 76730
rect 6818 76678 6832 76730
rect 6856 76678 6870 76730
rect 6870 76678 6882 76730
rect 6882 76678 6912 76730
rect 6936 76678 6946 76730
rect 6946 76678 6992 76730
rect 6696 76676 6752 76678
rect 6776 76676 6832 76678
rect 6856 76676 6912 76678
rect 6936 76676 6992 76678
rect 2722 76440 2778 76496
rect 5960 76186 6016 76188
rect 6040 76186 6096 76188
rect 6120 76186 6176 76188
rect 6200 76186 6256 76188
rect 5960 76134 6006 76186
rect 6006 76134 6016 76186
rect 6040 76134 6070 76186
rect 6070 76134 6082 76186
rect 6082 76134 6096 76186
rect 6120 76134 6134 76186
rect 6134 76134 6146 76186
rect 6146 76134 6176 76186
rect 6200 76134 6210 76186
rect 6210 76134 6256 76186
rect 5960 76132 6016 76134
rect 6040 76132 6096 76134
rect 6120 76132 6176 76134
rect 6200 76132 6256 76134
rect 2906 75780 2962 75816
rect 2906 75760 2908 75780
rect 2908 75760 2960 75780
rect 2960 75760 2962 75780
rect 7138 75796 7140 75816
rect 7140 75796 7192 75816
rect 7192 75796 7194 75816
rect 7138 75760 7194 75796
rect 6696 75642 6752 75644
rect 6776 75642 6832 75644
rect 6856 75642 6912 75644
rect 6936 75642 6992 75644
rect 6696 75590 6742 75642
rect 6742 75590 6752 75642
rect 6776 75590 6806 75642
rect 6806 75590 6818 75642
rect 6818 75590 6832 75642
rect 6856 75590 6870 75642
rect 6870 75590 6882 75642
rect 6882 75590 6912 75642
rect 6936 75590 6946 75642
rect 6946 75590 6992 75642
rect 6696 75588 6752 75590
rect 6776 75588 6832 75590
rect 6856 75588 6912 75590
rect 6936 75588 6992 75590
rect 5960 75098 6016 75100
rect 6040 75098 6096 75100
rect 6120 75098 6176 75100
rect 6200 75098 6256 75100
rect 5960 75046 6006 75098
rect 6006 75046 6016 75098
rect 6040 75046 6070 75098
rect 6070 75046 6082 75098
rect 6082 75046 6096 75098
rect 6120 75046 6134 75098
rect 6134 75046 6146 75098
rect 6146 75046 6176 75098
rect 6200 75046 6210 75098
rect 6210 75046 6256 75098
rect 5960 75044 6016 75046
rect 6040 75044 6096 75046
rect 6120 75044 6176 75046
rect 6200 75044 6256 75046
rect 5666 74536 5722 74592
rect 6696 74554 6752 74556
rect 6776 74554 6832 74556
rect 6856 74554 6912 74556
rect 6936 74554 6992 74556
rect 6696 74502 6742 74554
rect 6742 74502 6752 74554
rect 6776 74502 6806 74554
rect 6806 74502 6818 74554
rect 6818 74502 6832 74554
rect 6856 74502 6870 74554
rect 6870 74502 6882 74554
rect 6882 74502 6912 74554
rect 6936 74502 6946 74554
rect 6946 74502 6992 74554
rect 6696 74500 6752 74502
rect 6776 74500 6832 74502
rect 6856 74500 6912 74502
rect 6936 74500 6992 74502
rect 4378 74400 4434 74456
rect 5960 74010 6016 74012
rect 6040 74010 6096 74012
rect 6120 74010 6176 74012
rect 6200 74010 6256 74012
rect 5960 73958 6006 74010
rect 6006 73958 6016 74010
rect 6040 73958 6070 74010
rect 6070 73958 6082 74010
rect 6082 73958 6096 74010
rect 6120 73958 6134 74010
rect 6134 73958 6146 74010
rect 6146 73958 6176 74010
rect 6200 73958 6210 74010
rect 6210 73958 6256 74010
rect 5960 73956 6016 73958
rect 6040 73956 6096 73958
rect 6120 73956 6176 73958
rect 6200 73956 6256 73958
rect 6696 73466 6752 73468
rect 6776 73466 6832 73468
rect 6856 73466 6912 73468
rect 6936 73466 6992 73468
rect 6696 73414 6742 73466
rect 6742 73414 6752 73466
rect 6776 73414 6806 73466
rect 6806 73414 6818 73466
rect 6818 73414 6832 73466
rect 6856 73414 6870 73466
rect 6870 73414 6882 73466
rect 6882 73414 6912 73466
rect 6936 73414 6946 73466
rect 6946 73414 6992 73466
rect 6696 73412 6752 73414
rect 6776 73412 6832 73414
rect 6856 73412 6912 73414
rect 6936 73412 6992 73414
rect 7138 73312 7194 73368
rect 2906 73060 2962 73096
rect 2906 73040 2908 73060
rect 2908 73040 2960 73060
rect 2960 73040 2962 73060
rect 5960 72922 6016 72924
rect 6040 72922 6096 72924
rect 6120 72922 6176 72924
rect 6200 72922 6256 72924
rect 5960 72870 6006 72922
rect 6006 72870 6016 72922
rect 6040 72870 6070 72922
rect 6070 72870 6082 72922
rect 6082 72870 6096 72922
rect 6120 72870 6134 72922
rect 6134 72870 6146 72922
rect 6146 72870 6176 72922
rect 6200 72870 6210 72922
rect 6210 72870 6256 72922
rect 5960 72868 6016 72870
rect 6040 72868 6096 72870
rect 6120 72868 6176 72870
rect 6200 72868 6256 72870
rect 7138 72532 7140 72552
rect 7140 72532 7192 72552
rect 7192 72532 7194 72552
rect 7138 72496 7194 72532
rect 2906 72360 2962 72416
rect 6696 72378 6752 72380
rect 6776 72378 6832 72380
rect 6856 72378 6912 72380
rect 6936 72378 6992 72380
rect 6696 72326 6742 72378
rect 6742 72326 6752 72378
rect 6776 72326 6806 72378
rect 6806 72326 6818 72378
rect 6818 72326 6832 72378
rect 6856 72326 6870 72378
rect 6870 72326 6882 72378
rect 6882 72326 6912 72378
rect 6936 72326 6946 72378
rect 6946 72326 6992 72378
rect 6696 72324 6752 72326
rect 6776 72324 6832 72326
rect 6856 72324 6912 72326
rect 6936 72324 6992 72326
rect 5960 71834 6016 71836
rect 6040 71834 6096 71836
rect 6120 71834 6176 71836
rect 6200 71834 6256 71836
rect 5960 71782 6006 71834
rect 6006 71782 6016 71834
rect 6040 71782 6070 71834
rect 6070 71782 6082 71834
rect 6082 71782 6096 71834
rect 6120 71782 6134 71834
rect 6134 71782 6146 71834
rect 6146 71782 6176 71834
rect 6200 71782 6210 71834
rect 6210 71782 6256 71834
rect 5960 71780 6016 71782
rect 6040 71780 6096 71782
rect 6120 71780 6176 71782
rect 6200 71780 6256 71782
rect 7138 71444 7140 71464
rect 7140 71444 7192 71464
rect 7192 71444 7194 71464
rect 7138 71408 7194 71444
rect 6696 71290 6752 71292
rect 6776 71290 6832 71292
rect 6856 71290 6912 71292
rect 6936 71290 6992 71292
rect 6696 71238 6742 71290
rect 6742 71238 6752 71290
rect 6776 71238 6806 71290
rect 6806 71238 6818 71290
rect 6818 71238 6832 71290
rect 6856 71238 6870 71290
rect 6870 71238 6882 71290
rect 6882 71238 6912 71290
rect 6936 71238 6946 71290
rect 6946 71238 6992 71290
rect 6696 71236 6752 71238
rect 6776 71236 6832 71238
rect 6856 71236 6912 71238
rect 6936 71236 6992 71238
rect 2722 71000 2778 71056
rect 5960 70746 6016 70748
rect 6040 70746 6096 70748
rect 6120 70746 6176 70748
rect 6200 70746 6256 70748
rect 5960 70694 6006 70746
rect 6006 70694 6016 70746
rect 6040 70694 6070 70746
rect 6070 70694 6082 70746
rect 6082 70694 6096 70746
rect 6120 70694 6134 70746
rect 6134 70694 6146 70746
rect 6146 70694 6176 70746
rect 6200 70694 6210 70746
rect 6210 70694 6256 70746
rect 5960 70692 6016 70694
rect 6040 70692 6096 70694
rect 6120 70692 6176 70694
rect 6200 70692 6256 70694
rect 2906 70340 2962 70376
rect 2906 70320 2908 70340
rect 2908 70320 2960 70340
rect 2960 70320 2962 70340
rect 7138 70356 7140 70376
rect 7140 70356 7192 70376
rect 7192 70356 7194 70376
rect 7138 70320 7194 70356
rect 6696 70202 6752 70204
rect 6776 70202 6832 70204
rect 6856 70202 6912 70204
rect 6936 70202 6992 70204
rect 6696 70150 6742 70202
rect 6742 70150 6752 70202
rect 6776 70150 6806 70202
rect 6806 70150 6818 70202
rect 6818 70150 6832 70202
rect 6856 70150 6870 70202
rect 6870 70150 6882 70202
rect 6882 70150 6912 70202
rect 6936 70150 6946 70202
rect 6946 70150 6992 70202
rect 6696 70148 6752 70150
rect 6776 70148 6832 70150
rect 6856 70148 6912 70150
rect 6936 70148 6992 70150
rect 5960 69658 6016 69660
rect 6040 69658 6096 69660
rect 6120 69658 6176 69660
rect 6200 69658 6256 69660
rect 5960 69606 6006 69658
rect 6006 69606 6016 69658
rect 6040 69606 6070 69658
rect 6070 69606 6082 69658
rect 6082 69606 6096 69658
rect 6120 69606 6134 69658
rect 6134 69606 6146 69658
rect 6146 69606 6176 69658
rect 6200 69606 6210 69658
rect 6210 69606 6256 69658
rect 5960 69604 6016 69606
rect 6040 69604 6096 69606
rect 6120 69604 6176 69606
rect 6200 69604 6256 69606
rect 4378 68960 4434 69016
rect 6696 69114 6752 69116
rect 6776 69114 6832 69116
rect 6856 69114 6912 69116
rect 6936 69114 6992 69116
rect 6696 69062 6742 69114
rect 6742 69062 6752 69114
rect 6776 69062 6806 69114
rect 6806 69062 6818 69114
rect 6818 69062 6832 69114
rect 6856 69062 6870 69114
rect 6870 69062 6882 69114
rect 6882 69062 6912 69114
rect 6936 69062 6946 69114
rect 6946 69062 6992 69114
rect 6696 69060 6752 69062
rect 6776 69060 6832 69062
rect 6856 69060 6912 69062
rect 6936 69060 6992 69062
rect 5666 68824 5722 68880
rect 5960 68570 6016 68572
rect 6040 68570 6096 68572
rect 6120 68570 6176 68572
rect 6200 68570 6256 68572
rect 5960 68518 6006 68570
rect 6006 68518 6016 68570
rect 6040 68518 6070 68570
rect 6070 68518 6082 68570
rect 6082 68518 6096 68570
rect 6120 68518 6134 68570
rect 6134 68518 6146 68570
rect 6146 68518 6176 68570
rect 6200 68518 6210 68570
rect 6210 68518 6256 68570
rect 5960 68516 6016 68518
rect 6040 68516 6096 68518
rect 6120 68516 6176 68518
rect 6200 68516 6256 68518
rect 5666 68144 5722 68200
rect 6696 68026 6752 68028
rect 6776 68026 6832 68028
rect 6856 68026 6912 68028
rect 6936 68026 6992 68028
rect 6696 67974 6742 68026
rect 6742 67974 6752 68026
rect 6776 67974 6806 68026
rect 6806 67974 6818 68026
rect 6818 67974 6832 68026
rect 6856 67974 6870 68026
rect 6870 67974 6882 68026
rect 6882 67974 6912 68026
rect 6936 67974 6946 68026
rect 6946 67974 6992 68026
rect 6696 67972 6752 67974
rect 6776 67972 6832 67974
rect 6856 67972 6912 67974
rect 6936 67972 6992 67974
rect 2906 67620 2962 67656
rect 2906 67600 2908 67620
rect 2908 67600 2960 67620
rect 2960 67600 2962 67620
rect 5960 67482 6016 67484
rect 6040 67482 6096 67484
rect 6120 67482 6176 67484
rect 6200 67482 6256 67484
rect 5960 67430 6006 67482
rect 6006 67430 6016 67482
rect 6040 67430 6070 67482
rect 6070 67430 6082 67482
rect 6082 67430 6096 67482
rect 6120 67430 6134 67482
rect 6134 67430 6146 67482
rect 6146 67430 6176 67482
rect 6200 67430 6210 67482
rect 6210 67430 6256 67482
rect 5960 67428 6016 67430
rect 6040 67428 6096 67430
rect 6120 67428 6176 67430
rect 6200 67428 6256 67430
rect 7138 67092 7140 67112
rect 7140 67092 7192 67112
rect 7192 67092 7194 67112
rect 7138 67056 7194 67092
rect 2906 66920 2962 66976
rect 6696 66938 6752 66940
rect 6776 66938 6832 66940
rect 6856 66938 6912 66940
rect 6936 66938 6992 66940
rect 6696 66886 6742 66938
rect 6742 66886 6752 66938
rect 6776 66886 6806 66938
rect 6806 66886 6818 66938
rect 6818 66886 6832 66938
rect 6856 66886 6870 66938
rect 6870 66886 6882 66938
rect 6882 66886 6912 66938
rect 6936 66886 6946 66938
rect 6946 66886 6992 66938
rect 6696 66884 6752 66886
rect 6776 66884 6832 66886
rect 6856 66884 6912 66886
rect 6936 66884 6992 66886
rect 5960 66394 6016 66396
rect 6040 66394 6096 66396
rect 6120 66394 6176 66396
rect 6200 66394 6256 66396
rect 5960 66342 6006 66394
rect 6006 66342 6016 66394
rect 6040 66342 6070 66394
rect 6070 66342 6082 66394
rect 6082 66342 6096 66394
rect 6120 66342 6134 66394
rect 6134 66342 6146 66394
rect 6146 66342 6176 66394
rect 6200 66342 6210 66394
rect 6210 66342 6256 66394
rect 5960 66340 6016 66342
rect 6040 66340 6096 66342
rect 6120 66340 6176 66342
rect 6200 66340 6256 66342
rect 6696 65850 6752 65852
rect 6776 65850 6832 65852
rect 6856 65850 6912 65852
rect 6936 65850 6992 65852
rect 6696 65798 6742 65850
rect 6742 65798 6752 65850
rect 6776 65798 6806 65850
rect 6806 65798 6818 65850
rect 6818 65798 6832 65850
rect 6856 65798 6870 65850
rect 6870 65798 6882 65850
rect 6882 65798 6912 65850
rect 6936 65798 6946 65850
rect 6946 65798 6992 65850
rect 6696 65796 6752 65798
rect 6776 65796 6832 65798
rect 6856 65796 6912 65798
rect 6936 65796 6992 65798
rect 2906 65560 2962 65616
rect 5960 65306 6016 65308
rect 6040 65306 6096 65308
rect 6120 65306 6176 65308
rect 6200 65306 6256 65308
rect 5960 65254 6006 65306
rect 6006 65254 6016 65306
rect 6040 65254 6070 65306
rect 6070 65254 6082 65306
rect 6082 65254 6096 65306
rect 6120 65254 6134 65306
rect 6134 65254 6146 65306
rect 6146 65254 6176 65306
rect 6200 65254 6210 65306
rect 6210 65254 6256 65306
rect 5960 65252 6016 65254
rect 6040 65252 6096 65254
rect 6120 65252 6176 65254
rect 6200 65252 6256 65254
rect 2906 64900 2962 64936
rect 2906 64880 2908 64900
rect 2908 64880 2960 64900
rect 2960 64880 2962 64900
rect 6696 64762 6752 64764
rect 6776 64762 6832 64764
rect 6856 64762 6912 64764
rect 6936 64762 6992 64764
rect 6696 64710 6742 64762
rect 6742 64710 6752 64762
rect 6776 64710 6806 64762
rect 6806 64710 6818 64762
rect 6818 64710 6832 64762
rect 6856 64710 6870 64762
rect 6870 64710 6882 64762
rect 6882 64710 6912 64762
rect 6936 64710 6946 64762
rect 6946 64710 6992 64762
rect 6696 64708 6752 64710
rect 6776 64708 6832 64710
rect 6856 64708 6912 64710
rect 6936 64708 6992 64710
rect 5960 64218 6016 64220
rect 6040 64218 6096 64220
rect 6120 64218 6176 64220
rect 6200 64218 6256 64220
rect 5960 64166 6006 64218
rect 6006 64166 6016 64218
rect 6040 64166 6070 64218
rect 6070 64166 6082 64218
rect 6082 64166 6096 64218
rect 6120 64166 6134 64218
rect 6134 64166 6146 64218
rect 6146 64166 6176 64218
rect 6200 64166 6210 64218
rect 6210 64166 6256 64218
rect 5960 64164 6016 64166
rect 6040 64164 6096 64166
rect 6120 64164 6176 64166
rect 6200 64164 6256 64166
rect 6696 63674 6752 63676
rect 6776 63674 6832 63676
rect 6856 63674 6912 63676
rect 6936 63674 6992 63676
rect 6696 63622 6742 63674
rect 6742 63622 6752 63674
rect 6776 63622 6806 63674
rect 6806 63622 6818 63674
rect 6818 63622 6832 63674
rect 6856 63622 6870 63674
rect 6870 63622 6882 63674
rect 6882 63622 6912 63674
rect 6936 63622 6946 63674
rect 6946 63622 6992 63674
rect 6696 63620 6752 63622
rect 6776 63620 6832 63622
rect 6856 63620 6912 63622
rect 6936 63620 6992 63622
rect 5206 63520 5262 63576
rect 5960 63130 6016 63132
rect 6040 63130 6096 63132
rect 6120 63130 6176 63132
rect 6200 63130 6256 63132
rect 5960 63078 6006 63130
rect 6006 63078 6016 63130
rect 6040 63078 6070 63130
rect 6070 63078 6082 63130
rect 6082 63078 6096 63130
rect 6120 63078 6134 63130
rect 6134 63078 6146 63130
rect 6146 63078 6176 63130
rect 6200 63078 6210 63130
rect 6210 63078 6256 63130
rect 5960 63076 6016 63078
rect 6040 63076 6096 63078
rect 6120 63076 6176 63078
rect 6200 63076 6256 63078
rect 6696 62586 6752 62588
rect 6776 62586 6832 62588
rect 6856 62586 6912 62588
rect 6936 62586 6992 62588
rect 6696 62534 6742 62586
rect 6742 62534 6752 62586
rect 6776 62534 6806 62586
rect 6806 62534 6818 62586
rect 6818 62534 6832 62586
rect 6856 62534 6870 62586
rect 6870 62534 6882 62586
rect 6882 62534 6912 62586
rect 6936 62534 6946 62586
rect 6946 62534 6992 62586
rect 6696 62532 6752 62534
rect 6776 62532 6832 62534
rect 6856 62532 6912 62534
rect 6936 62532 6992 62534
rect 4930 62160 4986 62216
rect 5960 62042 6016 62044
rect 6040 62042 6096 62044
rect 6120 62042 6176 62044
rect 6200 62042 6256 62044
rect 5960 61990 6006 62042
rect 6006 61990 6016 62042
rect 6040 61990 6070 62042
rect 6070 61990 6082 62042
rect 6082 61990 6096 62042
rect 6120 61990 6134 62042
rect 6134 61990 6146 62042
rect 6146 61990 6176 62042
rect 6200 61990 6210 62042
rect 6210 61990 6256 62042
rect 5960 61988 6016 61990
rect 6040 61988 6096 61990
rect 6120 61988 6176 61990
rect 6200 61988 6256 61990
rect 2906 61480 2962 61536
rect 6696 61498 6752 61500
rect 6776 61498 6832 61500
rect 6856 61498 6912 61500
rect 6936 61498 6992 61500
rect 6696 61446 6742 61498
rect 6742 61446 6752 61498
rect 6776 61446 6806 61498
rect 6806 61446 6818 61498
rect 6818 61446 6832 61498
rect 6856 61446 6870 61498
rect 6870 61446 6882 61498
rect 6882 61446 6912 61498
rect 6936 61446 6946 61498
rect 6946 61446 6992 61498
rect 6696 61444 6752 61446
rect 6776 61444 6832 61446
rect 6856 61444 6912 61446
rect 6936 61444 6992 61446
rect 5960 60954 6016 60956
rect 6040 60954 6096 60956
rect 6120 60954 6176 60956
rect 6200 60954 6256 60956
rect 5960 60902 6006 60954
rect 6006 60902 6016 60954
rect 6040 60902 6070 60954
rect 6070 60902 6082 60954
rect 6082 60902 6096 60954
rect 6120 60902 6134 60954
rect 6134 60902 6146 60954
rect 6146 60902 6176 60954
rect 6200 60902 6210 60954
rect 6210 60902 6256 60954
rect 5960 60900 6016 60902
rect 6040 60900 6096 60902
rect 6120 60900 6176 60902
rect 6200 60900 6256 60902
rect 6696 60410 6752 60412
rect 6776 60410 6832 60412
rect 6856 60410 6912 60412
rect 6936 60410 6992 60412
rect 6696 60358 6742 60410
rect 6742 60358 6752 60410
rect 6776 60358 6806 60410
rect 6806 60358 6818 60410
rect 6818 60358 6832 60410
rect 6856 60358 6870 60410
rect 6870 60358 6882 60410
rect 6882 60358 6912 60410
rect 6936 60358 6946 60410
rect 6946 60358 6992 60410
rect 6696 60356 6752 60358
rect 6776 60356 6832 60358
rect 6856 60356 6912 60358
rect 6936 60356 6992 60358
rect 2906 60120 2962 60176
rect 5960 59866 6016 59868
rect 6040 59866 6096 59868
rect 6120 59866 6176 59868
rect 6200 59866 6256 59868
rect 5960 59814 6006 59866
rect 6006 59814 6016 59866
rect 6040 59814 6070 59866
rect 6070 59814 6082 59866
rect 6082 59814 6096 59866
rect 6120 59814 6134 59866
rect 6134 59814 6146 59866
rect 6146 59814 6176 59866
rect 6200 59814 6210 59866
rect 6210 59814 6256 59866
rect 5960 59812 6016 59814
rect 6040 59812 6096 59814
rect 6120 59812 6176 59814
rect 6200 59812 6256 59814
rect 5206 59476 5208 59496
rect 5208 59476 5260 59496
rect 5260 59476 5262 59496
rect 5206 59440 5262 59476
rect 6696 59322 6752 59324
rect 6776 59322 6832 59324
rect 6856 59322 6912 59324
rect 6936 59322 6992 59324
rect 6696 59270 6742 59322
rect 6742 59270 6752 59322
rect 6776 59270 6806 59322
rect 6806 59270 6818 59322
rect 6818 59270 6832 59322
rect 6856 59270 6870 59322
rect 6870 59270 6882 59322
rect 6882 59270 6912 59322
rect 6936 59270 6946 59322
rect 6946 59270 6992 59322
rect 6696 59268 6752 59270
rect 6776 59268 6832 59270
rect 6856 59268 6912 59270
rect 6936 59268 6992 59270
rect 5960 58778 6016 58780
rect 6040 58778 6096 58780
rect 6120 58778 6176 58780
rect 6200 58778 6256 58780
rect 5960 58726 6006 58778
rect 6006 58726 6016 58778
rect 6040 58726 6070 58778
rect 6070 58726 6082 58778
rect 6082 58726 6096 58778
rect 6120 58726 6134 58778
rect 6134 58726 6146 58778
rect 6146 58726 6176 58778
rect 6200 58726 6210 58778
rect 6210 58726 6256 58778
rect 5960 58724 6016 58726
rect 6040 58724 6096 58726
rect 6120 58724 6176 58726
rect 6200 58724 6256 58726
rect 5206 58080 5262 58136
rect 6696 58234 6752 58236
rect 6776 58234 6832 58236
rect 6856 58234 6912 58236
rect 6936 58234 6992 58236
rect 6696 58182 6742 58234
rect 6742 58182 6752 58234
rect 6776 58182 6806 58234
rect 6806 58182 6818 58234
rect 6818 58182 6832 58234
rect 6856 58182 6870 58234
rect 6870 58182 6882 58234
rect 6882 58182 6912 58234
rect 6936 58182 6946 58234
rect 6946 58182 6992 58234
rect 6696 58180 6752 58182
rect 6776 58180 6832 58182
rect 6856 58180 6912 58182
rect 6936 58180 6992 58182
rect 5390 57944 5446 58000
rect 5960 57690 6016 57692
rect 6040 57690 6096 57692
rect 6120 57690 6176 57692
rect 6200 57690 6256 57692
rect 5960 57638 6006 57690
rect 6006 57638 6016 57690
rect 6040 57638 6070 57690
rect 6070 57638 6082 57690
rect 6082 57638 6096 57690
rect 6120 57638 6134 57690
rect 6134 57638 6146 57690
rect 6146 57638 6176 57690
rect 6200 57638 6210 57690
rect 6210 57638 6256 57690
rect 5960 57636 6016 57638
rect 6040 57636 6096 57638
rect 6120 57636 6176 57638
rect 6200 57636 6256 57638
rect 6696 57146 6752 57148
rect 6776 57146 6832 57148
rect 6856 57146 6912 57148
rect 6936 57146 6992 57148
rect 6696 57094 6742 57146
rect 6742 57094 6752 57146
rect 6776 57094 6806 57146
rect 6806 57094 6818 57146
rect 6818 57094 6832 57146
rect 6856 57094 6870 57146
rect 6870 57094 6882 57146
rect 6882 57094 6912 57146
rect 6936 57094 6946 57146
rect 6946 57094 6992 57146
rect 6696 57092 6752 57094
rect 6776 57092 6832 57094
rect 6856 57092 6912 57094
rect 6936 57092 6992 57094
rect 4930 56720 4986 56776
rect 5960 56602 6016 56604
rect 6040 56602 6096 56604
rect 6120 56602 6176 56604
rect 6200 56602 6256 56604
rect 5960 56550 6006 56602
rect 6006 56550 6016 56602
rect 6040 56550 6070 56602
rect 6070 56550 6082 56602
rect 6082 56550 6096 56602
rect 6120 56550 6134 56602
rect 6134 56550 6146 56602
rect 6146 56550 6176 56602
rect 6200 56550 6210 56602
rect 6210 56550 6256 56602
rect 5960 56548 6016 56550
rect 6040 56548 6096 56550
rect 6120 56548 6176 56550
rect 6200 56548 6256 56550
rect 2906 56040 2962 56096
rect 6696 56058 6752 56060
rect 6776 56058 6832 56060
rect 6856 56058 6912 56060
rect 6936 56058 6992 56060
rect 6696 56006 6742 56058
rect 6742 56006 6752 56058
rect 6776 56006 6806 56058
rect 6806 56006 6818 56058
rect 6818 56006 6832 56058
rect 6856 56006 6870 56058
rect 6870 56006 6882 56058
rect 6882 56006 6912 56058
rect 6936 56006 6946 56058
rect 6946 56006 6992 56058
rect 6696 56004 6752 56006
rect 6776 56004 6832 56006
rect 6856 56004 6912 56006
rect 6936 56004 6992 56006
rect 5960 55514 6016 55516
rect 6040 55514 6096 55516
rect 6120 55514 6176 55516
rect 6200 55514 6256 55516
rect 5960 55462 6006 55514
rect 6006 55462 6016 55514
rect 6040 55462 6070 55514
rect 6070 55462 6082 55514
rect 6082 55462 6096 55514
rect 6120 55462 6134 55514
rect 6134 55462 6146 55514
rect 6146 55462 6176 55514
rect 6200 55462 6210 55514
rect 6210 55462 6256 55514
rect 5960 55460 6016 55462
rect 6040 55460 6096 55462
rect 6120 55460 6176 55462
rect 6200 55460 6256 55462
rect 6696 54970 6752 54972
rect 6776 54970 6832 54972
rect 6856 54970 6912 54972
rect 6936 54970 6992 54972
rect 6696 54918 6742 54970
rect 6742 54918 6752 54970
rect 6776 54918 6806 54970
rect 6806 54918 6818 54970
rect 6818 54918 6832 54970
rect 6856 54918 6870 54970
rect 6870 54918 6882 54970
rect 6882 54918 6912 54970
rect 6936 54918 6946 54970
rect 6946 54918 6992 54970
rect 6696 54916 6752 54918
rect 6776 54916 6832 54918
rect 6856 54916 6912 54918
rect 6936 54916 6992 54918
rect 2906 54680 2962 54736
rect 5960 54426 6016 54428
rect 6040 54426 6096 54428
rect 6120 54426 6176 54428
rect 6200 54426 6256 54428
rect 5960 54374 6006 54426
rect 6006 54374 6016 54426
rect 6040 54374 6070 54426
rect 6070 54374 6082 54426
rect 6082 54374 6096 54426
rect 6120 54374 6134 54426
rect 6134 54374 6146 54426
rect 6146 54374 6176 54426
rect 6200 54374 6210 54426
rect 6210 54374 6256 54426
rect 5960 54372 6016 54374
rect 6040 54372 6096 54374
rect 6120 54372 6176 54374
rect 6200 54372 6256 54374
rect 5114 54036 5116 54056
rect 5116 54036 5168 54056
rect 5168 54036 5170 54056
rect 5114 54000 5170 54036
rect 5666 54036 5668 54056
rect 5668 54036 5720 54056
rect 5720 54036 5722 54056
rect 5666 54000 5722 54036
rect 6696 53882 6752 53884
rect 6776 53882 6832 53884
rect 6856 53882 6912 53884
rect 6936 53882 6992 53884
rect 6696 53830 6742 53882
rect 6742 53830 6752 53882
rect 6776 53830 6806 53882
rect 6806 53830 6818 53882
rect 6818 53830 6832 53882
rect 6856 53830 6870 53882
rect 6870 53830 6882 53882
rect 6882 53830 6912 53882
rect 6936 53830 6946 53882
rect 6946 53830 6992 53882
rect 6696 53828 6752 53830
rect 6776 53828 6832 53830
rect 6856 53828 6912 53830
rect 6936 53828 6992 53830
rect 5960 53338 6016 53340
rect 6040 53338 6096 53340
rect 6120 53338 6176 53340
rect 6200 53338 6256 53340
rect 5960 53286 6006 53338
rect 6006 53286 6016 53338
rect 6040 53286 6070 53338
rect 6070 53286 6082 53338
rect 6082 53286 6096 53338
rect 6120 53286 6134 53338
rect 6134 53286 6146 53338
rect 6146 53286 6176 53338
rect 6200 53286 6210 53338
rect 6210 53286 6256 53338
rect 5960 53284 6016 53286
rect 6040 53284 6096 53286
rect 6120 53284 6176 53286
rect 6200 53284 6256 53286
rect 6696 52794 6752 52796
rect 6776 52794 6832 52796
rect 6856 52794 6912 52796
rect 6936 52794 6992 52796
rect 6696 52742 6742 52794
rect 6742 52742 6752 52794
rect 6776 52742 6806 52794
rect 6806 52742 6818 52794
rect 6818 52742 6832 52794
rect 6856 52742 6870 52794
rect 6870 52742 6882 52794
rect 6882 52742 6912 52794
rect 6936 52742 6946 52794
rect 6946 52742 6992 52794
rect 6696 52740 6752 52742
rect 6776 52740 6832 52742
rect 6856 52740 6912 52742
rect 6936 52740 6992 52742
rect 2906 52640 2962 52696
rect 5960 52250 6016 52252
rect 6040 52250 6096 52252
rect 6120 52250 6176 52252
rect 6200 52250 6256 52252
rect 5960 52198 6006 52250
rect 6006 52198 6016 52250
rect 6040 52198 6070 52250
rect 6070 52198 6082 52250
rect 6082 52198 6096 52250
rect 6120 52198 6134 52250
rect 6134 52198 6146 52250
rect 6146 52198 6176 52250
rect 6200 52198 6210 52250
rect 6210 52198 6256 52250
rect 5960 52196 6016 52198
rect 6040 52196 6096 52198
rect 6120 52196 6176 52198
rect 6200 52196 6256 52198
rect 6696 51706 6752 51708
rect 6776 51706 6832 51708
rect 6856 51706 6912 51708
rect 6936 51706 6992 51708
rect 6696 51654 6742 51706
rect 6742 51654 6752 51706
rect 6776 51654 6806 51706
rect 6806 51654 6818 51706
rect 6818 51654 6832 51706
rect 6856 51654 6870 51706
rect 6870 51654 6882 51706
rect 6882 51654 6912 51706
rect 6936 51654 6946 51706
rect 6946 51654 6992 51706
rect 6696 51652 6752 51654
rect 6776 51652 6832 51654
rect 6856 51652 6912 51654
rect 6936 51652 6992 51654
rect 2906 51280 2962 51336
rect 5960 51162 6016 51164
rect 6040 51162 6096 51164
rect 6120 51162 6176 51164
rect 6200 51162 6256 51164
rect 5960 51110 6006 51162
rect 6006 51110 6016 51162
rect 6040 51110 6070 51162
rect 6070 51110 6082 51162
rect 6082 51110 6096 51162
rect 6120 51110 6134 51162
rect 6134 51110 6146 51162
rect 6146 51110 6176 51162
rect 6200 51110 6210 51162
rect 6210 51110 6256 51162
rect 5960 51108 6016 51110
rect 6040 51108 6096 51110
rect 6120 51108 6176 51110
rect 6200 51108 6256 51110
rect 6696 50618 6752 50620
rect 6776 50618 6832 50620
rect 6856 50618 6912 50620
rect 6936 50618 6992 50620
rect 6696 50566 6742 50618
rect 6742 50566 6752 50618
rect 6776 50566 6806 50618
rect 6806 50566 6818 50618
rect 6818 50566 6832 50618
rect 6856 50566 6870 50618
rect 6870 50566 6882 50618
rect 6882 50566 6912 50618
rect 6936 50566 6946 50618
rect 6946 50566 6992 50618
rect 6696 50564 6752 50566
rect 6776 50564 6832 50566
rect 6856 50564 6912 50566
rect 6936 50564 6992 50566
rect 5960 50074 6016 50076
rect 6040 50074 6096 50076
rect 6120 50074 6176 50076
rect 6200 50074 6256 50076
rect 5960 50022 6006 50074
rect 6006 50022 6016 50074
rect 6040 50022 6070 50074
rect 6070 50022 6082 50074
rect 6082 50022 6096 50074
rect 6120 50022 6134 50074
rect 6134 50022 6146 50074
rect 6146 50022 6176 50074
rect 6200 50022 6210 50074
rect 6210 50022 6256 50074
rect 5960 50020 6016 50022
rect 6040 50020 6096 50022
rect 6120 50020 6176 50022
rect 6200 50020 6256 50022
rect 6696 49530 6752 49532
rect 6776 49530 6832 49532
rect 6856 49530 6912 49532
rect 6936 49530 6992 49532
rect 6696 49478 6742 49530
rect 6742 49478 6752 49530
rect 6776 49478 6806 49530
rect 6806 49478 6818 49530
rect 6818 49478 6832 49530
rect 6856 49478 6870 49530
rect 6870 49478 6882 49530
rect 6882 49478 6912 49530
rect 6936 49478 6946 49530
rect 6946 49478 6992 49530
rect 6696 49476 6752 49478
rect 6776 49476 6832 49478
rect 6856 49476 6912 49478
rect 6936 49476 6992 49478
rect 5960 48986 6016 48988
rect 6040 48986 6096 48988
rect 6120 48986 6176 48988
rect 6200 48986 6256 48988
rect 5960 48934 6006 48986
rect 6006 48934 6016 48986
rect 6040 48934 6070 48986
rect 6070 48934 6082 48986
rect 6082 48934 6096 48986
rect 6120 48934 6134 48986
rect 6134 48934 6146 48986
rect 6146 48934 6176 48986
rect 6200 48934 6210 48986
rect 6210 48934 6256 48986
rect 5960 48932 6016 48934
rect 6040 48932 6096 48934
rect 6120 48932 6176 48934
rect 6200 48932 6256 48934
rect 6696 48442 6752 48444
rect 6776 48442 6832 48444
rect 6856 48442 6912 48444
rect 6936 48442 6992 48444
rect 6696 48390 6742 48442
rect 6742 48390 6752 48442
rect 6776 48390 6806 48442
rect 6806 48390 6818 48442
rect 6818 48390 6832 48442
rect 6856 48390 6870 48442
rect 6870 48390 6882 48442
rect 6882 48390 6912 48442
rect 6936 48390 6946 48442
rect 6946 48390 6992 48442
rect 6696 48388 6752 48390
rect 6776 48388 6832 48390
rect 6856 48388 6912 48390
rect 6936 48388 6992 48390
rect 5960 47898 6016 47900
rect 6040 47898 6096 47900
rect 6120 47898 6176 47900
rect 6200 47898 6256 47900
rect 5960 47846 6006 47898
rect 6006 47846 6016 47898
rect 6040 47846 6070 47898
rect 6070 47846 6082 47898
rect 6082 47846 6096 47898
rect 6120 47846 6134 47898
rect 6134 47846 6146 47898
rect 6146 47846 6176 47898
rect 6200 47846 6210 47898
rect 6210 47846 6256 47898
rect 5960 47844 6016 47846
rect 6040 47844 6096 47846
rect 6120 47844 6176 47846
rect 6200 47844 6256 47846
rect 6696 47354 6752 47356
rect 6776 47354 6832 47356
rect 6856 47354 6912 47356
rect 6936 47354 6992 47356
rect 6696 47302 6742 47354
rect 6742 47302 6752 47354
rect 6776 47302 6806 47354
rect 6806 47302 6818 47354
rect 6818 47302 6832 47354
rect 6856 47302 6870 47354
rect 6870 47302 6882 47354
rect 6882 47302 6912 47354
rect 6936 47302 6946 47354
rect 6946 47302 6992 47354
rect 6696 47300 6752 47302
rect 6776 47300 6832 47302
rect 6856 47300 6912 47302
rect 6936 47300 6992 47302
rect 5960 46810 6016 46812
rect 6040 46810 6096 46812
rect 6120 46810 6176 46812
rect 6200 46810 6256 46812
rect 5960 46758 6006 46810
rect 6006 46758 6016 46810
rect 6040 46758 6070 46810
rect 6070 46758 6082 46810
rect 6082 46758 6096 46810
rect 6120 46758 6134 46810
rect 6134 46758 6146 46810
rect 6146 46758 6176 46810
rect 6200 46758 6210 46810
rect 6210 46758 6256 46810
rect 5960 46756 6016 46758
rect 6040 46756 6096 46758
rect 6120 46756 6176 46758
rect 6200 46756 6256 46758
rect 6696 46266 6752 46268
rect 6776 46266 6832 46268
rect 6856 46266 6912 46268
rect 6936 46266 6992 46268
rect 6696 46214 6742 46266
rect 6742 46214 6752 46266
rect 6776 46214 6806 46266
rect 6806 46214 6818 46266
rect 6818 46214 6832 46266
rect 6856 46214 6870 46266
rect 6870 46214 6882 46266
rect 6882 46214 6912 46266
rect 6936 46214 6946 46266
rect 6946 46214 6992 46266
rect 6696 46212 6752 46214
rect 6776 46212 6832 46214
rect 6856 46212 6912 46214
rect 6936 46212 6992 46214
rect 5960 45722 6016 45724
rect 6040 45722 6096 45724
rect 6120 45722 6176 45724
rect 6200 45722 6256 45724
rect 5960 45670 6006 45722
rect 6006 45670 6016 45722
rect 6040 45670 6070 45722
rect 6070 45670 6082 45722
rect 6082 45670 6096 45722
rect 6120 45670 6134 45722
rect 6134 45670 6146 45722
rect 6146 45670 6176 45722
rect 6200 45670 6210 45722
rect 6210 45670 6256 45722
rect 5960 45668 6016 45670
rect 6040 45668 6096 45670
rect 6120 45668 6176 45670
rect 6200 45668 6256 45670
rect 7230 65832 7286 65888
rect 7230 64744 7286 64800
rect 17728 87066 17784 87068
rect 17808 87066 17864 87068
rect 17888 87066 17944 87068
rect 17968 87066 18024 87068
rect 17728 87014 17774 87066
rect 17774 87014 17784 87066
rect 17808 87014 17838 87066
rect 17838 87014 17850 87066
rect 17850 87014 17864 87066
rect 17888 87014 17902 87066
rect 17902 87014 17914 87066
rect 17914 87014 17944 87066
rect 17968 87014 17978 87066
rect 17978 87014 18024 87066
rect 17728 87012 17784 87014
rect 17808 87012 17864 87014
rect 17888 87012 17944 87014
rect 17968 87012 18024 87014
rect 17728 85978 17784 85980
rect 17808 85978 17864 85980
rect 17888 85978 17944 85980
rect 17968 85978 18024 85980
rect 17728 85926 17774 85978
rect 17774 85926 17784 85978
rect 17808 85926 17838 85978
rect 17838 85926 17850 85978
rect 17850 85926 17864 85978
rect 17888 85926 17902 85978
rect 17902 85926 17914 85978
rect 17914 85926 17944 85978
rect 17968 85926 17978 85978
rect 17978 85926 18024 85978
rect 17728 85924 17784 85926
rect 17808 85924 17864 85926
rect 17888 85924 17944 85926
rect 17968 85924 18024 85926
rect 17728 84890 17784 84892
rect 17808 84890 17864 84892
rect 17888 84890 17944 84892
rect 17968 84890 18024 84892
rect 17728 84838 17774 84890
rect 17774 84838 17784 84890
rect 17808 84838 17838 84890
rect 17838 84838 17850 84890
rect 17850 84838 17864 84890
rect 17888 84838 17902 84890
rect 17902 84838 17914 84890
rect 17914 84838 17944 84890
rect 17968 84838 17978 84890
rect 17978 84838 18024 84890
rect 17728 84836 17784 84838
rect 17808 84836 17864 84838
rect 17888 84836 17944 84838
rect 17968 84836 18024 84838
rect 18388 86522 18444 86524
rect 18468 86522 18524 86524
rect 18548 86522 18604 86524
rect 18628 86522 18684 86524
rect 18388 86470 18434 86522
rect 18434 86470 18444 86522
rect 18468 86470 18498 86522
rect 18498 86470 18510 86522
rect 18510 86470 18524 86522
rect 18548 86470 18562 86522
rect 18562 86470 18574 86522
rect 18574 86470 18604 86522
rect 18628 86470 18638 86522
rect 18638 86470 18684 86522
rect 18388 86468 18444 86470
rect 18468 86468 18524 86470
rect 18548 86468 18604 86470
rect 18628 86468 18684 86470
rect 18388 85434 18444 85436
rect 18468 85434 18524 85436
rect 18548 85434 18604 85436
rect 18628 85434 18684 85436
rect 18388 85382 18434 85434
rect 18434 85382 18444 85434
rect 18468 85382 18498 85434
rect 18498 85382 18510 85434
rect 18510 85382 18524 85434
rect 18548 85382 18562 85434
rect 18562 85382 18574 85434
rect 18574 85382 18604 85434
rect 18628 85382 18638 85434
rect 18638 85382 18684 85434
rect 18388 85380 18444 85382
rect 18468 85380 18524 85382
rect 18548 85380 18604 85382
rect 18628 85380 18684 85382
rect 18388 84346 18444 84348
rect 18468 84346 18524 84348
rect 18548 84346 18604 84348
rect 18628 84346 18684 84348
rect 18388 84294 18434 84346
rect 18434 84294 18444 84346
rect 18468 84294 18498 84346
rect 18498 84294 18510 84346
rect 18510 84294 18524 84346
rect 18548 84294 18562 84346
rect 18562 84294 18574 84346
rect 18574 84294 18604 84346
rect 18628 84294 18638 84346
rect 18638 84294 18684 84346
rect 18388 84292 18444 84294
rect 18468 84292 18524 84294
rect 18548 84292 18604 84294
rect 18628 84292 18684 84294
rect 7230 62452 7286 62488
rect 7230 62432 7232 62452
rect 7232 62432 7284 62452
rect 7284 62432 7286 62452
rect 7230 61480 7286 61536
rect 7230 60392 7286 60448
rect 7230 59304 7286 59360
rect 7230 57012 7286 57048
rect 7230 56992 7232 57012
rect 7232 56992 7284 57012
rect 7284 56992 7286 57012
rect 7230 56040 7286 56096
rect 7230 54952 7286 55008
rect 7230 52776 7286 52832
rect 7230 51572 7286 51608
rect 7230 51552 7232 51572
rect 7232 51552 7284 51572
rect 7284 51552 7286 51572
rect 10542 82288 10598 82344
rect 36128 87066 36184 87068
rect 36208 87066 36264 87068
rect 36288 87066 36344 87068
rect 36368 87066 36424 87068
rect 36128 87014 36174 87066
rect 36174 87014 36184 87066
rect 36208 87014 36238 87066
rect 36238 87014 36250 87066
rect 36250 87014 36264 87066
rect 36288 87014 36302 87066
rect 36302 87014 36314 87066
rect 36314 87014 36344 87066
rect 36368 87014 36378 87066
rect 36378 87014 36424 87066
rect 36128 87012 36184 87014
rect 36208 87012 36264 87014
rect 36288 87012 36344 87014
rect 36368 87012 36424 87014
rect 36788 86522 36844 86524
rect 36868 86522 36924 86524
rect 36948 86522 37004 86524
rect 37028 86522 37084 86524
rect 36788 86470 36834 86522
rect 36834 86470 36844 86522
rect 36868 86470 36898 86522
rect 36898 86470 36910 86522
rect 36910 86470 36924 86522
rect 36948 86470 36962 86522
rect 36962 86470 36974 86522
rect 36974 86470 37004 86522
rect 37028 86470 37038 86522
rect 37038 86470 37084 86522
rect 36788 86468 36844 86470
rect 36868 86468 36924 86470
rect 36948 86468 37004 86470
rect 37028 86468 37084 86470
rect 36128 85978 36184 85980
rect 36208 85978 36264 85980
rect 36288 85978 36344 85980
rect 36368 85978 36424 85980
rect 36128 85926 36174 85978
rect 36174 85926 36184 85978
rect 36208 85926 36238 85978
rect 36238 85926 36250 85978
rect 36250 85926 36264 85978
rect 36288 85926 36302 85978
rect 36302 85926 36314 85978
rect 36314 85926 36344 85978
rect 36368 85926 36378 85978
rect 36378 85926 36424 85978
rect 36128 85924 36184 85926
rect 36208 85924 36264 85926
rect 36288 85924 36344 85926
rect 36368 85924 36424 85926
rect 36788 85434 36844 85436
rect 36868 85434 36924 85436
rect 36948 85434 37004 85436
rect 37028 85434 37084 85436
rect 36788 85382 36834 85434
rect 36834 85382 36844 85434
rect 36868 85382 36898 85434
rect 36898 85382 36910 85434
rect 36910 85382 36924 85434
rect 36948 85382 36962 85434
rect 36962 85382 36974 85434
rect 36974 85382 37004 85434
rect 37028 85382 37038 85434
rect 37038 85382 37084 85434
rect 36788 85380 36844 85382
rect 36868 85380 36924 85382
rect 36948 85380 37004 85382
rect 37028 85380 37084 85382
rect 36128 84890 36184 84892
rect 36208 84890 36264 84892
rect 36288 84890 36344 84892
rect 36368 84890 36424 84892
rect 36128 84838 36174 84890
rect 36174 84838 36184 84890
rect 36208 84838 36238 84890
rect 36238 84838 36250 84890
rect 36250 84838 36264 84890
rect 36288 84838 36302 84890
rect 36302 84838 36314 84890
rect 36314 84838 36344 84890
rect 36368 84838 36378 84890
rect 36378 84838 36424 84890
rect 36128 84836 36184 84838
rect 36208 84836 36264 84838
rect 36288 84836 36344 84838
rect 36368 84836 36424 84838
rect 36788 84346 36844 84348
rect 36868 84346 36924 84348
rect 36948 84346 37004 84348
rect 37028 84346 37084 84348
rect 36788 84294 36834 84346
rect 36834 84294 36844 84346
rect 36868 84294 36898 84346
rect 36898 84294 36910 84346
rect 36910 84294 36924 84346
rect 36948 84294 36962 84346
rect 36962 84294 36974 84346
rect 36974 84294 37004 84346
rect 37028 84294 37038 84346
rect 37038 84294 37084 84346
rect 36788 84292 36844 84294
rect 36868 84292 36924 84294
rect 36948 84292 37004 84294
rect 37028 84292 37084 84294
rect 55188 87610 55244 87612
rect 55268 87610 55324 87612
rect 55348 87610 55404 87612
rect 55428 87610 55484 87612
rect 55188 87558 55234 87610
rect 55234 87558 55244 87610
rect 55268 87558 55298 87610
rect 55298 87558 55310 87610
rect 55310 87558 55324 87610
rect 55348 87558 55362 87610
rect 55362 87558 55374 87610
rect 55374 87558 55404 87610
rect 55428 87558 55438 87610
rect 55438 87558 55484 87610
rect 55188 87556 55244 87558
rect 55268 87556 55324 87558
rect 55348 87556 55404 87558
rect 55428 87556 55484 87558
rect 73588 87610 73644 87612
rect 73668 87610 73724 87612
rect 73748 87610 73804 87612
rect 73828 87610 73884 87612
rect 73588 87558 73634 87610
rect 73634 87558 73644 87610
rect 73668 87558 73698 87610
rect 73698 87558 73710 87610
rect 73710 87558 73724 87610
rect 73748 87558 73762 87610
rect 73762 87558 73774 87610
rect 73774 87558 73804 87610
rect 73828 87558 73838 87610
rect 73838 87558 73884 87610
rect 73588 87556 73644 87558
rect 73668 87556 73724 87558
rect 73748 87556 73804 87558
rect 73828 87556 73884 87558
rect 9990 82016 10046 82072
rect 10542 82016 10598 82072
rect 9622 63588 9678 63644
rect 45962 50532 46018 50588
rect 45870 49444 45926 49500
rect 7138 45468 7140 45488
rect 7140 45468 7192 45488
rect 7192 45468 7194 45488
rect 7138 45432 7194 45468
rect 9990 45588 10046 45624
rect 9990 45568 9992 45588
rect 9992 45568 10044 45588
rect 10044 45568 10046 45588
rect 10542 45568 10598 45624
rect 12778 45432 12834 45488
rect 7506 45296 7562 45352
rect 11674 45296 11730 45352
rect 2906 45160 2962 45216
rect 6696 45178 6752 45180
rect 6776 45178 6832 45180
rect 6856 45178 6912 45180
rect 6936 45178 6992 45180
rect 6696 45126 6742 45178
rect 6742 45126 6752 45178
rect 6776 45126 6806 45178
rect 6806 45126 6818 45178
rect 6818 45126 6832 45178
rect 6856 45126 6870 45178
rect 6870 45126 6882 45178
rect 6882 45126 6912 45178
rect 6936 45126 6946 45178
rect 6946 45126 6992 45178
rect 6696 45124 6752 45126
rect 6776 45124 6832 45126
rect 6856 45124 6912 45126
rect 6936 45124 6992 45126
rect 5960 44634 6016 44636
rect 6040 44634 6096 44636
rect 6120 44634 6176 44636
rect 6200 44634 6256 44636
rect 5960 44582 6006 44634
rect 6006 44582 6016 44634
rect 6040 44582 6070 44634
rect 6070 44582 6082 44634
rect 6082 44582 6096 44634
rect 6120 44582 6134 44634
rect 6134 44582 6146 44634
rect 6146 44582 6176 44634
rect 6200 44582 6210 44634
rect 6210 44582 6256 44634
rect 7138 44616 7194 44672
rect 5960 44580 6016 44582
rect 6040 44580 6096 44582
rect 6120 44580 6176 44582
rect 6200 44580 6256 44582
rect 2906 44480 2962 44536
rect 6696 44090 6752 44092
rect 6776 44090 6832 44092
rect 6856 44090 6912 44092
rect 6936 44090 6992 44092
rect 6696 44038 6742 44090
rect 6742 44038 6752 44090
rect 6776 44038 6806 44090
rect 6806 44038 6818 44090
rect 6818 44038 6832 44090
rect 6856 44038 6870 44090
rect 6870 44038 6882 44090
rect 6882 44038 6912 44090
rect 6936 44038 6946 44090
rect 6946 44038 6992 44090
rect 6696 44036 6752 44038
rect 6776 44036 6832 44038
rect 6856 44036 6912 44038
rect 6936 44036 6992 44038
rect 2722 43800 2778 43856
rect 5960 43546 6016 43548
rect 6040 43546 6096 43548
rect 6120 43546 6176 43548
rect 6200 43546 6256 43548
rect 5960 43494 6006 43546
rect 6006 43494 6016 43546
rect 6040 43494 6070 43546
rect 6070 43494 6082 43546
rect 6082 43494 6096 43546
rect 6120 43494 6134 43546
rect 6134 43494 6146 43546
rect 6146 43494 6176 43546
rect 6200 43494 6210 43546
rect 6210 43494 6256 43546
rect 8150 43528 8206 43584
rect 5960 43492 6016 43494
rect 6040 43492 6096 43494
rect 6120 43492 6176 43494
rect 6200 43492 6256 43494
rect 6696 43002 6752 43004
rect 6776 43002 6832 43004
rect 6856 43002 6912 43004
rect 6936 43002 6992 43004
rect 6696 42950 6742 43002
rect 6742 42950 6752 43002
rect 6776 42950 6806 43002
rect 6806 42950 6818 43002
rect 6818 42950 6832 43002
rect 6856 42950 6870 43002
rect 6870 42950 6882 43002
rect 6882 42950 6912 43002
rect 6936 42950 6946 43002
rect 6946 42950 6992 43002
rect 6696 42948 6752 42950
rect 6776 42948 6832 42950
rect 6856 42948 6912 42950
rect 6936 42948 6992 42950
rect 2906 42440 2962 42496
rect 5960 42458 6016 42460
rect 6040 42458 6096 42460
rect 6120 42458 6176 42460
rect 6200 42458 6256 42460
rect 5960 42406 6006 42458
rect 6006 42406 6016 42458
rect 6040 42406 6070 42458
rect 6070 42406 6082 42458
rect 6082 42406 6096 42458
rect 6120 42406 6134 42458
rect 6134 42406 6146 42458
rect 6146 42406 6176 42458
rect 6200 42406 6210 42458
rect 6210 42406 6256 42458
rect 7138 42440 7194 42496
rect 5960 42404 6016 42406
rect 6040 42404 6096 42406
rect 6120 42404 6176 42406
rect 6200 42404 6256 42406
rect 6696 41914 6752 41916
rect 6776 41914 6832 41916
rect 6856 41914 6912 41916
rect 6936 41914 6992 41916
rect 6696 41862 6742 41914
rect 6742 41862 6752 41914
rect 6776 41862 6806 41914
rect 6806 41862 6818 41914
rect 6818 41862 6832 41914
rect 6856 41862 6870 41914
rect 6870 41862 6882 41914
rect 6882 41862 6912 41914
rect 6936 41862 6946 41914
rect 6946 41862 6992 41914
rect 6696 41860 6752 41862
rect 6776 41860 6832 41862
rect 6856 41860 6912 41862
rect 6936 41860 6992 41862
rect 5666 41488 5722 41544
rect 5960 41370 6016 41372
rect 6040 41370 6096 41372
rect 6120 41370 6176 41372
rect 6200 41370 6256 41372
rect 5960 41318 6006 41370
rect 6006 41318 6016 41370
rect 6040 41318 6070 41370
rect 6070 41318 6082 41370
rect 6082 41318 6096 41370
rect 6120 41318 6134 41370
rect 6134 41318 6146 41370
rect 6146 41318 6176 41370
rect 6200 41318 6210 41370
rect 6210 41318 6256 41370
rect 5960 41316 6016 41318
rect 6040 41316 6096 41318
rect 6120 41316 6176 41318
rect 6200 41316 6256 41318
rect 4378 41080 4434 41136
rect 6696 40826 6752 40828
rect 6776 40826 6832 40828
rect 6856 40826 6912 40828
rect 6936 40826 6992 40828
rect 6696 40774 6742 40826
rect 6742 40774 6752 40826
rect 6776 40774 6806 40826
rect 6806 40774 6818 40826
rect 6818 40774 6832 40826
rect 6856 40774 6870 40826
rect 6870 40774 6882 40826
rect 6882 40774 6912 40826
rect 6936 40774 6946 40826
rect 6946 40774 6992 40826
rect 6696 40772 6752 40774
rect 6776 40772 6832 40774
rect 6856 40772 6912 40774
rect 6936 40772 6992 40774
rect 2906 40420 2962 40456
rect 2906 40400 2908 40420
rect 2908 40400 2960 40420
rect 2960 40400 2962 40420
rect 5960 40282 6016 40284
rect 6040 40282 6096 40284
rect 6120 40282 6176 40284
rect 6200 40282 6256 40284
rect 5960 40230 6006 40282
rect 6006 40230 6016 40282
rect 6040 40230 6070 40282
rect 6070 40230 6082 40282
rect 6082 40230 6096 40282
rect 6120 40230 6134 40282
rect 6134 40230 6146 40282
rect 6146 40230 6176 40282
rect 6200 40230 6210 40282
rect 6210 40230 6256 40282
rect 7138 40264 7194 40320
rect 5960 40228 6016 40230
rect 6040 40228 6096 40230
rect 6120 40228 6176 40230
rect 6200 40228 6256 40230
rect 6696 39738 6752 39740
rect 6776 39738 6832 39740
rect 6856 39738 6912 39740
rect 6936 39738 6992 39740
rect 6696 39686 6742 39738
rect 6742 39686 6752 39738
rect 6776 39686 6806 39738
rect 6806 39686 6818 39738
rect 6818 39686 6832 39738
rect 6856 39686 6870 39738
rect 6870 39686 6882 39738
rect 6882 39686 6912 39738
rect 6936 39686 6946 39738
rect 6946 39686 6992 39738
rect 6696 39684 6752 39686
rect 6776 39684 6832 39686
rect 6856 39684 6912 39686
rect 6936 39684 6992 39686
rect 5960 39194 6016 39196
rect 6040 39194 6096 39196
rect 6120 39194 6176 39196
rect 6200 39194 6256 39196
rect 5960 39142 6006 39194
rect 6006 39142 6016 39194
rect 6040 39142 6070 39194
rect 6070 39142 6082 39194
rect 6082 39142 6096 39194
rect 6120 39142 6134 39194
rect 6134 39142 6146 39194
rect 6146 39142 6176 39194
rect 6200 39142 6210 39194
rect 6210 39142 6256 39194
rect 7138 39176 7194 39232
rect 5960 39140 6016 39142
rect 6040 39140 6096 39142
rect 6120 39140 6176 39142
rect 6200 39140 6256 39142
rect 2906 39040 2962 39096
rect 6696 38650 6752 38652
rect 6776 38650 6832 38652
rect 6856 38650 6912 38652
rect 6936 38650 6992 38652
rect 6696 38598 6742 38650
rect 6742 38598 6752 38650
rect 6776 38598 6806 38650
rect 6806 38598 6818 38650
rect 6818 38598 6832 38650
rect 6856 38598 6870 38650
rect 6870 38598 6882 38650
rect 6882 38598 6912 38650
rect 6936 38598 6946 38650
rect 6946 38598 6992 38650
rect 6696 38596 6752 38598
rect 6776 38596 6832 38598
rect 6856 38596 6912 38598
rect 6936 38596 6992 38598
rect 4378 38360 4434 38416
rect 5960 38106 6016 38108
rect 6040 38106 6096 38108
rect 6120 38106 6176 38108
rect 6200 38106 6256 38108
rect 5960 38054 6006 38106
rect 6006 38054 6016 38106
rect 6040 38054 6070 38106
rect 6070 38054 6082 38106
rect 6082 38054 6096 38106
rect 6120 38054 6134 38106
rect 6134 38054 6146 38106
rect 6146 38054 6176 38106
rect 6200 38054 6210 38106
rect 6210 38054 6256 38106
rect 7782 38088 7838 38144
rect 5960 38052 6016 38054
rect 6040 38052 6096 38054
rect 6120 38052 6176 38054
rect 6200 38052 6256 38054
rect 6696 37562 6752 37564
rect 6776 37562 6832 37564
rect 6856 37562 6912 37564
rect 6936 37562 6992 37564
rect 6696 37510 6742 37562
rect 6742 37510 6752 37562
rect 6776 37510 6806 37562
rect 6806 37510 6818 37562
rect 6818 37510 6832 37562
rect 6856 37510 6870 37562
rect 6870 37510 6882 37562
rect 6882 37510 6912 37562
rect 6936 37510 6946 37562
rect 6946 37510 6992 37562
rect 6696 37508 6752 37510
rect 6776 37508 6832 37510
rect 6856 37508 6912 37510
rect 6936 37508 6992 37510
rect 2906 37000 2962 37056
rect 5960 37018 6016 37020
rect 6040 37018 6096 37020
rect 6120 37018 6176 37020
rect 6200 37018 6256 37020
rect 5960 36966 6006 37018
rect 6006 36966 6016 37018
rect 6040 36966 6070 37018
rect 6070 36966 6082 37018
rect 6082 36966 6096 37018
rect 6120 36966 6134 37018
rect 6134 36966 6146 37018
rect 6146 36966 6176 37018
rect 6200 36966 6210 37018
rect 6210 36966 6256 37018
rect 7230 37000 7286 37056
rect 5960 36964 6016 36966
rect 6040 36964 6096 36966
rect 6120 36964 6176 36966
rect 6200 36964 6256 36966
rect 6696 36474 6752 36476
rect 6776 36474 6832 36476
rect 6856 36474 6912 36476
rect 6936 36474 6992 36476
rect 6696 36422 6742 36474
rect 6742 36422 6752 36474
rect 6776 36422 6806 36474
rect 6806 36422 6818 36474
rect 6818 36422 6832 36474
rect 6856 36422 6870 36474
rect 6870 36422 6882 36474
rect 6882 36422 6912 36474
rect 6936 36422 6946 36474
rect 6946 36422 6992 36474
rect 6696 36420 6752 36422
rect 6776 36420 6832 36422
rect 6856 36420 6912 36422
rect 6936 36420 6992 36422
rect 5666 36048 5722 36104
rect 5960 35930 6016 35932
rect 6040 35930 6096 35932
rect 6120 35930 6176 35932
rect 6200 35930 6256 35932
rect 5960 35878 6006 35930
rect 6006 35878 6016 35930
rect 6040 35878 6070 35930
rect 6070 35878 6082 35930
rect 6082 35878 6096 35930
rect 6120 35878 6134 35930
rect 6134 35878 6146 35930
rect 6146 35878 6176 35930
rect 6200 35878 6210 35930
rect 6210 35878 6256 35930
rect 5960 35876 6016 35878
rect 6040 35876 6096 35878
rect 6120 35876 6176 35878
rect 6200 35876 6256 35878
rect 4378 35640 4434 35696
rect 6696 35386 6752 35388
rect 6776 35386 6832 35388
rect 6856 35386 6912 35388
rect 6936 35386 6992 35388
rect 6696 35334 6742 35386
rect 6742 35334 6752 35386
rect 6776 35334 6806 35386
rect 6806 35334 6818 35386
rect 6818 35334 6832 35386
rect 6856 35334 6870 35386
rect 6870 35334 6882 35386
rect 6882 35334 6912 35386
rect 6936 35334 6946 35386
rect 6946 35334 6992 35386
rect 6696 35332 6752 35334
rect 6776 35332 6832 35334
rect 6856 35332 6912 35334
rect 6936 35332 6992 35334
rect 2906 34980 2962 35016
rect 2906 34960 2908 34980
rect 2908 34960 2960 34980
rect 2960 34960 2962 34980
rect 5960 34842 6016 34844
rect 6040 34842 6096 34844
rect 6120 34842 6176 34844
rect 6200 34842 6256 34844
rect 5960 34790 6006 34842
rect 6006 34790 6016 34842
rect 6040 34790 6070 34842
rect 6070 34790 6082 34842
rect 6082 34790 6096 34842
rect 6120 34790 6134 34842
rect 6134 34790 6146 34842
rect 6146 34790 6176 34842
rect 6200 34790 6210 34842
rect 6210 34790 6256 34842
rect 7230 34824 7286 34880
rect 5960 34788 6016 34790
rect 6040 34788 6096 34790
rect 6120 34788 6176 34790
rect 6200 34788 6256 34790
rect 6696 34298 6752 34300
rect 6776 34298 6832 34300
rect 6856 34298 6912 34300
rect 6936 34298 6992 34300
rect 6696 34246 6742 34298
rect 6742 34246 6752 34298
rect 6776 34246 6806 34298
rect 6806 34246 6818 34298
rect 6818 34246 6832 34298
rect 6856 34246 6870 34298
rect 6870 34246 6882 34298
rect 6882 34246 6912 34298
rect 6936 34246 6946 34298
rect 6946 34246 6992 34298
rect 6696 34244 6752 34246
rect 6776 34244 6832 34246
rect 6856 34244 6912 34246
rect 6936 34244 6992 34246
rect 5960 33754 6016 33756
rect 6040 33754 6096 33756
rect 6120 33754 6176 33756
rect 6200 33754 6256 33756
rect 5960 33702 6006 33754
rect 6006 33702 6016 33754
rect 6040 33702 6070 33754
rect 6070 33702 6082 33754
rect 6082 33702 6096 33754
rect 6120 33702 6134 33754
rect 6134 33702 6146 33754
rect 6146 33702 6176 33754
rect 6200 33702 6210 33754
rect 6210 33702 6256 33754
rect 7230 33736 7286 33792
rect 5960 33700 6016 33702
rect 6040 33700 6096 33702
rect 6120 33700 6176 33702
rect 6200 33700 6256 33702
rect 2906 33600 2962 33656
rect 6696 33210 6752 33212
rect 6776 33210 6832 33212
rect 6856 33210 6912 33212
rect 6936 33210 6992 33212
rect 6696 33158 6742 33210
rect 6742 33158 6752 33210
rect 6776 33158 6806 33210
rect 6806 33158 6818 33210
rect 6818 33158 6832 33210
rect 6856 33158 6870 33210
rect 6870 33158 6882 33210
rect 6882 33158 6912 33210
rect 6936 33158 6946 33210
rect 6946 33158 6992 33210
rect 6696 33156 6752 33158
rect 6776 33156 6832 33158
rect 6856 33156 6912 33158
rect 6936 33156 6992 33158
rect 4378 32920 4434 32976
rect 5666 32920 5722 32976
rect 5960 32666 6016 32668
rect 6040 32666 6096 32668
rect 6120 32666 6176 32668
rect 6200 32666 6256 32668
rect 5960 32614 6006 32666
rect 6006 32614 6016 32666
rect 6040 32614 6070 32666
rect 6070 32614 6082 32666
rect 6082 32614 6096 32666
rect 6120 32614 6134 32666
rect 6134 32614 6146 32666
rect 6146 32614 6176 32666
rect 6200 32614 6210 32666
rect 6210 32614 6256 32666
rect 5960 32612 6016 32614
rect 6040 32612 6096 32614
rect 6120 32612 6176 32614
rect 6200 32612 6256 32614
rect 6696 32122 6752 32124
rect 6776 32122 6832 32124
rect 6856 32122 6912 32124
rect 6936 32122 6992 32124
rect 6696 32070 6742 32122
rect 6742 32070 6752 32122
rect 6776 32070 6806 32122
rect 6806 32070 6818 32122
rect 6818 32070 6832 32122
rect 6856 32070 6870 32122
rect 6870 32070 6882 32122
rect 6882 32070 6912 32122
rect 6936 32070 6946 32122
rect 6946 32070 6992 32122
rect 6696 32068 6752 32070
rect 6776 32068 6832 32070
rect 6856 32068 6912 32070
rect 6936 32068 6992 32070
rect 2906 31560 2962 31616
rect 5960 31578 6016 31580
rect 6040 31578 6096 31580
rect 6120 31578 6176 31580
rect 6200 31578 6256 31580
rect 5960 31526 6006 31578
rect 6006 31526 6016 31578
rect 6040 31526 6070 31578
rect 6070 31526 6082 31578
rect 6082 31526 6096 31578
rect 6120 31526 6134 31578
rect 6134 31526 6146 31578
rect 6146 31526 6176 31578
rect 6200 31526 6210 31578
rect 6210 31526 6256 31578
rect 7230 31560 7286 31616
rect 5960 31524 6016 31526
rect 6040 31524 6096 31526
rect 6120 31524 6176 31526
rect 6200 31524 6256 31526
rect 6696 31034 6752 31036
rect 6776 31034 6832 31036
rect 6856 31034 6912 31036
rect 6936 31034 6992 31036
rect 6696 30982 6742 31034
rect 6742 30982 6752 31034
rect 6776 30982 6806 31034
rect 6806 30982 6818 31034
rect 6818 30982 6832 31034
rect 6856 30982 6870 31034
rect 6870 30982 6882 31034
rect 6882 30982 6912 31034
rect 6936 30982 6946 31034
rect 6946 30982 6992 31034
rect 6696 30980 6752 30982
rect 6776 30980 6832 30982
rect 6856 30980 6912 30982
rect 6936 30980 6992 30982
rect 5960 30490 6016 30492
rect 6040 30490 6096 30492
rect 6120 30490 6176 30492
rect 6200 30490 6256 30492
rect 5960 30438 6006 30490
rect 6006 30438 6016 30490
rect 6040 30438 6070 30490
rect 6070 30438 6082 30490
rect 6082 30438 6096 30490
rect 6120 30438 6134 30490
rect 6134 30438 6146 30490
rect 6146 30438 6176 30490
rect 6200 30438 6210 30490
rect 6210 30438 6256 30490
rect 5960 30436 6016 30438
rect 6040 30436 6096 30438
rect 6120 30436 6176 30438
rect 6200 30436 6256 30438
rect 4378 30200 4434 30256
rect 5666 30200 5722 30256
rect 6696 29946 6752 29948
rect 6776 29946 6832 29948
rect 6856 29946 6912 29948
rect 6936 29946 6992 29948
rect 6696 29894 6742 29946
rect 6742 29894 6752 29946
rect 6776 29894 6806 29946
rect 6806 29894 6818 29946
rect 6818 29894 6832 29946
rect 6856 29894 6870 29946
rect 6870 29894 6882 29946
rect 6882 29894 6912 29946
rect 6936 29894 6946 29946
rect 6946 29894 6992 29946
rect 6696 29892 6752 29894
rect 6776 29892 6832 29894
rect 6856 29892 6912 29894
rect 6936 29892 6992 29894
rect 2906 29520 2962 29576
rect 5960 29402 6016 29404
rect 6040 29402 6096 29404
rect 6120 29402 6176 29404
rect 6200 29402 6256 29404
rect 5960 29350 6006 29402
rect 6006 29350 6016 29402
rect 6040 29350 6070 29402
rect 6070 29350 6082 29402
rect 6082 29350 6096 29402
rect 6120 29350 6134 29402
rect 6134 29350 6146 29402
rect 6146 29350 6176 29402
rect 6200 29350 6210 29402
rect 6210 29350 6256 29402
rect 7230 29384 7286 29440
rect 5960 29348 6016 29350
rect 6040 29348 6096 29350
rect 6120 29348 6176 29350
rect 6200 29348 6256 29350
rect 6696 28858 6752 28860
rect 6776 28858 6832 28860
rect 6856 28858 6912 28860
rect 6936 28858 6992 28860
rect 6696 28806 6742 28858
rect 6742 28806 6752 28858
rect 6776 28806 6806 28858
rect 6806 28806 6818 28858
rect 6818 28806 6832 28858
rect 6856 28806 6870 28858
rect 6870 28806 6882 28858
rect 6882 28806 6912 28858
rect 6936 28806 6946 28858
rect 6946 28806 6992 28858
rect 6696 28804 6752 28806
rect 6776 28804 6832 28806
rect 6856 28804 6912 28806
rect 6936 28804 6992 28806
rect 5960 28314 6016 28316
rect 6040 28314 6096 28316
rect 6120 28314 6176 28316
rect 6200 28314 6256 28316
rect 5960 28262 6006 28314
rect 6006 28262 6016 28314
rect 6040 28262 6070 28314
rect 6070 28262 6082 28314
rect 6082 28262 6096 28314
rect 6120 28262 6134 28314
rect 6134 28262 6146 28314
rect 6146 28262 6176 28314
rect 6200 28262 6210 28314
rect 6210 28262 6256 28314
rect 7230 28296 7286 28352
rect 5960 28260 6016 28262
rect 6040 28260 6096 28262
rect 6120 28260 6176 28262
rect 6200 28260 6256 28262
rect 2906 28160 2962 28216
rect 6696 27770 6752 27772
rect 6776 27770 6832 27772
rect 6856 27770 6912 27772
rect 6936 27770 6992 27772
rect 6696 27718 6742 27770
rect 6742 27718 6752 27770
rect 6776 27718 6806 27770
rect 6806 27718 6818 27770
rect 6818 27718 6832 27770
rect 6856 27718 6870 27770
rect 6870 27718 6882 27770
rect 6882 27718 6912 27770
rect 6936 27718 6946 27770
rect 6946 27718 6992 27770
rect 6696 27716 6752 27718
rect 6776 27716 6832 27718
rect 6856 27716 6912 27718
rect 6936 27716 6992 27718
rect 5114 27480 5170 27536
rect 5390 27480 5446 27536
rect 5960 27226 6016 27228
rect 6040 27226 6096 27228
rect 6120 27226 6176 27228
rect 6200 27226 6256 27228
rect 5960 27174 6006 27226
rect 6006 27174 6016 27226
rect 6040 27174 6070 27226
rect 6070 27174 6082 27226
rect 6082 27174 6096 27226
rect 6120 27174 6134 27226
rect 6134 27174 6146 27226
rect 6146 27174 6176 27226
rect 6200 27174 6210 27226
rect 6210 27174 6256 27226
rect 5960 27172 6016 27174
rect 6040 27172 6096 27174
rect 6120 27172 6176 27174
rect 6200 27172 6256 27174
rect 6696 26682 6752 26684
rect 6776 26682 6832 26684
rect 6856 26682 6912 26684
rect 6936 26682 6992 26684
rect 6696 26630 6742 26682
rect 6742 26630 6752 26682
rect 6776 26630 6806 26682
rect 6806 26630 6818 26682
rect 6818 26630 6832 26682
rect 6856 26630 6870 26682
rect 6870 26630 6882 26682
rect 6882 26630 6912 26682
rect 6936 26630 6946 26682
rect 6946 26630 6992 26682
rect 6696 26628 6752 26630
rect 6776 26628 6832 26630
rect 6856 26628 6912 26630
rect 6936 26628 6992 26630
rect 2906 26120 2962 26176
rect 5960 26138 6016 26140
rect 6040 26138 6096 26140
rect 6120 26138 6176 26140
rect 6200 26138 6256 26140
rect 5960 26086 6006 26138
rect 6006 26086 6016 26138
rect 6040 26086 6070 26138
rect 6070 26086 6082 26138
rect 6082 26086 6096 26138
rect 6120 26086 6134 26138
rect 6134 26086 6146 26138
rect 6146 26086 6176 26138
rect 6200 26086 6210 26138
rect 6210 26086 6256 26138
rect 7138 26120 7194 26176
rect 5960 26084 6016 26086
rect 6040 26084 6096 26086
rect 6120 26084 6176 26086
rect 6200 26084 6256 26086
rect 6696 25594 6752 25596
rect 6776 25594 6832 25596
rect 6856 25594 6912 25596
rect 6936 25594 6992 25596
rect 6696 25542 6742 25594
rect 6742 25542 6752 25594
rect 6776 25542 6806 25594
rect 6806 25542 6818 25594
rect 6818 25542 6832 25594
rect 6856 25542 6870 25594
rect 6870 25542 6882 25594
rect 6882 25542 6912 25594
rect 6936 25542 6946 25594
rect 6946 25542 6992 25594
rect 6696 25540 6752 25542
rect 6776 25540 6832 25542
rect 6856 25540 6912 25542
rect 6936 25540 6992 25542
rect 5960 25050 6016 25052
rect 6040 25050 6096 25052
rect 6120 25050 6176 25052
rect 6200 25050 6256 25052
rect 5960 24998 6006 25050
rect 6006 24998 6016 25050
rect 6040 24998 6070 25050
rect 6070 24998 6082 25050
rect 6082 24998 6096 25050
rect 6120 24998 6134 25050
rect 6134 24998 6146 25050
rect 6146 24998 6176 25050
rect 6200 24998 6210 25050
rect 6210 24998 6256 25050
rect 7138 25032 7194 25088
rect 5960 24996 6016 24998
rect 6040 24996 6096 24998
rect 6120 24996 6176 24998
rect 6200 24996 6256 24998
rect 4930 24760 4986 24816
rect 6696 24506 6752 24508
rect 6776 24506 6832 24508
rect 6856 24506 6912 24508
rect 6936 24506 6992 24508
rect 6696 24454 6742 24506
rect 6742 24454 6752 24506
rect 6776 24454 6806 24506
rect 6806 24454 6818 24506
rect 6818 24454 6832 24506
rect 6856 24454 6870 24506
rect 6870 24454 6882 24506
rect 6882 24454 6912 24506
rect 6936 24454 6946 24506
rect 6946 24454 6992 24506
rect 6696 24452 6752 24454
rect 6776 24452 6832 24454
rect 6856 24452 6912 24454
rect 6936 24452 6992 24454
rect 2906 24080 2962 24136
rect 5960 23962 6016 23964
rect 6040 23962 6096 23964
rect 6120 23962 6176 23964
rect 6200 23962 6256 23964
rect 5960 23910 6006 23962
rect 6006 23910 6016 23962
rect 6040 23910 6070 23962
rect 6070 23910 6082 23962
rect 6082 23910 6096 23962
rect 6120 23910 6134 23962
rect 6134 23910 6146 23962
rect 6146 23910 6176 23962
rect 6200 23910 6210 23962
rect 6210 23910 6256 23962
rect 7138 23944 7194 24000
rect 5960 23908 6016 23910
rect 6040 23908 6096 23910
rect 6120 23908 6176 23910
rect 6200 23908 6256 23910
rect 6696 23418 6752 23420
rect 6776 23418 6832 23420
rect 6856 23418 6912 23420
rect 6936 23418 6992 23420
rect 6696 23366 6742 23418
rect 6742 23366 6752 23418
rect 6776 23366 6806 23418
rect 6806 23366 6818 23418
rect 6818 23366 6832 23418
rect 6856 23366 6870 23418
rect 6870 23366 6882 23418
rect 6882 23366 6912 23418
rect 6936 23366 6946 23418
rect 6946 23366 6992 23418
rect 6696 23364 6752 23366
rect 6776 23364 6832 23366
rect 6856 23364 6912 23366
rect 6936 23364 6992 23366
rect 5960 22874 6016 22876
rect 6040 22874 6096 22876
rect 6120 22874 6176 22876
rect 6200 22874 6256 22876
rect 5960 22822 6006 22874
rect 6006 22822 6016 22874
rect 6040 22822 6070 22874
rect 6070 22822 6082 22874
rect 6082 22822 6096 22874
rect 6120 22822 6134 22874
rect 6134 22822 6146 22874
rect 6146 22822 6176 22874
rect 6200 22822 6210 22874
rect 6210 22822 6256 22874
rect 7138 22856 7194 22912
rect 5960 22820 6016 22822
rect 6040 22820 6096 22822
rect 6120 22820 6176 22822
rect 6200 22820 6256 22822
rect 2906 22720 2962 22776
rect 6696 22330 6752 22332
rect 6776 22330 6832 22332
rect 6856 22330 6912 22332
rect 6936 22330 6992 22332
rect 6696 22278 6742 22330
rect 6742 22278 6752 22330
rect 6776 22278 6806 22330
rect 6806 22278 6818 22330
rect 6818 22278 6832 22330
rect 6856 22278 6870 22330
rect 6870 22278 6882 22330
rect 6882 22278 6912 22330
rect 6936 22278 6946 22330
rect 6946 22278 6992 22330
rect 6696 22276 6752 22278
rect 6776 22276 6832 22278
rect 6856 22276 6912 22278
rect 6936 22276 6992 22278
rect 4930 22040 4986 22096
rect 5960 21786 6016 21788
rect 6040 21786 6096 21788
rect 6120 21786 6176 21788
rect 6200 21786 6256 21788
rect 5960 21734 6006 21786
rect 6006 21734 6016 21786
rect 6040 21734 6070 21786
rect 6070 21734 6082 21786
rect 6082 21734 6096 21786
rect 6120 21734 6134 21786
rect 6134 21734 6146 21786
rect 6146 21734 6176 21786
rect 6200 21734 6210 21786
rect 6210 21734 6256 21786
rect 9162 21768 9218 21824
rect 5960 21732 6016 21734
rect 6040 21732 6096 21734
rect 6120 21732 6176 21734
rect 6200 21732 6256 21734
rect 6696 21242 6752 21244
rect 6776 21242 6832 21244
rect 6856 21242 6912 21244
rect 6936 21242 6992 21244
rect 6696 21190 6742 21242
rect 6742 21190 6752 21242
rect 6776 21190 6806 21242
rect 6806 21190 6818 21242
rect 6818 21190 6832 21242
rect 6856 21190 6870 21242
rect 6870 21190 6882 21242
rect 6882 21190 6912 21242
rect 6936 21190 6946 21242
rect 6946 21190 6992 21242
rect 6696 21188 6752 21190
rect 6776 21188 6832 21190
rect 6856 21188 6912 21190
rect 6936 21188 6992 21190
rect 5206 20680 5262 20736
rect 5960 20698 6016 20700
rect 6040 20698 6096 20700
rect 6120 20698 6176 20700
rect 6200 20698 6256 20700
rect 5960 20646 6006 20698
rect 6006 20646 6016 20698
rect 6040 20646 6070 20698
rect 6070 20646 6082 20698
rect 6082 20646 6096 20698
rect 6120 20646 6134 20698
rect 6134 20646 6146 20698
rect 6146 20646 6176 20698
rect 6200 20646 6210 20698
rect 6210 20646 6256 20698
rect 9254 20680 9310 20736
rect 5960 20644 6016 20646
rect 6040 20644 6096 20646
rect 6120 20644 6176 20646
rect 6200 20644 6256 20646
rect 6696 20154 6752 20156
rect 6776 20154 6832 20156
rect 6856 20154 6912 20156
rect 6936 20154 6992 20156
rect 6696 20102 6742 20154
rect 6742 20102 6752 20154
rect 6776 20102 6806 20154
rect 6806 20102 6818 20154
rect 6818 20102 6832 20154
rect 6856 20102 6870 20154
rect 6870 20102 6882 20154
rect 6882 20102 6912 20154
rect 6936 20102 6946 20154
rect 6946 20102 6992 20154
rect 6696 20100 6752 20102
rect 6776 20100 6832 20102
rect 6856 20100 6912 20102
rect 6936 20100 6992 20102
rect 5960 19610 6016 19612
rect 6040 19610 6096 19612
rect 6120 19610 6176 19612
rect 6200 19610 6256 19612
rect 5960 19558 6006 19610
rect 6006 19558 6016 19610
rect 6040 19558 6070 19610
rect 6070 19558 6082 19610
rect 6082 19558 6096 19610
rect 6120 19558 6134 19610
rect 6134 19558 6146 19610
rect 6146 19558 6176 19610
rect 6200 19558 6210 19610
rect 6210 19558 6256 19610
rect 7138 19592 7194 19648
rect 5960 19556 6016 19558
rect 6040 19556 6096 19558
rect 6120 19556 6176 19558
rect 6200 19556 6256 19558
rect 4930 19320 4986 19376
rect 6696 19066 6752 19068
rect 6776 19066 6832 19068
rect 6856 19066 6912 19068
rect 6936 19066 6992 19068
rect 6696 19014 6742 19066
rect 6742 19014 6752 19066
rect 6776 19014 6806 19066
rect 6806 19014 6818 19066
rect 6818 19014 6832 19066
rect 6856 19014 6870 19066
rect 6870 19014 6882 19066
rect 6882 19014 6912 19066
rect 6936 19014 6946 19066
rect 6946 19014 6992 19066
rect 6696 19012 6752 19014
rect 6776 19012 6832 19014
rect 6856 19012 6912 19014
rect 6936 19012 6992 19014
rect 2906 18640 2962 18696
rect 5960 18522 6016 18524
rect 6040 18522 6096 18524
rect 6120 18522 6176 18524
rect 6200 18522 6256 18524
rect 5960 18470 6006 18522
rect 6006 18470 6016 18522
rect 6040 18470 6070 18522
rect 6070 18470 6082 18522
rect 6082 18470 6096 18522
rect 6120 18470 6134 18522
rect 6134 18470 6146 18522
rect 6146 18470 6176 18522
rect 6200 18470 6210 18522
rect 6210 18470 6256 18522
rect 7138 18504 7194 18560
rect 5960 18468 6016 18470
rect 6040 18468 6096 18470
rect 6120 18468 6176 18470
rect 6200 18468 6256 18470
rect 6696 17978 6752 17980
rect 6776 17978 6832 17980
rect 6856 17978 6912 17980
rect 6936 17978 6992 17980
rect 6696 17926 6742 17978
rect 6742 17926 6752 17978
rect 6776 17926 6806 17978
rect 6806 17926 6818 17978
rect 6818 17926 6832 17978
rect 6856 17926 6870 17978
rect 6870 17926 6882 17978
rect 6882 17926 6912 17978
rect 6936 17926 6946 17978
rect 6946 17926 6992 17978
rect 6696 17924 6752 17926
rect 6776 17924 6832 17926
rect 6856 17924 6912 17926
rect 6936 17924 6992 17926
rect 5960 17434 6016 17436
rect 6040 17434 6096 17436
rect 6120 17434 6176 17436
rect 6200 17434 6256 17436
rect 5960 17382 6006 17434
rect 6006 17382 6016 17434
rect 6040 17382 6070 17434
rect 6070 17382 6082 17434
rect 6082 17382 6096 17434
rect 6120 17382 6134 17434
rect 6134 17382 6146 17434
rect 6146 17382 6176 17434
rect 6200 17382 6210 17434
rect 6210 17382 6256 17434
rect 7230 17416 7286 17472
rect 5960 17380 6016 17382
rect 6040 17380 6096 17382
rect 6120 17380 6176 17382
rect 6200 17380 6256 17382
rect 2906 17280 2962 17336
rect 6696 16890 6752 16892
rect 6776 16890 6832 16892
rect 6856 16890 6912 16892
rect 6936 16890 6992 16892
rect 6696 16838 6742 16890
rect 6742 16838 6752 16890
rect 6776 16838 6806 16890
rect 6806 16838 6818 16890
rect 6818 16838 6832 16890
rect 6856 16838 6870 16890
rect 6870 16838 6882 16890
rect 6882 16838 6912 16890
rect 6936 16838 6946 16890
rect 6946 16838 6992 16890
rect 6696 16836 6752 16838
rect 6776 16836 6832 16838
rect 6856 16836 6912 16838
rect 6936 16836 6992 16838
rect 5206 16600 5262 16656
rect 5390 16600 5446 16656
rect 5960 16346 6016 16348
rect 6040 16346 6096 16348
rect 6120 16346 6176 16348
rect 6200 16346 6256 16348
rect 5960 16294 6006 16346
rect 6006 16294 6016 16346
rect 6040 16294 6070 16346
rect 6070 16294 6082 16346
rect 6082 16294 6096 16346
rect 6120 16294 6134 16346
rect 6134 16294 6146 16346
rect 6146 16294 6176 16346
rect 6200 16294 6210 16346
rect 6210 16294 6256 16346
rect 5960 16292 6016 16294
rect 6040 16292 6096 16294
rect 6120 16292 6176 16294
rect 6200 16292 6256 16294
rect 6696 15802 6752 15804
rect 6776 15802 6832 15804
rect 6856 15802 6912 15804
rect 6936 15802 6992 15804
rect 6696 15750 6742 15802
rect 6742 15750 6752 15802
rect 6776 15750 6806 15802
rect 6806 15750 6818 15802
rect 6818 15750 6832 15802
rect 6856 15750 6870 15802
rect 6870 15750 6882 15802
rect 6882 15750 6912 15802
rect 6936 15750 6946 15802
rect 6946 15750 6992 15802
rect 6696 15748 6752 15750
rect 6776 15748 6832 15750
rect 6856 15748 6912 15750
rect 6936 15748 6992 15750
rect 5206 15240 5262 15296
rect 5960 15258 6016 15260
rect 6040 15258 6096 15260
rect 6120 15258 6176 15260
rect 6200 15258 6256 15260
rect 5960 15206 6006 15258
rect 6006 15206 6016 15258
rect 6040 15206 6070 15258
rect 6070 15206 6082 15258
rect 6082 15206 6096 15258
rect 6120 15206 6134 15258
rect 6134 15206 6146 15258
rect 6146 15206 6176 15258
rect 6200 15206 6210 15258
rect 6210 15206 6256 15258
rect 5960 15204 6016 15206
rect 6040 15204 6096 15206
rect 6120 15204 6176 15206
rect 6200 15204 6256 15206
rect 5666 14968 5722 15024
rect 6696 14714 6752 14716
rect 6776 14714 6832 14716
rect 6856 14714 6912 14716
rect 6936 14714 6992 14716
rect 6696 14662 6742 14714
rect 6742 14662 6752 14714
rect 6776 14662 6806 14714
rect 6806 14662 6818 14714
rect 6818 14662 6832 14714
rect 6856 14662 6870 14714
rect 6870 14662 6882 14714
rect 6882 14662 6912 14714
rect 6936 14662 6946 14714
rect 6946 14662 6992 14714
rect 6696 14660 6752 14662
rect 6776 14660 6832 14662
rect 6856 14660 6912 14662
rect 6936 14660 6992 14662
rect 5960 14170 6016 14172
rect 6040 14170 6096 14172
rect 6120 14170 6176 14172
rect 6200 14170 6256 14172
rect 5960 14118 6006 14170
rect 6006 14118 6016 14170
rect 6040 14118 6070 14170
rect 6070 14118 6082 14170
rect 6082 14118 6096 14170
rect 6120 14118 6134 14170
rect 6134 14118 6146 14170
rect 6146 14118 6176 14170
rect 6200 14118 6210 14170
rect 6210 14118 6256 14170
rect 5960 14116 6016 14118
rect 6040 14116 6096 14118
rect 6120 14116 6176 14118
rect 6200 14116 6256 14118
rect 6696 13626 6752 13628
rect 6776 13626 6832 13628
rect 6856 13626 6912 13628
rect 6936 13626 6992 13628
rect 6696 13574 6742 13626
rect 6742 13574 6752 13626
rect 6776 13574 6806 13626
rect 6806 13574 6818 13626
rect 6818 13574 6832 13626
rect 6856 13574 6870 13626
rect 6870 13574 6882 13626
rect 6882 13574 6912 13626
rect 6936 13574 6946 13626
rect 6946 13574 6992 13626
rect 6696 13572 6752 13574
rect 6776 13572 6832 13574
rect 6856 13572 6912 13574
rect 6936 13572 6992 13574
rect 46054 48356 46110 48412
rect 45962 14120 46018 14176
rect 5960 13082 6016 13084
rect 6040 13082 6096 13084
rect 6120 13082 6176 13084
rect 6200 13082 6256 13084
rect 5960 13030 6006 13082
rect 6006 13030 6016 13082
rect 6040 13030 6070 13082
rect 6070 13030 6082 13082
rect 6082 13030 6096 13082
rect 6120 13030 6134 13082
rect 6134 13030 6146 13082
rect 6146 13030 6176 13082
rect 6200 13030 6210 13082
rect 6210 13030 6256 13082
rect 5960 13028 6016 13030
rect 6040 13028 6096 13030
rect 6120 13028 6176 13030
rect 6200 13028 6256 13030
rect 45870 13032 45926 13088
rect 6696 12538 6752 12540
rect 6776 12538 6832 12540
rect 6856 12538 6912 12540
rect 6936 12538 6992 12540
rect 6696 12486 6742 12538
rect 6742 12486 6752 12538
rect 6776 12486 6806 12538
rect 6806 12486 6818 12538
rect 6818 12486 6832 12538
rect 6856 12486 6870 12538
rect 6870 12486 6882 12538
rect 6882 12486 6912 12538
rect 6936 12486 6946 12538
rect 6946 12486 6992 12538
rect 6696 12484 6752 12486
rect 6776 12484 6832 12486
rect 6856 12484 6912 12486
rect 6936 12484 6992 12486
rect 5960 11994 6016 11996
rect 6040 11994 6096 11996
rect 6120 11994 6176 11996
rect 6200 11994 6256 11996
rect 5960 11942 6006 11994
rect 6006 11942 6016 11994
rect 6040 11942 6070 11994
rect 6070 11942 6082 11994
rect 6082 11942 6096 11994
rect 6120 11942 6134 11994
rect 6134 11942 6146 11994
rect 6146 11942 6176 11994
rect 6200 11942 6210 11994
rect 6210 11942 6256 11994
rect 5960 11940 6016 11942
rect 6040 11940 6096 11942
rect 6120 11940 6176 11942
rect 6200 11940 6256 11942
rect 6696 11450 6752 11452
rect 6776 11450 6832 11452
rect 6856 11450 6912 11452
rect 6936 11450 6992 11452
rect 6696 11398 6742 11450
rect 6742 11398 6752 11450
rect 6776 11398 6806 11450
rect 6806 11398 6818 11450
rect 6818 11398 6832 11450
rect 6856 11398 6870 11450
rect 6870 11398 6882 11450
rect 6882 11398 6912 11450
rect 6936 11398 6946 11450
rect 6946 11398 6992 11450
rect 6696 11396 6752 11398
rect 6776 11396 6832 11398
rect 6856 11396 6912 11398
rect 6936 11396 6992 11398
rect 5960 10906 6016 10908
rect 6040 10906 6096 10908
rect 6120 10906 6176 10908
rect 6200 10906 6256 10908
rect 5960 10854 6006 10906
rect 6006 10854 6016 10906
rect 6040 10854 6070 10906
rect 6070 10854 6082 10906
rect 6082 10854 6096 10906
rect 6120 10854 6134 10906
rect 6134 10854 6146 10906
rect 6146 10854 6176 10906
rect 6200 10854 6210 10906
rect 6210 10854 6256 10906
rect 5960 10852 6016 10854
rect 6040 10852 6096 10854
rect 6120 10852 6176 10854
rect 6200 10852 6256 10854
rect 45870 10820 45926 10876
rect 6696 10362 6752 10364
rect 6776 10362 6832 10364
rect 6856 10362 6912 10364
rect 6936 10362 6992 10364
rect 6696 10310 6742 10362
rect 6742 10310 6752 10362
rect 6776 10310 6806 10362
rect 6806 10310 6818 10362
rect 6818 10310 6832 10362
rect 6856 10310 6870 10362
rect 6870 10310 6882 10362
rect 6882 10310 6912 10362
rect 6936 10310 6946 10362
rect 6946 10310 6992 10362
rect 6696 10308 6752 10310
rect 6776 10308 6832 10310
rect 6856 10308 6912 10310
rect 6936 10308 6992 10310
rect 5960 9818 6016 9820
rect 6040 9818 6096 9820
rect 6120 9818 6176 9820
rect 6200 9818 6256 9820
rect 5960 9766 6006 9818
rect 6006 9766 6016 9818
rect 6040 9766 6070 9818
rect 6070 9766 6082 9818
rect 6082 9766 6096 9818
rect 6120 9766 6134 9818
rect 6134 9766 6146 9818
rect 6146 9766 6176 9818
rect 6200 9766 6210 9818
rect 6210 9766 6256 9818
rect 5960 9764 6016 9766
rect 6040 9764 6096 9766
rect 6120 9764 6176 9766
rect 6200 9764 6256 9766
rect 6696 9274 6752 9276
rect 6776 9274 6832 9276
rect 6856 9274 6912 9276
rect 6936 9274 6992 9276
rect 6696 9222 6742 9274
rect 6742 9222 6752 9274
rect 6776 9222 6806 9274
rect 6806 9222 6818 9274
rect 6818 9222 6832 9274
rect 6856 9222 6870 9274
rect 6870 9222 6882 9274
rect 6882 9222 6912 9274
rect 6936 9222 6946 9274
rect 6946 9222 6992 9274
rect 6696 9220 6752 9222
rect 6776 9220 6832 9222
rect 6856 9220 6912 9222
rect 6936 9220 6992 9222
rect 5960 8730 6016 8732
rect 6040 8730 6096 8732
rect 6120 8730 6176 8732
rect 6200 8730 6256 8732
rect 5960 8678 6006 8730
rect 6006 8678 6016 8730
rect 6040 8678 6070 8730
rect 6070 8678 6082 8730
rect 6082 8678 6096 8730
rect 6120 8678 6134 8730
rect 6134 8678 6146 8730
rect 6146 8678 6176 8730
rect 6200 8678 6210 8730
rect 6210 8678 6256 8730
rect 5960 8676 6016 8678
rect 6040 8676 6096 8678
rect 6120 8676 6176 8678
rect 6200 8676 6256 8678
rect 6696 8186 6752 8188
rect 6776 8186 6832 8188
rect 6856 8186 6912 8188
rect 6936 8186 6992 8188
rect 6696 8134 6742 8186
rect 6742 8134 6752 8186
rect 6776 8134 6806 8186
rect 6806 8134 6818 8186
rect 6818 8134 6832 8186
rect 6856 8134 6870 8186
rect 6870 8134 6882 8186
rect 6882 8134 6912 8186
rect 6936 8134 6946 8186
rect 6946 8134 6992 8186
rect 6696 8132 6752 8134
rect 6776 8132 6832 8134
rect 6856 8132 6912 8134
rect 6936 8132 6992 8134
rect 5960 7642 6016 7644
rect 6040 7642 6096 7644
rect 6120 7642 6176 7644
rect 6200 7642 6256 7644
rect 5960 7590 6006 7642
rect 6006 7590 6016 7642
rect 6040 7590 6070 7642
rect 6070 7590 6082 7642
rect 6082 7590 6096 7642
rect 6120 7590 6134 7642
rect 6134 7590 6146 7642
rect 6146 7590 6176 7642
rect 6200 7590 6210 7642
rect 6210 7590 6256 7642
rect 5960 7588 6016 7590
rect 6040 7588 6096 7590
rect 6120 7588 6176 7590
rect 6200 7588 6256 7590
rect 6696 7098 6752 7100
rect 6776 7098 6832 7100
rect 6856 7098 6912 7100
rect 6936 7098 6992 7100
rect 6696 7046 6742 7098
rect 6742 7046 6752 7098
rect 6776 7046 6806 7098
rect 6806 7046 6818 7098
rect 6818 7046 6832 7098
rect 6856 7046 6870 7098
rect 6870 7046 6882 7098
rect 6882 7046 6912 7098
rect 6936 7046 6946 7098
rect 6946 7046 6992 7098
rect 6696 7044 6752 7046
rect 6776 7044 6832 7046
rect 6856 7044 6912 7046
rect 6936 7044 6992 7046
rect 17728 7642 17784 7644
rect 17808 7642 17864 7644
rect 17888 7642 17944 7644
rect 17968 7642 18024 7644
rect 17728 7590 17774 7642
rect 17774 7590 17784 7642
rect 17808 7590 17838 7642
rect 17838 7590 17850 7642
rect 17850 7590 17864 7642
rect 17888 7590 17902 7642
rect 17902 7590 17914 7642
rect 17914 7590 17944 7642
rect 17968 7590 17978 7642
rect 17978 7590 18024 7642
rect 17728 7588 17784 7590
rect 17808 7588 17864 7590
rect 17888 7588 17944 7590
rect 17968 7588 18024 7590
rect 17728 6554 17784 6556
rect 17808 6554 17864 6556
rect 17888 6554 17944 6556
rect 17968 6554 18024 6556
rect 17728 6502 17774 6554
rect 17774 6502 17784 6554
rect 17808 6502 17838 6554
rect 17838 6502 17850 6554
rect 17850 6502 17864 6554
rect 17888 6502 17902 6554
rect 17902 6502 17914 6554
rect 17914 6502 17944 6554
rect 17968 6502 17978 6554
rect 17978 6502 18024 6554
rect 17728 6500 17784 6502
rect 17808 6500 17864 6502
rect 17888 6500 17944 6502
rect 17968 6500 18024 6502
rect 17728 5466 17784 5468
rect 17808 5466 17864 5468
rect 17888 5466 17944 5468
rect 17968 5466 18024 5468
rect 17728 5414 17774 5466
rect 17774 5414 17784 5466
rect 17808 5414 17838 5466
rect 17838 5414 17850 5466
rect 17850 5414 17864 5466
rect 17888 5414 17902 5466
rect 17902 5414 17914 5466
rect 17914 5414 17944 5466
rect 17968 5414 17978 5466
rect 17978 5414 18024 5466
rect 17728 5412 17784 5414
rect 17808 5412 17864 5414
rect 17888 5412 17944 5414
rect 17968 5412 18024 5414
rect 18388 7098 18444 7100
rect 18468 7098 18524 7100
rect 18548 7098 18604 7100
rect 18628 7098 18684 7100
rect 18388 7046 18434 7098
rect 18434 7046 18444 7098
rect 18468 7046 18498 7098
rect 18498 7046 18510 7098
rect 18510 7046 18524 7098
rect 18548 7046 18562 7098
rect 18562 7046 18574 7098
rect 18574 7046 18604 7098
rect 18628 7046 18638 7098
rect 18638 7046 18684 7098
rect 18388 7044 18444 7046
rect 18468 7044 18524 7046
rect 18548 7044 18604 7046
rect 18628 7044 18684 7046
rect 18388 6010 18444 6012
rect 18468 6010 18524 6012
rect 18548 6010 18604 6012
rect 18628 6010 18684 6012
rect 18388 5958 18434 6010
rect 18434 5958 18444 6010
rect 18468 5958 18498 6010
rect 18498 5958 18510 6010
rect 18510 5958 18524 6010
rect 18548 5958 18562 6010
rect 18562 5958 18574 6010
rect 18574 5958 18604 6010
rect 18628 5958 18638 6010
rect 18638 5958 18684 6010
rect 18388 5956 18444 5958
rect 18468 5956 18524 5958
rect 18548 5956 18604 5958
rect 18628 5956 18684 5958
rect 36128 7642 36184 7644
rect 36208 7642 36264 7644
rect 36288 7642 36344 7644
rect 36368 7642 36424 7644
rect 36128 7590 36174 7642
rect 36174 7590 36184 7642
rect 36208 7590 36238 7642
rect 36238 7590 36250 7642
rect 36250 7590 36264 7642
rect 36288 7590 36302 7642
rect 36302 7590 36314 7642
rect 36314 7590 36344 7642
rect 36368 7590 36378 7642
rect 36378 7590 36424 7642
rect 36128 7588 36184 7590
rect 36208 7588 36264 7590
rect 36288 7588 36344 7590
rect 36368 7588 36424 7590
rect 36788 7098 36844 7100
rect 36868 7098 36924 7100
rect 36948 7098 37004 7100
rect 37028 7098 37084 7100
rect 36788 7046 36834 7098
rect 36834 7046 36844 7098
rect 36868 7046 36898 7098
rect 36898 7046 36910 7098
rect 36910 7046 36924 7098
rect 36948 7046 36962 7098
rect 36962 7046 36974 7098
rect 36974 7046 37004 7098
rect 37028 7046 37038 7098
rect 37038 7046 37084 7098
rect 36788 7044 36844 7046
rect 36868 7044 36924 7046
rect 36948 7044 37004 7046
rect 37028 7044 37084 7046
rect 36128 6554 36184 6556
rect 36208 6554 36264 6556
rect 36288 6554 36344 6556
rect 36368 6554 36424 6556
rect 36128 6502 36174 6554
rect 36174 6502 36184 6554
rect 36208 6502 36238 6554
rect 36238 6502 36250 6554
rect 36250 6502 36264 6554
rect 36288 6502 36302 6554
rect 36302 6502 36314 6554
rect 36314 6502 36344 6554
rect 36368 6502 36378 6554
rect 36378 6502 36424 6554
rect 36128 6500 36184 6502
rect 36208 6500 36264 6502
rect 36288 6500 36344 6502
rect 36368 6500 36424 6502
rect 36788 6010 36844 6012
rect 36868 6010 36924 6012
rect 36948 6010 37004 6012
rect 37028 6010 37084 6012
rect 36788 5958 36834 6010
rect 36834 5958 36844 6010
rect 36868 5958 36898 6010
rect 36898 5958 36910 6010
rect 36910 5958 36924 6010
rect 36948 5958 36962 6010
rect 36962 5958 36974 6010
rect 36974 5958 37004 6010
rect 37028 5958 37038 6010
rect 37038 5958 37084 6010
rect 36788 5956 36844 5958
rect 36868 5956 36924 5958
rect 36948 5956 37004 5958
rect 37028 5956 37084 5958
rect 36128 5466 36184 5468
rect 36208 5466 36264 5468
rect 36288 5466 36344 5468
rect 36368 5466 36424 5468
rect 36128 5414 36174 5466
rect 36174 5414 36184 5466
rect 36208 5414 36238 5466
rect 36238 5414 36250 5466
rect 36250 5414 36264 5466
rect 36288 5414 36302 5466
rect 36302 5414 36314 5466
rect 36314 5414 36344 5466
rect 36368 5414 36378 5466
rect 36378 5414 36424 5466
rect 36128 5412 36184 5414
rect 36208 5412 36264 5414
rect 36288 5412 36344 5414
rect 36368 5412 36424 5414
rect 46146 47268 46202 47324
rect 46146 13032 46202 13088
rect 46054 11944 46110 12000
rect 54528 87066 54584 87068
rect 54608 87066 54664 87068
rect 54688 87066 54744 87068
rect 54768 87066 54824 87068
rect 54528 87014 54574 87066
rect 54574 87014 54584 87066
rect 54608 87014 54638 87066
rect 54638 87014 54650 87066
rect 54650 87014 54664 87066
rect 54688 87014 54702 87066
rect 54702 87014 54714 87066
rect 54714 87014 54744 87066
rect 54768 87014 54778 87066
rect 54778 87014 54824 87066
rect 54528 87012 54584 87014
rect 54608 87012 54664 87014
rect 54688 87012 54744 87014
rect 54768 87012 54824 87014
rect 55188 86522 55244 86524
rect 55268 86522 55324 86524
rect 55348 86522 55404 86524
rect 55428 86522 55484 86524
rect 55188 86470 55234 86522
rect 55234 86470 55244 86522
rect 55268 86470 55298 86522
rect 55298 86470 55310 86522
rect 55310 86470 55324 86522
rect 55348 86470 55362 86522
rect 55362 86470 55374 86522
rect 55374 86470 55404 86522
rect 55428 86470 55438 86522
rect 55438 86470 55484 86522
rect 55188 86468 55244 86470
rect 55268 86468 55324 86470
rect 55348 86468 55404 86470
rect 55428 86468 55484 86470
rect 54528 85978 54584 85980
rect 54608 85978 54664 85980
rect 54688 85978 54744 85980
rect 54768 85978 54824 85980
rect 54528 85926 54574 85978
rect 54574 85926 54584 85978
rect 54608 85926 54638 85978
rect 54638 85926 54650 85978
rect 54650 85926 54664 85978
rect 54688 85926 54702 85978
rect 54702 85926 54714 85978
rect 54714 85926 54744 85978
rect 54768 85926 54778 85978
rect 54778 85926 54824 85978
rect 54528 85924 54584 85926
rect 54608 85924 54664 85926
rect 54688 85924 54744 85926
rect 54768 85924 54824 85926
rect 55188 85434 55244 85436
rect 55268 85434 55324 85436
rect 55348 85434 55404 85436
rect 55428 85434 55484 85436
rect 55188 85382 55234 85434
rect 55234 85382 55244 85434
rect 55268 85382 55298 85434
rect 55298 85382 55310 85434
rect 55310 85382 55324 85434
rect 55348 85382 55362 85434
rect 55362 85382 55374 85434
rect 55374 85382 55404 85434
rect 55428 85382 55438 85434
rect 55438 85382 55484 85434
rect 55188 85380 55244 85382
rect 55268 85380 55324 85382
rect 55348 85380 55404 85382
rect 55428 85380 55484 85382
rect 54528 84890 54584 84892
rect 54608 84890 54664 84892
rect 54688 84890 54744 84892
rect 54768 84890 54824 84892
rect 54528 84838 54574 84890
rect 54574 84838 54584 84890
rect 54608 84838 54638 84890
rect 54638 84838 54650 84890
rect 54650 84838 54664 84890
rect 54688 84838 54702 84890
rect 54702 84838 54714 84890
rect 54714 84838 54744 84890
rect 54768 84838 54778 84890
rect 54778 84838 54824 84890
rect 54528 84836 54584 84838
rect 54608 84836 54664 84838
rect 54688 84836 54744 84838
rect 54768 84836 54824 84838
rect 55188 84346 55244 84348
rect 55268 84346 55324 84348
rect 55348 84346 55404 84348
rect 55428 84346 55484 84348
rect 55188 84294 55234 84346
rect 55234 84294 55244 84346
rect 55268 84294 55298 84346
rect 55298 84294 55310 84346
rect 55310 84294 55324 84346
rect 55348 84294 55362 84346
rect 55362 84294 55374 84346
rect 55374 84294 55404 84346
rect 55428 84294 55438 84346
rect 55438 84294 55484 84346
rect 55188 84292 55244 84294
rect 55268 84292 55324 84294
rect 55348 84292 55404 84294
rect 55428 84292 55484 84294
rect 72928 87066 72984 87068
rect 73008 87066 73064 87068
rect 73088 87066 73144 87068
rect 73168 87066 73224 87068
rect 72928 87014 72974 87066
rect 72974 87014 72984 87066
rect 73008 87014 73038 87066
rect 73038 87014 73050 87066
rect 73050 87014 73064 87066
rect 73088 87014 73102 87066
rect 73102 87014 73114 87066
rect 73114 87014 73144 87066
rect 73168 87014 73178 87066
rect 73178 87014 73224 87066
rect 72928 87012 72984 87014
rect 73008 87012 73064 87014
rect 73088 87012 73144 87014
rect 73168 87012 73224 87014
rect 72928 85978 72984 85980
rect 73008 85978 73064 85980
rect 73088 85978 73144 85980
rect 73168 85978 73224 85980
rect 72928 85926 72974 85978
rect 72974 85926 72984 85978
rect 73008 85926 73038 85978
rect 73038 85926 73050 85978
rect 73050 85926 73064 85978
rect 73088 85926 73102 85978
rect 73102 85926 73114 85978
rect 73114 85926 73144 85978
rect 73168 85926 73178 85978
rect 73178 85926 73224 85978
rect 72928 85924 72984 85926
rect 73008 85924 73064 85926
rect 73088 85924 73144 85926
rect 73168 85924 73224 85926
rect 72928 84890 72984 84892
rect 73008 84890 73064 84892
rect 73088 84890 73144 84892
rect 73168 84890 73224 84892
rect 72928 84838 72974 84890
rect 72974 84838 72984 84890
rect 73008 84838 73038 84890
rect 73038 84838 73050 84890
rect 73050 84838 73064 84890
rect 73088 84838 73102 84890
rect 73102 84838 73114 84890
rect 73114 84838 73144 84890
rect 73168 84838 73178 84890
rect 73178 84838 73224 84890
rect 72928 84836 72984 84838
rect 73008 84836 73064 84838
rect 73088 84836 73144 84838
rect 73168 84836 73224 84838
rect 73588 86522 73644 86524
rect 73668 86522 73724 86524
rect 73748 86522 73804 86524
rect 73828 86522 73884 86524
rect 73588 86470 73634 86522
rect 73634 86470 73644 86522
rect 73668 86470 73698 86522
rect 73698 86470 73710 86522
rect 73710 86470 73724 86522
rect 73748 86470 73762 86522
rect 73762 86470 73774 86522
rect 73774 86470 73804 86522
rect 73828 86470 73838 86522
rect 73838 86470 73884 86522
rect 73588 86468 73644 86470
rect 73668 86468 73724 86470
rect 73748 86468 73804 86470
rect 73828 86468 73884 86470
rect 73588 85434 73644 85436
rect 73668 85434 73724 85436
rect 73748 85434 73804 85436
rect 73828 85434 73884 85436
rect 73588 85382 73634 85434
rect 73634 85382 73644 85434
rect 73668 85382 73698 85434
rect 73698 85382 73710 85434
rect 73710 85382 73724 85434
rect 73748 85382 73762 85434
rect 73762 85382 73774 85434
rect 73774 85382 73804 85434
rect 73828 85382 73838 85434
rect 73838 85382 73884 85434
rect 73588 85380 73644 85382
rect 73668 85380 73724 85382
rect 73748 85380 73804 85382
rect 73828 85380 73884 85382
rect 73588 84346 73644 84348
rect 73668 84346 73724 84348
rect 73748 84346 73804 84348
rect 73828 84346 73884 84348
rect 73588 84294 73634 84346
rect 73634 84294 73644 84346
rect 73668 84294 73698 84346
rect 73698 84294 73710 84346
rect 73710 84294 73724 84346
rect 73748 84294 73762 84346
rect 73762 84294 73774 84346
rect 73774 84294 73804 84346
rect 73828 84294 73838 84346
rect 73838 84294 73884 84346
rect 73588 84292 73644 84294
rect 73668 84292 73724 84294
rect 73748 84292 73804 84294
rect 73828 84292 73884 84294
rect 86552 84890 86608 84892
rect 86632 84890 86688 84892
rect 86712 84890 86768 84892
rect 86792 84890 86848 84892
rect 86552 84838 86598 84890
rect 86598 84838 86608 84890
rect 86632 84838 86662 84890
rect 86662 84838 86674 84890
rect 86674 84838 86688 84890
rect 86712 84838 86726 84890
rect 86726 84838 86738 84890
rect 86738 84838 86768 84890
rect 86792 84838 86802 84890
rect 86802 84838 86848 84890
rect 86552 84836 86608 84838
rect 86632 84836 86688 84838
rect 86712 84836 86768 84838
rect 86792 84836 86848 84838
rect 87288 84346 87344 84348
rect 87368 84346 87424 84348
rect 87448 84346 87504 84348
rect 87528 84346 87584 84348
rect 87288 84294 87334 84346
rect 87334 84294 87344 84346
rect 87368 84294 87398 84346
rect 87398 84294 87410 84346
rect 87410 84294 87424 84346
rect 87448 84294 87462 84346
rect 87462 84294 87474 84346
rect 87474 84294 87504 84346
rect 87528 84294 87538 84346
rect 87538 84294 87584 84346
rect 87288 84292 87344 84294
rect 87368 84292 87424 84294
rect 87448 84292 87504 84294
rect 87528 84292 87584 84294
rect 86552 83802 86608 83804
rect 86632 83802 86688 83804
rect 86712 83802 86768 83804
rect 86792 83802 86848 83804
rect 86552 83750 86598 83802
rect 86598 83750 86608 83802
rect 86632 83750 86662 83802
rect 86662 83750 86674 83802
rect 86674 83750 86688 83802
rect 86712 83750 86726 83802
rect 86726 83750 86738 83802
rect 86738 83750 86768 83802
rect 86792 83750 86802 83802
rect 86802 83750 86848 83802
rect 86552 83748 86608 83750
rect 86632 83748 86688 83750
rect 86712 83748 86768 83750
rect 86792 83748 86848 83750
rect 87288 83258 87344 83260
rect 87368 83258 87424 83260
rect 87448 83258 87504 83260
rect 87528 83258 87584 83260
rect 87288 83206 87334 83258
rect 87334 83206 87344 83258
rect 87368 83206 87398 83258
rect 87398 83206 87410 83258
rect 87410 83206 87424 83258
rect 87448 83206 87462 83258
rect 87462 83206 87474 83258
rect 87474 83206 87504 83258
rect 87528 83206 87538 83258
rect 87538 83206 87584 83258
rect 87288 83204 87344 83206
rect 87368 83204 87424 83206
rect 87448 83204 87504 83206
rect 87528 83204 87584 83206
rect 47066 45704 47122 45760
rect 47342 45704 47398 45760
rect 50178 45432 50234 45488
rect 49074 45296 49130 45352
rect 47342 45160 47398 45216
rect 47970 45160 48026 45216
rect 86552 82714 86608 82716
rect 86632 82714 86688 82716
rect 86712 82714 86768 82716
rect 86792 82714 86848 82716
rect 86552 82662 86598 82714
rect 86598 82662 86608 82714
rect 86632 82662 86662 82714
rect 86662 82662 86674 82714
rect 86674 82662 86688 82714
rect 86712 82662 86726 82714
rect 86726 82662 86738 82714
rect 86738 82662 86768 82714
rect 86792 82662 86802 82714
rect 86802 82662 86848 82714
rect 86552 82660 86608 82662
rect 86632 82660 86688 82662
rect 86712 82660 86768 82662
rect 86792 82660 86848 82662
rect 87288 82170 87344 82172
rect 87368 82170 87424 82172
rect 87448 82170 87504 82172
rect 87528 82170 87584 82172
rect 87288 82118 87334 82170
rect 87334 82118 87344 82170
rect 87368 82118 87398 82170
rect 87398 82118 87410 82170
rect 87410 82118 87424 82170
rect 87448 82118 87462 82170
rect 87462 82118 87474 82170
rect 87474 82118 87504 82170
rect 87528 82118 87538 82170
rect 87538 82118 87584 82170
rect 87288 82116 87344 82118
rect 87368 82116 87424 82118
rect 87448 82116 87504 82118
rect 87528 82116 87584 82118
rect 86552 81626 86608 81628
rect 86632 81626 86688 81628
rect 86712 81626 86768 81628
rect 86792 81626 86848 81628
rect 86552 81574 86598 81626
rect 86598 81574 86608 81626
rect 86632 81574 86662 81626
rect 86662 81574 86674 81626
rect 86674 81574 86688 81626
rect 86712 81574 86726 81626
rect 86726 81574 86738 81626
rect 86738 81574 86768 81626
rect 86792 81574 86802 81626
rect 86802 81574 86848 81626
rect 86552 81572 86608 81574
rect 86632 81572 86688 81574
rect 86712 81572 86768 81574
rect 86792 81572 86848 81574
rect 88374 81244 88376 81256
rect 88376 81244 88428 81256
rect 88428 81244 88430 81256
rect 88374 81200 88430 81244
rect 87288 81082 87344 81084
rect 87368 81082 87424 81084
rect 87448 81082 87504 81084
rect 87528 81082 87584 81084
rect 83498 80996 83554 81052
rect 87288 81030 87334 81082
rect 87334 81030 87344 81082
rect 87368 81030 87398 81082
rect 87398 81030 87410 81082
rect 87410 81030 87424 81082
rect 87448 81030 87462 81082
rect 87462 81030 87474 81082
rect 87474 81030 87504 81082
rect 87528 81030 87538 81082
rect 87538 81030 87584 81082
rect 87288 81028 87344 81030
rect 87368 81028 87424 81030
rect 87448 81028 87504 81030
rect 87528 81028 87584 81030
rect 86552 80538 86608 80540
rect 86632 80538 86688 80540
rect 86712 80538 86768 80540
rect 86792 80538 86848 80540
rect 86552 80486 86598 80538
rect 86598 80486 86608 80538
rect 86632 80486 86662 80538
rect 86662 80486 86674 80538
rect 86674 80486 86688 80538
rect 86712 80486 86726 80538
rect 86726 80486 86738 80538
rect 86738 80486 86768 80538
rect 86792 80486 86802 80538
rect 86802 80486 86848 80538
rect 86552 80484 86608 80486
rect 86632 80484 86688 80486
rect 86712 80484 86768 80486
rect 86792 80484 86848 80486
rect 87288 79994 87344 79996
rect 87368 79994 87424 79996
rect 87448 79994 87504 79996
rect 87528 79994 87584 79996
rect 83498 79908 83554 79964
rect 87288 79942 87334 79994
rect 87334 79942 87344 79994
rect 87368 79942 87398 79994
rect 87398 79942 87410 79994
rect 87410 79942 87424 79994
rect 87448 79942 87462 79994
rect 87462 79942 87474 79994
rect 87474 79942 87504 79994
rect 87528 79942 87538 79994
rect 87538 79942 87584 79994
rect 87288 79940 87344 79942
rect 87368 79940 87424 79942
rect 87448 79940 87504 79942
rect 87528 79940 87584 79942
rect 88282 79840 88338 79896
rect 86552 79450 86608 79452
rect 86632 79450 86688 79452
rect 86712 79450 86768 79452
rect 86792 79450 86848 79452
rect 86552 79398 86598 79450
rect 86598 79398 86608 79450
rect 86632 79398 86662 79450
rect 86662 79398 86674 79450
rect 86674 79398 86688 79450
rect 86712 79398 86726 79450
rect 86726 79398 86738 79450
rect 86738 79398 86768 79450
rect 86792 79398 86802 79450
rect 86802 79398 86848 79450
rect 86552 79396 86608 79398
rect 86632 79396 86688 79398
rect 86712 79396 86768 79398
rect 86792 79396 86848 79398
rect 87288 78906 87344 78908
rect 87368 78906 87424 78908
rect 87448 78906 87504 78908
rect 87528 78906 87584 78908
rect 87288 78854 87334 78906
rect 87334 78854 87344 78906
rect 87368 78854 87398 78906
rect 87398 78854 87410 78906
rect 87410 78854 87424 78906
rect 87448 78854 87462 78906
rect 87462 78854 87474 78906
rect 87474 78854 87504 78906
rect 87528 78854 87538 78906
rect 87538 78854 87584 78906
rect 87288 78852 87344 78854
rect 87368 78852 87424 78854
rect 87448 78852 87504 78854
rect 87528 78852 87584 78854
rect 88006 78616 88062 78672
rect 88282 78480 88338 78536
rect 86552 78362 86608 78364
rect 86632 78362 86688 78364
rect 86712 78362 86768 78364
rect 86792 78362 86848 78364
rect 86552 78310 86598 78362
rect 86598 78310 86608 78362
rect 86632 78310 86662 78362
rect 86662 78310 86674 78362
rect 86674 78310 86688 78362
rect 86712 78310 86726 78362
rect 86726 78310 86738 78362
rect 86738 78310 86768 78362
rect 86792 78310 86802 78362
rect 86802 78310 86848 78362
rect 86552 78308 86608 78310
rect 86632 78308 86688 78310
rect 86712 78308 86768 78310
rect 86792 78308 86848 78310
rect 87822 77956 87878 77992
rect 87822 77936 87824 77956
rect 87824 77936 87876 77956
rect 87876 77936 87878 77956
rect 87288 77818 87344 77820
rect 87368 77818 87424 77820
rect 87448 77818 87504 77820
rect 87528 77818 87584 77820
rect 87288 77766 87334 77818
rect 87334 77766 87344 77818
rect 87368 77766 87398 77818
rect 87398 77766 87410 77818
rect 87410 77766 87424 77818
rect 87448 77766 87462 77818
rect 87462 77766 87474 77818
rect 87474 77766 87504 77818
rect 87528 77766 87538 77818
rect 87538 77766 87584 77818
rect 88282 77800 88338 77856
rect 87288 77764 87344 77766
rect 87368 77764 87424 77766
rect 87448 77764 87504 77766
rect 87528 77764 87584 77766
rect 86552 77274 86608 77276
rect 86632 77274 86688 77276
rect 86712 77274 86768 77276
rect 86792 77274 86848 77276
rect 86552 77222 86598 77274
rect 86598 77222 86608 77274
rect 86632 77222 86662 77274
rect 86662 77222 86674 77274
rect 86674 77222 86688 77274
rect 86712 77222 86726 77274
rect 86726 77222 86738 77274
rect 86738 77222 86768 77274
rect 86792 77222 86802 77274
rect 86802 77222 86848 77274
rect 86552 77220 86608 77222
rect 86632 77220 86688 77222
rect 86712 77220 86768 77222
rect 86792 77220 86848 77222
rect 86626 76712 86682 76768
rect 87288 76730 87344 76732
rect 87368 76730 87424 76732
rect 87448 76730 87504 76732
rect 87528 76730 87584 76732
rect 87288 76678 87334 76730
rect 87334 76678 87344 76730
rect 87368 76678 87398 76730
rect 87398 76678 87410 76730
rect 87410 76678 87424 76730
rect 87448 76678 87462 76730
rect 87462 76678 87474 76730
rect 87474 76678 87504 76730
rect 87528 76678 87538 76730
rect 87538 76678 87584 76730
rect 87288 76676 87344 76678
rect 87368 76676 87424 76678
rect 87448 76676 87504 76678
rect 87528 76676 87584 76678
rect 88006 76440 88062 76496
rect 86552 76186 86608 76188
rect 86632 76186 86688 76188
rect 86712 76186 86768 76188
rect 86792 76186 86848 76188
rect 86552 76134 86598 76186
rect 86598 76134 86608 76186
rect 86632 76134 86662 76186
rect 86662 76134 86674 76186
rect 86674 76134 86688 76186
rect 86712 76134 86726 76186
rect 86726 76134 86738 76186
rect 86738 76134 86768 76186
rect 86792 76134 86802 76186
rect 86802 76134 86848 76186
rect 86552 76132 86608 76134
rect 86632 76132 86688 76134
rect 86712 76132 86768 76134
rect 86792 76132 86848 76134
rect 88466 75796 88468 75816
rect 88468 75796 88520 75816
rect 88520 75796 88522 75816
rect 88466 75760 88522 75796
rect 86902 75624 86958 75680
rect 87288 75642 87344 75644
rect 87368 75642 87424 75644
rect 87448 75642 87504 75644
rect 87528 75642 87584 75644
rect 87288 75590 87334 75642
rect 87334 75590 87344 75642
rect 87368 75590 87398 75642
rect 87398 75590 87410 75642
rect 87410 75590 87424 75642
rect 87448 75590 87462 75642
rect 87462 75590 87474 75642
rect 87474 75590 87504 75642
rect 87528 75590 87538 75642
rect 87538 75590 87584 75642
rect 87288 75588 87344 75590
rect 87368 75588 87424 75590
rect 87448 75588 87504 75590
rect 87528 75588 87584 75590
rect 86552 75098 86608 75100
rect 86632 75098 86688 75100
rect 86712 75098 86768 75100
rect 86792 75098 86848 75100
rect 86552 75046 86598 75098
rect 86598 75046 86608 75098
rect 86632 75046 86662 75098
rect 86662 75046 86674 75098
rect 86674 75046 86688 75098
rect 86712 75046 86726 75098
rect 86726 75046 86738 75098
rect 86738 75046 86768 75098
rect 86792 75046 86802 75098
rect 86802 75046 86848 75098
rect 86552 75044 86608 75046
rect 86632 75044 86688 75046
rect 86712 75044 86768 75046
rect 86792 75044 86848 75046
rect 84418 74536 84474 74592
rect 87288 74554 87344 74556
rect 87368 74554 87424 74556
rect 87448 74554 87504 74556
rect 87528 74554 87584 74556
rect 87288 74502 87334 74554
rect 87334 74502 87344 74554
rect 87368 74502 87398 74554
rect 87398 74502 87410 74554
rect 87410 74502 87424 74554
rect 87448 74502 87462 74554
rect 87462 74502 87474 74554
rect 87474 74502 87504 74554
rect 87528 74502 87538 74554
rect 87538 74502 87584 74554
rect 87288 74500 87344 74502
rect 87368 74500 87424 74502
rect 87448 74500 87504 74502
rect 87528 74500 87584 74502
rect 88558 74400 88614 74456
rect 86552 74010 86608 74012
rect 86632 74010 86688 74012
rect 86712 74010 86768 74012
rect 86792 74010 86848 74012
rect 86552 73958 86598 74010
rect 86598 73958 86608 74010
rect 86632 73958 86662 74010
rect 86662 73958 86674 74010
rect 86674 73958 86688 74010
rect 86712 73958 86726 74010
rect 86726 73958 86738 74010
rect 86738 73958 86768 74010
rect 86792 73958 86802 74010
rect 86802 73958 86848 74010
rect 86552 73956 86608 73958
rect 86632 73956 86688 73958
rect 86712 73956 86768 73958
rect 86792 73956 86848 73958
rect 87288 73466 87344 73468
rect 87368 73466 87424 73468
rect 87448 73466 87504 73468
rect 87528 73466 87584 73468
rect 87288 73414 87334 73466
rect 87334 73414 87344 73466
rect 87368 73414 87398 73466
rect 87398 73414 87410 73466
rect 87410 73414 87424 73466
rect 87448 73414 87462 73466
rect 87462 73414 87474 73466
rect 87474 73414 87504 73466
rect 87528 73414 87538 73466
rect 87538 73414 87584 73466
rect 87288 73412 87344 73414
rect 87368 73412 87424 73414
rect 87448 73412 87504 73414
rect 87528 73412 87584 73414
rect 88006 73196 88062 73232
rect 88006 73176 88008 73196
rect 88008 73176 88060 73196
rect 88060 73176 88062 73196
rect 88282 73040 88338 73096
rect 86552 72922 86608 72924
rect 86632 72922 86688 72924
rect 86712 72922 86768 72924
rect 86792 72922 86848 72924
rect 86552 72870 86598 72922
rect 86598 72870 86608 72922
rect 86632 72870 86662 72922
rect 86662 72870 86674 72922
rect 86674 72870 86688 72922
rect 86712 72870 86726 72922
rect 86726 72870 86738 72922
rect 86738 72870 86768 72922
rect 86792 72870 86802 72922
rect 86802 72870 86848 72922
rect 86552 72868 86608 72870
rect 86632 72868 86688 72870
rect 86712 72868 86768 72870
rect 86792 72868 86848 72870
rect 87178 72532 87180 72552
rect 87180 72532 87232 72552
rect 87232 72532 87234 72552
rect 87178 72496 87234 72532
rect 87288 72378 87344 72380
rect 87368 72378 87424 72380
rect 87448 72378 87504 72380
rect 87528 72378 87584 72380
rect 87288 72326 87334 72378
rect 87334 72326 87344 72378
rect 87368 72326 87398 72378
rect 87398 72326 87410 72378
rect 87410 72326 87424 72378
rect 87448 72326 87462 72378
rect 87462 72326 87474 72378
rect 87474 72326 87504 72378
rect 87528 72326 87538 72378
rect 87538 72326 87584 72378
rect 88282 72360 88338 72416
rect 87288 72324 87344 72326
rect 87368 72324 87424 72326
rect 87448 72324 87504 72326
rect 87528 72324 87584 72326
rect 86552 71834 86608 71836
rect 86632 71834 86688 71836
rect 86712 71834 86768 71836
rect 86792 71834 86848 71836
rect 86552 71782 86598 71834
rect 86598 71782 86608 71834
rect 86632 71782 86662 71834
rect 86662 71782 86674 71834
rect 86674 71782 86688 71834
rect 86712 71782 86726 71834
rect 86726 71782 86738 71834
rect 86738 71782 86768 71834
rect 86792 71782 86802 71834
rect 86802 71782 86848 71834
rect 86552 71780 86608 71782
rect 86632 71780 86688 71782
rect 86712 71780 86768 71782
rect 86792 71780 86848 71782
rect 86902 71272 86958 71328
rect 87288 71290 87344 71292
rect 87368 71290 87424 71292
rect 87448 71290 87504 71292
rect 87528 71290 87584 71292
rect 87288 71238 87334 71290
rect 87334 71238 87344 71290
rect 87368 71238 87398 71290
rect 87398 71238 87410 71290
rect 87410 71238 87424 71290
rect 87448 71238 87462 71290
rect 87462 71238 87474 71290
rect 87474 71238 87504 71290
rect 87528 71238 87538 71290
rect 87538 71238 87584 71290
rect 87288 71236 87344 71238
rect 87368 71236 87424 71238
rect 87448 71236 87504 71238
rect 87528 71236 87584 71238
rect 88282 71000 88338 71056
rect 86552 70746 86608 70748
rect 86632 70746 86688 70748
rect 86712 70746 86768 70748
rect 86792 70746 86848 70748
rect 86552 70694 86598 70746
rect 86598 70694 86608 70746
rect 86632 70694 86662 70746
rect 86662 70694 86674 70746
rect 86674 70694 86688 70746
rect 86712 70694 86726 70746
rect 86726 70694 86738 70746
rect 86738 70694 86768 70746
rect 86792 70694 86802 70746
rect 86802 70694 86848 70746
rect 86552 70692 86608 70694
rect 86632 70692 86688 70694
rect 86712 70692 86768 70694
rect 86792 70692 86848 70694
rect 88190 70320 88246 70376
rect 86902 70184 86958 70240
rect 87288 70202 87344 70204
rect 87368 70202 87424 70204
rect 87448 70202 87504 70204
rect 87528 70202 87584 70204
rect 87288 70150 87334 70202
rect 87334 70150 87344 70202
rect 87368 70150 87398 70202
rect 87398 70150 87410 70202
rect 87410 70150 87424 70202
rect 87448 70150 87462 70202
rect 87462 70150 87474 70202
rect 87474 70150 87504 70202
rect 87528 70150 87538 70202
rect 87538 70150 87584 70202
rect 87288 70148 87344 70150
rect 87368 70148 87424 70150
rect 87448 70148 87504 70150
rect 87528 70148 87584 70150
rect 86552 69658 86608 69660
rect 86632 69658 86688 69660
rect 86712 69658 86768 69660
rect 86792 69658 86848 69660
rect 86552 69606 86598 69658
rect 86598 69606 86608 69658
rect 86632 69606 86662 69658
rect 86662 69606 86674 69658
rect 86674 69606 86688 69658
rect 86712 69606 86726 69658
rect 86726 69606 86738 69658
rect 86738 69606 86768 69658
rect 86792 69606 86802 69658
rect 86802 69606 86848 69658
rect 86552 69604 86608 69606
rect 86632 69604 86688 69606
rect 86712 69604 86768 69606
rect 86792 69604 86848 69606
rect 86902 69096 86958 69152
rect 87288 69114 87344 69116
rect 87368 69114 87424 69116
rect 87448 69114 87504 69116
rect 87528 69114 87584 69116
rect 87288 69062 87334 69114
rect 87334 69062 87344 69114
rect 87368 69062 87398 69114
rect 87398 69062 87410 69114
rect 87410 69062 87424 69114
rect 87448 69062 87462 69114
rect 87462 69062 87474 69114
rect 87474 69062 87504 69114
rect 87528 69062 87538 69114
rect 87538 69062 87584 69114
rect 87288 69060 87344 69062
rect 87368 69060 87424 69062
rect 87448 69060 87504 69062
rect 87528 69060 87584 69062
rect 88558 68960 88614 69016
rect 86552 68570 86608 68572
rect 86632 68570 86688 68572
rect 86712 68570 86768 68572
rect 86792 68570 86848 68572
rect 86552 68518 86598 68570
rect 86598 68518 86608 68570
rect 86632 68518 86662 68570
rect 86662 68518 86674 68570
rect 86674 68518 86688 68570
rect 86712 68518 86726 68570
rect 86726 68518 86738 68570
rect 86738 68518 86768 68570
rect 86792 68518 86802 68570
rect 86802 68518 86848 68570
rect 86552 68516 86608 68518
rect 86632 68516 86688 68518
rect 86712 68516 86768 68518
rect 86792 68516 86848 68518
rect 87288 68026 87344 68028
rect 87368 68026 87424 68028
rect 87448 68026 87504 68028
rect 87528 68026 87584 68028
rect 87288 67974 87334 68026
rect 87334 67974 87344 68026
rect 87368 67974 87398 68026
rect 87398 67974 87410 68026
rect 87410 67974 87424 68026
rect 87448 67974 87462 68026
rect 87462 67974 87474 68026
rect 87474 67974 87504 68026
rect 87528 67974 87538 68026
rect 87538 67974 87584 68026
rect 87288 67972 87344 67974
rect 87368 67972 87424 67974
rect 87448 67972 87504 67974
rect 87528 67972 87584 67974
rect 84418 67872 84474 67928
rect 88282 67600 88338 67656
rect 86552 67482 86608 67484
rect 86632 67482 86688 67484
rect 86712 67482 86768 67484
rect 86792 67482 86848 67484
rect 86552 67430 86598 67482
rect 86598 67430 86608 67482
rect 86632 67430 86662 67482
rect 86662 67430 86674 67482
rect 86674 67430 86688 67482
rect 86712 67430 86726 67482
rect 86726 67430 86738 67482
rect 86738 67430 86768 67482
rect 86792 67430 86802 67482
rect 86802 67430 86848 67482
rect 86552 67428 86608 67430
rect 86632 67428 86688 67430
rect 86712 67428 86768 67430
rect 86792 67428 86848 67430
rect 86902 66920 86958 66976
rect 87288 66938 87344 66940
rect 87368 66938 87424 66940
rect 87448 66938 87504 66940
rect 87528 66938 87584 66940
rect 87288 66886 87334 66938
rect 87334 66886 87344 66938
rect 87368 66886 87398 66938
rect 87398 66886 87410 66938
rect 87410 66886 87424 66938
rect 87448 66886 87462 66938
rect 87462 66886 87474 66938
rect 87474 66886 87504 66938
rect 87528 66886 87538 66938
rect 87538 66886 87584 66938
rect 88282 66920 88338 66976
rect 87288 66884 87344 66886
rect 87368 66884 87424 66886
rect 87448 66884 87504 66886
rect 87528 66884 87584 66886
rect 86552 66394 86608 66396
rect 86632 66394 86688 66396
rect 86712 66394 86768 66396
rect 86792 66394 86848 66396
rect 86552 66342 86598 66394
rect 86598 66342 86608 66394
rect 86632 66342 86662 66394
rect 86662 66342 86674 66394
rect 86674 66342 86688 66394
rect 86712 66342 86726 66394
rect 86726 66342 86738 66394
rect 86738 66342 86768 66394
rect 86792 66342 86802 66394
rect 86802 66342 86848 66394
rect 86552 66340 86608 66342
rect 86632 66340 86688 66342
rect 86712 66340 86768 66342
rect 86792 66340 86848 66342
rect 87086 65832 87142 65888
rect 87288 65850 87344 65852
rect 87368 65850 87424 65852
rect 87448 65850 87504 65852
rect 87528 65850 87584 65852
rect 87288 65798 87334 65850
rect 87334 65798 87344 65850
rect 87368 65798 87398 65850
rect 87398 65798 87410 65850
rect 87410 65798 87424 65850
rect 87448 65798 87462 65850
rect 87462 65798 87474 65850
rect 87474 65798 87504 65850
rect 87528 65798 87538 65850
rect 87538 65798 87584 65850
rect 87288 65796 87344 65798
rect 87368 65796 87424 65798
rect 87448 65796 87504 65798
rect 87528 65796 87584 65798
rect 88190 65560 88246 65616
rect 86552 65306 86608 65308
rect 86632 65306 86688 65308
rect 86712 65306 86768 65308
rect 86792 65306 86848 65308
rect 86552 65254 86598 65306
rect 86598 65254 86608 65306
rect 86632 65254 86662 65306
rect 86662 65254 86674 65306
rect 86674 65254 86688 65306
rect 86712 65254 86726 65306
rect 86726 65254 86738 65306
rect 86738 65254 86768 65306
rect 86792 65254 86802 65306
rect 86802 65254 86848 65306
rect 86552 65252 86608 65254
rect 86632 65252 86688 65254
rect 86712 65252 86768 65254
rect 86792 65252 86848 65254
rect 88374 64900 88430 64936
rect 88374 64880 88376 64900
rect 88376 64880 88428 64900
rect 88428 64880 88430 64900
rect 87086 64744 87142 64800
rect 87288 64762 87344 64764
rect 87368 64762 87424 64764
rect 87448 64762 87504 64764
rect 87528 64762 87584 64764
rect 87288 64710 87334 64762
rect 87334 64710 87344 64762
rect 87368 64710 87398 64762
rect 87398 64710 87410 64762
rect 87410 64710 87424 64762
rect 87448 64710 87462 64762
rect 87462 64710 87474 64762
rect 87474 64710 87504 64762
rect 87528 64710 87538 64762
rect 87538 64710 87584 64762
rect 87288 64708 87344 64710
rect 87368 64708 87424 64710
rect 87448 64708 87504 64710
rect 87528 64708 87584 64710
rect 86552 64218 86608 64220
rect 86632 64218 86688 64220
rect 86712 64218 86768 64220
rect 86792 64218 86848 64220
rect 86552 64166 86598 64218
rect 86598 64166 86608 64218
rect 86632 64166 86662 64218
rect 86662 64166 86674 64218
rect 86674 64166 86688 64218
rect 86712 64166 86726 64218
rect 86726 64166 86738 64218
rect 86738 64166 86768 64218
rect 86792 64166 86802 64218
rect 86802 64166 86848 64218
rect 86552 64164 86608 64166
rect 86632 64164 86688 64166
rect 86712 64164 86768 64166
rect 86792 64164 86848 64166
rect 84418 63656 84474 63712
rect 87288 63674 87344 63676
rect 87368 63674 87424 63676
rect 87448 63674 87504 63676
rect 87528 63674 87584 63676
rect 87288 63622 87334 63674
rect 87334 63622 87344 63674
rect 87368 63622 87398 63674
rect 87398 63622 87410 63674
rect 87410 63622 87424 63674
rect 87448 63622 87462 63674
rect 87462 63622 87474 63674
rect 87474 63622 87504 63674
rect 87528 63622 87538 63674
rect 87538 63622 87584 63674
rect 87288 63620 87344 63622
rect 87368 63620 87424 63622
rect 87448 63620 87504 63622
rect 87528 63620 87584 63622
rect 88558 63520 88614 63576
rect 86552 63130 86608 63132
rect 86632 63130 86688 63132
rect 86712 63130 86768 63132
rect 86792 63130 86848 63132
rect 86552 63078 86598 63130
rect 86598 63078 86608 63130
rect 86632 63078 86662 63130
rect 86662 63078 86674 63130
rect 86674 63078 86688 63130
rect 86712 63078 86726 63130
rect 86726 63078 86738 63130
rect 86738 63078 86768 63130
rect 86792 63078 86802 63130
rect 86802 63078 86848 63130
rect 86552 63076 86608 63078
rect 86632 63076 86688 63078
rect 86712 63076 86768 63078
rect 86792 63076 86848 63078
rect 87288 62586 87344 62588
rect 87368 62586 87424 62588
rect 87448 62586 87504 62588
rect 87528 62586 87584 62588
rect 87288 62534 87334 62586
rect 87334 62534 87344 62586
rect 87368 62534 87398 62586
rect 87398 62534 87410 62586
rect 87410 62534 87424 62586
rect 87448 62534 87462 62586
rect 87462 62534 87474 62586
rect 87474 62534 87504 62586
rect 87528 62534 87538 62586
rect 87538 62534 87584 62586
rect 87288 62532 87344 62534
rect 87368 62532 87424 62534
rect 87448 62532 87504 62534
rect 87528 62532 87584 62534
rect 87086 62432 87142 62488
rect 88558 62160 88614 62216
rect 86552 62042 86608 62044
rect 86632 62042 86688 62044
rect 86712 62042 86768 62044
rect 86792 62042 86848 62044
rect 86552 61990 86598 62042
rect 86598 61990 86608 62042
rect 86632 61990 86662 62042
rect 86662 61990 86674 62042
rect 86674 61990 86688 62042
rect 86712 61990 86726 62042
rect 86726 61990 86738 62042
rect 86738 61990 86768 62042
rect 86792 61990 86802 62042
rect 86802 61990 86848 62042
rect 86552 61988 86608 61990
rect 86632 61988 86688 61990
rect 86712 61988 86768 61990
rect 86792 61988 86848 61990
rect 87086 61480 87142 61536
rect 87288 61498 87344 61500
rect 87368 61498 87424 61500
rect 87448 61498 87504 61500
rect 87528 61498 87584 61500
rect 87288 61446 87334 61498
rect 87334 61446 87344 61498
rect 87368 61446 87398 61498
rect 87398 61446 87410 61498
rect 87410 61446 87424 61498
rect 87448 61446 87462 61498
rect 87462 61446 87474 61498
rect 87474 61446 87504 61498
rect 87528 61446 87538 61498
rect 87538 61446 87584 61498
rect 88190 61480 88246 61536
rect 87288 61444 87344 61446
rect 87368 61444 87424 61446
rect 87448 61444 87504 61446
rect 87528 61444 87584 61446
rect 86552 60954 86608 60956
rect 86632 60954 86688 60956
rect 86712 60954 86768 60956
rect 86792 60954 86848 60956
rect 86552 60902 86598 60954
rect 86598 60902 86608 60954
rect 86632 60902 86662 60954
rect 86662 60902 86674 60954
rect 86674 60902 86688 60954
rect 86712 60902 86726 60954
rect 86726 60902 86738 60954
rect 86738 60902 86768 60954
rect 86792 60902 86802 60954
rect 86802 60902 86848 60954
rect 86552 60900 86608 60902
rect 86632 60900 86688 60902
rect 86712 60900 86768 60902
rect 86792 60900 86848 60902
rect 87086 60392 87142 60448
rect 87288 60410 87344 60412
rect 87368 60410 87424 60412
rect 87448 60410 87504 60412
rect 87528 60410 87584 60412
rect 87288 60358 87334 60410
rect 87334 60358 87344 60410
rect 87368 60358 87398 60410
rect 87398 60358 87410 60410
rect 87410 60358 87424 60410
rect 87448 60358 87462 60410
rect 87462 60358 87474 60410
rect 87474 60358 87504 60410
rect 87528 60358 87538 60410
rect 87538 60358 87584 60410
rect 87288 60356 87344 60358
rect 87368 60356 87424 60358
rect 87448 60356 87504 60358
rect 87528 60356 87584 60358
rect 88190 60120 88246 60176
rect 86552 59866 86608 59868
rect 86632 59866 86688 59868
rect 86712 59866 86768 59868
rect 86792 59866 86848 59868
rect 86552 59814 86598 59866
rect 86598 59814 86608 59866
rect 86632 59814 86662 59866
rect 86662 59814 86674 59866
rect 86674 59814 86688 59866
rect 86712 59814 86726 59866
rect 86726 59814 86738 59866
rect 86738 59814 86768 59866
rect 86792 59814 86802 59866
rect 86802 59814 86848 59866
rect 86552 59812 86608 59814
rect 86632 59812 86688 59814
rect 86712 59812 86768 59814
rect 86792 59812 86848 59814
rect 87638 59476 87640 59496
rect 87640 59476 87692 59496
rect 87692 59476 87694 59496
rect 87638 59440 87694 59476
rect 88374 59460 88430 59496
rect 88374 59440 88376 59460
rect 88376 59440 88428 59460
rect 88428 59440 88430 59460
rect 87288 59322 87344 59324
rect 87368 59322 87424 59324
rect 87448 59322 87504 59324
rect 87528 59322 87584 59324
rect 87288 59270 87334 59322
rect 87334 59270 87344 59322
rect 87368 59270 87398 59322
rect 87398 59270 87410 59322
rect 87410 59270 87424 59322
rect 87448 59270 87462 59322
rect 87462 59270 87474 59322
rect 87474 59270 87504 59322
rect 87528 59270 87538 59322
rect 87538 59270 87584 59322
rect 87288 59268 87344 59270
rect 87368 59268 87424 59270
rect 87448 59268 87504 59270
rect 87528 59268 87584 59270
rect 86552 58778 86608 58780
rect 86632 58778 86688 58780
rect 86712 58778 86768 58780
rect 86792 58778 86848 58780
rect 86552 58726 86598 58778
rect 86598 58726 86608 58778
rect 86632 58726 86662 58778
rect 86662 58726 86674 58778
rect 86674 58726 86688 58778
rect 86712 58726 86726 58778
rect 86726 58726 86738 58778
rect 86738 58726 86768 58778
rect 86792 58726 86802 58778
rect 86802 58726 86848 58778
rect 86552 58724 86608 58726
rect 86632 58724 86688 58726
rect 86712 58724 86768 58726
rect 86792 58724 86848 58726
rect 87288 58234 87344 58236
rect 87368 58234 87424 58236
rect 87448 58234 87504 58236
rect 87528 58234 87584 58236
rect 87288 58182 87334 58234
rect 87334 58182 87344 58234
rect 87368 58182 87398 58234
rect 87398 58182 87410 58234
rect 87410 58182 87424 58234
rect 87448 58182 87462 58234
rect 87462 58182 87474 58234
rect 87474 58182 87504 58234
rect 87528 58182 87538 58234
rect 87538 58182 87584 58234
rect 87288 58180 87344 58182
rect 87368 58180 87424 58182
rect 87448 58180 87504 58182
rect 87528 58180 87584 58182
rect 88558 58080 88614 58136
rect 88006 57944 88062 58000
rect 86552 57690 86608 57692
rect 86632 57690 86688 57692
rect 86712 57690 86768 57692
rect 86792 57690 86848 57692
rect 86552 57638 86598 57690
rect 86598 57638 86608 57690
rect 86632 57638 86662 57690
rect 86662 57638 86674 57690
rect 86674 57638 86688 57690
rect 86712 57638 86726 57690
rect 86726 57638 86738 57690
rect 86738 57638 86768 57690
rect 86792 57638 86802 57690
rect 86802 57638 86848 57690
rect 86552 57636 86608 57638
rect 86632 57636 86688 57638
rect 86712 57636 86768 57638
rect 86792 57636 86848 57638
rect 87288 57146 87344 57148
rect 87368 57146 87424 57148
rect 87448 57146 87504 57148
rect 87528 57146 87584 57148
rect 87288 57094 87334 57146
rect 87334 57094 87344 57146
rect 87368 57094 87398 57146
rect 87398 57094 87410 57146
rect 87410 57094 87424 57146
rect 87448 57094 87462 57146
rect 87462 57094 87474 57146
rect 87474 57094 87504 57146
rect 87528 57094 87538 57146
rect 87538 57094 87584 57146
rect 87288 57092 87344 57094
rect 87368 57092 87424 57094
rect 87448 57092 87504 57094
rect 87528 57092 87584 57094
rect 88006 56910 88062 56912
rect 88006 56858 88008 56910
rect 88008 56858 88060 56910
rect 88060 56858 88062 56910
rect 88006 56856 88062 56858
rect 88834 56720 88890 56776
rect 86552 56602 86608 56604
rect 86632 56602 86688 56604
rect 86712 56602 86768 56604
rect 86792 56602 86848 56604
rect 86552 56550 86598 56602
rect 86598 56550 86608 56602
rect 86632 56550 86662 56602
rect 86662 56550 86674 56602
rect 86674 56550 86688 56602
rect 86712 56550 86726 56602
rect 86726 56550 86738 56602
rect 86738 56550 86768 56602
rect 86792 56550 86802 56602
rect 86802 56550 86848 56602
rect 86552 56548 86608 56550
rect 86632 56548 86688 56550
rect 86712 56548 86768 56550
rect 86792 56548 86848 56550
rect 87086 56040 87142 56096
rect 87288 56058 87344 56060
rect 87368 56058 87424 56060
rect 87448 56058 87504 56060
rect 87528 56058 87584 56060
rect 87288 56006 87334 56058
rect 87334 56006 87344 56058
rect 87368 56006 87398 56058
rect 87398 56006 87410 56058
rect 87410 56006 87424 56058
rect 87448 56006 87462 56058
rect 87462 56006 87474 56058
rect 87474 56006 87504 56058
rect 87528 56006 87538 56058
rect 87538 56006 87584 56058
rect 88190 56040 88246 56096
rect 87288 56004 87344 56006
rect 87368 56004 87424 56006
rect 87448 56004 87504 56006
rect 87528 56004 87584 56006
rect 86552 55514 86608 55516
rect 86632 55514 86688 55516
rect 86712 55514 86768 55516
rect 86792 55514 86848 55516
rect 86552 55462 86598 55514
rect 86598 55462 86608 55514
rect 86632 55462 86662 55514
rect 86662 55462 86674 55514
rect 86674 55462 86688 55514
rect 86712 55462 86726 55514
rect 86726 55462 86738 55514
rect 86738 55462 86768 55514
rect 86792 55462 86802 55514
rect 86802 55462 86848 55514
rect 86552 55460 86608 55462
rect 86632 55460 86688 55462
rect 86712 55460 86768 55462
rect 86792 55460 86848 55462
rect 87086 54952 87142 55008
rect 87288 54970 87344 54972
rect 87368 54970 87424 54972
rect 87448 54970 87504 54972
rect 87528 54970 87584 54972
rect 87288 54918 87334 54970
rect 87334 54918 87344 54970
rect 87368 54918 87398 54970
rect 87398 54918 87410 54970
rect 87410 54918 87424 54970
rect 87448 54918 87462 54970
rect 87462 54918 87474 54970
rect 87474 54918 87504 54970
rect 87528 54918 87538 54970
rect 87538 54918 87584 54970
rect 87288 54916 87344 54918
rect 87368 54916 87424 54918
rect 87448 54916 87504 54918
rect 87528 54916 87584 54918
rect 88190 54680 88246 54736
rect 86552 54426 86608 54428
rect 86632 54426 86688 54428
rect 86712 54426 86768 54428
rect 86792 54426 86848 54428
rect 86552 54374 86598 54426
rect 86598 54374 86608 54426
rect 86632 54374 86662 54426
rect 86662 54374 86674 54426
rect 86674 54374 86688 54426
rect 86712 54374 86726 54426
rect 86726 54374 86738 54426
rect 86738 54374 86768 54426
rect 86792 54374 86802 54426
rect 86802 54374 86848 54426
rect 86552 54372 86608 54374
rect 86632 54372 86688 54374
rect 86712 54372 86768 54374
rect 86792 54372 86848 54374
rect 88650 54036 88652 54056
rect 88652 54036 88704 54056
rect 88704 54036 88706 54056
rect 88650 54000 88706 54036
rect 84418 53864 84474 53920
rect 87288 53882 87344 53884
rect 87368 53882 87424 53884
rect 87448 53882 87504 53884
rect 87528 53882 87584 53884
rect 87288 53830 87334 53882
rect 87334 53830 87344 53882
rect 87368 53830 87398 53882
rect 87398 53830 87410 53882
rect 87410 53830 87424 53882
rect 87448 53830 87462 53882
rect 87462 53830 87474 53882
rect 87474 53830 87504 53882
rect 87528 53830 87538 53882
rect 87538 53830 87584 53882
rect 87288 53828 87344 53830
rect 87368 53828 87424 53830
rect 87448 53828 87504 53830
rect 87528 53828 87584 53830
rect 86552 53338 86608 53340
rect 86632 53338 86688 53340
rect 86712 53338 86768 53340
rect 86792 53338 86848 53340
rect 86552 53286 86598 53338
rect 86598 53286 86608 53338
rect 86632 53286 86662 53338
rect 86662 53286 86674 53338
rect 86674 53286 86688 53338
rect 86712 53286 86726 53338
rect 86726 53286 86738 53338
rect 86738 53286 86768 53338
rect 86792 53286 86802 53338
rect 86802 53286 86848 53338
rect 86552 53284 86608 53286
rect 86632 53284 86688 53286
rect 86712 53284 86768 53286
rect 86792 53284 86848 53286
rect 87086 52776 87142 52832
rect 87288 52794 87344 52796
rect 87368 52794 87424 52796
rect 87448 52794 87504 52796
rect 87528 52794 87584 52796
rect 87288 52742 87334 52794
rect 87334 52742 87344 52794
rect 87368 52742 87398 52794
rect 87398 52742 87410 52794
rect 87410 52742 87424 52794
rect 87448 52742 87462 52794
rect 87462 52742 87474 52794
rect 87474 52742 87504 52794
rect 87528 52742 87538 52794
rect 87538 52742 87584 52794
rect 87288 52740 87344 52742
rect 87368 52740 87424 52742
rect 87448 52740 87504 52742
rect 87528 52740 87584 52742
rect 88282 52640 88338 52696
rect 86552 52250 86608 52252
rect 86632 52250 86688 52252
rect 86712 52250 86768 52252
rect 86792 52250 86848 52252
rect 86552 52198 86598 52250
rect 86598 52198 86608 52250
rect 86632 52198 86662 52250
rect 86662 52198 86674 52250
rect 86674 52198 86688 52250
rect 86712 52198 86726 52250
rect 86726 52198 86738 52250
rect 86738 52198 86768 52250
rect 86792 52198 86802 52250
rect 86802 52198 86848 52250
rect 86552 52196 86608 52198
rect 86632 52196 86688 52198
rect 86712 52196 86768 52198
rect 86792 52196 86848 52198
rect 87288 51706 87344 51708
rect 87368 51706 87424 51708
rect 87448 51706 87504 51708
rect 87528 51706 87584 51708
rect 87288 51654 87334 51706
rect 87334 51654 87344 51706
rect 87368 51654 87398 51706
rect 87398 51654 87410 51706
rect 87410 51654 87424 51706
rect 87448 51654 87462 51706
rect 87462 51654 87474 51706
rect 87474 51654 87504 51706
rect 87528 51654 87538 51706
rect 87538 51654 87584 51706
rect 87288 51652 87344 51654
rect 87368 51652 87424 51654
rect 87448 51652 87504 51654
rect 87528 51652 87584 51654
rect 85798 51552 85854 51608
rect 88190 51316 88192 51336
rect 88192 51316 88244 51336
rect 88244 51316 88246 51336
rect 88190 51280 88246 51316
rect 86552 51162 86608 51164
rect 86632 51162 86688 51164
rect 86712 51162 86768 51164
rect 86792 51162 86848 51164
rect 86552 51110 86598 51162
rect 86598 51110 86608 51162
rect 86632 51110 86662 51162
rect 86662 51110 86674 51162
rect 86674 51110 86688 51162
rect 86712 51110 86726 51162
rect 86726 51110 86738 51162
rect 86738 51110 86768 51162
rect 86792 51110 86802 51162
rect 86802 51110 86848 51162
rect 86552 51108 86608 51110
rect 86632 51108 86688 51110
rect 86712 51108 86768 51110
rect 86792 51108 86848 51110
rect 87288 50618 87344 50620
rect 87368 50618 87424 50620
rect 87448 50618 87504 50620
rect 87528 50618 87584 50620
rect 87288 50566 87334 50618
rect 87334 50566 87344 50618
rect 87368 50566 87398 50618
rect 87398 50566 87410 50618
rect 87410 50566 87424 50618
rect 87448 50566 87462 50618
rect 87462 50566 87474 50618
rect 87474 50566 87504 50618
rect 87528 50566 87538 50618
rect 87538 50566 87584 50618
rect 87288 50564 87344 50566
rect 87368 50564 87424 50566
rect 87448 50564 87504 50566
rect 87528 50564 87584 50566
rect 85430 50464 85486 50520
rect 85338 48288 85394 48344
rect 84418 38088 84474 38144
rect 84418 35912 84474 35968
rect 84418 32648 84474 32704
rect 84418 30472 84474 30528
rect 85246 27208 85302 27264
rect 84418 21768 84474 21824
rect 84418 20680 84474 20736
rect 84418 15240 84474 15296
rect 83682 14152 83738 14208
rect 83498 13032 83554 13088
rect 83498 11944 83554 12000
rect 46422 10888 46478 10944
rect 83314 10820 83370 10876
rect 54528 7642 54584 7644
rect 54608 7642 54664 7644
rect 54688 7642 54744 7644
rect 54768 7642 54824 7644
rect 54528 7590 54574 7642
rect 54574 7590 54584 7642
rect 54608 7590 54638 7642
rect 54638 7590 54650 7642
rect 54650 7590 54664 7642
rect 54688 7590 54702 7642
rect 54702 7590 54714 7642
rect 54714 7590 54744 7642
rect 54768 7590 54778 7642
rect 54778 7590 54824 7642
rect 54528 7588 54584 7590
rect 54608 7588 54664 7590
rect 54688 7588 54744 7590
rect 54768 7588 54824 7590
rect 54528 6554 54584 6556
rect 54608 6554 54664 6556
rect 54688 6554 54744 6556
rect 54768 6554 54824 6556
rect 54528 6502 54574 6554
rect 54574 6502 54584 6554
rect 54608 6502 54638 6554
rect 54638 6502 54650 6554
rect 54650 6502 54664 6554
rect 54688 6502 54702 6554
rect 54702 6502 54714 6554
rect 54714 6502 54744 6554
rect 54768 6502 54778 6554
rect 54778 6502 54824 6554
rect 54528 6500 54584 6502
rect 54608 6500 54664 6502
rect 54688 6500 54744 6502
rect 54768 6500 54824 6502
rect 54528 5466 54584 5468
rect 54608 5466 54664 5468
rect 54688 5466 54744 5468
rect 54768 5466 54824 5468
rect 54528 5414 54574 5466
rect 54574 5414 54584 5466
rect 54608 5414 54638 5466
rect 54638 5414 54650 5466
rect 54650 5414 54664 5466
rect 54688 5414 54702 5466
rect 54702 5414 54714 5466
rect 54714 5414 54744 5466
rect 54768 5414 54778 5466
rect 54778 5414 54824 5466
rect 54528 5412 54584 5414
rect 54608 5412 54664 5414
rect 54688 5412 54744 5414
rect 54768 5412 54824 5414
rect 55188 7098 55244 7100
rect 55268 7098 55324 7100
rect 55348 7098 55404 7100
rect 55428 7098 55484 7100
rect 55188 7046 55234 7098
rect 55234 7046 55244 7098
rect 55268 7046 55298 7098
rect 55298 7046 55310 7098
rect 55310 7046 55324 7098
rect 55348 7046 55362 7098
rect 55362 7046 55374 7098
rect 55374 7046 55404 7098
rect 55428 7046 55438 7098
rect 55438 7046 55484 7098
rect 55188 7044 55244 7046
rect 55268 7044 55324 7046
rect 55348 7044 55404 7046
rect 55428 7044 55484 7046
rect 55188 6010 55244 6012
rect 55268 6010 55324 6012
rect 55348 6010 55404 6012
rect 55428 6010 55484 6012
rect 55188 5958 55234 6010
rect 55234 5958 55244 6010
rect 55268 5958 55298 6010
rect 55298 5958 55310 6010
rect 55310 5958 55324 6010
rect 55348 5958 55362 6010
rect 55362 5958 55374 6010
rect 55374 5958 55404 6010
rect 55428 5958 55438 6010
rect 55438 5958 55484 6010
rect 55188 5956 55244 5958
rect 55268 5956 55324 5958
rect 55348 5956 55404 5958
rect 55428 5956 55484 5958
rect 72928 7642 72984 7644
rect 73008 7642 73064 7644
rect 73088 7642 73144 7644
rect 73168 7642 73224 7644
rect 72928 7590 72974 7642
rect 72974 7590 72984 7642
rect 73008 7590 73038 7642
rect 73038 7590 73050 7642
rect 73050 7590 73064 7642
rect 73088 7590 73102 7642
rect 73102 7590 73114 7642
rect 73114 7590 73144 7642
rect 73168 7590 73178 7642
rect 73178 7590 73224 7642
rect 72928 7588 72984 7590
rect 73008 7588 73064 7590
rect 73088 7588 73144 7590
rect 73168 7588 73224 7590
rect 72928 6554 72984 6556
rect 73008 6554 73064 6556
rect 73088 6554 73144 6556
rect 73168 6554 73224 6556
rect 72928 6502 72974 6554
rect 72974 6502 72984 6554
rect 73008 6502 73038 6554
rect 73038 6502 73050 6554
rect 73050 6502 73064 6554
rect 73088 6502 73102 6554
rect 73102 6502 73114 6554
rect 73114 6502 73144 6554
rect 73168 6502 73178 6554
rect 73178 6502 73224 6554
rect 72928 6500 72984 6502
rect 73008 6500 73064 6502
rect 73088 6500 73144 6502
rect 73168 6500 73224 6502
rect 72928 5466 72984 5468
rect 73008 5466 73064 5468
rect 73088 5466 73144 5468
rect 73168 5466 73224 5468
rect 72928 5414 72974 5466
rect 72974 5414 72984 5466
rect 73008 5414 73038 5466
rect 73038 5414 73050 5466
rect 73050 5414 73064 5466
rect 73088 5414 73102 5466
rect 73102 5414 73114 5466
rect 73114 5414 73144 5466
rect 73168 5414 73178 5466
rect 73178 5414 73224 5466
rect 72928 5412 72984 5414
rect 73008 5412 73064 5414
rect 73088 5412 73144 5414
rect 73168 5412 73224 5414
rect 73588 7098 73644 7100
rect 73668 7098 73724 7100
rect 73748 7098 73804 7100
rect 73828 7098 73884 7100
rect 73588 7046 73634 7098
rect 73634 7046 73644 7098
rect 73668 7046 73698 7098
rect 73698 7046 73710 7098
rect 73710 7046 73724 7098
rect 73748 7046 73762 7098
rect 73762 7046 73774 7098
rect 73774 7046 73804 7098
rect 73828 7046 73838 7098
rect 73838 7046 73884 7098
rect 73588 7044 73644 7046
rect 73668 7044 73724 7046
rect 73748 7044 73804 7046
rect 73828 7044 73884 7046
rect 73588 6010 73644 6012
rect 73668 6010 73724 6012
rect 73748 6010 73804 6012
rect 73828 6010 73884 6012
rect 73588 5958 73634 6010
rect 73634 5958 73644 6010
rect 73668 5958 73698 6010
rect 73698 5958 73710 6010
rect 73710 5958 73724 6010
rect 73748 5958 73762 6010
rect 73762 5958 73774 6010
rect 73774 5958 73804 6010
rect 73828 5958 73838 6010
rect 73838 5958 73884 6010
rect 73588 5956 73644 5958
rect 73668 5956 73724 5958
rect 73748 5956 73804 5958
rect 73828 5956 73884 5958
rect 86552 50074 86608 50076
rect 86632 50074 86688 50076
rect 86712 50074 86768 50076
rect 86792 50074 86848 50076
rect 86552 50022 86598 50074
rect 86598 50022 86608 50074
rect 86632 50022 86662 50074
rect 86662 50022 86674 50074
rect 86674 50022 86688 50074
rect 86712 50022 86726 50074
rect 86726 50022 86738 50074
rect 86738 50022 86768 50074
rect 86792 50022 86802 50074
rect 86802 50022 86848 50074
rect 86552 50020 86608 50022
rect 86632 50020 86688 50022
rect 86712 50020 86768 50022
rect 86792 50020 86848 50022
rect 87288 49530 87344 49532
rect 87368 49530 87424 49532
rect 87448 49530 87504 49532
rect 87528 49530 87584 49532
rect 87288 49478 87334 49530
rect 87334 49478 87344 49530
rect 87368 49478 87398 49530
rect 87398 49478 87410 49530
rect 87410 49478 87424 49530
rect 87448 49478 87462 49530
rect 87462 49478 87474 49530
rect 87474 49478 87504 49530
rect 87528 49478 87538 49530
rect 87538 49478 87584 49530
rect 87288 49476 87344 49478
rect 87368 49476 87424 49478
rect 87448 49476 87504 49478
rect 87528 49476 87584 49478
rect 85522 49376 85578 49432
rect 86552 48986 86608 48988
rect 86632 48986 86688 48988
rect 86712 48986 86768 48988
rect 86792 48986 86848 48988
rect 86552 48934 86598 48986
rect 86598 48934 86608 48986
rect 86632 48934 86662 48986
rect 86662 48934 86674 48986
rect 86674 48934 86688 48986
rect 86712 48934 86726 48986
rect 86726 48934 86738 48986
rect 86738 48934 86768 48986
rect 86792 48934 86802 48986
rect 86802 48934 86848 48986
rect 86552 48932 86608 48934
rect 86632 48932 86688 48934
rect 86712 48932 86768 48934
rect 86792 48932 86848 48934
rect 88190 48596 88192 48616
rect 88192 48596 88244 48616
rect 88244 48596 88246 48616
rect 88190 48560 88246 48596
rect 87288 48442 87344 48444
rect 87368 48442 87424 48444
rect 87448 48442 87504 48444
rect 87528 48442 87584 48444
rect 87288 48390 87334 48442
rect 87334 48390 87344 48442
rect 87368 48390 87398 48442
rect 87398 48390 87410 48442
rect 87410 48390 87424 48442
rect 87448 48390 87462 48442
rect 87462 48390 87474 48442
rect 87474 48390 87504 48442
rect 87528 48390 87538 48442
rect 87538 48390 87584 48442
rect 87288 48388 87344 48390
rect 87368 48388 87424 48390
rect 87448 48388 87504 48390
rect 87528 48388 87584 48390
rect 86552 47898 86608 47900
rect 86632 47898 86688 47900
rect 86712 47898 86768 47900
rect 86792 47898 86848 47900
rect 86552 47846 86598 47898
rect 86598 47846 86608 47898
rect 86632 47846 86662 47898
rect 86662 47846 86674 47898
rect 86674 47846 86688 47898
rect 86712 47846 86726 47898
rect 86726 47846 86738 47898
rect 86738 47846 86768 47898
rect 86792 47846 86802 47898
rect 86802 47846 86848 47898
rect 88190 47880 88246 47936
rect 86552 47844 86608 47846
rect 86632 47844 86688 47846
rect 86712 47844 86768 47846
rect 86792 47844 86848 47846
rect 85798 47336 85854 47392
rect 87288 47354 87344 47356
rect 87368 47354 87424 47356
rect 87448 47354 87504 47356
rect 87528 47354 87584 47356
rect 87288 47302 87334 47354
rect 87334 47302 87344 47354
rect 87368 47302 87398 47354
rect 87398 47302 87410 47354
rect 87410 47302 87424 47354
rect 87448 47302 87462 47354
rect 87462 47302 87474 47354
rect 87474 47302 87504 47354
rect 87528 47302 87538 47354
rect 87538 47302 87584 47354
rect 87288 47300 87344 47302
rect 87368 47300 87424 47302
rect 87448 47300 87504 47302
rect 87528 47300 87584 47302
rect 88190 47200 88246 47256
rect 86552 46810 86608 46812
rect 86632 46810 86688 46812
rect 86712 46810 86768 46812
rect 86792 46810 86848 46812
rect 86552 46758 86598 46810
rect 86598 46758 86608 46810
rect 86632 46758 86662 46810
rect 86662 46758 86674 46810
rect 86674 46758 86688 46810
rect 86712 46758 86726 46810
rect 86726 46758 86738 46810
rect 86738 46758 86768 46810
rect 86792 46758 86802 46810
rect 86802 46758 86848 46810
rect 86552 46756 86608 46758
rect 86632 46756 86688 46758
rect 86712 46756 86768 46758
rect 86792 46756 86848 46758
rect 88190 46520 88246 46576
rect 87288 46266 87344 46268
rect 87368 46266 87424 46268
rect 87448 46266 87504 46268
rect 87528 46266 87584 46268
rect 87288 46214 87334 46266
rect 87334 46214 87344 46266
rect 87368 46214 87398 46266
rect 87398 46214 87410 46266
rect 87410 46214 87424 46266
rect 87448 46214 87462 46266
rect 87462 46214 87474 46266
rect 87474 46214 87504 46266
rect 87528 46214 87538 46266
rect 87538 46214 87584 46266
rect 87288 46212 87344 46214
rect 87368 46212 87424 46214
rect 87448 46212 87504 46214
rect 87528 46212 87584 46214
rect 88190 45860 88246 45896
rect 88190 45840 88192 45860
rect 88192 45840 88244 45860
rect 88244 45840 88246 45860
rect 86552 45722 86608 45724
rect 86632 45722 86688 45724
rect 86712 45722 86768 45724
rect 86792 45722 86848 45724
rect 86552 45670 86598 45722
rect 86598 45670 86608 45722
rect 86632 45670 86662 45722
rect 86662 45670 86674 45722
rect 86674 45670 86688 45722
rect 86712 45670 86726 45722
rect 86726 45670 86738 45722
rect 86738 45670 86768 45722
rect 86792 45670 86802 45722
rect 86802 45670 86848 45722
rect 86552 45668 86608 45670
rect 86632 45668 86688 45670
rect 86712 45668 86768 45670
rect 86792 45668 86848 45670
rect 85982 45468 85984 45488
rect 85984 45468 86036 45488
rect 86036 45468 86038 45488
rect 85982 45432 86038 45468
rect 86166 45332 86168 45352
rect 86168 45332 86220 45352
rect 86220 45332 86222 45352
rect 86166 45296 86222 45332
rect 85614 45160 85670 45216
rect 87288 45178 87344 45180
rect 87368 45178 87424 45180
rect 87448 45178 87504 45180
rect 87528 45178 87584 45180
rect 87288 45126 87334 45178
rect 87334 45126 87344 45178
rect 87368 45126 87398 45178
rect 87398 45126 87410 45178
rect 87410 45126 87424 45178
rect 87448 45126 87462 45178
rect 87462 45126 87474 45178
rect 87474 45126 87504 45178
rect 87528 45126 87538 45178
rect 87538 45126 87584 45178
rect 88190 45160 88246 45216
rect 87288 45124 87344 45126
rect 87368 45124 87424 45126
rect 87448 45124 87504 45126
rect 87528 45124 87584 45126
rect 87178 44788 87180 44808
rect 87180 44788 87232 44808
rect 87232 44788 87234 44808
rect 87178 44752 87234 44788
rect 86552 44634 86608 44636
rect 86632 44634 86688 44636
rect 86712 44634 86768 44636
rect 86792 44634 86848 44636
rect 86552 44582 86598 44634
rect 86598 44582 86608 44634
rect 86632 44582 86662 44634
rect 86662 44582 86674 44634
rect 86674 44582 86688 44634
rect 86712 44582 86726 44634
rect 86726 44582 86738 44634
rect 86738 44582 86768 44634
rect 86792 44582 86802 44634
rect 86802 44582 86848 44634
rect 86552 44580 86608 44582
rect 86632 44580 86688 44582
rect 86712 44580 86768 44582
rect 86792 44580 86848 44582
rect 88282 44480 88338 44536
rect 87288 44090 87344 44092
rect 87368 44090 87424 44092
rect 87448 44090 87504 44092
rect 87528 44090 87584 44092
rect 87288 44038 87334 44090
rect 87334 44038 87344 44090
rect 87368 44038 87398 44090
rect 87398 44038 87410 44090
rect 87410 44038 87424 44090
rect 87448 44038 87462 44090
rect 87462 44038 87474 44090
rect 87474 44038 87504 44090
rect 87528 44038 87538 44090
rect 87538 44038 87584 44090
rect 87288 44036 87344 44038
rect 87368 44036 87424 44038
rect 87448 44036 87504 44038
rect 87528 44036 87584 44038
rect 88282 43800 88338 43856
rect 85798 43528 85854 43584
rect 86552 43546 86608 43548
rect 86632 43546 86688 43548
rect 86712 43546 86768 43548
rect 86792 43546 86848 43548
rect 86552 43494 86598 43546
rect 86598 43494 86608 43546
rect 86632 43494 86662 43546
rect 86662 43494 86674 43546
rect 86674 43494 86688 43546
rect 86712 43494 86726 43546
rect 86726 43494 86738 43546
rect 86738 43494 86768 43546
rect 86792 43494 86802 43546
rect 86802 43494 86848 43546
rect 86552 43492 86608 43494
rect 86632 43492 86688 43494
rect 86712 43492 86768 43494
rect 86792 43492 86848 43494
rect 87288 43002 87344 43004
rect 87368 43002 87424 43004
rect 87448 43002 87504 43004
rect 87528 43002 87584 43004
rect 87288 42950 87334 43002
rect 87334 42950 87344 43002
rect 87368 42950 87398 43002
rect 87398 42950 87410 43002
rect 87410 42950 87424 43002
rect 87448 42950 87462 43002
rect 87462 42950 87474 43002
rect 87474 42950 87504 43002
rect 87528 42950 87538 43002
rect 87538 42950 87584 43002
rect 87288 42948 87344 42950
rect 87368 42948 87424 42950
rect 87448 42948 87504 42950
rect 87528 42948 87584 42950
rect 86350 42440 86406 42496
rect 86552 42458 86608 42460
rect 86632 42458 86688 42460
rect 86712 42458 86768 42460
rect 86792 42458 86848 42460
rect 86552 42406 86598 42458
rect 86598 42406 86608 42458
rect 86632 42406 86662 42458
rect 86662 42406 86674 42458
rect 86674 42406 86688 42458
rect 86712 42406 86726 42458
rect 86726 42406 86738 42458
rect 86738 42406 86768 42458
rect 86792 42406 86802 42458
rect 86802 42406 86848 42458
rect 88282 42440 88338 42496
rect 86552 42404 86608 42406
rect 86632 42404 86688 42406
rect 86712 42404 86768 42406
rect 86792 42404 86848 42406
rect 87288 41914 87344 41916
rect 87368 41914 87424 41916
rect 87448 41914 87504 41916
rect 87528 41914 87584 41916
rect 87288 41862 87334 41914
rect 87334 41862 87344 41914
rect 87368 41862 87398 41914
rect 87398 41862 87410 41914
rect 87410 41862 87424 41914
rect 87448 41862 87462 41914
rect 87462 41862 87474 41914
rect 87474 41862 87504 41914
rect 87528 41862 87538 41914
rect 87538 41862 87584 41914
rect 87288 41860 87344 41862
rect 87368 41860 87424 41862
rect 87448 41860 87504 41862
rect 87528 41860 87584 41862
rect 87178 41488 87234 41544
rect 86552 41370 86608 41372
rect 86632 41370 86688 41372
rect 86712 41370 86768 41372
rect 86792 41370 86848 41372
rect 86552 41318 86598 41370
rect 86598 41318 86608 41370
rect 86632 41318 86662 41370
rect 86662 41318 86674 41370
rect 86674 41318 86688 41370
rect 86712 41318 86726 41370
rect 86726 41318 86738 41370
rect 86738 41318 86768 41370
rect 86792 41318 86802 41370
rect 86802 41318 86848 41370
rect 86552 41316 86608 41318
rect 86632 41316 86688 41318
rect 86712 41316 86768 41318
rect 86792 41316 86848 41318
rect 88282 41080 88338 41136
rect 87288 40826 87344 40828
rect 87368 40826 87424 40828
rect 87448 40826 87504 40828
rect 87528 40826 87584 40828
rect 87288 40774 87334 40826
rect 87334 40774 87344 40826
rect 87368 40774 87398 40826
rect 87398 40774 87410 40826
rect 87410 40774 87424 40826
rect 87448 40774 87462 40826
rect 87462 40774 87474 40826
rect 87474 40774 87504 40826
rect 87528 40774 87538 40826
rect 87538 40774 87584 40826
rect 87288 40772 87344 40774
rect 87368 40772 87424 40774
rect 87448 40772 87504 40774
rect 87528 40772 87584 40774
rect 87914 40400 87970 40456
rect 88282 40400 88338 40456
rect 86552 40282 86608 40284
rect 86632 40282 86688 40284
rect 86712 40282 86768 40284
rect 86792 40282 86848 40284
rect 86552 40230 86598 40282
rect 86598 40230 86608 40282
rect 86632 40230 86662 40282
rect 86662 40230 86674 40282
rect 86674 40230 86688 40282
rect 86712 40230 86726 40282
rect 86726 40230 86738 40282
rect 86738 40230 86768 40282
rect 86792 40230 86802 40282
rect 86802 40230 86848 40282
rect 86552 40228 86608 40230
rect 86632 40228 86688 40230
rect 86712 40228 86768 40230
rect 86792 40228 86848 40230
rect 87288 39738 87344 39740
rect 87368 39738 87424 39740
rect 87448 39738 87504 39740
rect 87528 39738 87584 39740
rect 87288 39686 87334 39738
rect 87334 39686 87344 39738
rect 87368 39686 87398 39738
rect 87398 39686 87410 39738
rect 87410 39686 87424 39738
rect 87448 39686 87462 39738
rect 87462 39686 87474 39738
rect 87474 39686 87504 39738
rect 87528 39686 87538 39738
rect 87538 39686 87584 39738
rect 87288 39684 87344 39686
rect 87368 39684 87424 39686
rect 87448 39684 87504 39686
rect 87528 39684 87584 39686
rect 87178 39348 87180 39368
rect 87180 39348 87232 39368
rect 87232 39348 87234 39368
rect 87178 39312 87234 39348
rect 86552 39194 86608 39196
rect 86632 39194 86688 39196
rect 86712 39194 86768 39196
rect 86792 39194 86848 39196
rect 86552 39142 86598 39194
rect 86598 39142 86608 39194
rect 86632 39142 86662 39194
rect 86662 39142 86674 39194
rect 86674 39142 86688 39194
rect 86712 39142 86726 39194
rect 86726 39142 86738 39194
rect 86738 39142 86768 39194
rect 86792 39142 86802 39194
rect 86802 39142 86848 39194
rect 86552 39140 86608 39142
rect 86632 39140 86688 39142
rect 86712 39140 86768 39142
rect 86792 39140 86848 39142
rect 88282 39040 88338 39096
rect 87288 38650 87344 38652
rect 87368 38650 87424 38652
rect 87448 38650 87504 38652
rect 87528 38650 87584 38652
rect 87288 38598 87334 38650
rect 87334 38598 87344 38650
rect 87368 38598 87398 38650
rect 87398 38598 87410 38650
rect 87410 38598 87424 38650
rect 87448 38598 87462 38650
rect 87462 38598 87474 38650
rect 87474 38598 87504 38650
rect 87528 38598 87538 38650
rect 87538 38598 87584 38650
rect 87288 38596 87344 38598
rect 87368 38596 87424 38598
rect 87448 38596 87504 38598
rect 87528 38596 87584 38598
rect 88282 38360 88338 38416
rect 86552 38106 86608 38108
rect 86632 38106 86688 38108
rect 86712 38106 86768 38108
rect 86792 38106 86848 38108
rect 86552 38054 86598 38106
rect 86598 38054 86608 38106
rect 86632 38054 86662 38106
rect 86662 38054 86674 38106
rect 86674 38054 86688 38106
rect 86712 38054 86726 38106
rect 86726 38054 86738 38106
rect 86738 38054 86768 38106
rect 86792 38054 86802 38106
rect 86802 38054 86848 38106
rect 86552 38052 86608 38054
rect 86632 38052 86688 38054
rect 86712 38052 86768 38054
rect 86792 38052 86848 38054
rect 87288 37562 87344 37564
rect 87368 37562 87424 37564
rect 87448 37562 87504 37564
rect 87528 37562 87584 37564
rect 87288 37510 87334 37562
rect 87334 37510 87344 37562
rect 87368 37510 87398 37562
rect 87398 37510 87410 37562
rect 87410 37510 87424 37562
rect 87448 37510 87462 37562
rect 87462 37510 87474 37562
rect 87474 37510 87504 37562
rect 87528 37510 87538 37562
rect 87538 37510 87584 37562
rect 87288 37508 87344 37510
rect 87368 37508 87424 37510
rect 87448 37508 87504 37510
rect 87528 37508 87584 37510
rect 86350 37000 86406 37056
rect 86552 37018 86608 37020
rect 86632 37018 86688 37020
rect 86712 37018 86768 37020
rect 86792 37018 86848 37020
rect 86552 36966 86598 37018
rect 86598 36966 86608 37018
rect 86632 36966 86662 37018
rect 86662 36966 86674 37018
rect 86674 36966 86688 37018
rect 86712 36966 86726 37018
rect 86726 36966 86738 37018
rect 86738 36966 86768 37018
rect 86792 36966 86802 37018
rect 86802 36966 86848 37018
rect 88282 37000 88338 37056
rect 86552 36964 86608 36966
rect 86632 36964 86688 36966
rect 86712 36964 86768 36966
rect 86792 36964 86848 36966
rect 87288 36474 87344 36476
rect 87368 36474 87424 36476
rect 87448 36474 87504 36476
rect 87528 36474 87584 36476
rect 87288 36422 87334 36474
rect 87334 36422 87344 36474
rect 87368 36422 87398 36474
rect 87398 36422 87410 36474
rect 87410 36422 87424 36474
rect 87448 36422 87462 36474
rect 87462 36422 87474 36474
rect 87474 36422 87504 36474
rect 87528 36422 87538 36474
rect 87538 36422 87584 36474
rect 87288 36420 87344 36422
rect 87368 36420 87424 36422
rect 87448 36420 87504 36422
rect 87528 36420 87584 36422
rect 86552 35930 86608 35932
rect 86632 35930 86688 35932
rect 86712 35930 86768 35932
rect 86792 35930 86848 35932
rect 86552 35878 86598 35930
rect 86598 35878 86608 35930
rect 86632 35878 86662 35930
rect 86662 35878 86674 35930
rect 86674 35878 86688 35930
rect 86712 35878 86726 35930
rect 86726 35878 86738 35930
rect 86738 35878 86768 35930
rect 86792 35878 86802 35930
rect 86802 35878 86848 35930
rect 86552 35876 86608 35878
rect 86632 35876 86688 35878
rect 86712 35876 86768 35878
rect 86792 35876 86848 35878
rect 88558 35640 88614 35696
rect 87288 35386 87344 35388
rect 87368 35386 87424 35388
rect 87448 35386 87504 35388
rect 87528 35386 87584 35388
rect 87288 35334 87334 35386
rect 87334 35334 87344 35386
rect 87368 35334 87398 35386
rect 87398 35334 87410 35386
rect 87410 35334 87424 35386
rect 87448 35334 87462 35386
rect 87462 35334 87474 35386
rect 87474 35334 87504 35386
rect 87528 35334 87538 35386
rect 87538 35334 87584 35386
rect 87288 35332 87344 35334
rect 87368 35332 87424 35334
rect 87448 35332 87504 35334
rect 87528 35332 87584 35334
rect 88282 34960 88338 35016
rect 86350 34824 86406 34880
rect 86552 34842 86608 34844
rect 86632 34842 86688 34844
rect 86712 34842 86768 34844
rect 86792 34842 86848 34844
rect 86552 34790 86598 34842
rect 86598 34790 86608 34842
rect 86632 34790 86662 34842
rect 86662 34790 86674 34842
rect 86674 34790 86688 34842
rect 86712 34790 86726 34842
rect 86726 34790 86738 34842
rect 86738 34790 86768 34842
rect 86792 34790 86802 34842
rect 86802 34790 86848 34842
rect 86552 34788 86608 34790
rect 86632 34788 86688 34790
rect 86712 34788 86768 34790
rect 86792 34788 86848 34790
rect 87288 34298 87344 34300
rect 87368 34298 87424 34300
rect 87448 34298 87504 34300
rect 87528 34298 87584 34300
rect 87288 34246 87334 34298
rect 87334 34246 87344 34298
rect 87368 34246 87398 34298
rect 87398 34246 87410 34298
rect 87410 34246 87424 34298
rect 87448 34246 87462 34298
rect 87462 34246 87474 34298
rect 87474 34246 87504 34298
rect 87528 34246 87538 34298
rect 87538 34246 87584 34298
rect 87288 34244 87344 34246
rect 87368 34244 87424 34246
rect 87448 34244 87504 34246
rect 87528 34244 87584 34246
rect 86350 33736 86406 33792
rect 86552 33754 86608 33756
rect 86632 33754 86688 33756
rect 86712 33754 86768 33756
rect 86792 33754 86848 33756
rect 86552 33702 86598 33754
rect 86598 33702 86608 33754
rect 86632 33702 86662 33754
rect 86662 33702 86674 33754
rect 86674 33702 86688 33754
rect 86712 33702 86726 33754
rect 86726 33702 86738 33754
rect 86738 33702 86768 33754
rect 86792 33702 86802 33754
rect 86802 33702 86848 33754
rect 86552 33700 86608 33702
rect 86632 33700 86688 33702
rect 86712 33700 86768 33702
rect 86792 33700 86848 33702
rect 88282 33600 88338 33656
rect 87288 33210 87344 33212
rect 87368 33210 87424 33212
rect 87448 33210 87504 33212
rect 87528 33210 87584 33212
rect 87288 33158 87334 33210
rect 87334 33158 87344 33210
rect 87368 33158 87398 33210
rect 87398 33158 87410 33210
rect 87410 33158 87424 33210
rect 87448 33158 87462 33210
rect 87462 33158 87474 33210
rect 87474 33158 87504 33210
rect 87528 33158 87538 33210
rect 87538 33158 87584 33210
rect 87288 33156 87344 33158
rect 87368 33156 87424 33158
rect 87448 33156 87504 33158
rect 87528 33156 87584 33158
rect 88558 32920 88614 32976
rect 86552 32666 86608 32668
rect 86632 32666 86688 32668
rect 86712 32666 86768 32668
rect 86792 32666 86848 32668
rect 86552 32614 86598 32666
rect 86598 32614 86608 32666
rect 86632 32614 86662 32666
rect 86662 32614 86674 32666
rect 86674 32614 86688 32666
rect 86712 32614 86726 32666
rect 86726 32614 86738 32666
rect 86738 32614 86768 32666
rect 86792 32614 86802 32666
rect 86802 32614 86848 32666
rect 86552 32612 86608 32614
rect 86632 32612 86688 32614
rect 86712 32612 86768 32614
rect 86792 32612 86848 32614
rect 87288 32122 87344 32124
rect 87368 32122 87424 32124
rect 87448 32122 87504 32124
rect 87528 32122 87584 32124
rect 87288 32070 87334 32122
rect 87334 32070 87344 32122
rect 87368 32070 87398 32122
rect 87398 32070 87410 32122
rect 87410 32070 87424 32122
rect 87448 32070 87462 32122
rect 87462 32070 87474 32122
rect 87474 32070 87504 32122
rect 87528 32070 87538 32122
rect 87538 32070 87584 32122
rect 87288 32068 87344 32070
rect 87368 32068 87424 32070
rect 87448 32068 87504 32070
rect 87528 32068 87584 32070
rect 86350 31560 86406 31616
rect 86552 31578 86608 31580
rect 86632 31578 86688 31580
rect 86712 31578 86768 31580
rect 86792 31578 86848 31580
rect 86552 31526 86598 31578
rect 86598 31526 86608 31578
rect 86632 31526 86662 31578
rect 86662 31526 86674 31578
rect 86674 31526 86688 31578
rect 86712 31526 86726 31578
rect 86726 31526 86738 31578
rect 86738 31526 86768 31578
rect 86792 31526 86802 31578
rect 86802 31526 86848 31578
rect 88282 31560 88338 31616
rect 86552 31524 86608 31526
rect 86632 31524 86688 31526
rect 86712 31524 86768 31526
rect 86792 31524 86848 31526
rect 87288 31034 87344 31036
rect 87368 31034 87424 31036
rect 87448 31034 87504 31036
rect 87528 31034 87584 31036
rect 87288 30982 87334 31034
rect 87334 30982 87344 31034
rect 87368 30982 87398 31034
rect 87398 30982 87410 31034
rect 87410 30982 87424 31034
rect 87448 30982 87462 31034
rect 87462 30982 87474 31034
rect 87474 30982 87504 31034
rect 87528 30982 87538 31034
rect 87538 30982 87584 31034
rect 87288 30980 87344 30982
rect 87368 30980 87424 30982
rect 87448 30980 87504 30982
rect 87528 30980 87584 30982
rect 86552 30490 86608 30492
rect 86632 30490 86688 30492
rect 86712 30490 86768 30492
rect 86792 30490 86848 30492
rect 86552 30438 86598 30490
rect 86598 30438 86608 30490
rect 86632 30438 86662 30490
rect 86662 30438 86674 30490
rect 86674 30438 86688 30490
rect 86712 30438 86726 30490
rect 86726 30438 86738 30490
rect 86738 30438 86768 30490
rect 86792 30438 86802 30490
rect 86802 30438 86848 30490
rect 86552 30436 86608 30438
rect 86632 30436 86688 30438
rect 86712 30436 86768 30438
rect 86792 30436 86848 30438
rect 88558 30200 88614 30256
rect 87288 29946 87344 29948
rect 87368 29946 87424 29948
rect 87448 29946 87504 29948
rect 87528 29946 87584 29948
rect 87288 29894 87334 29946
rect 87334 29894 87344 29946
rect 87368 29894 87398 29946
rect 87398 29894 87410 29946
rect 87410 29894 87424 29946
rect 87448 29894 87462 29946
rect 87462 29894 87474 29946
rect 87474 29894 87504 29946
rect 87528 29894 87538 29946
rect 87538 29894 87584 29946
rect 87288 29892 87344 29894
rect 87368 29892 87424 29894
rect 87448 29892 87504 29894
rect 87528 29892 87584 29894
rect 88282 29540 88338 29576
rect 88282 29520 88284 29540
rect 88284 29520 88336 29540
rect 88336 29520 88338 29540
rect 86350 29384 86406 29440
rect 86552 29402 86608 29404
rect 86632 29402 86688 29404
rect 86712 29402 86768 29404
rect 86792 29402 86848 29404
rect 86552 29350 86598 29402
rect 86598 29350 86608 29402
rect 86632 29350 86662 29402
rect 86662 29350 86674 29402
rect 86674 29350 86688 29402
rect 86712 29350 86726 29402
rect 86726 29350 86738 29402
rect 86738 29350 86768 29402
rect 86792 29350 86802 29402
rect 86802 29350 86848 29402
rect 86552 29348 86608 29350
rect 86632 29348 86688 29350
rect 86712 29348 86768 29350
rect 86792 29348 86848 29350
rect 87288 28858 87344 28860
rect 87368 28858 87424 28860
rect 87448 28858 87504 28860
rect 87528 28858 87584 28860
rect 87288 28806 87334 28858
rect 87334 28806 87344 28858
rect 87368 28806 87398 28858
rect 87398 28806 87410 28858
rect 87410 28806 87424 28858
rect 87448 28806 87462 28858
rect 87462 28806 87474 28858
rect 87474 28806 87504 28858
rect 87528 28806 87538 28858
rect 87538 28806 87584 28858
rect 87288 28804 87344 28806
rect 87368 28804 87424 28806
rect 87448 28804 87504 28806
rect 87528 28804 87584 28806
rect 86350 28296 86406 28352
rect 86552 28314 86608 28316
rect 86632 28314 86688 28316
rect 86712 28314 86768 28316
rect 86792 28314 86848 28316
rect 86552 28262 86598 28314
rect 86598 28262 86608 28314
rect 86632 28262 86662 28314
rect 86662 28262 86674 28314
rect 86674 28262 86688 28314
rect 86712 28262 86726 28314
rect 86726 28262 86738 28314
rect 86738 28262 86768 28314
rect 86792 28262 86802 28314
rect 86802 28262 86848 28314
rect 86552 28260 86608 28262
rect 86632 28260 86688 28262
rect 86712 28260 86768 28262
rect 86792 28260 86848 28262
rect 88190 28160 88246 28216
rect 87288 27770 87344 27772
rect 87368 27770 87424 27772
rect 87448 27770 87504 27772
rect 87528 27770 87584 27772
rect 87288 27718 87334 27770
rect 87334 27718 87344 27770
rect 87368 27718 87398 27770
rect 87398 27718 87410 27770
rect 87410 27718 87424 27770
rect 87448 27718 87462 27770
rect 87462 27718 87474 27770
rect 87474 27718 87504 27770
rect 87528 27718 87538 27770
rect 87538 27718 87584 27770
rect 87288 27716 87344 27718
rect 87368 27716 87424 27718
rect 87448 27716 87504 27718
rect 87528 27716 87584 27718
rect 88926 27480 88982 27536
rect 86552 27226 86608 27228
rect 86632 27226 86688 27228
rect 86712 27226 86768 27228
rect 86792 27226 86848 27228
rect 86552 27174 86598 27226
rect 86598 27174 86608 27226
rect 86632 27174 86662 27226
rect 86662 27174 86674 27226
rect 86674 27174 86688 27226
rect 86712 27174 86726 27226
rect 86726 27174 86738 27226
rect 86738 27174 86768 27226
rect 86792 27174 86802 27226
rect 86802 27174 86848 27226
rect 86552 27172 86608 27174
rect 86632 27172 86688 27174
rect 86712 27172 86768 27174
rect 86792 27172 86848 27174
rect 87288 26682 87344 26684
rect 87368 26682 87424 26684
rect 87448 26682 87504 26684
rect 87528 26682 87584 26684
rect 87288 26630 87334 26682
rect 87334 26630 87344 26682
rect 87368 26630 87398 26682
rect 87398 26630 87410 26682
rect 87410 26630 87424 26682
rect 87448 26630 87462 26682
rect 87462 26630 87474 26682
rect 87474 26630 87504 26682
rect 87528 26630 87538 26682
rect 87538 26630 87584 26682
rect 87288 26628 87344 26630
rect 87368 26628 87424 26630
rect 87448 26628 87504 26630
rect 87528 26628 87584 26630
rect 87730 26256 87786 26312
rect 86552 26138 86608 26140
rect 86632 26138 86688 26140
rect 86712 26138 86768 26140
rect 86792 26138 86848 26140
rect 86552 26086 86598 26138
rect 86598 26086 86608 26138
rect 86632 26086 86662 26138
rect 86662 26086 86674 26138
rect 86674 26086 86688 26138
rect 86712 26086 86726 26138
rect 86726 26086 86738 26138
rect 86738 26086 86768 26138
rect 86792 26086 86802 26138
rect 86802 26086 86848 26138
rect 88190 26120 88246 26176
rect 86552 26084 86608 26086
rect 86632 26084 86688 26086
rect 86712 26084 86768 26086
rect 86792 26084 86848 26086
rect 87288 25594 87344 25596
rect 87368 25594 87424 25596
rect 87448 25594 87504 25596
rect 87528 25594 87584 25596
rect 87288 25542 87334 25594
rect 87334 25542 87344 25594
rect 87368 25542 87398 25594
rect 87398 25542 87410 25594
rect 87410 25542 87424 25594
rect 87448 25542 87462 25594
rect 87462 25542 87474 25594
rect 87474 25542 87504 25594
rect 87528 25542 87538 25594
rect 87538 25542 87584 25594
rect 87288 25540 87344 25542
rect 87368 25540 87424 25542
rect 87448 25540 87504 25542
rect 87528 25540 87584 25542
rect 87730 25168 87786 25224
rect 86552 25050 86608 25052
rect 86632 25050 86688 25052
rect 86712 25050 86768 25052
rect 86792 25050 86848 25052
rect 86552 24998 86598 25050
rect 86598 24998 86608 25050
rect 86632 24998 86662 25050
rect 86662 24998 86674 25050
rect 86674 24998 86688 25050
rect 86712 24998 86726 25050
rect 86726 24998 86738 25050
rect 86738 24998 86768 25050
rect 86792 24998 86802 25050
rect 86802 24998 86848 25050
rect 86552 24996 86608 24998
rect 86632 24996 86688 24998
rect 86712 24996 86768 24998
rect 86792 24996 86848 24998
rect 88558 24760 88614 24816
rect 87288 24506 87344 24508
rect 87368 24506 87424 24508
rect 87448 24506 87504 24508
rect 87528 24506 87584 24508
rect 87288 24454 87334 24506
rect 87334 24454 87344 24506
rect 87368 24454 87398 24506
rect 87398 24454 87410 24506
rect 87410 24454 87424 24506
rect 87448 24454 87462 24506
rect 87462 24454 87474 24506
rect 87474 24454 87504 24506
rect 87528 24454 87538 24506
rect 87538 24454 87584 24506
rect 87288 24452 87344 24454
rect 87368 24452 87424 24454
rect 87448 24452 87504 24454
rect 87528 24452 87584 24454
rect 87730 24080 87786 24136
rect 88282 24100 88338 24136
rect 88282 24080 88284 24100
rect 88284 24080 88336 24100
rect 88336 24080 88338 24100
rect 86552 23962 86608 23964
rect 86632 23962 86688 23964
rect 86712 23962 86768 23964
rect 86792 23962 86848 23964
rect 86552 23910 86598 23962
rect 86598 23910 86608 23962
rect 86632 23910 86662 23962
rect 86662 23910 86674 23962
rect 86674 23910 86688 23962
rect 86712 23910 86726 23962
rect 86726 23910 86738 23962
rect 86738 23910 86768 23962
rect 86792 23910 86802 23962
rect 86802 23910 86848 23962
rect 86552 23908 86608 23910
rect 86632 23908 86688 23910
rect 86712 23908 86768 23910
rect 86792 23908 86848 23910
rect 87288 23418 87344 23420
rect 87368 23418 87424 23420
rect 87448 23418 87504 23420
rect 87528 23418 87584 23420
rect 87288 23366 87334 23418
rect 87334 23366 87344 23418
rect 87368 23366 87398 23418
rect 87398 23366 87410 23418
rect 87410 23366 87424 23418
rect 87448 23366 87462 23418
rect 87462 23366 87474 23418
rect 87474 23366 87504 23418
rect 87528 23366 87538 23418
rect 87538 23366 87584 23418
rect 87288 23364 87344 23366
rect 87368 23364 87424 23366
rect 87448 23364 87504 23366
rect 87528 23364 87584 23366
rect 86350 22856 86406 22912
rect 86552 22874 86608 22876
rect 86632 22874 86688 22876
rect 86712 22874 86768 22876
rect 86792 22874 86848 22876
rect 86552 22822 86598 22874
rect 86598 22822 86608 22874
rect 86632 22822 86662 22874
rect 86662 22822 86674 22874
rect 86674 22822 86688 22874
rect 86712 22822 86726 22874
rect 86726 22822 86738 22874
rect 86738 22822 86768 22874
rect 86792 22822 86802 22874
rect 86802 22822 86848 22874
rect 86552 22820 86608 22822
rect 86632 22820 86688 22822
rect 86712 22820 86768 22822
rect 86792 22820 86848 22822
rect 88282 22720 88338 22776
rect 87288 22330 87344 22332
rect 87368 22330 87424 22332
rect 87448 22330 87504 22332
rect 87528 22330 87584 22332
rect 87288 22278 87334 22330
rect 87334 22278 87344 22330
rect 87368 22278 87398 22330
rect 87398 22278 87410 22330
rect 87410 22278 87424 22330
rect 87448 22278 87462 22330
rect 87462 22278 87474 22330
rect 87474 22278 87504 22330
rect 87528 22278 87538 22330
rect 87538 22278 87584 22330
rect 87288 22276 87344 22278
rect 87368 22276 87424 22278
rect 87448 22276 87504 22278
rect 87528 22276 87584 22278
rect 88558 22040 88614 22096
rect 86552 21786 86608 21788
rect 86632 21786 86688 21788
rect 86712 21786 86768 21788
rect 86792 21786 86848 21788
rect 86552 21734 86598 21786
rect 86598 21734 86608 21786
rect 86632 21734 86662 21786
rect 86662 21734 86674 21786
rect 86674 21734 86688 21786
rect 86712 21734 86726 21786
rect 86726 21734 86738 21786
rect 86738 21734 86768 21786
rect 86792 21734 86802 21786
rect 86802 21734 86848 21786
rect 86552 21732 86608 21734
rect 86632 21732 86688 21734
rect 86712 21732 86768 21734
rect 86792 21732 86848 21734
rect 87288 21242 87344 21244
rect 87368 21242 87424 21244
rect 87448 21242 87504 21244
rect 87528 21242 87584 21244
rect 87288 21190 87334 21242
rect 87334 21190 87344 21242
rect 87368 21190 87398 21242
rect 87398 21190 87410 21242
rect 87410 21190 87424 21242
rect 87448 21190 87462 21242
rect 87462 21190 87474 21242
rect 87474 21190 87504 21242
rect 87528 21190 87538 21242
rect 87538 21190 87584 21242
rect 87288 21188 87344 21190
rect 87368 21188 87424 21190
rect 87448 21188 87504 21190
rect 87528 21188 87584 21190
rect 86552 20698 86608 20700
rect 86632 20698 86688 20700
rect 86712 20698 86768 20700
rect 86792 20698 86848 20700
rect 86552 20646 86598 20698
rect 86598 20646 86608 20698
rect 86632 20646 86662 20698
rect 86662 20646 86674 20698
rect 86674 20646 86688 20698
rect 86712 20646 86726 20698
rect 86726 20646 86738 20698
rect 86738 20646 86768 20698
rect 86792 20646 86802 20698
rect 86802 20646 86848 20698
rect 88558 20680 88614 20736
rect 86552 20644 86608 20646
rect 86632 20644 86688 20646
rect 86712 20644 86768 20646
rect 86792 20644 86848 20646
rect 87288 20154 87344 20156
rect 87368 20154 87424 20156
rect 87448 20154 87504 20156
rect 87528 20154 87584 20156
rect 87288 20102 87334 20154
rect 87334 20102 87344 20154
rect 87368 20102 87398 20154
rect 87398 20102 87410 20154
rect 87410 20102 87424 20154
rect 87448 20102 87462 20154
rect 87462 20102 87474 20154
rect 87474 20102 87504 20154
rect 87528 20102 87538 20154
rect 87538 20102 87584 20154
rect 87288 20100 87344 20102
rect 87368 20100 87424 20102
rect 87448 20100 87504 20102
rect 87528 20100 87584 20102
rect 87730 19728 87786 19784
rect 86552 19610 86608 19612
rect 86632 19610 86688 19612
rect 86712 19610 86768 19612
rect 86792 19610 86848 19612
rect 86552 19558 86598 19610
rect 86598 19558 86608 19610
rect 86632 19558 86662 19610
rect 86662 19558 86674 19610
rect 86674 19558 86688 19610
rect 86712 19558 86726 19610
rect 86726 19558 86738 19610
rect 86738 19558 86768 19610
rect 86792 19558 86802 19610
rect 86802 19558 86848 19610
rect 86552 19556 86608 19558
rect 86632 19556 86688 19558
rect 86712 19556 86768 19558
rect 86792 19556 86848 19558
rect 88558 19320 88614 19376
rect 87288 19066 87344 19068
rect 87368 19066 87424 19068
rect 87448 19066 87504 19068
rect 87528 19066 87584 19068
rect 87288 19014 87334 19066
rect 87334 19014 87344 19066
rect 87368 19014 87398 19066
rect 87398 19014 87410 19066
rect 87410 19014 87424 19066
rect 87448 19014 87462 19066
rect 87462 19014 87474 19066
rect 87474 19014 87504 19066
rect 87528 19014 87538 19066
rect 87538 19014 87584 19066
rect 87288 19012 87344 19014
rect 87368 19012 87424 19014
rect 87448 19012 87504 19014
rect 87528 19012 87584 19014
rect 87730 18640 87786 18696
rect 88282 18660 88338 18696
rect 88282 18640 88284 18660
rect 88284 18640 88336 18660
rect 88336 18640 88338 18660
rect 86552 18522 86608 18524
rect 86632 18522 86688 18524
rect 86712 18522 86768 18524
rect 86792 18522 86848 18524
rect 86552 18470 86598 18522
rect 86598 18470 86608 18522
rect 86632 18470 86662 18522
rect 86662 18470 86674 18522
rect 86674 18470 86688 18522
rect 86712 18470 86726 18522
rect 86726 18470 86738 18522
rect 86738 18470 86768 18522
rect 86792 18470 86802 18522
rect 86802 18470 86848 18522
rect 86552 18468 86608 18470
rect 86632 18468 86688 18470
rect 86712 18468 86768 18470
rect 86792 18468 86848 18470
rect 87288 17978 87344 17980
rect 87368 17978 87424 17980
rect 87448 17978 87504 17980
rect 87528 17978 87584 17980
rect 87288 17926 87334 17978
rect 87334 17926 87344 17978
rect 87368 17926 87398 17978
rect 87398 17926 87410 17978
rect 87410 17926 87424 17978
rect 87448 17926 87462 17978
rect 87462 17926 87474 17978
rect 87474 17926 87504 17978
rect 87528 17926 87538 17978
rect 87538 17926 87584 17978
rect 87288 17924 87344 17926
rect 87368 17924 87424 17926
rect 87448 17924 87504 17926
rect 87528 17924 87584 17926
rect 86350 17416 86406 17472
rect 86552 17434 86608 17436
rect 86632 17434 86688 17436
rect 86712 17434 86768 17436
rect 86792 17434 86848 17436
rect 86552 17382 86598 17434
rect 86598 17382 86608 17434
rect 86632 17382 86662 17434
rect 86662 17382 86674 17434
rect 86674 17382 86688 17434
rect 86712 17382 86726 17434
rect 86726 17382 86738 17434
rect 86738 17382 86768 17434
rect 86792 17382 86802 17434
rect 86802 17382 86848 17434
rect 86552 17380 86608 17382
rect 86632 17380 86688 17382
rect 86712 17380 86768 17382
rect 86792 17380 86848 17382
rect 88190 17280 88246 17336
rect 87288 16890 87344 16892
rect 87368 16890 87424 16892
rect 87448 16890 87504 16892
rect 87528 16890 87584 16892
rect 87288 16838 87334 16890
rect 87334 16838 87344 16890
rect 87368 16838 87398 16890
rect 87398 16838 87410 16890
rect 87410 16838 87424 16890
rect 87448 16838 87462 16890
rect 87462 16838 87474 16890
rect 87474 16838 87504 16890
rect 87528 16838 87538 16890
rect 87538 16838 87584 16890
rect 87288 16836 87344 16838
rect 87368 16836 87424 16838
rect 87448 16836 87504 16838
rect 87528 16836 87584 16838
rect 88558 16600 88614 16656
rect 88006 16464 88062 16520
rect 86552 16346 86608 16348
rect 86632 16346 86688 16348
rect 86712 16346 86768 16348
rect 86792 16346 86848 16348
rect 86552 16294 86598 16346
rect 86598 16294 86608 16346
rect 86632 16294 86662 16346
rect 86662 16294 86674 16346
rect 86674 16294 86688 16346
rect 86712 16294 86726 16346
rect 86726 16294 86738 16346
rect 86738 16294 86768 16346
rect 86792 16294 86802 16346
rect 86802 16294 86848 16346
rect 86552 16292 86608 16294
rect 86632 16292 86688 16294
rect 86712 16292 86768 16294
rect 86792 16292 86848 16294
rect 87288 15802 87344 15804
rect 87368 15802 87424 15804
rect 87448 15802 87504 15804
rect 87528 15802 87584 15804
rect 87288 15750 87334 15802
rect 87334 15750 87344 15802
rect 87368 15750 87398 15802
rect 87398 15750 87410 15802
rect 87410 15750 87424 15802
rect 87448 15750 87462 15802
rect 87462 15750 87474 15802
rect 87474 15750 87504 15802
rect 87528 15750 87538 15802
rect 87538 15750 87584 15802
rect 87288 15748 87344 15750
rect 87368 15748 87424 15750
rect 87448 15748 87504 15750
rect 87528 15748 87584 15750
rect 86552 15258 86608 15260
rect 86632 15258 86688 15260
rect 86712 15258 86768 15260
rect 86792 15258 86848 15260
rect 86552 15206 86598 15258
rect 86598 15206 86608 15258
rect 86632 15206 86662 15258
rect 86662 15206 86674 15258
rect 86674 15206 86688 15258
rect 86712 15206 86726 15258
rect 86726 15206 86738 15258
rect 86738 15206 86768 15258
rect 86792 15206 86802 15258
rect 86802 15206 86848 15258
rect 88558 15240 88614 15296
rect 86552 15204 86608 15206
rect 86632 15204 86688 15206
rect 86712 15204 86768 15206
rect 86792 15204 86848 15206
rect 87288 14714 87344 14716
rect 87368 14714 87424 14716
rect 87448 14714 87504 14716
rect 87528 14714 87584 14716
rect 87288 14662 87334 14714
rect 87334 14662 87344 14714
rect 87368 14662 87398 14714
rect 87398 14662 87410 14714
rect 87410 14662 87424 14714
rect 87448 14662 87462 14714
rect 87462 14662 87474 14714
rect 87474 14662 87504 14714
rect 87528 14662 87538 14714
rect 87538 14662 87584 14714
rect 87288 14660 87344 14662
rect 87368 14660 87424 14662
rect 87448 14660 87504 14662
rect 87528 14660 87584 14662
rect 88006 14560 88062 14616
rect 86552 14170 86608 14172
rect 86632 14170 86688 14172
rect 86712 14170 86768 14172
rect 86792 14170 86848 14172
rect 86552 14118 86598 14170
rect 86598 14118 86608 14170
rect 86632 14118 86662 14170
rect 86662 14118 86674 14170
rect 86674 14118 86688 14170
rect 86712 14118 86726 14170
rect 86726 14118 86738 14170
rect 86738 14118 86768 14170
rect 86792 14118 86802 14170
rect 86802 14118 86848 14170
rect 86552 14116 86608 14118
rect 86632 14116 86688 14118
rect 86712 14116 86768 14118
rect 86792 14116 86848 14118
rect 87288 13626 87344 13628
rect 87368 13626 87424 13628
rect 87448 13626 87504 13628
rect 87528 13626 87584 13628
rect 87288 13574 87334 13626
rect 87334 13574 87344 13626
rect 87368 13574 87398 13626
rect 87398 13574 87410 13626
rect 87410 13574 87424 13626
rect 87448 13574 87462 13626
rect 87462 13574 87474 13626
rect 87474 13574 87504 13626
rect 87528 13574 87538 13626
rect 87538 13574 87584 13626
rect 87288 13572 87344 13574
rect 87368 13572 87424 13574
rect 87448 13572 87504 13574
rect 87528 13572 87584 13574
rect 86552 13082 86608 13084
rect 86632 13082 86688 13084
rect 86712 13082 86768 13084
rect 86792 13082 86848 13084
rect 86552 13030 86598 13082
rect 86598 13030 86608 13082
rect 86632 13030 86662 13082
rect 86662 13030 86674 13082
rect 86674 13030 86688 13082
rect 86712 13030 86726 13082
rect 86726 13030 86738 13082
rect 86738 13030 86768 13082
rect 86792 13030 86802 13082
rect 86802 13030 86848 13082
rect 86552 13028 86608 13030
rect 86632 13028 86688 13030
rect 86712 13028 86768 13030
rect 86792 13028 86848 13030
rect 88190 13200 88246 13256
rect 87288 12538 87344 12540
rect 87368 12538 87424 12540
rect 87448 12538 87504 12540
rect 87528 12538 87584 12540
rect 87288 12486 87334 12538
rect 87334 12486 87344 12538
rect 87368 12486 87398 12538
rect 87398 12486 87410 12538
rect 87410 12486 87424 12538
rect 87448 12486 87462 12538
rect 87462 12486 87474 12538
rect 87474 12486 87504 12538
rect 87528 12486 87538 12538
rect 87538 12486 87584 12538
rect 88558 12520 88614 12576
rect 87288 12484 87344 12486
rect 87368 12484 87424 12486
rect 87448 12484 87504 12486
rect 87528 12484 87584 12486
rect 86552 11994 86608 11996
rect 86632 11994 86688 11996
rect 86712 11994 86768 11996
rect 86792 11994 86848 11996
rect 86552 11942 86598 11994
rect 86598 11942 86608 11994
rect 86632 11942 86662 11994
rect 86662 11942 86674 11994
rect 86674 11942 86688 11994
rect 86712 11942 86726 11994
rect 86726 11942 86738 11994
rect 86738 11942 86768 11994
rect 86792 11942 86802 11994
rect 86802 11942 86848 11994
rect 86552 11940 86608 11942
rect 86632 11940 86688 11942
rect 86712 11940 86768 11942
rect 86792 11940 86848 11942
rect 87288 11450 87344 11452
rect 87368 11450 87424 11452
rect 87448 11450 87504 11452
rect 87528 11450 87584 11452
rect 87288 11398 87334 11450
rect 87334 11398 87344 11450
rect 87368 11398 87398 11450
rect 87398 11398 87410 11450
rect 87410 11398 87424 11450
rect 87448 11398 87462 11450
rect 87462 11398 87474 11450
rect 87474 11398 87504 11450
rect 87528 11398 87538 11450
rect 87538 11398 87584 11450
rect 87288 11396 87344 11398
rect 87368 11396 87424 11398
rect 87448 11396 87504 11398
rect 87528 11396 87584 11398
rect 86552 10906 86608 10908
rect 86632 10906 86688 10908
rect 86712 10906 86768 10908
rect 86792 10906 86848 10908
rect 86552 10854 86598 10906
rect 86598 10854 86608 10906
rect 86632 10854 86662 10906
rect 86662 10854 86674 10906
rect 86674 10854 86688 10906
rect 86712 10854 86726 10906
rect 86726 10854 86738 10906
rect 86738 10854 86768 10906
rect 86792 10854 86802 10906
rect 86802 10854 86848 10906
rect 86552 10852 86608 10854
rect 86632 10852 86688 10854
rect 86712 10852 86768 10854
rect 86792 10852 86848 10854
rect 88374 10524 88376 10536
rect 88376 10524 88428 10536
rect 88428 10524 88430 10536
rect 88374 10480 88430 10524
rect 87288 10362 87344 10364
rect 87368 10362 87424 10364
rect 87448 10362 87504 10364
rect 87528 10362 87584 10364
rect 87288 10310 87334 10362
rect 87334 10310 87344 10362
rect 87368 10310 87398 10362
rect 87398 10310 87410 10362
rect 87410 10310 87424 10362
rect 87448 10310 87462 10362
rect 87462 10310 87474 10362
rect 87474 10310 87504 10362
rect 87528 10310 87538 10362
rect 87538 10310 87584 10362
rect 87288 10308 87344 10310
rect 87368 10308 87424 10310
rect 87448 10308 87504 10310
rect 87528 10308 87584 10310
rect 86552 9818 86608 9820
rect 86632 9818 86688 9820
rect 86712 9818 86768 9820
rect 86792 9818 86848 9820
rect 86552 9766 86598 9818
rect 86598 9766 86608 9818
rect 86632 9766 86662 9818
rect 86662 9766 86674 9818
rect 86674 9766 86688 9818
rect 86712 9766 86726 9818
rect 86726 9766 86738 9818
rect 86738 9766 86768 9818
rect 86792 9766 86802 9818
rect 86802 9766 86848 9818
rect 88558 9800 88614 9856
rect 86552 9764 86608 9766
rect 86632 9764 86688 9766
rect 86712 9764 86768 9766
rect 86792 9764 86848 9766
rect 87288 9274 87344 9276
rect 87368 9274 87424 9276
rect 87448 9274 87504 9276
rect 87528 9274 87584 9276
rect 87288 9222 87334 9274
rect 87334 9222 87344 9274
rect 87368 9222 87398 9274
rect 87398 9222 87410 9274
rect 87410 9222 87424 9274
rect 87448 9222 87462 9274
rect 87462 9222 87474 9274
rect 87474 9222 87504 9274
rect 87528 9222 87538 9274
rect 87538 9222 87584 9274
rect 87288 9220 87344 9222
rect 87368 9220 87424 9222
rect 87448 9220 87504 9222
rect 87528 9220 87584 9222
rect 86552 8730 86608 8732
rect 86632 8730 86688 8732
rect 86712 8730 86768 8732
rect 86792 8730 86848 8732
rect 86552 8678 86598 8730
rect 86598 8678 86608 8730
rect 86632 8678 86662 8730
rect 86662 8678 86674 8730
rect 86674 8678 86688 8730
rect 86712 8678 86726 8730
rect 86726 8678 86738 8730
rect 86738 8678 86768 8730
rect 86792 8678 86802 8730
rect 86802 8678 86848 8730
rect 86552 8676 86608 8678
rect 86632 8676 86688 8678
rect 86712 8676 86768 8678
rect 86792 8676 86848 8678
rect 87288 8186 87344 8188
rect 87368 8186 87424 8188
rect 87448 8186 87504 8188
rect 87528 8186 87584 8188
rect 87288 8134 87334 8186
rect 87334 8134 87344 8186
rect 87368 8134 87398 8186
rect 87398 8134 87410 8186
rect 87410 8134 87424 8186
rect 87448 8134 87462 8186
rect 87462 8134 87474 8186
rect 87474 8134 87504 8186
rect 87528 8134 87538 8186
rect 87538 8134 87584 8186
rect 87288 8132 87344 8134
rect 87368 8132 87424 8134
rect 87448 8132 87504 8134
rect 87528 8132 87584 8134
rect 86552 7642 86608 7644
rect 86632 7642 86688 7644
rect 86712 7642 86768 7644
rect 86792 7642 86848 7644
rect 86552 7590 86598 7642
rect 86598 7590 86608 7642
rect 86632 7590 86662 7642
rect 86662 7590 86674 7642
rect 86674 7590 86688 7642
rect 86712 7590 86726 7642
rect 86726 7590 86738 7642
rect 86738 7590 86768 7642
rect 86792 7590 86802 7642
rect 86802 7590 86848 7642
rect 86552 7588 86608 7590
rect 86632 7588 86688 7590
rect 86712 7588 86768 7590
rect 86792 7588 86848 7590
rect 87288 7098 87344 7100
rect 87368 7098 87424 7100
rect 87448 7098 87504 7100
rect 87528 7098 87584 7100
rect 87288 7046 87334 7098
rect 87334 7046 87344 7098
rect 87368 7046 87398 7098
rect 87398 7046 87410 7098
rect 87410 7046 87424 7098
rect 87448 7046 87462 7098
rect 87462 7046 87474 7098
rect 87474 7046 87504 7098
rect 87528 7046 87538 7098
rect 87538 7046 87584 7098
rect 87288 7044 87344 7046
rect 87368 7044 87424 7046
rect 87448 7044 87504 7046
rect 87528 7044 87584 7046
rect 18388 4922 18444 4924
rect 18468 4922 18524 4924
rect 18548 4922 18604 4924
rect 18628 4922 18684 4924
rect 18388 4870 18434 4922
rect 18434 4870 18444 4922
rect 18468 4870 18498 4922
rect 18498 4870 18510 4922
rect 18510 4870 18524 4922
rect 18548 4870 18562 4922
rect 18562 4870 18574 4922
rect 18574 4870 18604 4922
rect 18628 4870 18638 4922
rect 18638 4870 18684 4922
rect 18388 4868 18444 4870
rect 18468 4868 18524 4870
rect 18548 4868 18604 4870
rect 18628 4868 18684 4870
rect 36788 4922 36844 4924
rect 36868 4922 36924 4924
rect 36948 4922 37004 4924
rect 37028 4922 37084 4924
rect 36788 4870 36834 4922
rect 36834 4870 36844 4922
rect 36868 4870 36898 4922
rect 36898 4870 36910 4922
rect 36910 4870 36924 4922
rect 36948 4870 36962 4922
rect 36962 4870 36974 4922
rect 36974 4870 37004 4922
rect 37028 4870 37038 4922
rect 37038 4870 37084 4922
rect 36788 4868 36844 4870
rect 36868 4868 36924 4870
rect 36948 4868 37004 4870
rect 37028 4868 37084 4870
rect 55188 4922 55244 4924
rect 55268 4922 55324 4924
rect 55348 4922 55404 4924
rect 55428 4922 55484 4924
rect 55188 4870 55234 4922
rect 55234 4870 55244 4922
rect 55268 4870 55298 4922
rect 55298 4870 55310 4922
rect 55310 4870 55324 4922
rect 55348 4870 55362 4922
rect 55362 4870 55374 4922
rect 55374 4870 55404 4922
rect 55428 4870 55438 4922
rect 55438 4870 55484 4922
rect 55188 4868 55244 4870
rect 55268 4868 55324 4870
rect 55348 4868 55404 4870
rect 55428 4868 55484 4870
rect 73588 4922 73644 4924
rect 73668 4922 73724 4924
rect 73748 4922 73804 4924
rect 73828 4922 73884 4924
rect 73588 4870 73634 4922
rect 73634 4870 73644 4922
rect 73668 4870 73698 4922
rect 73698 4870 73710 4922
rect 73710 4870 73724 4922
rect 73748 4870 73762 4922
rect 73762 4870 73774 4922
rect 73774 4870 73804 4922
rect 73828 4870 73838 4922
rect 73838 4870 73884 4922
rect 73588 4868 73644 4870
rect 73668 4868 73724 4870
rect 73748 4868 73804 4870
rect 73828 4868 73884 4870
<< metal3 >>
rect 18378 87616 18694 87617
rect 18378 87552 18384 87616
rect 18448 87552 18464 87616
rect 18528 87552 18544 87616
rect 18608 87552 18624 87616
rect 18688 87552 18694 87616
rect 18378 87551 18694 87552
rect 36778 87616 37094 87617
rect 36778 87552 36784 87616
rect 36848 87552 36864 87616
rect 36928 87552 36944 87616
rect 37008 87552 37024 87616
rect 37088 87552 37094 87616
rect 36778 87551 37094 87552
rect 55178 87616 55494 87617
rect 55178 87552 55184 87616
rect 55248 87552 55264 87616
rect 55328 87552 55344 87616
rect 55408 87552 55424 87616
rect 55488 87552 55494 87616
rect 55178 87551 55494 87552
rect 73578 87616 73894 87617
rect 73578 87552 73584 87616
rect 73648 87552 73664 87616
rect 73728 87552 73744 87616
rect 73808 87552 73824 87616
rect 73888 87552 73894 87616
rect 73578 87551 73894 87552
rect 10302 87316 10308 87380
rect 10372 87378 10378 87380
rect 10721 87378 10787 87381
rect 10372 87376 10787 87378
rect 10372 87320 10726 87376
rect 10782 87320 10787 87376
rect 10372 87318 10787 87320
rect 10372 87316 10378 87318
rect 10721 87315 10787 87318
rect 17718 87072 18034 87073
rect 17718 87008 17724 87072
rect 17788 87008 17804 87072
rect 17868 87008 17884 87072
rect 17948 87008 17964 87072
rect 18028 87008 18034 87072
rect 17718 87007 18034 87008
rect 36118 87072 36434 87073
rect 36118 87008 36124 87072
rect 36188 87008 36204 87072
rect 36268 87008 36284 87072
rect 36348 87008 36364 87072
rect 36428 87008 36434 87072
rect 36118 87007 36434 87008
rect 54518 87072 54834 87073
rect 54518 87008 54524 87072
rect 54588 87008 54604 87072
rect 54668 87008 54684 87072
rect 54748 87008 54764 87072
rect 54828 87008 54834 87072
rect 54518 87007 54834 87008
rect 72918 87072 73234 87073
rect 72918 87008 72924 87072
rect 72988 87008 73004 87072
rect 73068 87008 73084 87072
rect 73148 87008 73164 87072
rect 73228 87008 73234 87072
rect 72918 87007 73234 87008
rect 18378 86528 18694 86529
rect 18378 86464 18384 86528
rect 18448 86464 18464 86528
rect 18528 86464 18544 86528
rect 18608 86464 18624 86528
rect 18688 86464 18694 86528
rect 18378 86463 18694 86464
rect 36778 86528 37094 86529
rect 36778 86464 36784 86528
rect 36848 86464 36864 86528
rect 36928 86464 36944 86528
rect 37008 86464 37024 86528
rect 37088 86464 37094 86528
rect 36778 86463 37094 86464
rect 55178 86528 55494 86529
rect 55178 86464 55184 86528
rect 55248 86464 55264 86528
rect 55328 86464 55344 86528
rect 55408 86464 55424 86528
rect 55488 86464 55494 86528
rect 55178 86463 55494 86464
rect 73578 86528 73894 86529
rect 73578 86464 73584 86528
rect 73648 86464 73664 86528
rect 73728 86464 73744 86528
rect 73808 86464 73824 86528
rect 73888 86464 73894 86528
rect 73578 86463 73894 86464
rect 17718 85984 18034 85985
rect 17718 85920 17724 85984
rect 17788 85920 17804 85984
rect 17868 85920 17884 85984
rect 17948 85920 17964 85984
rect 18028 85920 18034 85984
rect 17718 85919 18034 85920
rect 36118 85984 36434 85985
rect 36118 85920 36124 85984
rect 36188 85920 36204 85984
rect 36268 85920 36284 85984
rect 36348 85920 36364 85984
rect 36428 85920 36434 85984
rect 36118 85919 36434 85920
rect 54518 85984 54834 85985
rect 54518 85920 54524 85984
rect 54588 85920 54604 85984
rect 54668 85920 54684 85984
rect 54748 85920 54764 85984
rect 54828 85920 54834 85984
rect 54518 85919 54834 85920
rect 72918 85984 73234 85985
rect 72918 85920 72924 85984
rect 72988 85920 73004 85984
rect 73068 85920 73084 85984
rect 73148 85920 73164 85984
rect 73228 85920 73234 85984
rect 72918 85919 73234 85920
rect 18378 85440 18694 85441
rect 18378 85376 18384 85440
rect 18448 85376 18464 85440
rect 18528 85376 18544 85440
rect 18608 85376 18624 85440
rect 18688 85376 18694 85440
rect 18378 85375 18694 85376
rect 36778 85440 37094 85441
rect 36778 85376 36784 85440
rect 36848 85376 36864 85440
rect 36928 85376 36944 85440
rect 37008 85376 37024 85440
rect 37088 85376 37094 85440
rect 36778 85375 37094 85376
rect 55178 85440 55494 85441
rect 55178 85376 55184 85440
rect 55248 85376 55264 85440
rect 55328 85376 55344 85440
rect 55408 85376 55424 85440
rect 55488 85376 55494 85440
rect 55178 85375 55494 85376
rect 73578 85440 73894 85441
rect 73578 85376 73584 85440
rect 73648 85376 73664 85440
rect 73728 85376 73744 85440
rect 73808 85376 73824 85440
rect 73888 85376 73894 85440
rect 73578 85375 73894 85376
rect 5950 84896 6266 84897
rect 5950 84832 5956 84896
rect 6020 84832 6036 84896
rect 6100 84832 6116 84896
rect 6180 84832 6196 84896
rect 6260 84832 6266 84896
rect 5950 84831 6266 84832
rect 17718 84896 18034 84897
rect 17718 84832 17724 84896
rect 17788 84832 17804 84896
rect 17868 84832 17884 84896
rect 17948 84832 17964 84896
rect 18028 84832 18034 84896
rect 17718 84831 18034 84832
rect 36118 84896 36434 84897
rect 36118 84832 36124 84896
rect 36188 84832 36204 84896
rect 36268 84832 36284 84896
rect 36348 84832 36364 84896
rect 36428 84832 36434 84896
rect 36118 84831 36434 84832
rect 54518 84896 54834 84897
rect 54518 84832 54524 84896
rect 54588 84832 54604 84896
rect 54668 84832 54684 84896
rect 54748 84832 54764 84896
rect 54828 84832 54834 84896
rect 54518 84831 54834 84832
rect 72918 84896 73234 84897
rect 72918 84832 72924 84896
rect 72988 84832 73004 84896
rect 73068 84832 73084 84896
rect 73148 84832 73164 84896
rect 73228 84832 73234 84896
rect 72918 84831 73234 84832
rect 86542 84896 86858 84897
rect 86542 84832 86548 84896
rect 86612 84832 86628 84896
rect 86692 84832 86708 84896
rect 86772 84832 86788 84896
rect 86852 84832 86858 84896
rect 86542 84831 86858 84832
rect 6686 84352 7002 84353
rect 6686 84288 6692 84352
rect 6756 84288 6772 84352
rect 6836 84288 6852 84352
rect 6916 84288 6932 84352
rect 6996 84288 7002 84352
rect 6686 84287 7002 84288
rect 18378 84352 18694 84353
rect 18378 84288 18384 84352
rect 18448 84288 18464 84352
rect 18528 84288 18544 84352
rect 18608 84288 18624 84352
rect 18688 84288 18694 84352
rect 18378 84287 18694 84288
rect 36778 84352 37094 84353
rect 36778 84288 36784 84352
rect 36848 84288 36864 84352
rect 36928 84288 36944 84352
rect 37008 84288 37024 84352
rect 37088 84288 37094 84352
rect 36778 84287 37094 84288
rect 55178 84352 55494 84353
rect 55178 84288 55184 84352
rect 55248 84288 55264 84352
rect 55328 84288 55344 84352
rect 55408 84288 55424 84352
rect 55488 84288 55494 84352
rect 55178 84287 55494 84288
rect 73578 84352 73894 84353
rect 73578 84288 73584 84352
rect 73648 84288 73664 84352
rect 73728 84288 73744 84352
rect 73808 84288 73824 84352
rect 73888 84288 73894 84352
rect 73578 84287 73894 84288
rect 87278 84352 87594 84353
rect 87278 84288 87284 84352
rect 87348 84288 87364 84352
rect 87428 84288 87444 84352
rect 87508 84288 87524 84352
rect 87588 84288 87594 84352
rect 87278 84287 87594 84288
rect 5950 83808 6266 83809
rect 5950 83744 5956 83808
rect 6020 83744 6036 83808
rect 6100 83744 6116 83808
rect 6180 83744 6196 83808
rect 6260 83744 6266 83808
rect 5950 83743 6266 83744
rect 86542 83808 86858 83809
rect 86542 83744 86548 83808
rect 86612 83744 86628 83808
rect 86692 83744 86708 83808
rect 86772 83744 86788 83808
rect 86852 83744 86858 83808
rect 86542 83743 86858 83744
rect 6686 83264 7002 83265
rect 6686 83200 6692 83264
rect 6756 83200 6772 83264
rect 6836 83200 6852 83264
rect 6916 83200 6932 83264
rect 6996 83200 7002 83264
rect 6686 83199 7002 83200
rect 87278 83264 87594 83265
rect 87278 83200 87284 83264
rect 87348 83200 87364 83264
rect 87428 83200 87444 83264
rect 87508 83200 87524 83264
rect 87588 83200 87594 83264
rect 87278 83199 87594 83200
rect 5950 82720 6266 82721
rect 5950 82656 5956 82720
rect 6020 82656 6036 82720
rect 6100 82656 6116 82720
rect 6180 82656 6196 82720
rect 6260 82656 6266 82720
rect 5950 82655 6266 82656
rect 86542 82720 86858 82721
rect 86542 82656 86548 82720
rect 86612 82656 86628 82720
rect 86692 82656 86708 82720
rect 86772 82656 86788 82720
rect 86852 82656 86858 82720
rect 86542 82655 86858 82656
rect 10537 82346 10603 82349
rect 10494 82344 10603 82346
rect 10494 82288 10542 82344
rect 10598 82288 10603 82344
rect 10494 82283 10603 82288
rect 6686 82176 7002 82177
rect 6686 82112 6692 82176
rect 6756 82112 6772 82176
rect 6836 82112 6852 82176
rect 6916 82112 6932 82176
rect 6996 82112 7002 82176
rect 6686 82111 7002 82112
rect 10494 82077 10554 82283
rect 87278 82176 87594 82177
rect 87278 82112 87284 82176
rect 87348 82112 87364 82176
rect 87428 82112 87444 82176
rect 87508 82112 87524 82176
rect 87588 82112 87594 82176
rect 87278 82111 87594 82112
rect 9985 82074 10051 82077
rect 10494 82074 10603 82077
rect 9985 82072 10603 82074
rect 9985 82016 9990 82072
rect 10046 82016 10542 82072
rect 10598 82016 10603 82072
rect 9985 82014 10603 82016
rect 9985 82011 10051 82014
rect 10537 82011 10603 82014
rect 5950 81632 6266 81633
rect 5950 81568 5956 81632
rect 6020 81568 6036 81632
rect 6100 81568 6116 81632
rect 6180 81568 6196 81632
rect 6260 81568 6266 81632
rect 5950 81567 6266 81568
rect 86542 81632 86858 81633
rect 86542 81568 86548 81632
rect 86612 81568 86628 81632
rect 86692 81568 86708 81632
rect 86772 81568 86788 81632
rect 86852 81568 86858 81632
rect 86542 81567 86858 81568
rect 88369 81258 88435 81261
rect 89200 81258 90000 81288
rect 88369 81256 90000 81258
rect 88369 81200 88374 81256
rect 88430 81200 90000 81256
rect 88369 81198 90000 81200
rect 88369 81195 88435 81198
rect 89200 81168 90000 81198
rect 6686 81088 7002 81089
rect 6686 81024 6692 81088
rect 6756 81024 6772 81088
rect 6836 81024 6852 81088
rect 6916 81024 6932 81088
rect 6996 81024 7002 81088
rect 87278 81088 87594 81089
rect 6686 81023 7002 81024
rect 10302 80992 10308 81056
rect 10372 80992 10378 81056
rect 83493 81054 83559 81057
rect 45668 80994 46250 81054
rect 83020 81052 83559 81054
rect 83020 80996 83498 81052
rect 83554 80996 83559 81052
rect 87278 81024 87284 81088
rect 87348 81024 87364 81088
rect 87428 81024 87444 81088
rect 87508 81024 87524 81088
rect 87588 81024 87594 81088
rect 87278 81023 87594 81024
rect 83020 80994 83559 80996
rect 46190 80986 46250 80994
rect 83493 80991 83559 80994
rect 46190 80926 47508 80986
rect 5950 80544 6266 80545
rect 5950 80480 5956 80544
rect 6020 80480 6036 80544
rect 6100 80480 6116 80544
rect 6180 80480 6196 80544
rect 6260 80480 6266 80544
rect 5950 80479 6266 80480
rect 86542 80544 86858 80545
rect 86542 80480 86548 80544
rect 86612 80480 86628 80544
rect 86692 80480 86708 80544
rect 86772 80480 86788 80544
rect 86852 80480 86858 80544
rect 86542 80479 86858 80480
rect 7133 80170 7199 80173
rect 7133 80168 10186 80170
rect 7133 80112 7138 80168
rect 7194 80112 10186 80168
rect 7133 80110 10186 80112
rect 7133 80107 7199 80110
rect 6686 80000 7002 80001
rect 6686 79936 6692 80000
rect 6756 79936 6772 80000
rect 6836 79936 6852 80000
rect 6916 79936 6932 80000
rect 6996 79936 7002 80000
rect 10126 79936 10186 80110
rect 87278 80000 87594 80001
rect 83493 79966 83559 79969
rect 6686 79935 7002 79936
rect 1600 79898 2400 79928
rect 45668 79906 46250 79966
rect 83020 79964 83559 79966
rect 83020 79908 83498 79964
rect 83554 79908 83559 79964
rect 87278 79936 87284 80000
rect 87348 79936 87364 80000
rect 87428 79936 87444 80000
rect 87508 79936 87524 80000
rect 87588 79936 87594 80000
rect 87278 79935 87594 79936
rect 83020 79906 83559 79908
rect 2901 79898 2967 79901
rect 1600 79896 2967 79898
rect 1600 79840 2906 79896
rect 2962 79840 2967 79896
rect 1600 79838 2967 79840
rect 46190 79898 46250 79906
rect 83493 79903 83559 79906
rect 88277 79898 88343 79901
rect 89200 79898 90000 79928
rect 46190 79838 47508 79898
rect 88277 79896 90000 79898
rect 88277 79840 88282 79896
rect 88338 79840 90000 79896
rect 88277 79838 90000 79840
rect 1600 79808 2400 79838
rect 2901 79835 2967 79838
rect 88277 79835 88343 79838
rect 89200 79808 90000 79838
rect 5950 79456 6266 79457
rect 5950 79392 5956 79456
rect 6020 79392 6036 79456
rect 6100 79392 6116 79456
rect 6180 79392 6196 79456
rect 6260 79392 6266 79456
rect 5950 79391 6266 79392
rect 86542 79456 86858 79457
rect 86542 79392 86548 79456
rect 86612 79392 86628 79456
rect 86692 79392 86708 79456
rect 86772 79392 86788 79456
rect 86852 79392 86858 79456
rect 86542 79391 86858 79392
rect 6686 78912 7002 78913
rect 6686 78848 6692 78912
rect 6756 78848 6772 78912
rect 6836 78848 6852 78912
rect 6916 78848 6932 78912
rect 6996 78848 7002 78912
rect 87278 78912 87594 78913
rect 6686 78847 7002 78848
rect 45668 78818 46250 78878
rect 83020 78818 83602 78878
rect 87278 78848 87284 78912
rect 87348 78848 87364 78912
rect 87428 78848 87444 78912
rect 87508 78848 87524 78912
rect 87588 78848 87594 78912
rect 87278 78847 87594 78848
rect 7133 78810 7199 78813
rect 46190 78810 46250 78818
rect 83542 78810 83602 78818
rect 7133 78808 10156 78810
rect 7133 78752 7138 78808
rect 7194 78752 10156 78808
rect 7133 78750 10156 78752
rect 46190 78750 47508 78810
rect 83542 78750 85810 78810
rect 7133 78747 7199 78750
rect 85750 78674 85810 78750
rect 88001 78674 88067 78677
rect 85750 78672 88067 78674
rect 85750 78616 88006 78672
rect 88062 78616 88067 78672
rect 85750 78614 88067 78616
rect 88001 78611 88067 78614
rect 1600 78538 2400 78568
rect 2901 78538 2967 78541
rect 1600 78536 2967 78538
rect 1600 78480 2906 78536
rect 2962 78480 2967 78536
rect 1600 78478 2967 78480
rect 1600 78448 2400 78478
rect 2901 78475 2967 78478
rect 88277 78538 88343 78541
rect 89200 78538 90000 78568
rect 88277 78536 90000 78538
rect 88277 78480 88282 78536
rect 88338 78480 90000 78536
rect 88277 78478 90000 78480
rect 88277 78475 88343 78478
rect 89200 78448 90000 78478
rect 5950 78368 6266 78369
rect 5950 78304 5956 78368
rect 6020 78304 6036 78368
rect 6100 78304 6116 78368
rect 6180 78304 6196 78368
rect 6260 78304 6266 78368
rect 5950 78303 6266 78304
rect 86542 78368 86858 78369
rect 86542 78304 86548 78368
rect 86612 78304 86628 78368
rect 86692 78304 86708 78368
rect 86772 78304 86788 78368
rect 86852 78304 86858 78368
rect 86542 78303 86858 78304
rect 7133 77994 7199 77997
rect 87817 77994 87883 77997
rect 7133 77992 10186 77994
rect 7133 77936 7138 77992
rect 7194 77936 10186 77992
rect 7133 77934 10186 77936
rect 7133 77931 7199 77934
rect 1600 77858 2400 77888
rect 2901 77858 2967 77861
rect 1600 77856 2967 77858
rect 1600 77800 2906 77856
rect 2962 77800 2967 77856
rect 1600 77798 2967 77800
rect 1600 77768 2400 77798
rect 2901 77795 2967 77798
rect 6686 77824 7002 77825
rect 6686 77760 6692 77824
rect 6756 77760 6772 77824
rect 6836 77760 6852 77824
rect 6916 77760 6932 77824
rect 6996 77760 7002 77824
rect 10126 77760 10186 77934
rect 85750 77992 87883 77994
rect 85750 77936 87822 77992
rect 87878 77936 87883 77992
rect 85750 77934 87883 77936
rect 85750 77858 85810 77934
rect 87817 77931 87883 77934
rect 83542 77798 85810 77858
rect 88277 77858 88343 77861
rect 89200 77858 90000 77888
rect 88277 77856 90000 77858
rect 87278 77824 87594 77825
rect 83542 77790 83602 77798
rect 6686 77759 7002 77760
rect 45668 77730 46250 77790
rect 83020 77730 83602 77790
rect 87278 77760 87284 77824
rect 87348 77760 87364 77824
rect 87428 77760 87444 77824
rect 87508 77760 87524 77824
rect 87588 77760 87594 77824
rect 88277 77800 88282 77856
rect 88338 77800 90000 77856
rect 88277 77798 90000 77800
rect 88277 77795 88343 77798
rect 89200 77768 90000 77798
rect 87278 77759 87594 77760
rect 46190 77722 46250 77730
rect 46190 77662 47508 77722
rect 5950 77280 6266 77281
rect 5950 77216 5956 77280
rect 6020 77216 6036 77280
rect 6100 77216 6116 77280
rect 6180 77216 6196 77280
rect 6260 77216 6266 77280
rect 5950 77215 6266 77216
rect 86542 77280 86858 77281
rect 86542 77216 86548 77280
rect 86612 77216 86628 77280
rect 86692 77216 86708 77280
rect 86772 77216 86788 77280
rect 86852 77216 86858 77280
rect 86542 77215 86858 77216
rect 7133 76906 7199 76909
rect 7133 76904 10186 76906
rect 7133 76848 7138 76904
rect 7194 76848 10186 76904
rect 7133 76846 10186 76848
rect 7133 76843 7199 76846
rect 6686 76736 7002 76737
rect 6686 76672 6692 76736
rect 6756 76672 6772 76736
rect 6836 76672 6852 76736
rect 6916 76672 6932 76736
rect 6996 76672 7002 76736
rect 10126 76672 10186 76846
rect 86621 76770 86687 76773
rect 83542 76768 86687 76770
rect 83542 76712 86626 76768
rect 86682 76712 86687 76768
rect 83542 76710 86687 76712
rect 83542 76702 83602 76710
rect 86621 76707 86687 76710
rect 87278 76736 87594 76737
rect 6686 76671 7002 76672
rect 45668 76642 46250 76702
rect 83020 76642 83602 76702
rect 87278 76672 87284 76736
rect 87348 76672 87364 76736
rect 87428 76672 87444 76736
rect 87508 76672 87524 76736
rect 87588 76672 87594 76736
rect 87278 76671 87594 76672
rect 46190 76634 46250 76642
rect 46190 76574 47508 76634
rect 1600 76498 2400 76528
rect 2717 76498 2783 76501
rect 1600 76496 2783 76498
rect 1600 76440 2722 76496
rect 2778 76440 2783 76496
rect 1600 76438 2783 76440
rect 1600 76408 2400 76438
rect 2717 76435 2783 76438
rect 88001 76498 88067 76501
rect 89200 76498 90000 76528
rect 88001 76496 90000 76498
rect 88001 76440 88006 76496
rect 88062 76440 90000 76496
rect 88001 76438 90000 76440
rect 88001 76435 88067 76438
rect 89200 76408 90000 76438
rect 5950 76192 6266 76193
rect 5950 76128 5956 76192
rect 6020 76128 6036 76192
rect 6100 76128 6116 76192
rect 6180 76128 6196 76192
rect 6260 76128 6266 76192
rect 5950 76127 6266 76128
rect 86542 76192 86858 76193
rect 86542 76128 86548 76192
rect 86612 76128 86628 76192
rect 86692 76128 86708 76192
rect 86772 76128 86788 76192
rect 86852 76128 86858 76192
rect 86542 76127 86858 76128
rect 1600 75818 2400 75848
rect 2901 75818 2967 75821
rect 1600 75816 2967 75818
rect 1600 75760 2906 75816
rect 2962 75760 2967 75816
rect 1600 75758 2967 75760
rect 1600 75728 2400 75758
rect 2901 75755 2967 75758
rect 7133 75818 7199 75821
rect 88461 75818 88527 75821
rect 89200 75818 90000 75848
rect 7133 75816 10186 75818
rect 7133 75760 7138 75816
rect 7194 75760 10186 75816
rect 7133 75758 10186 75760
rect 7133 75755 7199 75758
rect 6686 75648 7002 75649
rect 6686 75584 6692 75648
rect 6756 75584 6772 75648
rect 6836 75584 6852 75648
rect 6916 75584 6932 75648
rect 6996 75584 7002 75648
rect 10126 75584 10186 75758
rect 88461 75816 90000 75818
rect 88461 75760 88466 75816
rect 88522 75760 90000 75816
rect 88461 75758 90000 75760
rect 88461 75755 88527 75758
rect 89200 75728 90000 75758
rect 86897 75682 86963 75685
rect 83542 75680 86963 75682
rect 83542 75624 86902 75680
rect 86958 75624 86963 75680
rect 83542 75622 86963 75624
rect 83542 75614 83602 75622
rect 86897 75619 86963 75622
rect 87278 75648 87594 75649
rect 6686 75583 7002 75584
rect 45668 75554 46250 75614
rect 83020 75554 83602 75614
rect 87278 75584 87284 75648
rect 87348 75584 87364 75648
rect 87428 75584 87444 75648
rect 87508 75584 87524 75648
rect 87588 75584 87594 75648
rect 87278 75583 87594 75584
rect 46190 75546 46250 75554
rect 46190 75486 47508 75546
rect 5950 75104 6266 75105
rect 5950 75040 5956 75104
rect 6020 75040 6036 75104
rect 6100 75040 6116 75104
rect 6180 75040 6196 75104
rect 6260 75040 6266 75104
rect 5950 75039 6266 75040
rect 86542 75104 86858 75105
rect 86542 75040 86548 75104
rect 86612 75040 86628 75104
rect 86692 75040 86708 75104
rect 86772 75040 86788 75104
rect 86852 75040 86858 75104
rect 86542 75039 86858 75040
rect 6446 74670 10186 74730
rect 5661 74594 5727 74597
rect 6446 74594 6506 74670
rect 5661 74592 6506 74594
rect 5661 74536 5666 74592
rect 5722 74536 6506 74592
rect 5661 74534 6506 74536
rect 6686 74560 7002 74561
rect 5661 74531 5727 74534
rect 6686 74496 6692 74560
rect 6756 74496 6772 74560
rect 6836 74496 6852 74560
rect 6916 74496 6932 74560
rect 6996 74496 7002 74560
rect 10126 74496 10186 74670
rect 84413 74594 84479 74597
rect 83358 74592 84479 74594
rect 83358 74536 84418 74592
rect 84474 74536 84479 74592
rect 83358 74534 84479 74536
rect 83358 74526 83418 74534
rect 84413 74531 84479 74534
rect 87278 74560 87594 74561
rect 6686 74495 7002 74496
rect 1600 74458 2400 74488
rect 45668 74466 46250 74526
rect 83020 74466 83418 74526
rect 87278 74496 87284 74560
rect 87348 74496 87364 74560
rect 87428 74496 87444 74560
rect 87508 74496 87524 74560
rect 87588 74496 87594 74560
rect 87278 74495 87594 74496
rect 4373 74458 4439 74461
rect 1600 74456 4439 74458
rect 1600 74400 4378 74456
rect 4434 74400 4439 74456
rect 1600 74398 4439 74400
rect 46190 74458 46250 74466
rect 88553 74458 88619 74461
rect 89200 74458 90000 74488
rect 46190 74398 47508 74458
rect 88553 74456 90000 74458
rect 88553 74400 88558 74456
rect 88614 74400 90000 74456
rect 88553 74398 90000 74400
rect 1600 74368 2400 74398
rect 4373 74395 4439 74398
rect 88553 74395 88619 74398
rect 89200 74368 90000 74398
rect 5950 74016 6266 74017
rect 5950 73952 5956 74016
rect 6020 73952 6036 74016
rect 6100 73952 6116 74016
rect 6180 73952 6196 74016
rect 6260 73952 6266 74016
rect 5950 73951 6266 73952
rect 86542 74016 86858 74017
rect 86542 73952 86548 74016
rect 86612 73952 86628 74016
rect 86692 73952 86708 74016
rect 86772 73952 86788 74016
rect 86852 73952 86858 74016
rect 86542 73951 86858 73952
rect 6686 73472 7002 73473
rect 6686 73408 6692 73472
rect 6756 73408 6772 73472
rect 6836 73408 6852 73472
rect 6916 73408 6932 73472
rect 6996 73408 7002 73472
rect 87278 73472 87594 73473
rect 6686 73407 7002 73408
rect 45668 73378 46066 73438
rect 83020 73378 83418 73438
rect 87278 73408 87284 73472
rect 87348 73408 87364 73472
rect 87428 73408 87444 73472
rect 87508 73408 87524 73472
rect 87588 73408 87594 73472
rect 87278 73407 87594 73408
rect 7133 73370 7199 73373
rect 46006 73370 46066 73378
rect 83358 73370 83418 73378
rect 7133 73368 10156 73370
rect 7133 73312 7138 73368
rect 7194 73312 10156 73368
rect 7133 73310 10156 73312
rect 46006 73310 47508 73370
rect 83358 73310 85810 73370
rect 7133 73307 7199 73310
rect 85750 73234 85810 73310
rect 88001 73234 88067 73237
rect 85750 73232 88067 73234
rect 85750 73176 88006 73232
rect 88062 73176 88067 73232
rect 85750 73174 88067 73176
rect 88001 73171 88067 73174
rect 1600 73098 2400 73128
rect 2901 73098 2967 73101
rect 1600 73096 2967 73098
rect 1600 73040 2906 73096
rect 2962 73040 2967 73096
rect 1600 73038 2967 73040
rect 1600 73008 2400 73038
rect 2901 73035 2967 73038
rect 88277 73098 88343 73101
rect 89200 73098 90000 73128
rect 88277 73096 90000 73098
rect 88277 73040 88282 73096
rect 88338 73040 90000 73096
rect 88277 73038 90000 73040
rect 88277 73035 88343 73038
rect 89200 73008 90000 73038
rect 5950 72928 6266 72929
rect 5950 72864 5956 72928
rect 6020 72864 6036 72928
rect 6100 72864 6116 72928
rect 6180 72864 6196 72928
rect 6260 72864 6266 72928
rect 5950 72863 6266 72864
rect 86542 72928 86858 72929
rect 86542 72864 86548 72928
rect 86612 72864 86628 72928
rect 86692 72864 86708 72928
rect 86772 72864 86788 72928
rect 86852 72864 86858 72928
rect 86542 72863 86858 72864
rect 7133 72554 7199 72557
rect 87173 72554 87239 72557
rect 7133 72552 10186 72554
rect 7133 72496 7138 72552
rect 7194 72496 10186 72552
rect 7133 72494 10186 72496
rect 7133 72491 7199 72494
rect 1600 72418 2400 72448
rect 2901 72418 2967 72421
rect 1600 72416 2967 72418
rect 1600 72360 2906 72416
rect 2962 72360 2967 72416
rect 1600 72358 2967 72360
rect 1600 72328 2400 72358
rect 2901 72355 2967 72358
rect 6686 72384 7002 72385
rect 6686 72320 6692 72384
rect 6756 72320 6772 72384
rect 6836 72320 6852 72384
rect 6916 72320 6932 72384
rect 6996 72320 7002 72384
rect 10126 72320 10186 72494
rect 85750 72552 87239 72554
rect 85750 72496 87178 72552
rect 87234 72496 87239 72552
rect 85750 72494 87239 72496
rect 85750 72418 85810 72494
rect 87173 72491 87239 72494
rect 83542 72358 85810 72418
rect 88277 72418 88343 72421
rect 89200 72418 90000 72448
rect 88277 72416 90000 72418
rect 87278 72384 87594 72385
rect 83542 72350 83602 72358
rect 6686 72319 7002 72320
rect 45668 72290 46250 72350
rect 83020 72290 83602 72350
rect 87278 72320 87284 72384
rect 87348 72320 87364 72384
rect 87428 72320 87444 72384
rect 87508 72320 87524 72384
rect 87588 72320 87594 72384
rect 88277 72360 88282 72416
rect 88338 72360 90000 72416
rect 88277 72358 90000 72360
rect 88277 72355 88343 72358
rect 89200 72328 90000 72358
rect 87278 72319 87594 72320
rect 46190 72282 46250 72290
rect 46190 72222 47508 72282
rect 5950 71840 6266 71841
rect 5950 71776 5956 71840
rect 6020 71776 6036 71840
rect 6100 71776 6116 71840
rect 6180 71776 6196 71840
rect 6260 71776 6266 71840
rect 5950 71775 6266 71776
rect 86542 71840 86858 71841
rect 86542 71776 86548 71840
rect 86612 71776 86628 71840
rect 86692 71776 86708 71840
rect 86772 71776 86788 71840
rect 86852 71776 86858 71840
rect 86542 71775 86858 71776
rect 7133 71466 7199 71469
rect 7133 71464 10186 71466
rect 7133 71408 7138 71464
rect 7194 71408 10186 71464
rect 7133 71406 10186 71408
rect 7133 71403 7199 71406
rect 6686 71296 7002 71297
rect 6686 71232 6692 71296
rect 6756 71232 6772 71296
rect 6836 71232 6852 71296
rect 6916 71232 6932 71296
rect 6996 71232 7002 71296
rect 10126 71232 10186 71406
rect 86897 71330 86963 71333
rect 83542 71328 86963 71330
rect 83542 71272 86902 71328
rect 86958 71272 86963 71328
rect 83542 71270 86963 71272
rect 83542 71262 83602 71270
rect 86897 71267 86963 71270
rect 87278 71296 87594 71297
rect 6686 71231 7002 71232
rect 45668 71202 46250 71262
rect 83020 71202 83602 71262
rect 87278 71232 87284 71296
rect 87348 71232 87364 71296
rect 87428 71232 87444 71296
rect 87508 71232 87524 71296
rect 87588 71232 87594 71296
rect 87278 71231 87594 71232
rect 46190 71194 46250 71202
rect 46190 71134 47508 71194
rect 1600 71058 2400 71088
rect 2717 71058 2783 71061
rect 1600 71056 2783 71058
rect 1600 71000 2722 71056
rect 2778 71000 2783 71056
rect 1600 70998 2783 71000
rect 1600 70968 2400 70998
rect 2717 70995 2783 70998
rect 88277 71058 88343 71061
rect 89200 71058 90000 71088
rect 88277 71056 90000 71058
rect 88277 71000 88282 71056
rect 88338 71000 90000 71056
rect 88277 70998 90000 71000
rect 88277 70995 88343 70998
rect 89200 70968 90000 70998
rect 5950 70752 6266 70753
rect 5950 70688 5956 70752
rect 6020 70688 6036 70752
rect 6100 70688 6116 70752
rect 6180 70688 6196 70752
rect 6260 70688 6266 70752
rect 5950 70687 6266 70688
rect 86542 70752 86858 70753
rect 86542 70688 86548 70752
rect 86612 70688 86628 70752
rect 86692 70688 86708 70752
rect 86772 70688 86788 70752
rect 86852 70688 86858 70752
rect 86542 70687 86858 70688
rect 1600 70378 2400 70408
rect 2901 70378 2967 70381
rect 1600 70376 2967 70378
rect 1600 70320 2906 70376
rect 2962 70320 2967 70376
rect 1600 70318 2967 70320
rect 1600 70288 2400 70318
rect 2901 70315 2967 70318
rect 7133 70378 7199 70381
rect 88185 70378 88251 70381
rect 89200 70378 90000 70408
rect 7133 70376 10186 70378
rect 7133 70320 7138 70376
rect 7194 70320 10186 70376
rect 7133 70318 10186 70320
rect 7133 70315 7199 70318
rect 6686 70208 7002 70209
rect 6686 70144 6692 70208
rect 6756 70144 6772 70208
rect 6836 70144 6852 70208
rect 6916 70144 6932 70208
rect 6996 70144 7002 70208
rect 10126 70144 10186 70318
rect 88185 70376 90000 70378
rect 88185 70320 88190 70376
rect 88246 70320 90000 70376
rect 88185 70318 90000 70320
rect 88185 70315 88251 70318
rect 89200 70288 90000 70318
rect 86897 70242 86963 70245
rect 83542 70240 86963 70242
rect 83542 70184 86902 70240
rect 86958 70184 86963 70240
rect 83542 70182 86963 70184
rect 83542 70174 83602 70182
rect 86897 70179 86963 70182
rect 87278 70208 87594 70209
rect 6686 70143 7002 70144
rect 45668 70114 46250 70174
rect 83020 70114 83602 70174
rect 87278 70144 87284 70208
rect 87348 70144 87364 70208
rect 87428 70144 87444 70208
rect 87508 70144 87524 70208
rect 87588 70144 87594 70208
rect 87278 70143 87594 70144
rect 46190 70106 46250 70114
rect 46190 70046 47508 70106
rect 5950 69664 6266 69665
rect 5950 69600 5956 69664
rect 6020 69600 6036 69664
rect 6100 69600 6116 69664
rect 6180 69600 6196 69664
rect 6260 69600 6266 69664
rect 5950 69599 6266 69600
rect 86542 69664 86858 69665
rect 86542 69600 86548 69664
rect 86612 69600 86628 69664
rect 86692 69600 86708 69664
rect 86772 69600 86788 69664
rect 86852 69600 86858 69664
rect 86542 69599 86858 69600
rect 86897 69154 86963 69157
rect 83542 69152 86963 69154
rect 6686 69120 7002 69121
rect 6686 69056 6692 69120
rect 6756 69056 6772 69120
rect 6836 69056 6852 69120
rect 6916 69056 6932 69120
rect 6996 69056 7002 69120
rect 83542 69096 86902 69152
rect 86958 69096 86963 69152
rect 83542 69094 86963 69096
rect 83542 69086 83602 69094
rect 86897 69091 86963 69094
rect 87278 69120 87594 69121
rect 6686 69055 7002 69056
rect 1600 69018 2400 69048
rect 45668 69026 46250 69086
rect 83020 69026 83602 69086
rect 87278 69056 87284 69120
rect 87348 69056 87364 69120
rect 87428 69056 87444 69120
rect 87508 69056 87524 69120
rect 87588 69056 87594 69120
rect 87278 69055 87594 69056
rect 4373 69018 4439 69021
rect 1600 69016 4439 69018
rect 1600 68960 4378 69016
rect 4434 68960 4439 69016
rect 46190 69018 46250 69026
rect 88553 69018 88619 69021
rect 89200 69018 90000 69048
rect 1600 68958 4439 68960
rect 1600 68928 2400 68958
rect 4373 68955 4439 68958
rect 5661 68882 5727 68885
rect 10126 68882 10186 68988
rect 46190 68958 47508 69018
rect 88553 69016 90000 69018
rect 88553 68960 88558 69016
rect 88614 68960 90000 69016
rect 88553 68958 90000 68960
rect 88553 68955 88619 68958
rect 89200 68928 90000 68958
rect 5661 68880 10186 68882
rect 5661 68824 5666 68880
rect 5722 68824 10186 68880
rect 5661 68822 10186 68824
rect 5661 68819 5727 68822
rect 5950 68576 6266 68577
rect 5950 68512 5956 68576
rect 6020 68512 6036 68576
rect 6100 68512 6116 68576
rect 6180 68512 6196 68576
rect 6260 68512 6266 68576
rect 5950 68511 6266 68512
rect 86542 68576 86858 68577
rect 86542 68512 86548 68576
rect 86612 68512 86628 68576
rect 86692 68512 86708 68576
rect 86772 68512 86788 68576
rect 86852 68512 86858 68576
rect 86542 68511 86858 68512
rect 5661 68202 5727 68205
rect 5661 68200 10186 68202
rect 5661 68144 5666 68200
rect 5722 68144 10186 68200
rect 5661 68142 10186 68144
rect 5661 68139 5727 68142
rect 6686 68032 7002 68033
rect 6686 67968 6692 68032
rect 6756 67968 6772 68032
rect 6836 67968 6852 68032
rect 6916 67968 6932 68032
rect 6996 67968 7002 68032
rect 10126 67968 10186 68142
rect 87278 68032 87594 68033
rect 6686 67967 7002 67968
rect 45668 67938 46250 67998
rect 83020 67938 83418 67998
rect 87278 67968 87284 68032
rect 87348 67968 87364 68032
rect 87428 67968 87444 68032
rect 87508 67968 87524 68032
rect 87588 67968 87594 68032
rect 87278 67967 87594 67968
rect 46190 67930 46250 67938
rect 83358 67930 83418 67938
rect 84413 67930 84479 67933
rect 46190 67870 47508 67930
rect 83358 67928 84479 67930
rect 83358 67872 84418 67928
rect 84474 67872 84479 67928
rect 83358 67870 84479 67872
rect 84413 67867 84479 67870
rect 1600 67658 2400 67688
rect 2901 67658 2967 67661
rect 1600 67656 2967 67658
rect 1600 67600 2906 67656
rect 2962 67600 2967 67656
rect 1600 67598 2967 67600
rect 1600 67568 2400 67598
rect 2901 67595 2967 67598
rect 88277 67658 88343 67661
rect 89200 67658 90000 67688
rect 88277 67656 90000 67658
rect 88277 67600 88282 67656
rect 88338 67600 90000 67656
rect 88277 67598 90000 67600
rect 88277 67595 88343 67598
rect 89200 67568 90000 67598
rect 5950 67488 6266 67489
rect 5950 67424 5956 67488
rect 6020 67424 6036 67488
rect 6100 67424 6116 67488
rect 6180 67424 6196 67488
rect 6260 67424 6266 67488
rect 5950 67423 6266 67424
rect 86542 67488 86858 67489
rect 86542 67424 86548 67488
rect 86612 67424 86628 67488
rect 86692 67424 86708 67488
rect 86772 67424 86788 67488
rect 86852 67424 86858 67488
rect 86542 67423 86858 67424
rect 7133 67114 7199 67117
rect 7133 67112 10186 67114
rect 7133 67056 7138 67112
rect 7194 67056 10186 67112
rect 7133 67054 10186 67056
rect 7133 67051 7199 67054
rect 1600 66978 2400 67008
rect 2901 66978 2967 66981
rect 1600 66976 2967 66978
rect 1600 66920 2906 66976
rect 2962 66920 2967 66976
rect 1600 66918 2967 66920
rect 1600 66888 2400 66918
rect 2901 66915 2967 66918
rect 6686 66944 7002 66945
rect 6686 66880 6692 66944
rect 6756 66880 6772 66944
rect 6836 66880 6852 66944
rect 6916 66880 6932 66944
rect 6996 66880 7002 66944
rect 10126 66880 10186 67054
rect 86897 66978 86963 66981
rect 83542 66976 86963 66978
rect 83542 66920 86902 66976
rect 86958 66920 86963 66976
rect 88277 66978 88343 66981
rect 89200 66978 90000 67008
rect 88277 66976 90000 66978
rect 83542 66918 86963 66920
rect 83542 66910 83602 66918
rect 86897 66915 86963 66918
rect 87278 66944 87594 66945
rect 6686 66879 7002 66880
rect 45668 66850 46250 66910
rect 83020 66850 83602 66910
rect 87278 66880 87284 66944
rect 87348 66880 87364 66944
rect 87428 66880 87444 66944
rect 87508 66880 87524 66944
rect 87588 66880 87594 66944
rect 88277 66920 88282 66976
rect 88338 66920 90000 66976
rect 88277 66918 90000 66920
rect 88277 66915 88343 66918
rect 89200 66888 90000 66918
rect 87278 66879 87594 66880
rect 46190 66842 46250 66850
rect 46190 66782 47508 66842
rect 5950 66400 6266 66401
rect 5950 66336 5956 66400
rect 6020 66336 6036 66400
rect 6100 66336 6116 66400
rect 6180 66336 6196 66400
rect 6260 66336 6266 66400
rect 5950 66335 6266 66336
rect 86542 66400 86858 66401
rect 86542 66336 86548 66400
rect 86612 66336 86628 66400
rect 86692 66336 86708 66400
rect 86772 66336 86788 66400
rect 86852 66336 86858 66400
rect 86542 66335 86858 66336
rect 7225 65890 7291 65893
rect 87081 65890 87147 65893
rect 7225 65888 10186 65890
rect 6686 65856 7002 65857
rect 6686 65792 6692 65856
rect 6756 65792 6772 65856
rect 6836 65792 6852 65856
rect 6916 65792 6932 65856
rect 6996 65792 7002 65856
rect 7225 65832 7230 65888
rect 7286 65832 10186 65888
rect 7225 65830 10186 65832
rect 7225 65827 7291 65830
rect 10126 65792 10186 65830
rect 83542 65888 87147 65890
rect 83542 65832 87086 65888
rect 87142 65832 87147 65888
rect 83542 65830 87147 65832
rect 83542 65822 83602 65830
rect 87081 65827 87147 65830
rect 87278 65856 87594 65857
rect 6686 65791 7002 65792
rect 45668 65762 46250 65822
rect 83020 65762 83602 65822
rect 87278 65792 87284 65856
rect 87348 65792 87364 65856
rect 87428 65792 87444 65856
rect 87508 65792 87524 65856
rect 87588 65792 87594 65856
rect 87278 65791 87594 65792
rect 46190 65754 46250 65762
rect 46190 65694 47508 65754
rect 1600 65618 2400 65648
rect 2901 65618 2967 65621
rect 1600 65616 2967 65618
rect 1600 65560 2906 65616
rect 2962 65560 2967 65616
rect 1600 65558 2967 65560
rect 1600 65528 2400 65558
rect 2901 65555 2967 65558
rect 88185 65618 88251 65621
rect 89200 65618 90000 65648
rect 88185 65616 90000 65618
rect 88185 65560 88190 65616
rect 88246 65560 90000 65616
rect 88185 65558 90000 65560
rect 88185 65555 88251 65558
rect 89200 65528 90000 65558
rect 5950 65312 6266 65313
rect 5950 65248 5956 65312
rect 6020 65248 6036 65312
rect 6100 65248 6116 65312
rect 6180 65248 6196 65312
rect 6260 65248 6266 65312
rect 5950 65247 6266 65248
rect 86542 65312 86858 65313
rect 86542 65248 86548 65312
rect 86612 65248 86628 65312
rect 86692 65248 86708 65312
rect 86772 65248 86788 65312
rect 86852 65248 86858 65312
rect 86542 65247 86858 65248
rect 1600 64938 2400 64968
rect 2901 64938 2967 64941
rect 1600 64936 2967 64938
rect 1600 64880 2906 64936
rect 2962 64880 2967 64936
rect 1600 64878 2967 64880
rect 1600 64848 2400 64878
rect 2901 64875 2967 64878
rect 88369 64938 88435 64941
rect 89200 64938 90000 64968
rect 88369 64936 90000 64938
rect 88369 64880 88374 64936
rect 88430 64880 90000 64936
rect 88369 64878 90000 64880
rect 88369 64875 88435 64878
rect 89200 64848 90000 64878
rect 7225 64802 7291 64805
rect 87081 64802 87147 64805
rect 7225 64800 10186 64802
rect 6686 64768 7002 64769
rect 6686 64704 6692 64768
rect 6756 64704 6772 64768
rect 6836 64704 6852 64768
rect 6916 64704 6932 64768
rect 6996 64704 7002 64768
rect 7225 64744 7230 64800
rect 7286 64744 10186 64800
rect 7225 64742 10186 64744
rect 7225 64739 7291 64742
rect 10126 64704 10186 64742
rect 83542 64800 87147 64802
rect 83542 64744 87086 64800
rect 87142 64744 87147 64800
rect 83542 64742 87147 64744
rect 83542 64734 83602 64742
rect 87081 64739 87147 64742
rect 87278 64768 87594 64769
rect 6686 64703 7002 64704
rect 45668 64674 46250 64734
rect 83020 64674 83602 64734
rect 87278 64704 87284 64768
rect 87348 64704 87364 64768
rect 87428 64704 87444 64768
rect 87508 64704 87524 64768
rect 87588 64704 87594 64768
rect 87278 64703 87594 64704
rect 46190 64666 46250 64674
rect 46190 64606 47508 64666
rect 5950 64224 6266 64225
rect 5950 64160 5956 64224
rect 6020 64160 6036 64224
rect 6100 64160 6116 64224
rect 6180 64160 6196 64224
rect 6260 64160 6266 64224
rect 5950 64159 6266 64160
rect 86542 64224 86858 64225
rect 86542 64160 86548 64224
rect 86612 64160 86628 64224
rect 86692 64160 86708 64224
rect 86772 64160 86788 64224
rect 86852 64160 86858 64224
rect 86542 64159 86858 64160
rect 84413 63714 84479 63717
rect 83358 63712 84479 63714
rect 6686 63680 7002 63681
rect 6686 63616 6692 63680
rect 6756 63616 6772 63680
rect 6836 63616 6852 63680
rect 6916 63616 6932 63680
rect 6996 63616 7002 63680
rect 83358 63656 84418 63712
rect 84474 63656 84479 63712
rect 83358 63654 84479 63656
rect 6686 63615 7002 63616
rect 9617 63646 9683 63649
rect 83358 63646 83418 63654
rect 84413 63651 84479 63654
rect 87278 63680 87594 63681
rect 9617 63644 10156 63646
rect 1600 63578 2400 63608
rect 9617 63588 9622 63644
rect 9678 63588 10156 63644
rect 9617 63586 10156 63588
rect 45668 63586 46250 63646
rect 83020 63586 83418 63646
rect 87278 63616 87284 63680
rect 87348 63616 87364 63680
rect 87428 63616 87444 63680
rect 87508 63616 87524 63680
rect 87588 63616 87594 63680
rect 87278 63615 87594 63616
rect 9617 63583 9683 63586
rect 5201 63578 5267 63581
rect 1600 63576 5267 63578
rect 1600 63520 5206 63576
rect 5262 63520 5267 63576
rect 1600 63518 5267 63520
rect 46190 63578 46250 63586
rect 88553 63578 88619 63581
rect 89200 63578 90000 63608
rect 46190 63518 47508 63578
rect 88553 63576 90000 63578
rect 88553 63520 88558 63576
rect 88614 63520 90000 63576
rect 88553 63518 90000 63520
rect 1600 63488 2400 63518
rect 5201 63515 5267 63518
rect 88553 63515 88619 63518
rect 89200 63488 90000 63518
rect 5950 63136 6266 63137
rect 5950 63072 5956 63136
rect 6020 63072 6036 63136
rect 6100 63072 6116 63136
rect 6180 63072 6196 63136
rect 6260 63072 6266 63136
rect 5950 63071 6266 63072
rect 86542 63136 86858 63137
rect 86542 63072 86548 63136
rect 86612 63072 86628 63136
rect 86692 63072 86708 63136
rect 86772 63072 86788 63136
rect 86852 63072 86858 63136
rect 86542 63071 86858 63072
rect 6686 62592 7002 62593
rect 6686 62528 6692 62592
rect 6756 62528 6772 62592
rect 6836 62528 6852 62592
rect 6916 62528 6932 62592
rect 6996 62528 7002 62592
rect 87278 62592 87594 62593
rect 6686 62527 7002 62528
rect 45668 62498 46250 62558
rect 83020 62498 83602 62558
rect 87278 62528 87284 62592
rect 87348 62528 87364 62592
rect 87428 62528 87444 62592
rect 87508 62528 87524 62592
rect 87588 62528 87594 62592
rect 87278 62527 87594 62528
rect 7225 62490 7291 62493
rect 46190 62490 46250 62498
rect 83542 62490 83602 62498
rect 87081 62490 87147 62493
rect 7225 62488 10156 62490
rect 7225 62432 7230 62488
rect 7286 62432 10156 62488
rect 7225 62430 10156 62432
rect 46190 62430 47508 62490
rect 83542 62488 87147 62490
rect 83542 62432 87086 62488
rect 87142 62432 87147 62488
rect 83542 62430 87147 62432
rect 7225 62427 7291 62430
rect 87081 62427 87147 62430
rect 1600 62218 2400 62248
rect 4925 62218 4991 62221
rect 1600 62216 4991 62218
rect 1600 62160 4930 62216
rect 4986 62160 4991 62216
rect 1600 62158 4991 62160
rect 1600 62128 2400 62158
rect 4925 62155 4991 62158
rect 88553 62218 88619 62221
rect 89200 62218 90000 62248
rect 88553 62216 90000 62218
rect 88553 62160 88558 62216
rect 88614 62160 90000 62216
rect 88553 62158 90000 62160
rect 88553 62155 88619 62158
rect 89200 62128 90000 62158
rect 5950 62048 6266 62049
rect 5950 61984 5956 62048
rect 6020 61984 6036 62048
rect 6100 61984 6116 62048
rect 6180 61984 6196 62048
rect 6260 61984 6266 62048
rect 5950 61983 6266 61984
rect 86542 62048 86858 62049
rect 86542 61984 86548 62048
rect 86612 61984 86628 62048
rect 86692 61984 86708 62048
rect 86772 61984 86788 62048
rect 86852 61984 86858 62048
rect 86542 61983 86858 61984
rect 1600 61538 2400 61568
rect 2901 61538 2967 61541
rect 1600 61536 2967 61538
rect 1600 61480 2906 61536
rect 2962 61480 2967 61536
rect 7225 61538 7291 61541
rect 87081 61538 87147 61541
rect 7225 61536 10186 61538
rect 1600 61478 2967 61480
rect 1600 61448 2400 61478
rect 2901 61475 2967 61478
rect 6686 61504 7002 61505
rect 6686 61440 6692 61504
rect 6756 61440 6772 61504
rect 6836 61440 6852 61504
rect 6916 61440 6932 61504
rect 6996 61440 7002 61504
rect 7225 61480 7230 61536
rect 7286 61480 10186 61536
rect 7225 61478 10186 61480
rect 7225 61475 7291 61478
rect 10126 61440 10186 61478
rect 83542 61536 87147 61538
rect 83542 61480 87086 61536
rect 87142 61480 87147 61536
rect 88185 61538 88251 61541
rect 89200 61538 90000 61568
rect 88185 61536 90000 61538
rect 83542 61478 87147 61480
rect 83542 61470 83602 61478
rect 87081 61475 87147 61478
rect 87278 61504 87594 61505
rect 6686 61439 7002 61440
rect 45668 61410 46250 61470
rect 83020 61410 83602 61470
rect 87278 61440 87284 61504
rect 87348 61440 87364 61504
rect 87428 61440 87444 61504
rect 87508 61440 87524 61504
rect 87588 61440 87594 61504
rect 88185 61480 88190 61536
rect 88246 61480 90000 61536
rect 88185 61478 90000 61480
rect 88185 61475 88251 61478
rect 89200 61448 90000 61478
rect 87278 61439 87594 61440
rect 46190 61402 46250 61410
rect 46190 61342 47508 61402
rect 5950 60960 6266 60961
rect 5950 60896 5956 60960
rect 6020 60896 6036 60960
rect 6100 60896 6116 60960
rect 6180 60896 6196 60960
rect 6260 60896 6266 60960
rect 5950 60895 6266 60896
rect 86542 60960 86858 60961
rect 86542 60896 86548 60960
rect 86612 60896 86628 60960
rect 86692 60896 86708 60960
rect 86772 60896 86788 60960
rect 86852 60896 86858 60960
rect 86542 60895 86858 60896
rect 7225 60450 7291 60453
rect 87081 60450 87147 60453
rect 7225 60448 10186 60450
rect 6686 60416 7002 60417
rect 6686 60352 6692 60416
rect 6756 60352 6772 60416
rect 6836 60352 6852 60416
rect 6916 60352 6932 60416
rect 6996 60352 7002 60416
rect 7225 60392 7230 60448
rect 7286 60392 10186 60448
rect 7225 60390 10186 60392
rect 7225 60387 7291 60390
rect 10126 60352 10186 60390
rect 83542 60448 87147 60450
rect 83542 60392 87086 60448
rect 87142 60392 87147 60448
rect 83542 60390 87147 60392
rect 83542 60382 83602 60390
rect 87081 60387 87147 60390
rect 87278 60416 87594 60417
rect 6686 60351 7002 60352
rect 45668 60322 46250 60382
rect 83020 60322 83602 60382
rect 87278 60352 87284 60416
rect 87348 60352 87364 60416
rect 87428 60352 87444 60416
rect 87508 60352 87524 60416
rect 87588 60352 87594 60416
rect 87278 60351 87594 60352
rect 46190 60314 46250 60322
rect 46190 60254 47508 60314
rect 1600 60178 2400 60208
rect 2901 60178 2967 60181
rect 1600 60176 2967 60178
rect 1600 60120 2906 60176
rect 2962 60120 2967 60176
rect 1600 60118 2967 60120
rect 1600 60088 2400 60118
rect 2901 60115 2967 60118
rect 88185 60178 88251 60181
rect 89200 60178 90000 60208
rect 88185 60176 90000 60178
rect 88185 60120 88190 60176
rect 88246 60120 90000 60176
rect 88185 60118 90000 60120
rect 88185 60115 88251 60118
rect 89200 60088 90000 60118
rect 5950 59872 6266 59873
rect 5950 59808 5956 59872
rect 6020 59808 6036 59872
rect 6100 59808 6116 59872
rect 6180 59808 6196 59872
rect 6260 59808 6266 59872
rect 5950 59807 6266 59808
rect 86542 59872 86858 59873
rect 86542 59808 86548 59872
rect 86612 59808 86628 59872
rect 86692 59808 86708 59872
rect 86772 59808 86788 59872
rect 86852 59808 86858 59872
rect 86542 59807 86858 59808
rect 1600 59498 2400 59528
rect 5201 59498 5267 59501
rect 87633 59498 87699 59501
rect 1600 59496 5267 59498
rect 1600 59440 5206 59496
rect 5262 59440 5267 59496
rect 1600 59438 5267 59440
rect 1600 59408 2400 59438
rect 5201 59435 5267 59438
rect 85750 59496 87699 59498
rect 85750 59440 87638 59496
rect 87694 59440 87699 59496
rect 85750 59438 87699 59440
rect 7225 59362 7291 59365
rect 85750 59362 85810 59438
rect 87633 59435 87699 59438
rect 88369 59498 88435 59501
rect 89200 59498 90000 59528
rect 88369 59496 90000 59498
rect 88369 59440 88374 59496
rect 88430 59440 90000 59496
rect 88369 59438 90000 59440
rect 88369 59435 88435 59438
rect 89200 59408 90000 59438
rect 7225 59360 10186 59362
rect 6686 59328 7002 59329
rect 6686 59264 6692 59328
rect 6756 59264 6772 59328
rect 6836 59264 6852 59328
rect 6916 59264 6932 59328
rect 6996 59264 7002 59328
rect 7225 59304 7230 59360
rect 7286 59304 10186 59360
rect 7225 59302 10186 59304
rect 7225 59299 7291 59302
rect 10126 59264 10186 59302
rect 83542 59302 85810 59362
rect 87278 59328 87594 59329
rect 83542 59294 83602 59302
rect 6686 59263 7002 59264
rect 45668 59234 46250 59294
rect 83020 59234 83602 59294
rect 87278 59264 87284 59328
rect 87348 59264 87364 59328
rect 87428 59264 87444 59328
rect 87508 59264 87524 59328
rect 87588 59264 87594 59328
rect 87278 59263 87594 59264
rect 46190 59226 46250 59234
rect 46190 59166 47508 59226
rect 5950 58784 6266 58785
rect 5950 58720 5956 58784
rect 6020 58720 6036 58784
rect 6100 58720 6116 58784
rect 6180 58720 6196 58784
rect 6260 58720 6266 58784
rect 5950 58719 6266 58720
rect 86542 58784 86858 58785
rect 86542 58720 86548 58784
rect 86612 58720 86628 58784
rect 86692 58720 86708 58784
rect 86772 58720 86788 58784
rect 86852 58720 86858 58784
rect 86542 58719 86858 58720
rect 6686 58240 7002 58241
rect 6686 58176 6692 58240
rect 6756 58176 6772 58240
rect 6836 58176 6852 58240
rect 6916 58176 6932 58240
rect 6996 58176 7002 58240
rect 87278 58240 87594 58241
rect 6686 58175 7002 58176
rect 1600 58138 2400 58168
rect 45668 58146 46250 58206
rect 83020 58146 83602 58206
rect 87278 58176 87284 58240
rect 87348 58176 87364 58240
rect 87428 58176 87444 58240
rect 87508 58176 87524 58240
rect 87588 58176 87594 58240
rect 87278 58175 87594 58176
rect 5201 58138 5267 58141
rect 1600 58136 5267 58138
rect 1600 58080 5206 58136
rect 5262 58080 5267 58136
rect 46190 58138 46250 58146
rect 83542 58138 83602 58146
rect 88553 58138 88619 58141
rect 89200 58138 90000 58168
rect 1600 58078 5267 58080
rect 1600 58048 2400 58078
rect 5201 58075 5267 58078
rect 5385 58002 5451 58005
rect 10126 58002 10186 58108
rect 46190 58078 47508 58138
rect 83542 58078 85810 58138
rect 5385 58000 10186 58002
rect 5385 57944 5390 58000
rect 5446 57944 10186 58000
rect 5385 57942 10186 57944
rect 85750 58002 85810 58078
rect 88553 58136 90000 58138
rect 88553 58080 88558 58136
rect 88614 58080 90000 58136
rect 88553 58078 90000 58080
rect 88553 58075 88619 58078
rect 89200 58048 90000 58078
rect 88001 58002 88067 58005
rect 85750 58000 88067 58002
rect 85750 57944 88006 58000
rect 88062 57944 88067 58000
rect 85750 57942 88067 57944
rect 5385 57939 5451 57942
rect 88001 57939 88067 57942
rect 5950 57696 6266 57697
rect 5950 57632 5956 57696
rect 6020 57632 6036 57696
rect 6100 57632 6116 57696
rect 6180 57632 6196 57696
rect 6260 57632 6266 57696
rect 5950 57631 6266 57632
rect 86542 57696 86858 57697
rect 86542 57632 86548 57696
rect 86612 57632 86628 57696
rect 86692 57632 86708 57696
rect 86772 57632 86788 57696
rect 86852 57632 86858 57696
rect 86542 57631 86858 57632
rect 6686 57152 7002 57153
rect 6686 57088 6692 57152
rect 6756 57088 6772 57152
rect 6836 57088 6852 57152
rect 6916 57088 6932 57152
rect 6996 57088 7002 57152
rect 87278 57152 87594 57153
rect 6686 57087 7002 57088
rect 45668 57058 46250 57118
rect 83020 57058 83602 57118
rect 87278 57088 87284 57152
rect 87348 57088 87364 57152
rect 87428 57088 87444 57152
rect 87508 57088 87524 57152
rect 87588 57088 87594 57152
rect 87278 57087 87594 57088
rect 7225 57050 7291 57053
rect 46190 57050 46250 57058
rect 83542 57050 83602 57058
rect 7225 57048 10156 57050
rect 7225 56992 7230 57048
rect 7286 56992 10156 57048
rect 7225 56990 10156 56992
rect 46190 56990 47508 57050
rect 83542 56990 85810 57050
rect 7225 56987 7291 56990
rect 85750 56914 85810 56990
rect 88001 56914 88067 56917
rect 85750 56912 88067 56914
rect 85750 56856 88006 56912
rect 88062 56856 88067 56912
rect 85750 56854 88067 56856
rect 88001 56851 88067 56854
rect 1600 56778 2400 56808
rect 4925 56778 4991 56781
rect 1600 56776 4991 56778
rect 1600 56720 4930 56776
rect 4986 56720 4991 56776
rect 1600 56718 4991 56720
rect 1600 56688 2400 56718
rect 4925 56715 4991 56718
rect 88829 56778 88895 56781
rect 89200 56778 90000 56808
rect 88829 56776 90000 56778
rect 88829 56720 88834 56776
rect 88890 56720 90000 56776
rect 88829 56718 90000 56720
rect 88829 56715 88895 56718
rect 89200 56688 90000 56718
rect 5950 56608 6266 56609
rect 5950 56544 5956 56608
rect 6020 56544 6036 56608
rect 6100 56544 6116 56608
rect 6180 56544 6196 56608
rect 6260 56544 6266 56608
rect 5950 56543 6266 56544
rect 86542 56608 86858 56609
rect 86542 56544 86548 56608
rect 86612 56544 86628 56608
rect 86692 56544 86708 56608
rect 86772 56544 86788 56608
rect 86852 56544 86858 56608
rect 86542 56543 86858 56544
rect 1600 56098 2400 56128
rect 2901 56098 2967 56101
rect 1600 56096 2967 56098
rect 1600 56040 2906 56096
rect 2962 56040 2967 56096
rect 7225 56098 7291 56101
rect 87081 56098 87147 56101
rect 7225 56096 10186 56098
rect 1600 56038 2967 56040
rect 1600 56008 2400 56038
rect 2901 56035 2967 56038
rect 6686 56064 7002 56065
rect 6686 56000 6692 56064
rect 6756 56000 6772 56064
rect 6836 56000 6852 56064
rect 6916 56000 6932 56064
rect 6996 56000 7002 56064
rect 7225 56040 7230 56096
rect 7286 56040 10186 56096
rect 7225 56038 10186 56040
rect 7225 56035 7291 56038
rect 10126 56000 10186 56038
rect 83542 56096 87147 56098
rect 83542 56040 87086 56096
rect 87142 56040 87147 56096
rect 88185 56098 88251 56101
rect 89200 56098 90000 56128
rect 88185 56096 90000 56098
rect 83542 56038 87147 56040
rect 83542 56030 83602 56038
rect 87081 56035 87147 56038
rect 87278 56064 87594 56065
rect 6686 55999 7002 56000
rect 45668 55970 46250 56030
rect 83020 55970 83602 56030
rect 87278 56000 87284 56064
rect 87348 56000 87364 56064
rect 87428 56000 87444 56064
rect 87508 56000 87524 56064
rect 87588 56000 87594 56064
rect 88185 56040 88190 56096
rect 88246 56040 90000 56096
rect 88185 56038 90000 56040
rect 88185 56035 88251 56038
rect 89200 56008 90000 56038
rect 87278 55999 87594 56000
rect 46190 55962 46250 55970
rect 46190 55902 47508 55962
rect 5950 55520 6266 55521
rect 5950 55456 5956 55520
rect 6020 55456 6036 55520
rect 6100 55456 6116 55520
rect 6180 55456 6196 55520
rect 6260 55456 6266 55520
rect 5950 55455 6266 55456
rect 86542 55520 86858 55521
rect 86542 55456 86548 55520
rect 86612 55456 86628 55520
rect 86692 55456 86708 55520
rect 86772 55456 86788 55520
rect 86852 55456 86858 55520
rect 86542 55455 86858 55456
rect 7225 55010 7291 55013
rect 87081 55010 87147 55013
rect 7225 55008 10186 55010
rect 6686 54976 7002 54977
rect 6686 54912 6692 54976
rect 6756 54912 6772 54976
rect 6836 54912 6852 54976
rect 6916 54912 6932 54976
rect 6996 54912 7002 54976
rect 7225 54952 7230 55008
rect 7286 54952 10186 55008
rect 7225 54950 10186 54952
rect 7225 54947 7291 54950
rect 10126 54912 10186 54950
rect 83542 55008 87147 55010
rect 83542 54952 87086 55008
rect 87142 54952 87147 55008
rect 83542 54950 87147 54952
rect 83542 54942 83602 54950
rect 87081 54947 87147 54950
rect 87278 54976 87594 54977
rect 6686 54911 7002 54912
rect 45668 54882 46250 54942
rect 83020 54882 83602 54942
rect 87278 54912 87284 54976
rect 87348 54912 87364 54976
rect 87428 54912 87444 54976
rect 87508 54912 87524 54976
rect 87588 54912 87594 54976
rect 87278 54911 87594 54912
rect 46190 54874 46250 54882
rect 46190 54814 47508 54874
rect 1600 54738 2400 54768
rect 2901 54738 2967 54741
rect 1600 54736 2967 54738
rect 1600 54680 2906 54736
rect 2962 54680 2967 54736
rect 1600 54678 2967 54680
rect 1600 54648 2400 54678
rect 2901 54675 2967 54678
rect 88185 54738 88251 54741
rect 89200 54738 90000 54768
rect 88185 54736 90000 54738
rect 88185 54680 88190 54736
rect 88246 54680 90000 54736
rect 88185 54678 90000 54680
rect 88185 54675 88251 54678
rect 89200 54648 90000 54678
rect 5950 54432 6266 54433
rect 5950 54368 5956 54432
rect 6020 54368 6036 54432
rect 6100 54368 6116 54432
rect 6180 54368 6196 54432
rect 6260 54368 6266 54432
rect 5950 54367 6266 54368
rect 86542 54432 86858 54433
rect 86542 54368 86548 54432
rect 86612 54368 86628 54432
rect 86692 54368 86708 54432
rect 86772 54368 86788 54432
rect 86852 54368 86858 54432
rect 86542 54367 86858 54368
rect 1600 54058 2400 54088
rect 5109 54058 5175 54061
rect 1600 54056 5175 54058
rect 1600 54000 5114 54056
rect 5170 54000 5175 54056
rect 1600 53998 5175 54000
rect 1600 53968 2400 53998
rect 5109 53995 5175 53998
rect 5661 54058 5727 54061
rect 88645 54058 88711 54061
rect 89200 54058 90000 54088
rect 5661 54056 10186 54058
rect 5661 54000 5666 54056
rect 5722 54000 10186 54056
rect 5661 53998 10186 54000
rect 5661 53995 5727 53998
rect 6686 53888 7002 53889
rect 6686 53824 6692 53888
rect 6756 53824 6772 53888
rect 6836 53824 6852 53888
rect 6916 53824 6932 53888
rect 6996 53824 7002 53888
rect 10126 53824 10186 53998
rect 88645 54056 90000 54058
rect 88645 54000 88650 54056
rect 88706 54000 90000 54056
rect 88645 53998 90000 54000
rect 88645 53995 88711 53998
rect 89200 53968 90000 53998
rect 84413 53922 84479 53925
rect 83358 53920 84479 53922
rect 83358 53864 84418 53920
rect 84474 53864 84479 53920
rect 83358 53862 84479 53864
rect 83358 53854 83418 53862
rect 84413 53859 84479 53862
rect 87278 53888 87594 53889
rect 6686 53823 7002 53824
rect 45668 53794 46250 53854
rect 83020 53794 83418 53854
rect 87278 53824 87284 53888
rect 87348 53824 87364 53888
rect 87428 53824 87444 53888
rect 87508 53824 87524 53888
rect 87588 53824 87594 53888
rect 87278 53823 87594 53824
rect 46190 53786 46250 53794
rect 46190 53726 47508 53786
rect 5950 53344 6266 53345
rect 5950 53280 5956 53344
rect 6020 53280 6036 53344
rect 6100 53280 6116 53344
rect 6180 53280 6196 53344
rect 6260 53280 6266 53344
rect 5950 53279 6266 53280
rect 86542 53344 86858 53345
rect 86542 53280 86548 53344
rect 86612 53280 86628 53344
rect 86692 53280 86708 53344
rect 86772 53280 86788 53344
rect 86852 53280 86858 53344
rect 86542 53279 86858 53280
rect 7225 52834 7291 52837
rect 87081 52834 87147 52837
rect 7225 52832 10186 52834
rect 6686 52800 7002 52801
rect 6686 52736 6692 52800
rect 6756 52736 6772 52800
rect 6836 52736 6852 52800
rect 6916 52736 6932 52800
rect 6996 52736 7002 52800
rect 7225 52776 7230 52832
rect 7286 52776 10186 52832
rect 7225 52774 10186 52776
rect 7225 52771 7291 52774
rect 10126 52736 10186 52774
rect 83542 52832 87147 52834
rect 83542 52776 87086 52832
rect 87142 52776 87147 52832
rect 83542 52774 87147 52776
rect 83542 52766 83602 52774
rect 87081 52771 87147 52774
rect 87278 52800 87594 52801
rect 6686 52735 7002 52736
rect 1600 52698 2400 52728
rect 45668 52706 46066 52766
rect 83020 52706 83602 52766
rect 87278 52736 87284 52800
rect 87348 52736 87364 52800
rect 87428 52736 87444 52800
rect 87508 52736 87524 52800
rect 87588 52736 87594 52800
rect 87278 52735 87594 52736
rect 2901 52698 2967 52701
rect 1600 52696 2967 52698
rect 1600 52640 2906 52696
rect 2962 52640 2967 52696
rect 1600 52638 2967 52640
rect 46006 52698 46066 52706
rect 88277 52698 88343 52701
rect 89200 52698 90000 52728
rect 46006 52638 47508 52698
rect 88277 52696 90000 52698
rect 88277 52640 88282 52696
rect 88338 52640 90000 52696
rect 88277 52638 90000 52640
rect 1600 52608 2400 52638
rect 2901 52635 2967 52638
rect 88277 52635 88343 52638
rect 89200 52608 90000 52638
rect 5950 52256 6266 52257
rect 5950 52192 5956 52256
rect 6020 52192 6036 52256
rect 6100 52192 6116 52256
rect 6180 52192 6196 52256
rect 6260 52192 6266 52256
rect 5950 52191 6266 52192
rect 86542 52256 86858 52257
rect 86542 52192 86548 52256
rect 86612 52192 86628 52256
rect 86692 52192 86708 52256
rect 86772 52192 86788 52256
rect 86852 52192 86858 52256
rect 86542 52191 86858 52192
rect 6686 51712 7002 51713
rect 6686 51648 6692 51712
rect 6756 51648 6772 51712
rect 6836 51648 6852 51712
rect 6916 51648 6932 51712
rect 6996 51648 7002 51712
rect 87278 51712 87594 51713
rect 6686 51647 7002 51648
rect 45668 51618 46250 51678
rect 83020 51618 83418 51678
rect 87278 51648 87284 51712
rect 87348 51648 87364 51712
rect 87428 51648 87444 51712
rect 87508 51648 87524 51712
rect 87588 51648 87594 51712
rect 87278 51647 87594 51648
rect 7225 51610 7291 51613
rect 46190 51610 46250 51618
rect 83358 51610 83418 51618
rect 85793 51610 85859 51613
rect 7225 51608 10156 51610
rect 7225 51552 7230 51608
rect 7286 51552 10156 51608
rect 7225 51550 10156 51552
rect 46190 51550 47508 51610
rect 83358 51608 85859 51610
rect 83358 51552 85798 51608
rect 85854 51552 85859 51608
rect 83358 51550 85859 51552
rect 7225 51547 7291 51550
rect 85793 51547 85859 51550
rect 1600 51338 2400 51368
rect 2901 51338 2967 51341
rect 1600 51336 2967 51338
rect 1600 51280 2906 51336
rect 2962 51280 2967 51336
rect 1600 51278 2967 51280
rect 1600 51248 2400 51278
rect 2901 51275 2967 51278
rect 88185 51338 88251 51341
rect 89200 51338 90000 51368
rect 88185 51336 90000 51338
rect 88185 51280 88190 51336
rect 88246 51280 90000 51336
rect 88185 51278 90000 51280
rect 88185 51275 88251 51278
rect 89200 51248 90000 51278
rect 5950 51168 6266 51169
rect 5950 51104 5956 51168
rect 6020 51104 6036 51168
rect 6100 51104 6116 51168
rect 6180 51104 6196 51168
rect 6260 51104 6266 51168
rect 5950 51103 6266 51104
rect 86542 51168 86858 51169
rect 86542 51104 86548 51168
rect 86612 51104 86628 51168
rect 86692 51104 86708 51168
rect 86772 51104 86788 51168
rect 86852 51104 86858 51168
rect 86542 51103 86858 51104
rect 6686 50624 7002 50625
rect 6686 50560 6692 50624
rect 6756 50560 6772 50624
rect 6836 50560 6852 50624
rect 6916 50560 6932 50624
rect 6996 50560 7002 50624
rect 87278 50624 87594 50625
rect 45957 50590 46023 50593
rect 6686 50559 7002 50560
rect 45668 50588 46023 50590
rect 45668 50532 45962 50588
rect 46018 50532 46023 50588
rect 45668 50530 46023 50532
rect 83020 50530 83418 50590
rect 87278 50560 87284 50624
rect 87348 50560 87364 50624
rect 87428 50560 87444 50624
rect 87508 50560 87524 50624
rect 87588 50560 87594 50624
rect 87278 50559 87594 50560
rect 45957 50527 46023 50530
rect 83358 50522 83418 50530
rect 85425 50522 85491 50525
rect 83358 50520 85491 50522
rect 83358 50464 85430 50520
rect 85486 50464 85491 50520
rect 83358 50462 85491 50464
rect 85425 50459 85491 50462
rect 5950 50080 6266 50081
rect 5950 50016 5956 50080
rect 6020 50016 6036 50080
rect 6100 50016 6116 50080
rect 6180 50016 6196 50080
rect 6260 50016 6266 50080
rect 5950 50015 6266 50016
rect 86542 50080 86858 50081
rect 86542 50016 86548 50080
rect 86612 50016 86628 50080
rect 86692 50016 86708 50080
rect 86772 50016 86788 50080
rect 86852 50016 86858 50080
rect 86542 50015 86858 50016
rect 6686 49536 7002 49537
rect 6686 49472 6692 49536
rect 6756 49472 6772 49536
rect 6836 49472 6852 49536
rect 6916 49472 6932 49536
rect 6996 49472 7002 49536
rect 87278 49536 87594 49537
rect 45865 49502 45931 49505
rect 6686 49471 7002 49472
rect 45668 49500 45931 49502
rect 45668 49444 45870 49500
rect 45926 49444 45931 49500
rect 45668 49442 45931 49444
rect 83020 49442 83418 49502
rect 87278 49472 87284 49536
rect 87348 49472 87364 49536
rect 87428 49472 87444 49536
rect 87508 49472 87524 49536
rect 87588 49472 87594 49536
rect 87278 49471 87594 49472
rect 45865 49439 45931 49442
rect 83358 49434 83418 49442
rect 85517 49434 85583 49437
rect 83358 49432 85583 49434
rect 83358 49376 85522 49432
rect 85578 49376 85583 49432
rect 83358 49374 85583 49376
rect 85517 49371 85583 49374
rect 5950 48992 6266 48993
rect 5950 48928 5956 48992
rect 6020 48928 6036 48992
rect 6100 48928 6116 48992
rect 6180 48928 6196 48992
rect 6260 48928 6266 48992
rect 5950 48927 6266 48928
rect 86542 48992 86858 48993
rect 86542 48928 86548 48992
rect 86612 48928 86628 48992
rect 86692 48928 86708 48992
rect 86772 48928 86788 48992
rect 86852 48928 86858 48992
rect 86542 48927 86858 48928
rect 88185 48618 88251 48621
rect 89200 48618 90000 48648
rect 88185 48616 90000 48618
rect 88185 48560 88190 48616
rect 88246 48560 90000 48616
rect 88185 48558 90000 48560
rect 88185 48555 88251 48558
rect 89200 48528 90000 48558
rect 6686 48448 7002 48449
rect 6686 48384 6692 48448
rect 6756 48384 6772 48448
rect 6836 48384 6852 48448
rect 6916 48384 6932 48448
rect 6996 48384 7002 48448
rect 87278 48448 87594 48449
rect 46049 48414 46115 48417
rect 6686 48383 7002 48384
rect 45668 48412 46115 48414
rect 45668 48356 46054 48412
rect 46110 48356 46115 48412
rect 45668 48354 46115 48356
rect 83020 48354 83418 48414
rect 87278 48384 87284 48448
rect 87348 48384 87364 48448
rect 87428 48384 87444 48448
rect 87508 48384 87524 48448
rect 87588 48384 87594 48448
rect 87278 48383 87594 48384
rect 46049 48351 46115 48354
rect 83358 48346 83418 48354
rect 85333 48346 85399 48349
rect 83358 48344 85399 48346
rect 83358 48288 85338 48344
rect 85394 48288 85399 48344
rect 83358 48286 85399 48288
rect 85333 48283 85399 48286
rect 88185 47938 88251 47941
rect 89200 47938 90000 47968
rect 88185 47936 90000 47938
rect 5950 47904 6266 47905
rect 5950 47840 5956 47904
rect 6020 47840 6036 47904
rect 6100 47840 6116 47904
rect 6180 47840 6196 47904
rect 6260 47840 6266 47904
rect 5950 47839 6266 47840
rect 86542 47904 86858 47905
rect 86542 47840 86548 47904
rect 86612 47840 86628 47904
rect 86692 47840 86708 47904
rect 86772 47840 86788 47904
rect 86852 47840 86858 47904
rect 88185 47880 88190 47936
rect 88246 47880 90000 47936
rect 88185 47878 90000 47880
rect 88185 47875 88251 47878
rect 89200 47848 90000 47878
rect 86542 47839 86858 47840
rect 85793 47394 85859 47397
rect 83358 47392 85859 47394
rect 6686 47360 7002 47361
rect 6686 47296 6692 47360
rect 6756 47296 6772 47360
rect 6836 47296 6852 47360
rect 6916 47296 6932 47360
rect 6996 47296 7002 47360
rect 83358 47336 85798 47392
rect 85854 47336 85859 47392
rect 83358 47334 85859 47336
rect 46141 47326 46207 47329
rect 83358 47326 83418 47334
rect 85793 47331 85859 47334
rect 87278 47360 87594 47361
rect 6686 47295 7002 47296
rect 45668 47324 46207 47326
rect 45668 47268 46146 47324
rect 46202 47268 46207 47324
rect 45668 47266 46207 47268
rect 83020 47266 83418 47326
rect 87278 47296 87284 47360
rect 87348 47296 87364 47360
rect 87428 47296 87444 47360
rect 87508 47296 87524 47360
rect 87588 47296 87594 47360
rect 87278 47295 87594 47296
rect 46141 47263 46207 47266
rect 88185 47258 88251 47261
rect 89200 47258 90000 47288
rect 88185 47256 90000 47258
rect 88185 47200 88190 47256
rect 88246 47200 90000 47256
rect 88185 47198 90000 47200
rect 88185 47195 88251 47198
rect 89200 47168 90000 47198
rect 5950 46816 6266 46817
rect 5950 46752 5956 46816
rect 6020 46752 6036 46816
rect 6100 46752 6116 46816
rect 6180 46752 6196 46816
rect 6260 46752 6266 46816
rect 5950 46751 6266 46752
rect 86542 46816 86858 46817
rect 86542 46752 86548 46816
rect 86612 46752 86628 46816
rect 86692 46752 86708 46816
rect 86772 46752 86788 46816
rect 86852 46752 86858 46816
rect 86542 46751 86858 46752
rect 88185 46578 88251 46581
rect 89200 46578 90000 46608
rect 88185 46576 90000 46578
rect 88185 46520 88190 46576
rect 88246 46520 90000 46576
rect 88185 46518 90000 46520
rect 88185 46515 88251 46518
rect 89200 46488 90000 46518
rect 6686 46272 7002 46273
rect 6686 46208 6692 46272
rect 6756 46208 6772 46272
rect 6836 46208 6852 46272
rect 6916 46208 6932 46272
rect 6996 46208 7002 46272
rect 6686 46207 7002 46208
rect 87278 46272 87594 46273
rect 87278 46208 87284 46272
rect 87348 46208 87364 46272
rect 87428 46208 87444 46272
rect 87508 46208 87524 46272
rect 87588 46208 87594 46272
rect 87278 46207 87594 46208
rect 88185 45898 88251 45901
rect 89200 45898 90000 45928
rect 88185 45896 90000 45898
rect 88185 45840 88190 45896
rect 88246 45840 90000 45896
rect 88185 45838 90000 45840
rect 88185 45835 88251 45838
rect 89200 45808 90000 45838
rect 47061 45762 47127 45765
rect 47337 45762 47403 45765
rect 47061 45760 47403 45762
rect 5950 45728 6266 45729
rect 5950 45664 5956 45728
rect 6020 45664 6036 45728
rect 6100 45664 6116 45728
rect 6180 45664 6196 45728
rect 6260 45664 6266 45728
rect 47061 45704 47066 45760
rect 47122 45704 47342 45760
rect 47398 45704 47403 45760
rect 47061 45702 47403 45704
rect 47061 45699 47127 45702
rect 47337 45699 47403 45702
rect 86542 45728 86858 45729
rect 5950 45663 6266 45664
rect 86542 45664 86548 45728
rect 86612 45664 86628 45728
rect 86692 45664 86708 45728
rect 86772 45664 86788 45728
rect 86852 45664 86858 45728
rect 86542 45663 86858 45664
rect 9985 45626 10051 45629
rect 10537 45626 10603 45629
rect 9985 45624 10603 45626
rect 9985 45568 9990 45624
rect 10046 45568 10542 45624
rect 10598 45568 10603 45624
rect 9985 45566 10603 45568
rect 9985 45563 10051 45566
rect 10537 45563 10603 45566
rect 7133 45490 7199 45493
rect 12773 45490 12839 45493
rect 50173 45490 50239 45493
rect 85977 45490 86043 45493
rect 7133 45488 86043 45490
rect 7133 45432 7138 45488
rect 7194 45432 12778 45488
rect 12834 45432 50178 45488
rect 50234 45432 85982 45488
rect 86038 45432 86043 45488
rect 7133 45430 86043 45432
rect 7133 45427 7199 45430
rect 12773 45427 12839 45430
rect 50173 45427 50239 45430
rect 85977 45427 86043 45430
rect 7501 45354 7567 45357
rect 11669 45354 11735 45357
rect 49069 45354 49135 45357
rect 86161 45354 86227 45357
rect 7501 45352 27850 45354
rect 7501 45296 7506 45352
rect 7562 45296 11674 45352
rect 11730 45296 27850 45352
rect 7501 45294 27850 45296
rect 7501 45291 7567 45294
rect 11669 45291 11735 45294
rect 1600 45218 2400 45248
rect 2901 45218 2967 45221
rect 1600 45216 2967 45218
rect 1600 45160 2906 45216
rect 2962 45160 2967 45216
rect 27790 45218 27850 45294
rect 47110 45352 86227 45354
rect 47110 45296 49074 45352
rect 49130 45296 86166 45352
rect 86222 45296 86227 45352
rect 47110 45294 86227 45296
rect 47110 45218 47170 45294
rect 49069 45291 49135 45294
rect 86161 45291 86227 45294
rect 1600 45158 2967 45160
rect 1600 45128 2400 45158
rect 2901 45155 2967 45158
rect 6686 45184 7002 45185
rect 6686 45120 6692 45184
rect 6756 45120 6772 45184
rect 6836 45120 6852 45184
rect 6916 45120 6932 45184
rect 6996 45120 7002 45184
rect 27790 45158 47170 45218
rect 47337 45218 47403 45221
rect 47965 45218 48031 45221
rect 85609 45218 85675 45221
rect 47337 45216 85675 45218
rect 47337 45160 47342 45216
rect 47398 45160 47970 45216
rect 48026 45160 85614 45216
rect 85670 45160 85675 45216
rect 88185 45218 88251 45221
rect 89200 45218 90000 45248
rect 88185 45216 90000 45218
rect 47337 45158 85675 45160
rect 47337 45155 47403 45158
rect 47965 45155 48031 45158
rect 85609 45155 85675 45158
rect 87278 45184 87594 45185
rect 6686 45119 7002 45120
rect 87278 45120 87284 45184
rect 87348 45120 87364 45184
rect 87428 45120 87444 45184
rect 87508 45120 87524 45184
rect 87588 45120 87594 45184
rect 88185 45160 88190 45216
rect 88246 45160 90000 45216
rect 88185 45158 90000 45160
rect 88185 45155 88251 45158
rect 89200 45128 90000 45158
rect 87278 45119 87594 45120
rect 87173 44810 87239 44813
rect 85198 44808 87239 44810
rect 85198 44752 87178 44808
rect 87234 44752 87239 44808
rect 85198 44750 87239 44752
rect 7133 44674 7199 44677
rect 85198 44674 85258 44750
rect 87173 44747 87239 44750
rect 7133 44672 10156 44674
rect 5950 44640 6266 44641
rect 5950 44576 5956 44640
rect 6020 44576 6036 44640
rect 6100 44576 6116 44640
rect 6180 44576 6196 44640
rect 6260 44576 6266 44640
rect 7133 44616 7138 44672
rect 7194 44616 10156 44672
rect 7133 44614 10156 44616
rect 45668 44614 47508 44674
rect 83020 44614 85258 44674
rect 86542 44640 86858 44641
rect 7133 44611 7199 44614
rect 5950 44575 6266 44576
rect 86542 44576 86548 44640
rect 86612 44576 86628 44640
rect 86692 44576 86708 44640
rect 86772 44576 86788 44640
rect 86852 44576 86858 44640
rect 86542 44575 86858 44576
rect 1600 44538 2400 44568
rect 2901 44538 2967 44541
rect 1600 44536 2967 44538
rect 1600 44480 2906 44536
rect 2962 44480 2967 44536
rect 1600 44478 2967 44480
rect 1600 44448 2400 44478
rect 2901 44475 2967 44478
rect 88277 44538 88343 44541
rect 89200 44538 90000 44568
rect 88277 44536 90000 44538
rect 88277 44480 88282 44536
rect 88338 44480 90000 44536
rect 88277 44478 90000 44480
rect 88277 44475 88343 44478
rect 89200 44448 90000 44478
rect 6686 44096 7002 44097
rect 6686 44032 6692 44096
rect 6756 44032 6772 44096
rect 6836 44032 6852 44096
rect 6916 44032 6932 44096
rect 6996 44032 7002 44096
rect 6686 44031 7002 44032
rect 87278 44096 87594 44097
rect 87278 44032 87284 44096
rect 87348 44032 87364 44096
rect 87428 44032 87444 44096
rect 87508 44032 87524 44096
rect 87588 44032 87594 44096
rect 87278 44031 87594 44032
rect 1600 43858 2400 43888
rect 2717 43858 2783 43861
rect 1600 43856 2783 43858
rect 1600 43800 2722 43856
rect 2778 43800 2783 43856
rect 1600 43798 2783 43800
rect 1600 43768 2400 43798
rect 2717 43795 2783 43798
rect 88277 43858 88343 43861
rect 89200 43858 90000 43888
rect 88277 43856 90000 43858
rect 88277 43800 88282 43856
rect 88338 43800 90000 43856
rect 88277 43798 90000 43800
rect 88277 43795 88343 43798
rect 89200 43768 90000 43798
rect 8145 43586 8211 43589
rect 85793 43586 85859 43589
rect 8145 43584 10156 43586
rect 5950 43552 6266 43553
rect 5950 43488 5956 43552
rect 6020 43488 6036 43552
rect 6100 43488 6116 43552
rect 6180 43488 6196 43552
rect 6260 43488 6266 43552
rect 8145 43528 8150 43584
rect 8206 43528 10156 43584
rect 46144 43554 47508 43586
rect 83542 43584 85859 43586
rect 83542 43554 85798 43584
rect 8145 43526 10156 43528
rect 45668 43526 47508 43554
rect 83020 43528 85798 43554
rect 85854 43528 85859 43584
rect 83020 43526 85859 43528
rect 8145 43523 8211 43526
rect 45668 43494 46204 43526
rect 83020 43494 83602 43526
rect 85793 43523 85859 43526
rect 86542 43552 86858 43553
rect 5950 43487 6266 43488
rect 86542 43488 86548 43552
rect 86612 43488 86628 43552
rect 86692 43488 86708 43552
rect 86772 43488 86788 43552
rect 86852 43488 86858 43552
rect 86542 43487 86858 43488
rect 6686 43008 7002 43009
rect 6686 42944 6692 43008
rect 6756 42944 6772 43008
rect 6836 42944 6852 43008
rect 6916 42944 6932 43008
rect 6996 42944 7002 43008
rect 6686 42943 7002 42944
rect 87278 43008 87594 43009
rect 87278 42944 87284 43008
rect 87348 42944 87364 43008
rect 87428 42944 87444 43008
rect 87508 42944 87524 43008
rect 87588 42944 87594 43008
rect 87278 42943 87594 42944
rect 1600 42498 2400 42528
rect 2901 42498 2967 42501
rect 1600 42496 2967 42498
rect 1600 42440 2906 42496
rect 2962 42440 2967 42496
rect 7133 42498 7199 42501
rect 86345 42498 86411 42501
rect 7133 42496 10156 42498
rect 1600 42438 2967 42440
rect 1600 42408 2400 42438
rect 2901 42435 2967 42438
rect 5950 42464 6266 42465
rect 5950 42400 5956 42464
rect 6020 42400 6036 42464
rect 6100 42400 6116 42464
rect 6180 42400 6196 42464
rect 6260 42400 6266 42464
rect 7133 42440 7138 42496
rect 7194 42440 10156 42496
rect 46144 42466 47508 42498
rect 83542 42496 86411 42498
rect 83542 42466 86350 42496
rect 7133 42438 10156 42440
rect 45668 42438 47508 42466
rect 83020 42440 86350 42466
rect 86406 42440 86411 42496
rect 88277 42498 88343 42501
rect 89200 42498 90000 42528
rect 88277 42496 90000 42498
rect 83020 42438 86411 42440
rect 7133 42435 7199 42438
rect 45668 42406 46204 42438
rect 83020 42406 83602 42438
rect 86345 42435 86411 42438
rect 86542 42464 86858 42465
rect 5950 42399 6266 42400
rect 86542 42400 86548 42464
rect 86612 42400 86628 42464
rect 86692 42400 86708 42464
rect 86772 42400 86788 42464
rect 86852 42400 86858 42464
rect 88277 42440 88282 42496
rect 88338 42440 90000 42496
rect 88277 42438 90000 42440
rect 88277 42435 88343 42438
rect 89200 42408 90000 42438
rect 86542 42399 86858 42400
rect 6686 41920 7002 41921
rect 6686 41856 6692 41920
rect 6756 41856 6772 41920
rect 6836 41856 6852 41920
rect 6916 41856 6932 41920
rect 6996 41856 7002 41920
rect 6686 41855 7002 41856
rect 87278 41920 87594 41921
rect 87278 41856 87284 41920
rect 87348 41856 87364 41920
rect 87428 41856 87444 41920
rect 87508 41856 87524 41920
rect 87588 41856 87594 41920
rect 87278 41855 87594 41856
rect 5661 41546 5727 41549
rect 87173 41546 87239 41549
rect 5661 41544 10186 41546
rect 5661 41488 5666 41544
rect 5722 41488 10186 41544
rect 5661 41486 10186 41488
rect 5661 41483 5727 41486
rect 10126 41380 10186 41486
rect 85750 41544 87239 41546
rect 85750 41488 87178 41544
rect 87234 41488 87239 41544
rect 85750 41486 87239 41488
rect 85750 41410 85810 41486
rect 87173 41483 87239 41486
rect 46144 41378 47508 41410
rect 83542 41378 85810 41410
rect 5950 41376 6266 41377
rect 5950 41312 5956 41376
rect 6020 41312 6036 41376
rect 6100 41312 6116 41376
rect 6180 41312 6196 41376
rect 6260 41312 6266 41376
rect 45668 41350 47508 41378
rect 83020 41350 85810 41378
rect 86542 41376 86858 41377
rect 45668 41318 46204 41350
rect 83020 41318 83602 41350
rect 5950 41311 6266 41312
rect 86542 41312 86548 41376
rect 86612 41312 86628 41376
rect 86692 41312 86708 41376
rect 86772 41312 86788 41376
rect 86852 41312 86858 41376
rect 86542 41311 86858 41312
rect 1600 41138 2400 41168
rect 4373 41138 4439 41141
rect 1600 41136 4439 41138
rect 1600 41080 4378 41136
rect 4434 41080 4439 41136
rect 1600 41078 4439 41080
rect 1600 41048 2400 41078
rect 4373 41075 4439 41078
rect 88277 41138 88343 41141
rect 89200 41138 90000 41168
rect 88277 41136 90000 41138
rect 88277 41080 88282 41136
rect 88338 41080 90000 41136
rect 88277 41078 90000 41080
rect 88277 41075 88343 41078
rect 89200 41048 90000 41078
rect 6686 40832 7002 40833
rect 6686 40768 6692 40832
rect 6756 40768 6772 40832
rect 6836 40768 6852 40832
rect 6916 40768 6932 40832
rect 6996 40768 7002 40832
rect 6686 40767 7002 40768
rect 87278 40832 87594 40833
rect 87278 40768 87284 40832
rect 87348 40768 87364 40832
rect 87428 40768 87444 40832
rect 87508 40768 87524 40832
rect 87588 40768 87594 40832
rect 87278 40767 87594 40768
rect 1600 40458 2400 40488
rect 2901 40458 2967 40461
rect 87909 40458 87975 40461
rect 1600 40456 2967 40458
rect 1600 40400 2906 40456
rect 2962 40400 2967 40456
rect 1600 40398 2967 40400
rect 1600 40368 2400 40398
rect 2901 40395 2967 40398
rect 85750 40456 87975 40458
rect 85750 40400 87914 40456
rect 87970 40400 87975 40456
rect 85750 40398 87975 40400
rect 7133 40322 7199 40325
rect 85750 40322 85810 40398
rect 87909 40395 87975 40398
rect 88277 40458 88343 40461
rect 89200 40458 90000 40488
rect 88277 40456 90000 40458
rect 88277 40400 88282 40456
rect 88338 40400 90000 40456
rect 88277 40398 90000 40400
rect 88277 40395 88343 40398
rect 89200 40368 90000 40398
rect 7133 40320 10156 40322
rect 5950 40288 6266 40289
rect 5950 40224 5956 40288
rect 6020 40224 6036 40288
rect 6100 40224 6116 40288
rect 6180 40224 6196 40288
rect 6260 40224 6266 40288
rect 7133 40264 7138 40320
rect 7194 40264 10156 40320
rect 46144 40290 47508 40322
rect 83542 40290 85810 40322
rect 7133 40262 10156 40264
rect 45668 40262 47508 40290
rect 83020 40262 85810 40290
rect 86542 40288 86858 40289
rect 7133 40259 7199 40262
rect 45668 40230 46204 40262
rect 83020 40230 83602 40262
rect 5950 40223 6266 40224
rect 86542 40224 86548 40288
rect 86612 40224 86628 40288
rect 86692 40224 86708 40288
rect 86772 40224 86788 40288
rect 86852 40224 86858 40288
rect 86542 40223 86858 40224
rect 6686 39744 7002 39745
rect 6686 39680 6692 39744
rect 6756 39680 6772 39744
rect 6836 39680 6852 39744
rect 6916 39680 6932 39744
rect 6996 39680 7002 39744
rect 6686 39679 7002 39680
rect 87278 39744 87594 39745
rect 87278 39680 87284 39744
rect 87348 39680 87364 39744
rect 87428 39680 87444 39744
rect 87508 39680 87524 39744
rect 87588 39680 87594 39744
rect 87278 39679 87594 39680
rect 87173 39370 87239 39373
rect 85750 39368 87239 39370
rect 85750 39312 87178 39368
rect 87234 39312 87239 39368
rect 85750 39310 87239 39312
rect 7133 39234 7199 39237
rect 85750 39234 85810 39310
rect 87173 39307 87239 39310
rect 7133 39232 10156 39234
rect 5950 39200 6266 39201
rect 5950 39136 5956 39200
rect 6020 39136 6036 39200
rect 6100 39136 6116 39200
rect 6180 39136 6196 39200
rect 6260 39136 6266 39200
rect 7133 39176 7138 39232
rect 7194 39176 10156 39232
rect 46144 39202 47508 39234
rect 83542 39202 85810 39234
rect 7133 39174 10156 39176
rect 45668 39174 47508 39202
rect 83020 39174 85810 39202
rect 86542 39200 86858 39201
rect 7133 39171 7199 39174
rect 45668 39142 46204 39174
rect 83020 39142 83602 39174
rect 5950 39135 6266 39136
rect 86542 39136 86548 39200
rect 86612 39136 86628 39200
rect 86692 39136 86708 39200
rect 86772 39136 86788 39200
rect 86852 39136 86858 39200
rect 86542 39135 86858 39136
rect 1600 39098 2400 39128
rect 2901 39098 2967 39101
rect 1600 39096 2967 39098
rect 1600 39040 2906 39096
rect 2962 39040 2967 39096
rect 1600 39038 2967 39040
rect 1600 39008 2400 39038
rect 2901 39035 2967 39038
rect 88277 39098 88343 39101
rect 89200 39098 90000 39128
rect 88277 39096 90000 39098
rect 88277 39040 88282 39096
rect 88338 39040 90000 39096
rect 88277 39038 90000 39040
rect 88277 39035 88343 39038
rect 89200 39008 90000 39038
rect 6686 38656 7002 38657
rect 6686 38592 6692 38656
rect 6756 38592 6772 38656
rect 6836 38592 6852 38656
rect 6916 38592 6932 38656
rect 6996 38592 7002 38656
rect 6686 38591 7002 38592
rect 87278 38656 87594 38657
rect 87278 38592 87284 38656
rect 87348 38592 87364 38656
rect 87428 38592 87444 38656
rect 87508 38592 87524 38656
rect 87588 38592 87594 38656
rect 87278 38591 87594 38592
rect 1600 38418 2400 38448
rect 4373 38418 4439 38421
rect 1600 38416 4439 38418
rect 1600 38360 4378 38416
rect 4434 38360 4439 38416
rect 1600 38358 4439 38360
rect 1600 38328 2400 38358
rect 4373 38355 4439 38358
rect 88277 38418 88343 38421
rect 89200 38418 90000 38448
rect 88277 38416 90000 38418
rect 88277 38360 88282 38416
rect 88338 38360 90000 38416
rect 88277 38358 90000 38360
rect 88277 38355 88343 38358
rect 89200 38328 90000 38358
rect 7777 38146 7843 38149
rect 84413 38146 84479 38149
rect 7777 38144 10156 38146
rect 5950 38112 6266 38113
rect 5950 38048 5956 38112
rect 6020 38048 6036 38112
rect 6100 38048 6116 38112
rect 6180 38048 6196 38112
rect 6260 38048 6266 38112
rect 7777 38088 7782 38144
rect 7838 38088 10156 38144
rect 46144 38114 47508 38146
rect 83542 38144 84479 38146
rect 83542 38114 84418 38144
rect 7777 38086 10156 38088
rect 45668 38086 47508 38114
rect 83020 38088 84418 38114
rect 84474 38088 84479 38144
rect 83020 38086 84479 38088
rect 7777 38083 7843 38086
rect 45668 38054 46204 38086
rect 83020 38054 83602 38086
rect 84413 38083 84479 38086
rect 86542 38112 86858 38113
rect 5950 38047 6266 38048
rect 86542 38048 86548 38112
rect 86612 38048 86628 38112
rect 86692 38048 86708 38112
rect 86772 38048 86788 38112
rect 86852 38048 86858 38112
rect 86542 38047 86858 38048
rect 6686 37568 7002 37569
rect 6686 37504 6692 37568
rect 6756 37504 6772 37568
rect 6836 37504 6852 37568
rect 6916 37504 6932 37568
rect 6996 37504 7002 37568
rect 6686 37503 7002 37504
rect 87278 37568 87594 37569
rect 87278 37504 87284 37568
rect 87348 37504 87364 37568
rect 87428 37504 87444 37568
rect 87508 37504 87524 37568
rect 87588 37504 87594 37568
rect 87278 37503 87594 37504
rect 1600 37058 2400 37088
rect 2901 37058 2967 37061
rect 1600 37056 2967 37058
rect 1600 37000 2906 37056
rect 2962 37000 2967 37056
rect 7225 37058 7291 37061
rect 86345 37058 86411 37061
rect 7225 37056 10156 37058
rect 1600 36998 2967 37000
rect 1600 36968 2400 36998
rect 2901 36995 2967 36998
rect 5950 37024 6266 37025
rect 5950 36960 5956 37024
rect 6020 36960 6036 37024
rect 6100 36960 6116 37024
rect 6180 36960 6196 37024
rect 6260 36960 6266 37024
rect 7225 37000 7230 37056
rect 7286 37000 10156 37056
rect 46006 37026 47508 37058
rect 83542 37056 86411 37058
rect 83542 37026 86350 37056
rect 7225 36998 10156 37000
rect 45668 36998 47508 37026
rect 83020 37000 86350 37026
rect 86406 37000 86411 37056
rect 88277 37058 88343 37061
rect 89200 37058 90000 37088
rect 88277 37056 90000 37058
rect 83020 36998 86411 37000
rect 7225 36995 7291 36998
rect 45668 36966 46066 36998
rect 83020 36966 83602 36998
rect 86345 36995 86411 36998
rect 86542 37024 86858 37025
rect 5950 36959 6266 36960
rect 86542 36960 86548 37024
rect 86612 36960 86628 37024
rect 86692 36960 86708 37024
rect 86772 36960 86788 37024
rect 86852 36960 86858 37024
rect 88277 37000 88282 37056
rect 88338 37000 90000 37056
rect 88277 36998 90000 37000
rect 88277 36995 88343 36998
rect 89200 36968 90000 36998
rect 86542 36959 86858 36960
rect 6686 36480 7002 36481
rect 6686 36416 6692 36480
rect 6756 36416 6772 36480
rect 6836 36416 6852 36480
rect 6916 36416 6932 36480
rect 6996 36416 7002 36480
rect 6686 36415 7002 36416
rect 87278 36480 87594 36481
rect 87278 36416 87284 36480
rect 87348 36416 87364 36480
rect 87428 36416 87444 36480
rect 87508 36416 87524 36480
rect 87588 36416 87594 36480
rect 87278 36415 87594 36416
rect 5661 36106 5727 36109
rect 5661 36104 10186 36106
rect 5661 36048 5666 36104
rect 5722 36048 10186 36104
rect 5661 36046 10186 36048
rect 5661 36043 5727 36046
rect 10126 35940 10186 36046
rect 84413 35970 84479 35973
rect 46006 35938 47508 35970
rect 83542 35968 84479 35970
rect 83542 35938 84418 35968
rect 5950 35936 6266 35937
rect 5950 35872 5956 35936
rect 6020 35872 6036 35936
rect 6100 35872 6116 35936
rect 6180 35872 6196 35936
rect 6260 35872 6266 35936
rect 45668 35910 47508 35938
rect 83020 35912 84418 35938
rect 84474 35912 84479 35968
rect 83020 35910 84479 35912
rect 45668 35878 46066 35910
rect 83020 35878 83602 35910
rect 84413 35907 84479 35910
rect 86542 35936 86858 35937
rect 5950 35871 6266 35872
rect 86542 35872 86548 35936
rect 86612 35872 86628 35936
rect 86692 35872 86708 35936
rect 86772 35872 86788 35936
rect 86852 35872 86858 35936
rect 86542 35871 86858 35872
rect 1600 35698 2400 35728
rect 4373 35698 4439 35701
rect 1600 35696 4439 35698
rect 1600 35640 4378 35696
rect 4434 35640 4439 35696
rect 1600 35638 4439 35640
rect 1600 35608 2400 35638
rect 4373 35635 4439 35638
rect 88553 35698 88619 35701
rect 89200 35698 90000 35728
rect 88553 35696 90000 35698
rect 88553 35640 88558 35696
rect 88614 35640 90000 35696
rect 88553 35638 90000 35640
rect 88553 35635 88619 35638
rect 89200 35608 90000 35638
rect 6686 35392 7002 35393
rect 6686 35328 6692 35392
rect 6756 35328 6772 35392
rect 6836 35328 6852 35392
rect 6916 35328 6932 35392
rect 6996 35328 7002 35392
rect 6686 35327 7002 35328
rect 87278 35392 87594 35393
rect 87278 35328 87284 35392
rect 87348 35328 87364 35392
rect 87428 35328 87444 35392
rect 87508 35328 87524 35392
rect 87588 35328 87594 35392
rect 87278 35327 87594 35328
rect 1600 35018 2400 35048
rect 2901 35018 2967 35021
rect 1600 35016 2967 35018
rect 1600 34960 2906 35016
rect 2962 34960 2967 35016
rect 1600 34958 2967 34960
rect 1600 34928 2400 34958
rect 2901 34955 2967 34958
rect 88277 35018 88343 35021
rect 89200 35018 90000 35048
rect 88277 35016 90000 35018
rect 88277 34960 88282 35016
rect 88338 34960 90000 35016
rect 88277 34958 90000 34960
rect 88277 34955 88343 34958
rect 89200 34928 90000 34958
rect 7225 34882 7291 34885
rect 86345 34882 86411 34885
rect 7225 34880 10156 34882
rect 5950 34848 6266 34849
rect 5950 34784 5956 34848
rect 6020 34784 6036 34848
rect 6100 34784 6116 34848
rect 6180 34784 6196 34848
rect 6260 34784 6266 34848
rect 7225 34824 7230 34880
rect 7286 34824 10156 34880
rect 46006 34850 47508 34882
rect 83542 34880 86411 34882
rect 83542 34850 86350 34880
rect 7225 34822 10156 34824
rect 45668 34822 47508 34850
rect 83020 34824 86350 34850
rect 86406 34824 86411 34880
rect 83020 34822 86411 34824
rect 7225 34819 7291 34822
rect 45668 34790 46066 34822
rect 83020 34790 83602 34822
rect 86345 34819 86411 34822
rect 86542 34848 86858 34849
rect 5950 34783 6266 34784
rect 86542 34784 86548 34848
rect 86612 34784 86628 34848
rect 86692 34784 86708 34848
rect 86772 34784 86788 34848
rect 86852 34784 86858 34848
rect 86542 34783 86858 34784
rect 6686 34304 7002 34305
rect 6686 34240 6692 34304
rect 6756 34240 6772 34304
rect 6836 34240 6852 34304
rect 6916 34240 6932 34304
rect 6996 34240 7002 34304
rect 6686 34239 7002 34240
rect 87278 34304 87594 34305
rect 87278 34240 87284 34304
rect 87348 34240 87364 34304
rect 87428 34240 87444 34304
rect 87508 34240 87524 34304
rect 87588 34240 87594 34304
rect 87278 34239 87594 34240
rect 7225 33794 7291 33797
rect 86345 33794 86411 33797
rect 7225 33792 10156 33794
rect 5950 33760 6266 33761
rect 5950 33696 5956 33760
rect 6020 33696 6036 33760
rect 6100 33696 6116 33760
rect 6180 33696 6196 33760
rect 6260 33696 6266 33760
rect 7225 33736 7230 33792
rect 7286 33736 10156 33792
rect 46006 33762 47508 33794
rect 83542 33792 86411 33794
rect 83542 33762 86350 33792
rect 7225 33734 10156 33736
rect 45668 33734 47508 33762
rect 83020 33736 86350 33762
rect 86406 33736 86411 33792
rect 83020 33734 86411 33736
rect 7225 33731 7291 33734
rect 45668 33702 46066 33734
rect 83020 33702 83602 33734
rect 86345 33731 86411 33734
rect 86542 33760 86858 33761
rect 5950 33695 6266 33696
rect 86542 33696 86548 33760
rect 86612 33696 86628 33760
rect 86692 33696 86708 33760
rect 86772 33696 86788 33760
rect 86852 33696 86858 33760
rect 86542 33695 86858 33696
rect 1600 33658 2400 33688
rect 2901 33658 2967 33661
rect 1600 33656 2967 33658
rect 1600 33600 2906 33656
rect 2962 33600 2967 33656
rect 1600 33598 2967 33600
rect 1600 33568 2400 33598
rect 2901 33595 2967 33598
rect 88277 33658 88343 33661
rect 89200 33658 90000 33688
rect 88277 33656 90000 33658
rect 88277 33600 88282 33656
rect 88338 33600 90000 33656
rect 88277 33598 90000 33600
rect 88277 33595 88343 33598
rect 89200 33568 90000 33598
rect 6686 33216 7002 33217
rect 6686 33152 6692 33216
rect 6756 33152 6772 33216
rect 6836 33152 6852 33216
rect 6916 33152 6932 33216
rect 6996 33152 7002 33216
rect 6686 33151 7002 33152
rect 87278 33216 87594 33217
rect 87278 33152 87284 33216
rect 87348 33152 87364 33216
rect 87428 33152 87444 33216
rect 87508 33152 87524 33216
rect 87588 33152 87594 33216
rect 87278 33151 87594 33152
rect 1600 32978 2400 33008
rect 4373 32978 4439 32981
rect 1600 32976 4439 32978
rect 1600 32920 4378 32976
rect 4434 32920 4439 32976
rect 1600 32918 4439 32920
rect 1600 32888 2400 32918
rect 4373 32915 4439 32918
rect 5661 32978 5727 32981
rect 88553 32978 88619 32981
rect 89200 32978 90000 33008
rect 5661 32976 10186 32978
rect 5661 32920 5666 32976
rect 5722 32920 10186 32976
rect 5661 32918 10186 32920
rect 5661 32915 5727 32918
rect 10126 32676 10186 32918
rect 88553 32976 90000 32978
rect 88553 32920 88558 32976
rect 88614 32920 90000 32976
rect 88553 32918 90000 32920
rect 88553 32915 88619 32918
rect 89200 32888 90000 32918
rect 84413 32706 84479 32709
rect 46006 32674 47508 32706
rect 83542 32704 84479 32706
rect 83542 32674 84418 32704
rect 5950 32672 6266 32673
rect 5950 32608 5956 32672
rect 6020 32608 6036 32672
rect 6100 32608 6116 32672
rect 6180 32608 6196 32672
rect 6260 32608 6266 32672
rect 45668 32646 47508 32674
rect 83020 32648 84418 32674
rect 84474 32648 84479 32704
rect 83020 32646 84479 32648
rect 45668 32614 46066 32646
rect 83020 32614 83602 32646
rect 84413 32643 84479 32646
rect 86542 32672 86858 32673
rect 5950 32607 6266 32608
rect 86542 32608 86548 32672
rect 86612 32608 86628 32672
rect 86692 32608 86708 32672
rect 86772 32608 86788 32672
rect 86852 32608 86858 32672
rect 86542 32607 86858 32608
rect 6686 32128 7002 32129
rect 6686 32064 6692 32128
rect 6756 32064 6772 32128
rect 6836 32064 6852 32128
rect 6916 32064 6932 32128
rect 6996 32064 7002 32128
rect 6686 32063 7002 32064
rect 87278 32128 87594 32129
rect 87278 32064 87284 32128
rect 87348 32064 87364 32128
rect 87428 32064 87444 32128
rect 87508 32064 87524 32128
rect 87588 32064 87594 32128
rect 87278 32063 87594 32064
rect 1600 31618 2400 31648
rect 2901 31618 2967 31621
rect 1600 31616 2967 31618
rect 1600 31560 2906 31616
rect 2962 31560 2967 31616
rect 7225 31618 7291 31621
rect 86345 31618 86411 31621
rect 7225 31616 10156 31618
rect 1600 31558 2967 31560
rect 1600 31528 2400 31558
rect 2901 31555 2967 31558
rect 5950 31584 6266 31585
rect 5950 31520 5956 31584
rect 6020 31520 6036 31584
rect 6100 31520 6116 31584
rect 6180 31520 6196 31584
rect 6260 31520 6266 31584
rect 7225 31560 7230 31616
rect 7286 31560 10156 31616
rect 46006 31586 47508 31618
rect 83542 31616 86411 31618
rect 83542 31586 86350 31616
rect 7225 31558 10156 31560
rect 45668 31558 47508 31586
rect 83020 31560 86350 31586
rect 86406 31560 86411 31616
rect 88277 31618 88343 31621
rect 89200 31618 90000 31648
rect 88277 31616 90000 31618
rect 83020 31558 86411 31560
rect 7225 31555 7291 31558
rect 45668 31526 46066 31558
rect 83020 31526 83602 31558
rect 86345 31555 86411 31558
rect 86542 31584 86858 31585
rect 5950 31519 6266 31520
rect 86542 31520 86548 31584
rect 86612 31520 86628 31584
rect 86692 31520 86708 31584
rect 86772 31520 86788 31584
rect 86852 31520 86858 31584
rect 88277 31560 88282 31616
rect 88338 31560 90000 31616
rect 88277 31558 90000 31560
rect 88277 31555 88343 31558
rect 89200 31528 90000 31558
rect 86542 31519 86858 31520
rect 6686 31040 7002 31041
rect 6686 30976 6692 31040
rect 6756 30976 6772 31040
rect 6836 30976 6852 31040
rect 6916 30976 6932 31040
rect 6996 30976 7002 31040
rect 6686 30975 7002 30976
rect 87278 31040 87594 31041
rect 87278 30976 87284 31040
rect 87348 30976 87364 31040
rect 87428 30976 87444 31040
rect 87508 30976 87524 31040
rect 87588 30976 87594 31040
rect 87278 30975 87594 30976
rect 84413 30530 84479 30533
rect 46006 30498 47508 30530
rect 83542 30528 84479 30530
rect 83542 30498 84418 30528
rect 5950 30496 6266 30497
rect 5950 30432 5956 30496
rect 6020 30432 6036 30496
rect 6100 30432 6116 30496
rect 6180 30432 6196 30496
rect 6260 30432 6266 30496
rect 45668 30470 47508 30498
rect 83020 30472 84418 30498
rect 84474 30472 84479 30528
rect 83020 30470 84479 30472
rect 45668 30438 46066 30470
rect 83020 30438 83602 30470
rect 84413 30467 84479 30470
rect 86542 30496 86858 30497
rect 86542 30432 86548 30496
rect 86612 30432 86628 30496
rect 86692 30432 86708 30496
rect 86772 30432 86788 30496
rect 86852 30432 86858 30496
rect 5950 30431 6266 30432
rect 1600 30258 2400 30288
rect 4373 30258 4439 30261
rect 1600 30256 4439 30258
rect 1600 30200 4378 30256
rect 4434 30200 4439 30256
rect 1600 30198 4439 30200
rect 1600 30168 2400 30198
rect 4373 30195 4439 30198
rect 5661 30258 5727 30261
rect 10126 30258 10186 30432
rect 86542 30431 86858 30432
rect 5661 30256 10186 30258
rect 5661 30200 5666 30256
rect 5722 30200 10186 30256
rect 5661 30198 10186 30200
rect 88553 30258 88619 30261
rect 89200 30258 90000 30288
rect 88553 30256 90000 30258
rect 88553 30200 88558 30256
rect 88614 30200 90000 30256
rect 88553 30198 90000 30200
rect 5661 30195 5727 30198
rect 88553 30195 88619 30198
rect 89200 30168 90000 30198
rect 6686 29952 7002 29953
rect 6686 29888 6692 29952
rect 6756 29888 6772 29952
rect 6836 29888 6852 29952
rect 6916 29888 6932 29952
rect 6996 29888 7002 29952
rect 6686 29887 7002 29888
rect 87278 29952 87594 29953
rect 87278 29888 87284 29952
rect 87348 29888 87364 29952
rect 87428 29888 87444 29952
rect 87508 29888 87524 29952
rect 87588 29888 87594 29952
rect 87278 29887 87594 29888
rect 1600 29578 2400 29608
rect 2901 29578 2967 29581
rect 1600 29576 2967 29578
rect 1600 29520 2906 29576
rect 2962 29520 2967 29576
rect 1600 29518 2967 29520
rect 1600 29488 2400 29518
rect 2901 29515 2967 29518
rect 88277 29578 88343 29581
rect 89200 29578 90000 29608
rect 88277 29576 90000 29578
rect 88277 29520 88282 29576
rect 88338 29520 90000 29576
rect 88277 29518 90000 29520
rect 88277 29515 88343 29518
rect 89200 29488 90000 29518
rect 7225 29442 7291 29445
rect 86345 29442 86411 29445
rect 7225 29440 10156 29442
rect 5950 29408 6266 29409
rect 5950 29344 5956 29408
rect 6020 29344 6036 29408
rect 6100 29344 6116 29408
rect 6180 29344 6196 29408
rect 6260 29344 6266 29408
rect 7225 29384 7230 29440
rect 7286 29384 10156 29440
rect 46006 29410 47508 29442
rect 83542 29440 86411 29442
rect 83542 29410 86350 29440
rect 7225 29382 10156 29384
rect 45668 29382 47508 29410
rect 83020 29384 86350 29410
rect 86406 29384 86411 29440
rect 83020 29382 86411 29384
rect 7225 29379 7291 29382
rect 45668 29350 46066 29382
rect 83020 29350 83602 29382
rect 86345 29379 86411 29382
rect 86542 29408 86858 29409
rect 5950 29343 6266 29344
rect 86542 29344 86548 29408
rect 86612 29344 86628 29408
rect 86692 29344 86708 29408
rect 86772 29344 86788 29408
rect 86852 29344 86858 29408
rect 86542 29343 86858 29344
rect 6686 28864 7002 28865
rect 6686 28800 6692 28864
rect 6756 28800 6772 28864
rect 6836 28800 6852 28864
rect 6916 28800 6932 28864
rect 6996 28800 7002 28864
rect 6686 28799 7002 28800
rect 87278 28864 87594 28865
rect 87278 28800 87284 28864
rect 87348 28800 87364 28864
rect 87428 28800 87444 28864
rect 87508 28800 87524 28864
rect 87588 28800 87594 28864
rect 87278 28799 87594 28800
rect 7225 28354 7291 28357
rect 86345 28354 86411 28357
rect 7225 28352 10156 28354
rect 5950 28320 6266 28321
rect 5950 28256 5956 28320
rect 6020 28256 6036 28320
rect 6100 28256 6116 28320
rect 6180 28256 6196 28320
rect 6260 28256 6266 28320
rect 7225 28296 7230 28352
rect 7286 28296 10156 28352
rect 46006 28322 47508 28354
rect 83542 28352 86411 28354
rect 83542 28322 86350 28352
rect 7225 28294 10156 28296
rect 45668 28294 47508 28322
rect 83020 28296 86350 28322
rect 86406 28296 86411 28352
rect 83020 28294 86411 28296
rect 7225 28291 7291 28294
rect 45668 28262 46066 28294
rect 83020 28262 83602 28294
rect 86345 28291 86411 28294
rect 86542 28320 86858 28321
rect 5950 28255 6266 28256
rect 86542 28256 86548 28320
rect 86612 28256 86628 28320
rect 86692 28256 86708 28320
rect 86772 28256 86788 28320
rect 86852 28256 86858 28320
rect 86542 28255 86858 28256
rect 1600 28218 2400 28248
rect 2901 28218 2967 28221
rect 1600 28216 2967 28218
rect 1600 28160 2906 28216
rect 2962 28160 2967 28216
rect 1600 28158 2967 28160
rect 1600 28128 2400 28158
rect 2901 28155 2967 28158
rect 88185 28218 88251 28221
rect 89200 28218 90000 28248
rect 88185 28216 90000 28218
rect 88185 28160 88190 28216
rect 88246 28160 90000 28216
rect 88185 28158 90000 28160
rect 88185 28155 88251 28158
rect 89200 28128 90000 28158
rect 6686 27776 7002 27777
rect 6686 27712 6692 27776
rect 6756 27712 6772 27776
rect 6836 27712 6852 27776
rect 6916 27712 6932 27776
rect 6996 27712 7002 27776
rect 6686 27711 7002 27712
rect 87278 27776 87594 27777
rect 87278 27712 87284 27776
rect 87348 27712 87364 27776
rect 87428 27712 87444 27776
rect 87508 27712 87524 27776
rect 87588 27712 87594 27776
rect 87278 27711 87594 27712
rect 1600 27538 2400 27568
rect 5109 27538 5175 27541
rect 1600 27536 5175 27538
rect 1600 27480 5114 27536
rect 5170 27480 5175 27536
rect 1600 27478 5175 27480
rect 1600 27448 2400 27478
rect 5109 27475 5175 27478
rect 5385 27538 5451 27541
rect 88921 27538 88987 27541
rect 89200 27538 90000 27568
rect 5385 27536 10186 27538
rect 5385 27480 5390 27536
rect 5446 27480 10186 27536
rect 5385 27478 10186 27480
rect 5385 27475 5451 27478
rect 10126 27236 10186 27478
rect 88921 27536 90000 27538
rect 88921 27480 88926 27536
rect 88982 27480 90000 27536
rect 88921 27478 90000 27480
rect 88921 27475 88987 27478
rect 89200 27448 90000 27478
rect 85241 27266 85307 27269
rect 46006 27234 47508 27266
rect 83542 27264 85307 27266
rect 83542 27234 85246 27264
rect 5950 27232 6266 27233
rect 5950 27168 5956 27232
rect 6020 27168 6036 27232
rect 6100 27168 6116 27232
rect 6180 27168 6196 27232
rect 6260 27168 6266 27232
rect 45668 27206 47508 27234
rect 83020 27208 85246 27234
rect 85302 27208 85307 27264
rect 83020 27206 85307 27208
rect 45668 27174 46066 27206
rect 83020 27174 83602 27206
rect 85241 27203 85307 27206
rect 86542 27232 86858 27233
rect 5950 27167 6266 27168
rect 86542 27168 86548 27232
rect 86612 27168 86628 27232
rect 86692 27168 86708 27232
rect 86772 27168 86788 27232
rect 86852 27168 86858 27232
rect 86542 27167 86858 27168
rect 6686 26688 7002 26689
rect 6686 26624 6692 26688
rect 6756 26624 6772 26688
rect 6836 26624 6852 26688
rect 6916 26624 6932 26688
rect 6996 26624 7002 26688
rect 6686 26623 7002 26624
rect 87278 26688 87594 26689
rect 87278 26624 87284 26688
rect 87348 26624 87364 26688
rect 87428 26624 87444 26688
rect 87508 26624 87524 26688
rect 87588 26624 87594 26688
rect 87278 26623 87594 26624
rect 87725 26314 87791 26317
rect 85750 26312 87791 26314
rect 85750 26256 87730 26312
rect 87786 26256 87791 26312
rect 85750 26254 87791 26256
rect 1600 26178 2400 26208
rect 2901 26178 2967 26181
rect 1600 26176 2967 26178
rect 1600 26120 2906 26176
rect 2962 26120 2967 26176
rect 7133 26178 7199 26181
rect 85750 26178 85810 26254
rect 87725 26251 87791 26254
rect 7133 26176 10156 26178
rect 1600 26118 2967 26120
rect 1600 26088 2400 26118
rect 2901 26115 2967 26118
rect 5950 26144 6266 26145
rect 5950 26080 5956 26144
rect 6020 26080 6036 26144
rect 6100 26080 6116 26144
rect 6180 26080 6196 26144
rect 6260 26080 6266 26144
rect 7133 26120 7138 26176
rect 7194 26120 10156 26176
rect 46006 26146 47508 26178
rect 83542 26146 85810 26178
rect 7133 26118 10156 26120
rect 45668 26118 47508 26146
rect 83020 26118 85810 26146
rect 88185 26178 88251 26181
rect 89200 26178 90000 26208
rect 88185 26176 90000 26178
rect 86542 26144 86858 26145
rect 7133 26115 7199 26118
rect 45668 26086 46066 26118
rect 83020 26086 83602 26118
rect 5950 26079 6266 26080
rect 86542 26080 86548 26144
rect 86612 26080 86628 26144
rect 86692 26080 86708 26144
rect 86772 26080 86788 26144
rect 86852 26080 86858 26144
rect 88185 26120 88190 26176
rect 88246 26120 90000 26176
rect 88185 26118 90000 26120
rect 88185 26115 88251 26118
rect 89200 26088 90000 26118
rect 86542 26079 86858 26080
rect 6686 25600 7002 25601
rect 6686 25536 6692 25600
rect 6756 25536 6772 25600
rect 6836 25536 6852 25600
rect 6916 25536 6932 25600
rect 6996 25536 7002 25600
rect 6686 25535 7002 25536
rect 87278 25600 87594 25601
rect 87278 25536 87284 25600
rect 87348 25536 87364 25600
rect 87428 25536 87444 25600
rect 87508 25536 87524 25600
rect 87588 25536 87594 25600
rect 87278 25535 87594 25536
rect 87725 25226 87791 25229
rect 85750 25224 87791 25226
rect 85750 25168 87730 25224
rect 87786 25168 87791 25224
rect 85750 25166 87791 25168
rect 7133 25090 7199 25093
rect 85750 25090 85810 25166
rect 87725 25163 87791 25166
rect 7133 25088 10156 25090
rect 5950 25056 6266 25057
rect 5950 24992 5956 25056
rect 6020 24992 6036 25056
rect 6100 24992 6116 25056
rect 6180 24992 6196 25056
rect 6260 24992 6266 25056
rect 7133 25032 7138 25088
rect 7194 25032 10156 25088
rect 46006 25058 47508 25090
rect 83358 25058 85810 25090
rect 7133 25030 10156 25032
rect 45668 25030 47508 25058
rect 83020 25030 85810 25058
rect 86542 25056 86858 25057
rect 7133 25027 7199 25030
rect 45668 24998 46066 25030
rect 83020 24998 83418 25030
rect 5950 24991 6266 24992
rect 86542 24992 86548 25056
rect 86612 24992 86628 25056
rect 86692 24992 86708 25056
rect 86772 24992 86788 25056
rect 86852 24992 86858 25056
rect 86542 24991 86858 24992
rect 1600 24818 2400 24848
rect 4925 24818 4991 24821
rect 1600 24816 4991 24818
rect 1600 24760 4930 24816
rect 4986 24760 4991 24816
rect 1600 24758 4991 24760
rect 1600 24728 2400 24758
rect 4925 24755 4991 24758
rect 88553 24818 88619 24821
rect 89200 24818 90000 24848
rect 88553 24816 90000 24818
rect 88553 24760 88558 24816
rect 88614 24760 90000 24816
rect 88553 24758 90000 24760
rect 88553 24755 88619 24758
rect 89200 24728 90000 24758
rect 6686 24512 7002 24513
rect 6686 24448 6692 24512
rect 6756 24448 6772 24512
rect 6836 24448 6852 24512
rect 6916 24448 6932 24512
rect 6996 24448 7002 24512
rect 6686 24447 7002 24448
rect 87278 24512 87594 24513
rect 87278 24448 87284 24512
rect 87348 24448 87364 24512
rect 87428 24448 87444 24512
rect 87508 24448 87524 24512
rect 87588 24448 87594 24512
rect 87278 24447 87594 24448
rect 1600 24138 2400 24168
rect 2901 24138 2967 24141
rect 87725 24138 87791 24141
rect 1600 24136 2967 24138
rect 1600 24080 2906 24136
rect 2962 24080 2967 24136
rect 1600 24078 2967 24080
rect 1600 24048 2400 24078
rect 2901 24075 2967 24078
rect 85750 24136 87791 24138
rect 85750 24080 87730 24136
rect 87786 24080 87791 24136
rect 85750 24078 87791 24080
rect 7133 24002 7199 24005
rect 85750 24002 85810 24078
rect 87725 24075 87791 24078
rect 88277 24138 88343 24141
rect 89200 24138 90000 24168
rect 88277 24136 90000 24138
rect 88277 24080 88282 24136
rect 88338 24080 90000 24136
rect 88277 24078 90000 24080
rect 88277 24075 88343 24078
rect 89200 24048 90000 24078
rect 7133 24000 10156 24002
rect 5950 23968 6266 23969
rect 5950 23904 5956 23968
rect 6020 23904 6036 23968
rect 6100 23904 6116 23968
rect 6180 23904 6196 23968
rect 6260 23904 6266 23968
rect 7133 23944 7138 24000
rect 7194 23944 10156 24000
rect 46006 23970 47508 24002
rect 83542 23970 85810 24002
rect 7133 23942 10156 23944
rect 45668 23942 47508 23970
rect 83020 23942 85810 23970
rect 86542 23968 86858 23969
rect 7133 23939 7199 23942
rect 45668 23910 46066 23942
rect 83020 23910 83602 23942
rect 5950 23903 6266 23904
rect 86542 23904 86548 23968
rect 86612 23904 86628 23968
rect 86692 23904 86708 23968
rect 86772 23904 86788 23968
rect 86852 23904 86858 23968
rect 86542 23903 86858 23904
rect 6686 23424 7002 23425
rect 6686 23360 6692 23424
rect 6756 23360 6772 23424
rect 6836 23360 6852 23424
rect 6916 23360 6932 23424
rect 6996 23360 7002 23424
rect 6686 23359 7002 23360
rect 87278 23424 87594 23425
rect 87278 23360 87284 23424
rect 87348 23360 87364 23424
rect 87428 23360 87444 23424
rect 87508 23360 87524 23424
rect 87588 23360 87594 23424
rect 87278 23359 87594 23360
rect 7133 22914 7199 22917
rect 86345 22914 86411 22917
rect 7133 22912 10156 22914
rect 5950 22880 6266 22881
rect 5950 22816 5956 22880
rect 6020 22816 6036 22880
rect 6100 22816 6116 22880
rect 6180 22816 6196 22880
rect 6260 22816 6266 22880
rect 7133 22856 7138 22912
rect 7194 22856 10156 22912
rect 46006 22882 47508 22914
rect 83542 22912 86411 22914
rect 83542 22882 86350 22912
rect 7133 22854 10156 22856
rect 45668 22854 47508 22882
rect 83020 22856 86350 22882
rect 86406 22856 86411 22912
rect 83020 22854 86411 22856
rect 7133 22851 7199 22854
rect 45668 22822 46066 22854
rect 83020 22822 83602 22854
rect 86345 22851 86411 22854
rect 86542 22880 86858 22881
rect 5950 22815 6266 22816
rect 86542 22816 86548 22880
rect 86612 22816 86628 22880
rect 86692 22816 86708 22880
rect 86772 22816 86788 22880
rect 86852 22816 86858 22880
rect 86542 22815 86858 22816
rect 1600 22778 2400 22808
rect 2901 22778 2967 22781
rect 1600 22776 2967 22778
rect 1600 22720 2906 22776
rect 2962 22720 2967 22776
rect 1600 22718 2967 22720
rect 1600 22688 2400 22718
rect 2901 22715 2967 22718
rect 88277 22778 88343 22781
rect 89200 22778 90000 22808
rect 88277 22776 90000 22778
rect 88277 22720 88282 22776
rect 88338 22720 90000 22776
rect 88277 22718 90000 22720
rect 88277 22715 88343 22718
rect 89200 22688 90000 22718
rect 6686 22336 7002 22337
rect 6686 22272 6692 22336
rect 6756 22272 6772 22336
rect 6836 22272 6852 22336
rect 6916 22272 6932 22336
rect 6996 22272 7002 22336
rect 6686 22271 7002 22272
rect 87278 22336 87594 22337
rect 87278 22272 87284 22336
rect 87348 22272 87364 22336
rect 87428 22272 87444 22336
rect 87508 22272 87524 22336
rect 87588 22272 87594 22336
rect 87278 22271 87594 22272
rect 1600 22098 2400 22128
rect 4925 22098 4991 22101
rect 1600 22096 4991 22098
rect 1600 22040 4930 22096
rect 4986 22040 4991 22096
rect 1600 22038 4991 22040
rect 1600 22008 2400 22038
rect 4925 22035 4991 22038
rect 88553 22098 88619 22101
rect 89200 22098 90000 22128
rect 88553 22096 90000 22098
rect 88553 22040 88558 22096
rect 88614 22040 90000 22096
rect 88553 22038 90000 22040
rect 88553 22035 88619 22038
rect 89200 22008 90000 22038
rect 9157 21826 9223 21829
rect 84413 21826 84479 21829
rect 9157 21824 10156 21826
rect 5950 21792 6266 21793
rect 5950 21728 5956 21792
rect 6020 21728 6036 21792
rect 6100 21728 6116 21792
rect 6180 21728 6196 21792
rect 6260 21728 6266 21792
rect 9157 21768 9162 21824
rect 9218 21768 10156 21824
rect 46006 21794 47508 21826
rect 83542 21824 84479 21826
rect 83542 21794 84418 21824
rect 9157 21766 10156 21768
rect 45668 21766 47508 21794
rect 83020 21768 84418 21794
rect 84474 21768 84479 21824
rect 83020 21766 84479 21768
rect 9157 21763 9223 21766
rect 45668 21734 46066 21766
rect 83020 21734 83602 21766
rect 84413 21763 84479 21766
rect 86542 21792 86858 21793
rect 5950 21727 6266 21728
rect 86542 21728 86548 21792
rect 86612 21728 86628 21792
rect 86692 21728 86708 21792
rect 86772 21728 86788 21792
rect 86852 21728 86858 21792
rect 86542 21727 86858 21728
rect 6686 21248 7002 21249
rect 6686 21184 6692 21248
rect 6756 21184 6772 21248
rect 6836 21184 6852 21248
rect 6916 21184 6932 21248
rect 6996 21184 7002 21248
rect 6686 21183 7002 21184
rect 87278 21248 87594 21249
rect 87278 21184 87284 21248
rect 87348 21184 87364 21248
rect 87428 21184 87444 21248
rect 87508 21184 87524 21248
rect 87588 21184 87594 21248
rect 87278 21183 87594 21184
rect 1600 20738 2400 20768
rect 5201 20738 5267 20741
rect 1600 20736 5267 20738
rect 1600 20680 5206 20736
rect 5262 20680 5267 20736
rect 9249 20738 9315 20741
rect 84413 20738 84479 20741
rect 9249 20736 10156 20738
rect 1600 20678 5267 20680
rect 1600 20648 2400 20678
rect 5201 20675 5267 20678
rect 5950 20704 6266 20705
rect 5950 20640 5956 20704
rect 6020 20640 6036 20704
rect 6100 20640 6116 20704
rect 6180 20640 6196 20704
rect 6260 20640 6266 20704
rect 9249 20680 9254 20736
rect 9310 20680 10156 20736
rect 46006 20706 47508 20738
rect 83542 20736 84479 20738
rect 83542 20706 84418 20736
rect 9249 20678 10156 20680
rect 45668 20678 47508 20706
rect 83020 20680 84418 20706
rect 84474 20680 84479 20736
rect 88553 20738 88619 20741
rect 89200 20738 90000 20768
rect 88553 20736 90000 20738
rect 83020 20678 84479 20680
rect 9249 20675 9315 20678
rect 45668 20646 46066 20678
rect 83020 20646 83602 20678
rect 84413 20675 84479 20678
rect 86542 20704 86858 20705
rect 5950 20639 6266 20640
rect 86542 20640 86548 20704
rect 86612 20640 86628 20704
rect 86692 20640 86708 20704
rect 86772 20640 86788 20704
rect 86852 20640 86858 20704
rect 88553 20680 88558 20736
rect 88614 20680 90000 20736
rect 88553 20678 90000 20680
rect 88553 20675 88619 20678
rect 89200 20648 90000 20678
rect 86542 20639 86858 20640
rect 6686 20160 7002 20161
rect 6686 20096 6692 20160
rect 6756 20096 6772 20160
rect 6836 20096 6852 20160
rect 6916 20096 6932 20160
rect 6996 20096 7002 20160
rect 6686 20095 7002 20096
rect 87278 20160 87594 20161
rect 87278 20096 87284 20160
rect 87348 20096 87364 20160
rect 87428 20096 87444 20160
rect 87508 20096 87524 20160
rect 87588 20096 87594 20160
rect 87278 20095 87594 20096
rect 87725 19786 87791 19789
rect 85750 19784 87791 19786
rect 85750 19728 87730 19784
rect 87786 19728 87791 19784
rect 85750 19726 87791 19728
rect 7133 19650 7199 19653
rect 85750 19650 85810 19726
rect 87725 19723 87791 19726
rect 7133 19648 10156 19650
rect 5950 19616 6266 19617
rect 5950 19552 5956 19616
rect 6020 19552 6036 19616
rect 6100 19552 6116 19616
rect 6180 19552 6196 19616
rect 6260 19552 6266 19616
rect 7133 19592 7138 19648
rect 7194 19592 10156 19648
rect 46006 19618 47508 19650
rect 83542 19618 85810 19650
rect 7133 19590 10156 19592
rect 45668 19590 47508 19618
rect 83020 19590 85810 19618
rect 86542 19616 86858 19617
rect 7133 19587 7199 19590
rect 45668 19558 46066 19590
rect 83020 19558 83602 19590
rect 5950 19551 6266 19552
rect 86542 19552 86548 19616
rect 86612 19552 86628 19616
rect 86692 19552 86708 19616
rect 86772 19552 86788 19616
rect 86852 19552 86858 19616
rect 86542 19551 86858 19552
rect 1600 19378 2400 19408
rect 4925 19378 4991 19381
rect 1600 19376 4991 19378
rect 1600 19320 4930 19376
rect 4986 19320 4991 19376
rect 1600 19318 4991 19320
rect 1600 19288 2400 19318
rect 4925 19315 4991 19318
rect 88553 19378 88619 19381
rect 89200 19378 90000 19408
rect 88553 19376 90000 19378
rect 88553 19320 88558 19376
rect 88614 19320 90000 19376
rect 88553 19318 90000 19320
rect 88553 19315 88619 19318
rect 89200 19288 90000 19318
rect 6686 19072 7002 19073
rect 6686 19008 6692 19072
rect 6756 19008 6772 19072
rect 6836 19008 6852 19072
rect 6916 19008 6932 19072
rect 6996 19008 7002 19072
rect 6686 19007 7002 19008
rect 87278 19072 87594 19073
rect 87278 19008 87284 19072
rect 87348 19008 87364 19072
rect 87428 19008 87444 19072
rect 87508 19008 87524 19072
rect 87588 19008 87594 19072
rect 87278 19007 87594 19008
rect 1600 18698 2400 18728
rect 2901 18698 2967 18701
rect 87725 18698 87791 18701
rect 1600 18696 2967 18698
rect 1600 18640 2906 18696
rect 2962 18640 2967 18696
rect 1600 18638 2967 18640
rect 1600 18608 2400 18638
rect 2901 18635 2967 18638
rect 85750 18696 87791 18698
rect 85750 18640 87730 18696
rect 87786 18640 87791 18696
rect 85750 18638 87791 18640
rect 7133 18562 7199 18565
rect 85750 18562 85810 18638
rect 87725 18635 87791 18638
rect 88277 18698 88343 18701
rect 89200 18698 90000 18728
rect 88277 18696 90000 18698
rect 88277 18640 88282 18696
rect 88338 18640 90000 18696
rect 88277 18638 90000 18640
rect 88277 18635 88343 18638
rect 89200 18608 90000 18638
rect 7133 18560 10156 18562
rect 5950 18528 6266 18529
rect 5950 18464 5956 18528
rect 6020 18464 6036 18528
rect 6100 18464 6116 18528
rect 6180 18464 6196 18528
rect 6260 18464 6266 18528
rect 7133 18504 7138 18560
rect 7194 18504 10156 18560
rect 46006 18530 47508 18562
rect 83542 18530 85810 18562
rect 7133 18502 10156 18504
rect 45668 18502 47508 18530
rect 83020 18502 85810 18530
rect 86542 18528 86858 18529
rect 7133 18499 7199 18502
rect 45668 18470 46066 18502
rect 83020 18470 83602 18502
rect 5950 18463 6266 18464
rect 86542 18464 86548 18528
rect 86612 18464 86628 18528
rect 86692 18464 86708 18528
rect 86772 18464 86788 18528
rect 86852 18464 86858 18528
rect 86542 18463 86858 18464
rect 6686 17984 7002 17985
rect 6686 17920 6692 17984
rect 6756 17920 6772 17984
rect 6836 17920 6852 17984
rect 6916 17920 6932 17984
rect 6996 17920 7002 17984
rect 6686 17919 7002 17920
rect 87278 17984 87594 17985
rect 87278 17920 87284 17984
rect 87348 17920 87364 17984
rect 87428 17920 87444 17984
rect 87508 17920 87524 17984
rect 87588 17920 87594 17984
rect 87278 17919 87594 17920
rect 7225 17474 7291 17477
rect 86345 17474 86411 17477
rect 7225 17472 10156 17474
rect 5950 17440 6266 17441
rect 5950 17376 5956 17440
rect 6020 17376 6036 17440
rect 6100 17376 6116 17440
rect 6180 17376 6196 17440
rect 6260 17376 6266 17440
rect 7225 17416 7230 17472
rect 7286 17416 10156 17472
rect 46006 17442 47508 17474
rect 83542 17472 86411 17474
rect 83542 17442 86350 17472
rect 7225 17414 10156 17416
rect 45668 17414 47508 17442
rect 83020 17416 86350 17442
rect 86406 17416 86411 17472
rect 83020 17414 86411 17416
rect 7225 17411 7291 17414
rect 45668 17382 46066 17414
rect 83020 17382 83602 17414
rect 86345 17411 86411 17414
rect 86542 17440 86858 17441
rect 5950 17375 6266 17376
rect 86542 17376 86548 17440
rect 86612 17376 86628 17440
rect 86692 17376 86708 17440
rect 86772 17376 86788 17440
rect 86852 17376 86858 17440
rect 86542 17375 86858 17376
rect 1600 17338 2400 17368
rect 2901 17338 2967 17341
rect 1600 17336 2967 17338
rect 1600 17280 2906 17336
rect 2962 17280 2967 17336
rect 1600 17278 2967 17280
rect 1600 17248 2400 17278
rect 2901 17275 2967 17278
rect 88185 17338 88251 17341
rect 89200 17338 90000 17368
rect 88185 17336 90000 17338
rect 88185 17280 88190 17336
rect 88246 17280 90000 17336
rect 88185 17278 90000 17280
rect 88185 17275 88251 17278
rect 89200 17248 90000 17278
rect 6686 16896 7002 16897
rect 6686 16832 6692 16896
rect 6756 16832 6772 16896
rect 6836 16832 6852 16896
rect 6916 16832 6932 16896
rect 6996 16832 7002 16896
rect 6686 16831 7002 16832
rect 87278 16896 87594 16897
rect 87278 16832 87284 16896
rect 87348 16832 87364 16896
rect 87428 16832 87444 16896
rect 87508 16832 87524 16896
rect 87588 16832 87594 16896
rect 87278 16831 87594 16832
rect 1600 16658 2400 16688
rect 5201 16658 5267 16661
rect 1600 16656 5267 16658
rect 1600 16600 5206 16656
rect 5262 16600 5267 16656
rect 1600 16598 5267 16600
rect 1600 16568 2400 16598
rect 5201 16595 5267 16598
rect 5385 16658 5451 16661
rect 88553 16658 88619 16661
rect 89200 16658 90000 16688
rect 5385 16656 10186 16658
rect 5385 16600 5390 16656
rect 5446 16600 10186 16656
rect 5385 16598 10186 16600
rect 5385 16595 5451 16598
rect 10126 16356 10186 16598
rect 88553 16656 90000 16658
rect 88553 16600 88558 16656
rect 88614 16600 90000 16656
rect 88553 16598 90000 16600
rect 88553 16595 88619 16598
rect 89200 16568 90000 16598
rect 88001 16522 88067 16525
rect 85750 16520 88067 16522
rect 85750 16464 88006 16520
rect 88062 16464 88067 16520
rect 85750 16462 88067 16464
rect 85750 16386 85810 16462
rect 88001 16459 88067 16462
rect 46006 16354 47508 16386
rect 83542 16354 85810 16386
rect 5950 16352 6266 16353
rect 5950 16288 5956 16352
rect 6020 16288 6036 16352
rect 6100 16288 6116 16352
rect 6180 16288 6196 16352
rect 6260 16288 6266 16352
rect 45668 16326 47508 16354
rect 83020 16326 85810 16354
rect 86542 16352 86858 16353
rect 45668 16294 46066 16326
rect 83020 16294 83602 16326
rect 5950 16287 6266 16288
rect 86542 16288 86548 16352
rect 86612 16288 86628 16352
rect 86692 16288 86708 16352
rect 86772 16288 86788 16352
rect 86852 16288 86858 16352
rect 86542 16287 86858 16288
rect 6686 15808 7002 15809
rect 6686 15744 6692 15808
rect 6756 15744 6772 15808
rect 6836 15744 6852 15808
rect 6916 15744 6932 15808
rect 6996 15744 7002 15808
rect 6686 15743 7002 15744
rect 87278 15808 87594 15809
rect 87278 15744 87284 15808
rect 87348 15744 87364 15808
rect 87428 15744 87444 15808
rect 87508 15744 87524 15808
rect 87588 15744 87594 15808
rect 87278 15743 87594 15744
rect 1600 15298 2400 15328
rect 5201 15298 5267 15301
rect 84413 15298 84479 15301
rect 1600 15296 5267 15298
rect 1600 15240 5206 15296
rect 5262 15240 5267 15296
rect 46006 15266 47508 15298
rect 83542 15296 84479 15298
rect 83542 15266 84418 15296
rect 1600 15238 5267 15240
rect 1600 15208 2400 15238
rect 5201 15235 5267 15238
rect 5950 15264 6266 15265
rect 5950 15200 5956 15264
rect 6020 15200 6036 15264
rect 6100 15200 6116 15264
rect 6180 15200 6196 15264
rect 6260 15200 6266 15264
rect 45668 15238 47508 15266
rect 83020 15240 84418 15266
rect 84474 15240 84479 15296
rect 88553 15298 88619 15301
rect 89200 15298 90000 15328
rect 88553 15296 90000 15298
rect 83020 15238 84479 15240
rect 45668 15206 46066 15238
rect 83020 15206 83602 15238
rect 84413 15235 84479 15238
rect 86542 15264 86858 15265
rect 86542 15200 86548 15264
rect 86612 15200 86628 15264
rect 86692 15200 86708 15264
rect 86772 15200 86788 15264
rect 86852 15200 86858 15264
rect 88553 15240 88558 15296
rect 88614 15240 90000 15296
rect 88553 15238 90000 15240
rect 88553 15235 88619 15238
rect 89200 15208 90000 15238
rect 5950 15199 6266 15200
rect 5661 15026 5727 15029
rect 10126 15026 10186 15200
rect 86542 15199 86858 15200
rect 5661 15024 10186 15026
rect 5661 14968 5666 15024
rect 5722 14968 10186 15024
rect 5661 14966 10186 14968
rect 5661 14963 5727 14966
rect 6686 14720 7002 14721
rect 6686 14656 6692 14720
rect 6756 14656 6772 14720
rect 6836 14656 6852 14720
rect 6916 14656 6932 14720
rect 6996 14656 7002 14720
rect 6686 14655 7002 14656
rect 87278 14720 87594 14721
rect 87278 14656 87284 14720
rect 87348 14656 87364 14720
rect 87428 14656 87444 14720
rect 87508 14656 87524 14720
rect 87588 14656 87594 14720
rect 87278 14655 87594 14656
rect 88001 14618 88067 14621
rect 89200 14618 90000 14648
rect 88001 14616 90000 14618
rect 88001 14560 88006 14616
rect 88062 14560 90000 14616
rect 88001 14558 90000 14560
rect 88001 14555 88067 14558
rect 89200 14528 90000 14558
rect 83677 14210 83743 14213
rect 83542 14208 83743 14210
rect 45957 14178 46023 14181
rect 83542 14178 83682 14208
rect 5950 14176 6266 14177
rect 5950 14112 5956 14176
rect 6020 14112 6036 14176
rect 6100 14112 6116 14176
rect 6180 14112 6196 14176
rect 6260 14112 6266 14176
rect 45668 14176 46023 14178
rect 45668 14120 45962 14176
rect 46018 14120 46023 14176
rect 45668 14118 46023 14120
rect 83020 14152 83682 14178
rect 83738 14152 83743 14208
rect 83020 14150 83743 14152
rect 83020 14118 83602 14150
rect 83677 14147 83743 14150
rect 86542 14176 86858 14177
rect 45957 14115 46023 14118
rect 5950 14111 6266 14112
rect 86542 14112 86548 14176
rect 86612 14112 86628 14176
rect 86692 14112 86708 14176
rect 86772 14112 86788 14176
rect 86852 14112 86858 14176
rect 86542 14111 86858 14112
rect 6686 13632 7002 13633
rect 6686 13568 6692 13632
rect 6756 13568 6772 13632
rect 6836 13568 6852 13632
rect 6916 13568 6932 13632
rect 6996 13568 7002 13632
rect 6686 13567 7002 13568
rect 87278 13632 87594 13633
rect 87278 13568 87284 13632
rect 87348 13568 87364 13632
rect 87428 13568 87444 13632
rect 87508 13568 87524 13632
rect 87588 13568 87594 13632
rect 87278 13567 87594 13568
rect 88185 13258 88251 13261
rect 89200 13258 90000 13288
rect 88185 13256 90000 13258
rect 88185 13200 88190 13256
rect 88246 13200 90000 13256
rect 88185 13198 90000 13200
rect 88185 13195 88251 13198
rect 89200 13168 90000 13198
rect 45865 13090 45931 13093
rect 46141 13090 46207 13093
rect 83493 13090 83559 13093
rect 5950 13088 6266 13089
rect 5950 13024 5956 13088
rect 6020 13024 6036 13088
rect 6100 13024 6116 13088
rect 6180 13024 6196 13088
rect 6260 13024 6266 13088
rect 45668 13088 46207 13090
rect 45668 13032 45870 13088
rect 45926 13032 46146 13088
rect 46202 13032 46207 13088
rect 45668 13030 46207 13032
rect 83020 13088 83559 13090
rect 83020 13032 83498 13088
rect 83554 13032 83559 13088
rect 83020 13030 83559 13032
rect 45865 13027 45931 13030
rect 46141 13027 46207 13030
rect 83493 13027 83559 13030
rect 86542 13088 86858 13089
rect 5950 13023 6266 13024
rect 86542 13024 86548 13088
rect 86612 13024 86628 13088
rect 86692 13024 86708 13088
rect 86772 13024 86788 13088
rect 86852 13024 86858 13088
rect 86542 13023 86858 13024
rect 88553 12578 88619 12581
rect 89200 12578 90000 12608
rect 88553 12576 90000 12578
rect 6686 12544 7002 12545
rect 6686 12480 6692 12544
rect 6756 12480 6772 12544
rect 6836 12480 6852 12544
rect 6916 12480 6932 12544
rect 6996 12480 7002 12544
rect 6686 12479 7002 12480
rect 87278 12544 87594 12545
rect 87278 12480 87284 12544
rect 87348 12480 87364 12544
rect 87428 12480 87444 12544
rect 87508 12480 87524 12544
rect 87588 12480 87594 12544
rect 88553 12520 88558 12576
rect 88614 12520 90000 12576
rect 88553 12518 90000 12520
rect 88553 12515 88619 12518
rect 89200 12488 90000 12518
rect 87278 12479 87594 12480
rect 46049 12002 46115 12005
rect 83493 12002 83559 12005
rect 5950 12000 6266 12001
rect 5950 11936 5956 12000
rect 6020 11936 6036 12000
rect 6100 11936 6116 12000
rect 6180 11936 6196 12000
rect 6260 11936 6266 12000
rect 45668 12000 46115 12002
rect 45668 11944 46054 12000
rect 46110 11944 46115 12000
rect 45668 11942 46115 11944
rect 83020 12000 83559 12002
rect 83020 11944 83498 12000
rect 83554 11944 83559 12000
rect 83020 11942 83559 11944
rect 46049 11939 46115 11942
rect 83493 11939 83559 11942
rect 86542 12000 86858 12001
rect 5950 11935 6266 11936
rect 86542 11936 86548 12000
rect 86612 11936 86628 12000
rect 86692 11936 86708 12000
rect 86772 11936 86788 12000
rect 86852 11936 86858 12000
rect 86542 11935 86858 11936
rect 6686 11456 7002 11457
rect 6686 11392 6692 11456
rect 6756 11392 6772 11456
rect 6836 11392 6852 11456
rect 6916 11392 6932 11456
rect 6996 11392 7002 11456
rect 6686 11391 7002 11392
rect 87278 11456 87594 11457
rect 87278 11392 87284 11456
rect 87348 11392 87364 11456
rect 87428 11392 87444 11456
rect 87508 11392 87524 11456
rect 87588 11392 87594 11456
rect 87278 11391 87594 11392
rect 46417 10946 46483 10949
rect 46190 10944 46483 10946
rect 5950 10912 6266 10913
rect 5950 10848 5956 10912
rect 6020 10848 6036 10912
rect 6100 10848 6116 10912
rect 6180 10848 6196 10912
rect 6260 10848 6266 10912
rect 46190 10888 46422 10944
rect 46478 10888 46483 10944
rect 46190 10886 46483 10888
rect 45865 10878 45931 10881
rect 46190 10878 46250 10886
rect 46417 10883 46483 10886
rect 86542 10912 86858 10913
rect 83309 10878 83375 10881
rect 5950 10847 6266 10848
rect 45668 10876 46250 10878
rect 45668 10820 45870 10876
rect 45926 10820 46250 10876
rect 45668 10818 46250 10820
rect 83020 10876 83375 10878
rect 83020 10820 83314 10876
rect 83370 10820 83375 10876
rect 86542 10848 86548 10912
rect 86612 10848 86628 10912
rect 86692 10848 86708 10912
rect 86772 10848 86788 10912
rect 86852 10848 86858 10912
rect 86542 10847 86858 10848
rect 83020 10818 83375 10820
rect 45865 10815 45931 10818
rect 83309 10815 83375 10818
rect 88369 10538 88435 10541
rect 89200 10538 90000 10568
rect 88369 10536 90000 10538
rect 88369 10480 88374 10536
rect 88430 10480 90000 10536
rect 88369 10478 90000 10480
rect 88369 10475 88435 10478
rect 89200 10448 90000 10478
rect 6686 10368 7002 10369
rect 6686 10304 6692 10368
rect 6756 10304 6772 10368
rect 6836 10304 6852 10368
rect 6916 10304 6932 10368
rect 6996 10304 7002 10368
rect 6686 10303 7002 10304
rect 87278 10368 87594 10369
rect 87278 10304 87284 10368
rect 87348 10304 87364 10368
rect 87428 10304 87444 10368
rect 87508 10304 87524 10368
rect 87588 10304 87594 10368
rect 87278 10303 87594 10304
rect 88553 9858 88619 9861
rect 89200 9858 90000 9888
rect 88553 9856 90000 9858
rect 5950 9824 6266 9825
rect 5950 9760 5956 9824
rect 6020 9760 6036 9824
rect 6100 9760 6116 9824
rect 6180 9760 6196 9824
rect 6260 9760 6266 9824
rect 5950 9759 6266 9760
rect 86542 9824 86858 9825
rect 86542 9760 86548 9824
rect 86612 9760 86628 9824
rect 86692 9760 86708 9824
rect 86772 9760 86788 9824
rect 86852 9760 86858 9824
rect 88553 9800 88558 9856
rect 88614 9800 90000 9856
rect 88553 9798 90000 9800
rect 88553 9795 88619 9798
rect 89200 9768 90000 9798
rect 86542 9759 86858 9760
rect 6686 9280 7002 9281
rect 6686 9216 6692 9280
rect 6756 9216 6772 9280
rect 6836 9216 6852 9280
rect 6916 9216 6932 9280
rect 6996 9216 7002 9280
rect 6686 9215 7002 9216
rect 87278 9280 87594 9281
rect 87278 9216 87284 9280
rect 87348 9216 87364 9280
rect 87428 9216 87444 9280
rect 87508 9216 87524 9280
rect 87588 9216 87594 9280
rect 87278 9215 87594 9216
rect 5950 8736 6266 8737
rect 5950 8672 5956 8736
rect 6020 8672 6036 8736
rect 6100 8672 6116 8736
rect 6180 8672 6196 8736
rect 6260 8672 6266 8736
rect 5950 8671 6266 8672
rect 86542 8736 86858 8737
rect 86542 8672 86548 8736
rect 86612 8672 86628 8736
rect 86692 8672 86708 8736
rect 86772 8672 86788 8736
rect 86852 8672 86858 8736
rect 86542 8671 86858 8672
rect 6686 8192 7002 8193
rect 6686 8128 6692 8192
rect 6756 8128 6772 8192
rect 6836 8128 6852 8192
rect 6916 8128 6932 8192
rect 6996 8128 7002 8192
rect 6686 8127 7002 8128
rect 87278 8192 87594 8193
rect 87278 8128 87284 8192
rect 87348 8128 87364 8192
rect 87428 8128 87444 8192
rect 87508 8128 87524 8192
rect 87588 8128 87594 8192
rect 87278 8127 87594 8128
rect 5950 7648 6266 7649
rect 5950 7584 5956 7648
rect 6020 7584 6036 7648
rect 6100 7584 6116 7648
rect 6180 7584 6196 7648
rect 6260 7584 6266 7648
rect 5950 7583 6266 7584
rect 17718 7648 18034 7649
rect 17718 7584 17724 7648
rect 17788 7584 17804 7648
rect 17868 7584 17884 7648
rect 17948 7584 17964 7648
rect 18028 7584 18034 7648
rect 17718 7583 18034 7584
rect 36118 7648 36434 7649
rect 36118 7584 36124 7648
rect 36188 7584 36204 7648
rect 36268 7584 36284 7648
rect 36348 7584 36364 7648
rect 36428 7584 36434 7648
rect 36118 7583 36434 7584
rect 54518 7648 54834 7649
rect 54518 7584 54524 7648
rect 54588 7584 54604 7648
rect 54668 7584 54684 7648
rect 54748 7584 54764 7648
rect 54828 7584 54834 7648
rect 54518 7583 54834 7584
rect 72918 7648 73234 7649
rect 72918 7584 72924 7648
rect 72988 7584 73004 7648
rect 73068 7584 73084 7648
rect 73148 7584 73164 7648
rect 73228 7584 73234 7648
rect 72918 7583 73234 7584
rect 86542 7648 86858 7649
rect 86542 7584 86548 7648
rect 86612 7584 86628 7648
rect 86692 7584 86708 7648
rect 86772 7584 86788 7648
rect 86852 7584 86858 7648
rect 86542 7583 86858 7584
rect 6686 7104 7002 7105
rect 6686 7040 6692 7104
rect 6756 7040 6772 7104
rect 6836 7040 6852 7104
rect 6916 7040 6932 7104
rect 6996 7040 7002 7104
rect 6686 7039 7002 7040
rect 18378 7104 18694 7105
rect 18378 7040 18384 7104
rect 18448 7040 18464 7104
rect 18528 7040 18544 7104
rect 18608 7040 18624 7104
rect 18688 7040 18694 7104
rect 18378 7039 18694 7040
rect 36778 7104 37094 7105
rect 36778 7040 36784 7104
rect 36848 7040 36864 7104
rect 36928 7040 36944 7104
rect 37008 7040 37024 7104
rect 37088 7040 37094 7104
rect 36778 7039 37094 7040
rect 55178 7104 55494 7105
rect 55178 7040 55184 7104
rect 55248 7040 55264 7104
rect 55328 7040 55344 7104
rect 55408 7040 55424 7104
rect 55488 7040 55494 7104
rect 55178 7039 55494 7040
rect 73578 7104 73894 7105
rect 73578 7040 73584 7104
rect 73648 7040 73664 7104
rect 73728 7040 73744 7104
rect 73808 7040 73824 7104
rect 73888 7040 73894 7104
rect 73578 7039 73894 7040
rect 87278 7104 87594 7105
rect 87278 7040 87284 7104
rect 87348 7040 87364 7104
rect 87428 7040 87444 7104
rect 87508 7040 87524 7104
rect 87588 7040 87594 7104
rect 87278 7039 87594 7040
rect 17718 6560 18034 6561
rect 17718 6496 17724 6560
rect 17788 6496 17804 6560
rect 17868 6496 17884 6560
rect 17948 6496 17964 6560
rect 18028 6496 18034 6560
rect 17718 6495 18034 6496
rect 36118 6560 36434 6561
rect 36118 6496 36124 6560
rect 36188 6496 36204 6560
rect 36268 6496 36284 6560
rect 36348 6496 36364 6560
rect 36428 6496 36434 6560
rect 36118 6495 36434 6496
rect 54518 6560 54834 6561
rect 54518 6496 54524 6560
rect 54588 6496 54604 6560
rect 54668 6496 54684 6560
rect 54748 6496 54764 6560
rect 54828 6496 54834 6560
rect 54518 6495 54834 6496
rect 72918 6560 73234 6561
rect 72918 6496 72924 6560
rect 72988 6496 73004 6560
rect 73068 6496 73084 6560
rect 73148 6496 73164 6560
rect 73228 6496 73234 6560
rect 72918 6495 73234 6496
rect 18378 6016 18694 6017
rect 18378 5952 18384 6016
rect 18448 5952 18464 6016
rect 18528 5952 18544 6016
rect 18608 5952 18624 6016
rect 18688 5952 18694 6016
rect 18378 5951 18694 5952
rect 36778 6016 37094 6017
rect 36778 5952 36784 6016
rect 36848 5952 36864 6016
rect 36928 5952 36944 6016
rect 37008 5952 37024 6016
rect 37088 5952 37094 6016
rect 36778 5951 37094 5952
rect 55178 6016 55494 6017
rect 55178 5952 55184 6016
rect 55248 5952 55264 6016
rect 55328 5952 55344 6016
rect 55408 5952 55424 6016
rect 55488 5952 55494 6016
rect 55178 5951 55494 5952
rect 73578 6016 73894 6017
rect 73578 5952 73584 6016
rect 73648 5952 73664 6016
rect 73728 5952 73744 6016
rect 73808 5952 73824 6016
rect 73888 5952 73894 6016
rect 73578 5951 73894 5952
rect 17718 5472 18034 5473
rect 17718 5408 17724 5472
rect 17788 5408 17804 5472
rect 17868 5408 17884 5472
rect 17948 5408 17964 5472
rect 18028 5408 18034 5472
rect 17718 5407 18034 5408
rect 36118 5472 36434 5473
rect 36118 5408 36124 5472
rect 36188 5408 36204 5472
rect 36268 5408 36284 5472
rect 36348 5408 36364 5472
rect 36428 5408 36434 5472
rect 36118 5407 36434 5408
rect 54518 5472 54834 5473
rect 54518 5408 54524 5472
rect 54588 5408 54604 5472
rect 54668 5408 54684 5472
rect 54748 5408 54764 5472
rect 54828 5408 54834 5472
rect 54518 5407 54834 5408
rect 72918 5472 73234 5473
rect 72918 5408 72924 5472
rect 72988 5408 73004 5472
rect 73068 5408 73084 5472
rect 73148 5408 73164 5472
rect 73228 5408 73234 5472
rect 72918 5407 73234 5408
rect 18378 4928 18694 4929
rect 18378 4864 18384 4928
rect 18448 4864 18464 4928
rect 18528 4864 18544 4928
rect 18608 4864 18624 4928
rect 18688 4864 18694 4928
rect 18378 4863 18694 4864
rect 36778 4928 37094 4929
rect 36778 4864 36784 4928
rect 36848 4864 36864 4928
rect 36928 4864 36944 4928
rect 37008 4864 37024 4928
rect 37088 4864 37094 4928
rect 36778 4863 37094 4864
rect 55178 4928 55494 4929
rect 55178 4864 55184 4928
rect 55248 4864 55264 4928
rect 55328 4864 55344 4928
rect 55408 4864 55424 4928
rect 55488 4864 55494 4928
rect 55178 4863 55494 4864
rect 73578 4928 73894 4929
rect 73578 4864 73584 4928
rect 73648 4864 73664 4928
rect 73728 4864 73744 4928
rect 73808 4864 73824 4928
rect 73888 4864 73894 4928
rect 73578 4863 73894 4864
<< via3 >>
rect 18384 87612 18448 87616
rect 18384 87556 18388 87612
rect 18388 87556 18444 87612
rect 18444 87556 18448 87612
rect 18384 87552 18448 87556
rect 18464 87612 18528 87616
rect 18464 87556 18468 87612
rect 18468 87556 18524 87612
rect 18524 87556 18528 87612
rect 18464 87552 18528 87556
rect 18544 87612 18608 87616
rect 18544 87556 18548 87612
rect 18548 87556 18604 87612
rect 18604 87556 18608 87612
rect 18544 87552 18608 87556
rect 18624 87612 18688 87616
rect 18624 87556 18628 87612
rect 18628 87556 18684 87612
rect 18684 87556 18688 87612
rect 18624 87552 18688 87556
rect 36784 87612 36848 87616
rect 36784 87556 36788 87612
rect 36788 87556 36844 87612
rect 36844 87556 36848 87612
rect 36784 87552 36848 87556
rect 36864 87612 36928 87616
rect 36864 87556 36868 87612
rect 36868 87556 36924 87612
rect 36924 87556 36928 87612
rect 36864 87552 36928 87556
rect 36944 87612 37008 87616
rect 36944 87556 36948 87612
rect 36948 87556 37004 87612
rect 37004 87556 37008 87612
rect 36944 87552 37008 87556
rect 37024 87612 37088 87616
rect 37024 87556 37028 87612
rect 37028 87556 37084 87612
rect 37084 87556 37088 87612
rect 37024 87552 37088 87556
rect 55184 87612 55248 87616
rect 55184 87556 55188 87612
rect 55188 87556 55244 87612
rect 55244 87556 55248 87612
rect 55184 87552 55248 87556
rect 55264 87612 55328 87616
rect 55264 87556 55268 87612
rect 55268 87556 55324 87612
rect 55324 87556 55328 87612
rect 55264 87552 55328 87556
rect 55344 87612 55408 87616
rect 55344 87556 55348 87612
rect 55348 87556 55404 87612
rect 55404 87556 55408 87612
rect 55344 87552 55408 87556
rect 55424 87612 55488 87616
rect 55424 87556 55428 87612
rect 55428 87556 55484 87612
rect 55484 87556 55488 87612
rect 55424 87552 55488 87556
rect 73584 87612 73648 87616
rect 73584 87556 73588 87612
rect 73588 87556 73644 87612
rect 73644 87556 73648 87612
rect 73584 87552 73648 87556
rect 73664 87612 73728 87616
rect 73664 87556 73668 87612
rect 73668 87556 73724 87612
rect 73724 87556 73728 87612
rect 73664 87552 73728 87556
rect 73744 87612 73808 87616
rect 73744 87556 73748 87612
rect 73748 87556 73804 87612
rect 73804 87556 73808 87612
rect 73744 87552 73808 87556
rect 73824 87612 73888 87616
rect 73824 87556 73828 87612
rect 73828 87556 73884 87612
rect 73884 87556 73888 87612
rect 73824 87552 73888 87556
rect 10308 87316 10372 87380
rect 17724 87068 17788 87072
rect 17724 87012 17728 87068
rect 17728 87012 17784 87068
rect 17784 87012 17788 87068
rect 17724 87008 17788 87012
rect 17804 87068 17868 87072
rect 17804 87012 17808 87068
rect 17808 87012 17864 87068
rect 17864 87012 17868 87068
rect 17804 87008 17868 87012
rect 17884 87068 17948 87072
rect 17884 87012 17888 87068
rect 17888 87012 17944 87068
rect 17944 87012 17948 87068
rect 17884 87008 17948 87012
rect 17964 87068 18028 87072
rect 17964 87012 17968 87068
rect 17968 87012 18024 87068
rect 18024 87012 18028 87068
rect 17964 87008 18028 87012
rect 36124 87068 36188 87072
rect 36124 87012 36128 87068
rect 36128 87012 36184 87068
rect 36184 87012 36188 87068
rect 36124 87008 36188 87012
rect 36204 87068 36268 87072
rect 36204 87012 36208 87068
rect 36208 87012 36264 87068
rect 36264 87012 36268 87068
rect 36204 87008 36268 87012
rect 36284 87068 36348 87072
rect 36284 87012 36288 87068
rect 36288 87012 36344 87068
rect 36344 87012 36348 87068
rect 36284 87008 36348 87012
rect 36364 87068 36428 87072
rect 36364 87012 36368 87068
rect 36368 87012 36424 87068
rect 36424 87012 36428 87068
rect 36364 87008 36428 87012
rect 54524 87068 54588 87072
rect 54524 87012 54528 87068
rect 54528 87012 54584 87068
rect 54584 87012 54588 87068
rect 54524 87008 54588 87012
rect 54604 87068 54668 87072
rect 54604 87012 54608 87068
rect 54608 87012 54664 87068
rect 54664 87012 54668 87068
rect 54604 87008 54668 87012
rect 54684 87068 54748 87072
rect 54684 87012 54688 87068
rect 54688 87012 54744 87068
rect 54744 87012 54748 87068
rect 54684 87008 54748 87012
rect 54764 87068 54828 87072
rect 54764 87012 54768 87068
rect 54768 87012 54824 87068
rect 54824 87012 54828 87068
rect 54764 87008 54828 87012
rect 72924 87068 72988 87072
rect 72924 87012 72928 87068
rect 72928 87012 72984 87068
rect 72984 87012 72988 87068
rect 72924 87008 72988 87012
rect 73004 87068 73068 87072
rect 73004 87012 73008 87068
rect 73008 87012 73064 87068
rect 73064 87012 73068 87068
rect 73004 87008 73068 87012
rect 73084 87068 73148 87072
rect 73084 87012 73088 87068
rect 73088 87012 73144 87068
rect 73144 87012 73148 87068
rect 73084 87008 73148 87012
rect 73164 87068 73228 87072
rect 73164 87012 73168 87068
rect 73168 87012 73224 87068
rect 73224 87012 73228 87068
rect 73164 87008 73228 87012
rect 18384 86524 18448 86528
rect 18384 86468 18388 86524
rect 18388 86468 18444 86524
rect 18444 86468 18448 86524
rect 18384 86464 18448 86468
rect 18464 86524 18528 86528
rect 18464 86468 18468 86524
rect 18468 86468 18524 86524
rect 18524 86468 18528 86524
rect 18464 86464 18528 86468
rect 18544 86524 18608 86528
rect 18544 86468 18548 86524
rect 18548 86468 18604 86524
rect 18604 86468 18608 86524
rect 18544 86464 18608 86468
rect 18624 86524 18688 86528
rect 18624 86468 18628 86524
rect 18628 86468 18684 86524
rect 18684 86468 18688 86524
rect 18624 86464 18688 86468
rect 36784 86524 36848 86528
rect 36784 86468 36788 86524
rect 36788 86468 36844 86524
rect 36844 86468 36848 86524
rect 36784 86464 36848 86468
rect 36864 86524 36928 86528
rect 36864 86468 36868 86524
rect 36868 86468 36924 86524
rect 36924 86468 36928 86524
rect 36864 86464 36928 86468
rect 36944 86524 37008 86528
rect 36944 86468 36948 86524
rect 36948 86468 37004 86524
rect 37004 86468 37008 86524
rect 36944 86464 37008 86468
rect 37024 86524 37088 86528
rect 37024 86468 37028 86524
rect 37028 86468 37084 86524
rect 37084 86468 37088 86524
rect 37024 86464 37088 86468
rect 55184 86524 55248 86528
rect 55184 86468 55188 86524
rect 55188 86468 55244 86524
rect 55244 86468 55248 86524
rect 55184 86464 55248 86468
rect 55264 86524 55328 86528
rect 55264 86468 55268 86524
rect 55268 86468 55324 86524
rect 55324 86468 55328 86524
rect 55264 86464 55328 86468
rect 55344 86524 55408 86528
rect 55344 86468 55348 86524
rect 55348 86468 55404 86524
rect 55404 86468 55408 86524
rect 55344 86464 55408 86468
rect 55424 86524 55488 86528
rect 55424 86468 55428 86524
rect 55428 86468 55484 86524
rect 55484 86468 55488 86524
rect 55424 86464 55488 86468
rect 73584 86524 73648 86528
rect 73584 86468 73588 86524
rect 73588 86468 73644 86524
rect 73644 86468 73648 86524
rect 73584 86464 73648 86468
rect 73664 86524 73728 86528
rect 73664 86468 73668 86524
rect 73668 86468 73724 86524
rect 73724 86468 73728 86524
rect 73664 86464 73728 86468
rect 73744 86524 73808 86528
rect 73744 86468 73748 86524
rect 73748 86468 73804 86524
rect 73804 86468 73808 86524
rect 73744 86464 73808 86468
rect 73824 86524 73888 86528
rect 73824 86468 73828 86524
rect 73828 86468 73884 86524
rect 73884 86468 73888 86524
rect 73824 86464 73888 86468
rect 17724 85980 17788 85984
rect 17724 85924 17728 85980
rect 17728 85924 17784 85980
rect 17784 85924 17788 85980
rect 17724 85920 17788 85924
rect 17804 85980 17868 85984
rect 17804 85924 17808 85980
rect 17808 85924 17864 85980
rect 17864 85924 17868 85980
rect 17804 85920 17868 85924
rect 17884 85980 17948 85984
rect 17884 85924 17888 85980
rect 17888 85924 17944 85980
rect 17944 85924 17948 85980
rect 17884 85920 17948 85924
rect 17964 85980 18028 85984
rect 17964 85924 17968 85980
rect 17968 85924 18024 85980
rect 18024 85924 18028 85980
rect 17964 85920 18028 85924
rect 36124 85980 36188 85984
rect 36124 85924 36128 85980
rect 36128 85924 36184 85980
rect 36184 85924 36188 85980
rect 36124 85920 36188 85924
rect 36204 85980 36268 85984
rect 36204 85924 36208 85980
rect 36208 85924 36264 85980
rect 36264 85924 36268 85980
rect 36204 85920 36268 85924
rect 36284 85980 36348 85984
rect 36284 85924 36288 85980
rect 36288 85924 36344 85980
rect 36344 85924 36348 85980
rect 36284 85920 36348 85924
rect 36364 85980 36428 85984
rect 36364 85924 36368 85980
rect 36368 85924 36424 85980
rect 36424 85924 36428 85980
rect 36364 85920 36428 85924
rect 54524 85980 54588 85984
rect 54524 85924 54528 85980
rect 54528 85924 54584 85980
rect 54584 85924 54588 85980
rect 54524 85920 54588 85924
rect 54604 85980 54668 85984
rect 54604 85924 54608 85980
rect 54608 85924 54664 85980
rect 54664 85924 54668 85980
rect 54604 85920 54668 85924
rect 54684 85980 54748 85984
rect 54684 85924 54688 85980
rect 54688 85924 54744 85980
rect 54744 85924 54748 85980
rect 54684 85920 54748 85924
rect 54764 85980 54828 85984
rect 54764 85924 54768 85980
rect 54768 85924 54824 85980
rect 54824 85924 54828 85980
rect 54764 85920 54828 85924
rect 72924 85980 72988 85984
rect 72924 85924 72928 85980
rect 72928 85924 72984 85980
rect 72984 85924 72988 85980
rect 72924 85920 72988 85924
rect 73004 85980 73068 85984
rect 73004 85924 73008 85980
rect 73008 85924 73064 85980
rect 73064 85924 73068 85980
rect 73004 85920 73068 85924
rect 73084 85980 73148 85984
rect 73084 85924 73088 85980
rect 73088 85924 73144 85980
rect 73144 85924 73148 85980
rect 73084 85920 73148 85924
rect 73164 85980 73228 85984
rect 73164 85924 73168 85980
rect 73168 85924 73224 85980
rect 73224 85924 73228 85980
rect 73164 85920 73228 85924
rect 18384 85436 18448 85440
rect 18384 85380 18388 85436
rect 18388 85380 18444 85436
rect 18444 85380 18448 85436
rect 18384 85376 18448 85380
rect 18464 85436 18528 85440
rect 18464 85380 18468 85436
rect 18468 85380 18524 85436
rect 18524 85380 18528 85436
rect 18464 85376 18528 85380
rect 18544 85436 18608 85440
rect 18544 85380 18548 85436
rect 18548 85380 18604 85436
rect 18604 85380 18608 85436
rect 18544 85376 18608 85380
rect 18624 85436 18688 85440
rect 18624 85380 18628 85436
rect 18628 85380 18684 85436
rect 18684 85380 18688 85436
rect 18624 85376 18688 85380
rect 36784 85436 36848 85440
rect 36784 85380 36788 85436
rect 36788 85380 36844 85436
rect 36844 85380 36848 85436
rect 36784 85376 36848 85380
rect 36864 85436 36928 85440
rect 36864 85380 36868 85436
rect 36868 85380 36924 85436
rect 36924 85380 36928 85436
rect 36864 85376 36928 85380
rect 36944 85436 37008 85440
rect 36944 85380 36948 85436
rect 36948 85380 37004 85436
rect 37004 85380 37008 85436
rect 36944 85376 37008 85380
rect 37024 85436 37088 85440
rect 37024 85380 37028 85436
rect 37028 85380 37084 85436
rect 37084 85380 37088 85436
rect 37024 85376 37088 85380
rect 55184 85436 55248 85440
rect 55184 85380 55188 85436
rect 55188 85380 55244 85436
rect 55244 85380 55248 85436
rect 55184 85376 55248 85380
rect 55264 85436 55328 85440
rect 55264 85380 55268 85436
rect 55268 85380 55324 85436
rect 55324 85380 55328 85436
rect 55264 85376 55328 85380
rect 55344 85436 55408 85440
rect 55344 85380 55348 85436
rect 55348 85380 55404 85436
rect 55404 85380 55408 85436
rect 55344 85376 55408 85380
rect 55424 85436 55488 85440
rect 55424 85380 55428 85436
rect 55428 85380 55484 85436
rect 55484 85380 55488 85436
rect 55424 85376 55488 85380
rect 73584 85436 73648 85440
rect 73584 85380 73588 85436
rect 73588 85380 73644 85436
rect 73644 85380 73648 85436
rect 73584 85376 73648 85380
rect 73664 85436 73728 85440
rect 73664 85380 73668 85436
rect 73668 85380 73724 85436
rect 73724 85380 73728 85436
rect 73664 85376 73728 85380
rect 73744 85436 73808 85440
rect 73744 85380 73748 85436
rect 73748 85380 73804 85436
rect 73804 85380 73808 85436
rect 73744 85376 73808 85380
rect 73824 85436 73888 85440
rect 73824 85380 73828 85436
rect 73828 85380 73884 85436
rect 73884 85380 73888 85436
rect 73824 85376 73888 85380
rect 5956 84892 6020 84896
rect 5956 84836 5960 84892
rect 5960 84836 6016 84892
rect 6016 84836 6020 84892
rect 5956 84832 6020 84836
rect 6036 84892 6100 84896
rect 6036 84836 6040 84892
rect 6040 84836 6096 84892
rect 6096 84836 6100 84892
rect 6036 84832 6100 84836
rect 6116 84892 6180 84896
rect 6116 84836 6120 84892
rect 6120 84836 6176 84892
rect 6176 84836 6180 84892
rect 6116 84832 6180 84836
rect 6196 84892 6260 84896
rect 6196 84836 6200 84892
rect 6200 84836 6256 84892
rect 6256 84836 6260 84892
rect 6196 84832 6260 84836
rect 17724 84892 17788 84896
rect 17724 84836 17728 84892
rect 17728 84836 17784 84892
rect 17784 84836 17788 84892
rect 17724 84832 17788 84836
rect 17804 84892 17868 84896
rect 17804 84836 17808 84892
rect 17808 84836 17864 84892
rect 17864 84836 17868 84892
rect 17804 84832 17868 84836
rect 17884 84892 17948 84896
rect 17884 84836 17888 84892
rect 17888 84836 17944 84892
rect 17944 84836 17948 84892
rect 17884 84832 17948 84836
rect 17964 84892 18028 84896
rect 17964 84836 17968 84892
rect 17968 84836 18024 84892
rect 18024 84836 18028 84892
rect 17964 84832 18028 84836
rect 36124 84892 36188 84896
rect 36124 84836 36128 84892
rect 36128 84836 36184 84892
rect 36184 84836 36188 84892
rect 36124 84832 36188 84836
rect 36204 84892 36268 84896
rect 36204 84836 36208 84892
rect 36208 84836 36264 84892
rect 36264 84836 36268 84892
rect 36204 84832 36268 84836
rect 36284 84892 36348 84896
rect 36284 84836 36288 84892
rect 36288 84836 36344 84892
rect 36344 84836 36348 84892
rect 36284 84832 36348 84836
rect 36364 84892 36428 84896
rect 36364 84836 36368 84892
rect 36368 84836 36424 84892
rect 36424 84836 36428 84892
rect 36364 84832 36428 84836
rect 54524 84892 54588 84896
rect 54524 84836 54528 84892
rect 54528 84836 54584 84892
rect 54584 84836 54588 84892
rect 54524 84832 54588 84836
rect 54604 84892 54668 84896
rect 54604 84836 54608 84892
rect 54608 84836 54664 84892
rect 54664 84836 54668 84892
rect 54604 84832 54668 84836
rect 54684 84892 54748 84896
rect 54684 84836 54688 84892
rect 54688 84836 54744 84892
rect 54744 84836 54748 84892
rect 54684 84832 54748 84836
rect 54764 84892 54828 84896
rect 54764 84836 54768 84892
rect 54768 84836 54824 84892
rect 54824 84836 54828 84892
rect 54764 84832 54828 84836
rect 72924 84892 72988 84896
rect 72924 84836 72928 84892
rect 72928 84836 72984 84892
rect 72984 84836 72988 84892
rect 72924 84832 72988 84836
rect 73004 84892 73068 84896
rect 73004 84836 73008 84892
rect 73008 84836 73064 84892
rect 73064 84836 73068 84892
rect 73004 84832 73068 84836
rect 73084 84892 73148 84896
rect 73084 84836 73088 84892
rect 73088 84836 73144 84892
rect 73144 84836 73148 84892
rect 73084 84832 73148 84836
rect 73164 84892 73228 84896
rect 73164 84836 73168 84892
rect 73168 84836 73224 84892
rect 73224 84836 73228 84892
rect 73164 84832 73228 84836
rect 86548 84892 86612 84896
rect 86548 84836 86552 84892
rect 86552 84836 86608 84892
rect 86608 84836 86612 84892
rect 86548 84832 86612 84836
rect 86628 84892 86692 84896
rect 86628 84836 86632 84892
rect 86632 84836 86688 84892
rect 86688 84836 86692 84892
rect 86628 84832 86692 84836
rect 86708 84892 86772 84896
rect 86708 84836 86712 84892
rect 86712 84836 86768 84892
rect 86768 84836 86772 84892
rect 86708 84832 86772 84836
rect 86788 84892 86852 84896
rect 86788 84836 86792 84892
rect 86792 84836 86848 84892
rect 86848 84836 86852 84892
rect 86788 84832 86852 84836
rect 6692 84348 6756 84352
rect 6692 84292 6696 84348
rect 6696 84292 6752 84348
rect 6752 84292 6756 84348
rect 6692 84288 6756 84292
rect 6772 84348 6836 84352
rect 6772 84292 6776 84348
rect 6776 84292 6832 84348
rect 6832 84292 6836 84348
rect 6772 84288 6836 84292
rect 6852 84348 6916 84352
rect 6852 84292 6856 84348
rect 6856 84292 6912 84348
rect 6912 84292 6916 84348
rect 6852 84288 6916 84292
rect 6932 84348 6996 84352
rect 6932 84292 6936 84348
rect 6936 84292 6992 84348
rect 6992 84292 6996 84348
rect 6932 84288 6996 84292
rect 18384 84348 18448 84352
rect 18384 84292 18388 84348
rect 18388 84292 18444 84348
rect 18444 84292 18448 84348
rect 18384 84288 18448 84292
rect 18464 84348 18528 84352
rect 18464 84292 18468 84348
rect 18468 84292 18524 84348
rect 18524 84292 18528 84348
rect 18464 84288 18528 84292
rect 18544 84348 18608 84352
rect 18544 84292 18548 84348
rect 18548 84292 18604 84348
rect 18604 84292 18608 84348
rect 18544 84288 18608 84292
rect 18624 84348 18688 84352
rect 18624 84292 18628 84348
rect 18628 84292 18684 84348
rect 18684 84292 18688 84348
rect 18624 84288 18688 84292
rect 36784 84348 36848 84352
rect 36784 84292 36788 84348
rect 36788 84292 36844 84348
rect 36844 84292 36848 84348
rect 36784 84288 36848 84292
rect 36864 84348 36928 84352
rect 36864 84292 36868 84348
rect 36868 84292 36924 84348
rect 36924 84292 36928 84348
rect 36864 84288 36928 84292
rect 36944 84348 37008 84352
rect 36944 84292 36948 84348
rect 36948 84292 37004 84348
rect 37004 84292 37008 84348
rect 36944 84288 37008 84292
rect 37024 84348 37088 84352
rect 37024 84292 37028 84348
rect 37028 84292 37084 84348
rect 37084 84292 37088 84348
rect 37024 84288 37088 84292
rect 55184 84348 55248 84352
rect 55184 84292 55188 84348
rect 55188 84292 55244 84348
rect 55244 84292 55248 84348
rect 55184 84288 55248 84292
rect 55264 84348 55328 84352
rect 55264 84292 55268 84348
rect 55268 84292 55324 84348
rect 55324 84292 55328 84348
rect 55264 84288 55328 84292
rect 55344 84348 55408 84352
rect 55344 84292 55348 84348
rect 55348 84292 55404 84348
rect 55404 84292 55408 84348
rect 55344 84288 55408 84292
rect 55424 84348 55488 84352
rect 55424 84292 55428 84348
rect 55428 84292 55484 84348
rect 55484 84292 55488 84348
rect 55424 84288 55488 84292
rect 73584 84348 73648 84352
rect 73584 84292 73588 84348
rect 73588 84292 73644 84348
rect 73644 84292 73648 84348
rect 73584 84288 73648 84292
rect 73664 84348 73728 84352
rect 73664 84292 73668 84348
rect 73668 84292 73724 84348
rect 73724 84292 73728 84348
rect 73664 84288 73728 84292
rect 73744 84348 73808 84352
rect 73744 84292 73748 84348
rect 73748 84292 73804 84348
rect 73804 84292 73808 84348
rect 73744 84288 73808 84292
rect 73824 84348 73888 84352
rect 73824 84292 73828 84348
rect 73828 84292 73884 84348
rect 73884 84292 73888 84348
rect 73824 84288 73888 84292
rect 87284 84348 87348 84352
rect 87284 84292 87288 84348
rect 87288 84292 87344 84348
rect 87344 84292 87348 84348
rect 87284 84288 87348 84292
rect 87364 84348 87428 84352
rect 87364 84292 87368 84348
rect 87368 84292 87424 84348
rect 87424 84292 87428 84348
rect 87364 84288 87428 84292
rect 87444 84348 87508 84352
rect 87444 84292 87448 84348
rect 87448 84292 87504 84348
rect 87504 84292 87508 84348
rect 87444 84288 87508 84292
rect 87524 84348 87588 84352
rect 87524 84292 87528 84348
rect 87528 84292 87584 84348
rect 87584 84292 87588 84348
rect 87524 84288 87588 84292
rect 5956 83804 6020 83808
rect 5956 83748 5960 83804
rect 5960 83748 6016 83804
rect 6016 83748 6020 83804
rect 5956 83744 6020 83748
rect 6036 83804 6100 83808
rect 6036 83748 6040 83804
rect 6040 83748 6096 83804
rect 6096 83748 6100 83804
rect 6036 83744 6100 83748
rect 6116 83804 6180 83808
rect 6116 83748 6120 83804
rect 6120 83748 6176 83804
rect 6176 83748 6180 83804
rect 6116 83744 6180 83748
rect 6196 83804 6260 83808
rect 6196 83748 6200 83804
rect 6200 83748 6256 83804
rect 6256 83748 6260 83804
rect 6196 83744 6260 83748
rect 86548 83804 86612 83808
rect 86548 83748 86552 83804
rect 86552 83748 86608 83804
rect 86608 83748 86612 83804
rect 86548 83744 86612 83748
rect 86628 83804 86692 83808
rect 86628 83748 86632 83804
rect 86632 83748 86688 83804
rect 86688 83748 86692 83804
rect 86628 83744 86692 83748
rect 86708 83804 86772 83808
rect 86708 83748 86712 83804
rect 86712 83748 86768 83804
rect 86768 83748 86772 83804
rect 86708 83744 86772 83748
rect 86788 83804 86852 83808
rect 86788 83748 86792 83804
rect 86792 83748 86848 83804
rect 86848 83748 86852 83804
rect 86788 83744 86852 83748
rect 6692 83260 6756 83264
rect 6692 83204 6696 83260
rect 6696 83204 6752 83260
rect 6752 83204 6756 83260
rect 6692 83200 6756 83204
rect 6772 83260 6836 83264
rect 6772 83204 6776 83260
rect 6776 83204 6832 83260
rect 6832 83204 6836 83260
rect 6772 83200 6836 83204
rect 6852 83260 6916 83264
rect 6852 83204 6856 83260
rect 6856 83204 6912 83260
rect 6912 83204 6916 83260
rect 6852 83200 6916 83204
rect 6932 83260 6996 83264
rect 6932 83204 6936 83260
rect 6936 83204 6992 83260
rect 6992 83204 6996 83260
rect 6932 83200 6996 83204
rect 87284 83260 87348 83264
rect 87284 83204 87288 83260
rect 87288 83204 87344 83260
rect 87344 83204 87348 83260
rect 87284 83200 87348 83204
rect 87364 83260 87428 83264
rect 87364 83204 87368 83260
rect 87368 83204 87424 83260
rect 87424 83204 87428 83260
rect 87364 83200 87428 83204
rect 87444 83260 87508 83264
rect 87444 83204 87448 83260
rect 87448 83204 87504 83260
rect 87504 83204 87508 83260
rect 87444 83200 87508 83204
rect 87524 83260 87588 83264
rect 87524 83204 87528 83260
rect 87528 83204 87584 83260
rect 87584 83204 87588 83260
rect 87524 83200 87588 83204
rect 5956 82716 6020 82720
rect 5956 82660 5960 82716
rect 5960 82660 6016 82716
rect 6016 82660 6020 82716
rect 5956 82656 6020 82660
rect 6036 82716 6100 82720
rect 6036 82660 6040 82716
rect 6040 82660 6096 82716
rect 6096 82660 6100 82716
rect 6036 82656 6100 82660
rect 6116 82716 6180 82720
rect 6116 82660 6120 82716
rect 6120 82660 6176 82716
rect 6176 82660 6180 82716
rect 6116 82656 6180 82660
rect 6196 82716 6260 82720
rect 6196 82660 6200 82716
rect 6200 82660 6256 82716
rect 6256 82660 6260 82716
rect 6196 82656 6260 82660
rect 86548 82716 86612 82720
rect 86548 82660 86552 82716
rect 86552 82660 86608 82716
rect 86608 82660 86612 82716
rect 86548 82656 86612 82660
rect 86628 82716 86692 82720
rect 86628 82660 86632 82716
rect 86632 82660 86688 82716
rect 86688 82660 86692 82716
rect 86628 82656 86692 82660
rect 86708 82716 86772 82720
rect 86708 82660 86712 82716
rect 86712 82660 86768 82716
rect 86768 82660 86772 82716
rect 86708 82656 86772 82660
rect 86788 82716 86852 82720
rect 86788 82660 86792 82716
rect 86792 82660 86848 82716
rect 86848 82660 86852 82716
rect 86788 82656 86852 82660
rect 6692 82172 6756 82176
rect 6692 82116 6696 82172
rect 6696 82116 6752 82172
rect 6752 82116 6756 82172
rect 6692 82112 6756 82116
rect 6772 82172 6836 82176
rect 6772 82116 6776 82172
rect 6776 82116 6832 82172
rect 6832 82116 6836 82172
rect 6772 82112 6836 82116
rect 6852 82172 6916 82176
rect 6852 82116 6856 82172
rect 6856 82116 6912 82172
rect 6912 82116 6916 82172
rect 6852 82112 6916 82116
rect 6932 82172 6996 82176
rect 6932 82116 6936 82172
rect 6936 82116 6992 82172
rect 6992 82116 6996 82172
rect 6932 82112 6996 82116
rect 87284 82172 87348 82176
rect 87284 82116 87288 82172
rect 87288 82116 87344 82172
rect 87344 82116 87348 82172
rect 87284 82112 87348 82116
rect 87364 82172 87428 82176
rect 87364 82116 87368 82172
rect 87368 82116 87424 82172
rect 87424 82116 87428 82172
rect 87364 82112 87428 82116
rect 87444 82172 87508 82176
rect 87444 82116 87448 82172
rect 87448 82116 87504 82172
rect 87504 82116 87508 82172
rect 87444 82112 87508 82116
rect 87524 82172 87588 82176
rect 87524 82116 87528 82172
rect 87528 82116 87584 82172
rect 87584 82116 87588 82172
rect 87524 82112 87588 82116
rect 5956 81628 6020 81632
rect 5956 81572 5960 81628
rect 5960 81572 6016 81628
rect 6016 81572 6020 81628
rect 5956 81568 6020 81572
rect 6036 81628 6100 81632
rect 6036 81572 6040 81628
rect 6040 81572 6096 81628
rect 6096 81572 6100 81628
rect 6036 81568 6100 81572
rect 6116 81628 6180 81632
rect 6116 81572 6120 81628
rect 6120 81572 6176 81628
rect 6176 81572 6180 81628
rect 6116 81568 6180 81572
rect 6196 81628 6260 81632
rect 6196 81572 6200 81628
rect 6200 81572 6256 81628
rect 6256 81572 6260 81628
rect 6196 81568 6260 81572
rect 86548 81628 86612 81632
rect 86548 81572 86552 81628
rect 86552 81572 86608 81628
rect 86608 81572 86612 81628
rect 86548 81568 86612 81572
rect 86628 81628 86692 81632
rect 86628 81572 86632 81628
rect 86632 81572 86688 81628
rect 86688 81572 86692 81628
rect 86628 81568 86692 81572
rect 86708 81628 86772 81632
rect 86708 81572 86712 81628
rect 86712 81572 86768 81628
rect 86768 81572 86772 81628
rect 86708 81568 86772 81572
rect 86788 81628 86852 81632
rect 86788 81572 86792 81628
rect 86792 81572 86848 81628
rect 86848 81572 86852 81628
rect 86788 81568 86852 81572
rect 6692 81084 6756 81088
rect 6692 81028 6696 81084
rect 6696 81028 6752 81084
rect 6752 81028 6756 81084
rect 6692 81024 6756 81028
rect 6772 81084 6836 81088
rect 6772 81028 6776 81084
rect 6776 81028 6832 81084
rect 6832 81028 6836 81084
rect 6772 81024 6836 81028
rect 6852 81084 6916 81088
rect 6852 81028 6856 81084
rect 6856 81028 6912 81084
rect 6912 81028 6916 81084
rect 6852 81024 6916 81028
rect 6932 81084 6996 81088
rect 6932 81028 6936 81084
rect 6936 81028 6992 81084
rect 6992 81028 6996 81084
rect 6932 81024 6996 81028
rect 10308 80992 10372 81056
rect 87284 81084 87348 81088
rect 87284 81028 87288 81084
rect 87288 81028 87344 81084
rect 87344 81028 87348 81084
rect 87284 81024 87348 81028
rect 87364 81084 87428 81088
rect 87364 81028 87368 81084
rect 87368 81028 87424 81084
rect 87424 81028 87428 81084
rect 87364 81024 87428 81028
rect 87444 81084 87508 81088
rect 87444 81028 87448 81084
rect 87448 81028 87504 81084
rect 87504 81028 87508 81084
rect 87444 81024 87508 81028
rect 87524 81084 87588 81088
rect 87524 81028 87528 81084
rect 87528 81028 87584 81084
rect 87584 81028 87588 81084
rect 87524 81024 87588 81028
rect 5956 80540 6020 80544
rect 5956 80484 5960 80540
rect 5960 80484 6016 80540
rect 6016 80484 6020 80540
rect 5956 80480 6020 80484
rect 6036 80540 6100 80544
rect 6036 80484 6040 80540
rect 6040 80484 6096 80540
rect 6096 80484 6100 80540
rect 6036 80480 6100 80484
rect 6116 80540 6180 80544
rect 6116 80484 6120 80540
rect 6120 80484 6176 80540
rect 6176 80484 6180 80540
rect 6116 80480 6180 80484
rect 6196 80540 6260 80544
rect 6196 80484 6200 80540
rect 6200 80484 6256 80540
rect 6256 80484 6260 80540
rect 6196 80480 6260 80484
rect 86548 80540 86612 80544
rect 86548 80484 86552 80540
rect 86552 80484 86608 80540
rect 86608 80484 86612 80540
rect 86548 80480 86612 80484
rect 86628 80540 86692 80544
rect 86628 80484 86632 80540
rect 86632 80484 86688 80540
rect 86688 80484 86692 80540
rect 86628 80480 86692 80484
rect 86708 80540 86772 80544
rect 86708 80484 86712 80540
rect 86712 80484 86768 80540
rect 86768 80484 86772 80540
rect 86708 80480 86772 80484
rect 86788 80540 86852 80544
rect 86788 80484 86792 80540
rect 86792 80484 86848 80540
rect 86848 80484 86852 80540
rect 86788 80480 86852 80484
rect 6692 79996 6756 80000
rect 6692 79940 6696 79996
rect 6696 79940 6752 79996
rect 6752 79940 6756 79996
rect 6692 79936 6756 79940
rect 6772 79996 6836 80000
rect 6772 79940 6776 79996
rect 6776 79940 6832 79996
rect 6832 79940 6836 79996
rect 6772 79936 6836 79940
rect 6852 79996 6916 80000
rect 6852 79940 6856 79996
rect 6856 79940 6912 79996
rect 6912 79940 6916 79996
rect 6852 79936 6916 79940
rect 6932 79996 6996 80000
rect 6932 79940 6936 79996
rect 6936 79940 6992 79996
rect 6992 79940 6996 79996
rect 6932 79936 6996 79940
rect 87284 79996 87348 80000
rect 87284 79940 87288 79996
rect 87288 79940 87344 79996
rect 87344 79940 87348 79996
rect 87284 79936 87348 79940
rect 87364 79996 87428 80000
rect 87364 79940 87368 79996
rect 87368 79940 87424 79996
rect 87424 79940 87428 79996
rect 87364 79936 87428 79940
rect 87444 79996 87508 80000
rect 87444 79940 87448 79996
rect 87448 79940 87504 79996
rect 87504 79940 87508 79996
rect 87444 79936 87508 79940
rect 87524 79996 87588 80000
rect 87524 79940 87528 79996
rect 87528 79940 87584 79996
rect 87584 79940 87588 79996
rect 87524 79936 87588 79940
rect 5956 79452 6020 79456
rect 5956 79396 5960 79452
rect 5960 79396 6016 79452
rect 6016 79396 6020 79452
rect 5956 79392 6020 79396
rect 6036 79452 6100 79456
rect 6036 79396 6040 79452
rect 6040 79396 6096 79452
rect 6096 79396 6100 79452
rect 6036 79392 6100 79396
rect 6116 79452 6180 79456
rect 6116 79396 6120 79452
rect 6120 79396 6176 79452
rect 6176 79396 6180 79452
rect 6116 79392 6180 79396
rect 6196 79452 6260 79456
rect 6196 79396 6200 79452
rect 6200 79396 6256 79452
rect 6256 79396 6260 79452
rect 6196 79392 6260 79396
rect 86548 79452 86612 79456
rect 86548 79396 86552 79452
rect 86552 79396 86608 79452
rect 86608 79396 86612 79452
rect 86548 79392 86612 79396
rect 86628 79452 86692 79456
rect 86628 79396 86632 79452
rect 86632 79396 86688 79452
rect 86688 79396 86692 79452
rect 86628 79392 86692 79396
rect 86708 79452 86772 79456
rect 86708 79396 86712 79452
rect 86712 79396 86768 79452
rect 86768 79396 86772 79452
rect 86708 79392 86772 79396
rect 86788 79452 86852 79456
rect 86788 79396 86792 79452
rect 86792 79396 86848 79452
rect 86848 79396 86852 79452
rect 86788 79392 86852 79396
rect 6692 78908 6756 78912
rect 6692 78852 6696 78908
rect 6696 78852 6752 78908
rect 6752 78852 6756 78908
rect 6692 78848 6756 78852
rect 6772 78908 6836 78912
rect 6772 78852 6776 78908
rect 6776 78852 6832 78908
rect 6832 78852 6836 78908
rect 6772 78848 6836 78852
rect 6852 78908 6916 78912
rect 6852 78852 6856 78908
rect 6856 78852 6912 78908
rect 6912 78852 6916 78908
rect 6852 78848 6916 78852
rect 6932 78908 6996 78912
rect 6932 78852 6936 78908
rect 6936 78852 6992 78908
rect 6992 78852 6996 78908
rect 6932 78848 6996 78852
rect 87284 78908 87348 78912
rect 87284 78852 87288 78908
rect 87288 78852 87344 78908
rect 87344 78852 87348 78908
rect 87284 78848 87348 78852
rect 87364 78908 87428 78912
rect 87364 78852 87368 78908
rect 87368 78852 87424 78908
rect 87424 78852 87428 78908
rect 87364 78848 87428 78852
rect 87444 78908 87508 78912
rect 87444 78852 87448 78908
rect 87448 78852 87504 78908
rect 87504 78852 87508 78908
rect 87444 78848 87508 78852
rect 87524 78908 87588 78912
rect 87524 78852 87528 78908
rect 87528 78852 87584 78908
rect 87584 78852 87588 78908
rect 87524 78848 87588 78852
rect 5956 78364 6020 78368
rect 5956 78308 5960 78364
rect 5960 78308 6016 78364
rect 6016 78308 6020 78364
rect 5956 78304 6020 78308
rect 6036 78364 6100 78368
rect 6036 78308 6040 78364
rect 6040 78308 6096 78364
rect 6096 78308 6100 78364
rect 6036 78304 6100 78308
rect 6116 78364 6180 78368
rect 6116 78308 6120 78364
rect 6120 78308 6176 78364
rect 6176 78308 6180 78364
rect 6116 78304 6180 78308
rect 6196 78364 6260 78368
rect 6196 78308 6200 78364
rect 6200 78308 6256 78364
rect 6256 78308 6260 78364
rect 6196 78304 6260 78308
rect 86548 78364 86612 78368
rect 86548 78308 86552 78364
rect 86552 78308 86608 78364
rect 86608 78308 86612 78364
rect 86548 78304 86612 78308
rect 86628 78364 86692 78368
rect 86628 78308 86632 78364
rect 86632 78308 86688 78364
rect 86688 78308 86692 78364
rect 86628 78304 86692 78308
rect 86708 78364 86772 78368
rect 86708 78308 86712 78364
rect 86712 78308 86768 78364
rect 86768 78308 86772 78364
rect 86708 78304 86772 78308
rect 86788 78364 86852 78368
rect 86788 78308 86792 78364
rect 86792 78308 86848 78364
rect 86848 78308 86852 78364
rect 86788 78304 86852 78308
rect 6692 77820 6756 77824
rect 6692 77764 6696 77820
rect 6696 77764 6752 77820
rect 6752 77764 6756 77820
rect 6692 77760 6756 77764
rect 6772 77820 6836 77824
rect 6772 77764 6776 77820
rect 6776 77764 6832 77820
rect 6832 77764 6836 77820
rect 6772 77760 6836 77764
rect 6852 77820 6916 77824
rect 6852 77764 6856 77820
rect 6856 77764 6912 77820
rect 6912 77764 6916 77820
rect 6852 77760 6916 77764
rect 6932 77820 6996 77824
rect 6932 77764 6936 77820
rect 6936 77764 6992 77820
rect 6992 77764 6996 77820
rect 6932 77760 6996 77764
rect 87284 77820 87348 77824
rect 87284 77764 87288 77820
rect 87288 77764 87344 77820
rect 87344 77764 87348 77820
rect 87284 77760 87348 77764
rect 87364 77820 87428 77824
rect 87364 77764 87368 77820
rect 87368 77764 87424 77820
rect 87424 77764 87428 77820
rect 87364 77760 87428 77764
rect 87444 77820 87508 77824
rect 87444 77764 87448 77820
rect 87448 77764 87504 77820
rect 87504 77764 87508 77820
rect 87444 77760 87508 77764
rect 87524 77820 87588 77824
rect 87524 77764 87528 77820
rect 87528 77764 87584 77820
rect 87584 77764 87588 77820
rect 87524 77760 87588 77764
rect 5956 77276 6020 77280
rect 5956 77220 5960 77276
rect 5960 77220 6016 77276
rect 6016 77220 6020 77276
rect 5956 77216 6020 77220
rect 6036 77276 6100 77280
rect 6036 77220 6040 77276
rect 6040 77220 6096 77276
rect 6096 77220 6100 77276
rect 6036 77216 6100 77220
rect 6116 77276 6180 77280
rect 6116 77220 6120 77276
rect 6120 77220 6176 77276
rect 6176 77220 6180 77276
rect 6116 77216 6180 77220
rect 6196 77276 6260 77280
rect 6196 77220 6200 77276
rect 6200 77220 6256 77276
rect 6256 77220 6260 77276
rect 6196 77216 6260 77220
rect 86548 77276 86612 77280
rect 86548 77220 86552 77276
rect 86552 77220 86608 77276
rect 86608 77220 86612 77276
rect 86548 77216 86612 77220
rect 86628 77276 86692 77280
rect 86628 77220 86632 77276
rect 86632 77220 86688 77276
rect 86688 77220 86692 77276
rect 86628 77216 86692 77220
rect 86708 77276 86772 77280
rect 86708 77220 86712 77276
rect 86712 77220 86768 77276
rect 86768 77220 86772 77276
rect 86708 77216 86772 77220
rect 86788 77276 86852 77280
rect 86788 77220 86792 77276
rect 86792 77220 86848 77276
rect 86848 77220 86852 77276
rect 86788 77216 86852 77220
rect 6692 76732 6756 76736
rect 6692 76676 6696 76732
rect 6696 76676 6752 76732
rect 6752 76676 6756 76732
rect 6692 76672 6756 76676
rect 6772 76732 6836 76736
rect 6772 76676 6776 76732
rect 6776 76676 6832 76732
rect 6832 76676 6836 76732
rect 6772 76672 6836 76676
rect 6852 76732 6916 76736
rect 6852 76676 6856 76732
rect 6856 76676 6912 76732
rect 6912 76676 6916 76732
rect 6852 76672 6916 76676
rect 6932 76732 6996 76736
rect 6932 76676 6936 76732
rect 6936 76676 6992 76732
rect 6992 76676 6996 76732
rect 6932 76672 6996 76676
rect 87284 76732 87348 76736
rect 87284 76676 87288 76732
rect 87288 76676 87344 76732
rect 87344 76676 87348 76732
rect 87284 76672 87348 76676
rect 87364 76732 87428 76736
rect 87364 76676 87368 76732
rect 87368 76676 87424 76732
rect 87424 76676 87428 76732
rect 87364 76672 87428 76676
rect 87444 76732 87508 76736
rect 87444 76676 87448 76732
rect 87448 76676 87504 76732
rect 87504 76676 87508 76732
rect 87444 76672 87508 76676
rect 87524 76732 87588 76736
rect 87524 76676 87528 76732
rect 87528 76676 87584 76732
rect 87584 76676 87588 76732
rect 87524 76672 87588 76676
rect 5956 76188 6020 76192
rect 5956 76132 5960 76188
rect 5960 76132 6016 76188
rect 6016 76132 6020 76188
rect 5956 76128 6020 76132
rect 6036 76188 6100 76192
rect 6036 76132 6040 76188
rect 6040 76132 6096 76188
rect 6096 76132 6100 76188
rect 6036 76128 6100 76132
rect 6116 76188 6180 76192
rect 6116 76132 6120 76188
rect 6120 76132 6176 76188
rect 6176 76132 6180 76188
rect 6116 76128 6180 76132
rect 6196 76188 6260 76192
rect 6196 76132 6200 76188
rect 6200 76132 6256 76188
rect 6256 76132 6260 76188
rect 6196 76128 6260 76132
rect 86548 76188 86612 76192
rect 86548 76132 86552 76188
rect 86552 76132 86608 76188
rect 86608 76132 86612 76188
rect 86548 76128 86612 76132
rect 86628 76188 86692 76192
rect 86628 76132 86632 76188
rect 86632 76132 86688 76188
rect 86688 76132 86692 76188
rect 86628 76128 86692 76132
rect 86708 76188 86772 76192
rect 86708 76132 86712 76188
rect 86712 76132 86768 76188
rect 86768 76132 86772 76188
rect 86708 76128 86772 76132
rect 86788 76188 86852 76192
rect 86788 76132 86792 76188
rect 86792 76132 86848 76188
rect 86848 76132 86852 76188
rect 86788 76128 86852 76132
rect 6692 75644 6756 75648
rect 6692 75588 6696 75644
rect 6696 75588 6752 75644
rect 6752 75588 6756 75644
rect 6692 75584 6756 75588
rect 6772 75644 6836 75648
rect 6772 75588 6776 75644
rect 6776 75588 6832 75644
rect 6832 75588 6836 75644
rect 6772 75584 6836 75588
rect 6852 75644 6916 75648
rect 6852 75588 6856 75644
rect 6856 75588 6912 75644
rect 6912 75588 6916 75644
rect 6852 75584 6916 75588
rect 6932 75644 6996 75648
rect 6932 75588 6936 75644
rect 6936 75588 6992 75644
rect 6992 75588 6996 75644
rect 6932 75584 6996 75588
rect 87284 75644 87348 75648
rect 87284 75588 87288 75644
rect 87288 75588 87344 75644
rect 87344 75588 87348 75644
rect 87284 75584 87348 75588
rect 87364 75644 87428 75648
rect 87364 75588 87368 75644
rect 87368 75588 87424 75644
rect 87424 75588 87428 75644
rect 87364 75584 87428 75588
rect 87444 75644 87508 75648
rect 87444 75588 87448 75644
rect 87448 75588 87504 75644
rect 87504 75588 87508 75644
rect 87444 75584 87508 75588
rect 87524 75644 87588 75648
rect 87524 75588 87528 75644
rect 87528 75588 87584 75644
rect 87584 75588 87588 75644
rect 87524 75584 87588 75588
rect 5956 75100 6020 75104
rect 5956 75044 5960 75100
rect 5960 75044 6016 75100
rect 6016 75044 6020 75100
rect 5956 75040 6020 75044
rect 6036 75100 6100 75104
rect 6036 75044 6040 75100
rect 6040 75044 6096 75100
rect 6096 75044 6100 75100
rect 6036 75040 6100 75044
rect 6116 75100 6180 75104
rect 6116 75044 6120 75100
rect 6120 75044 6176 75100
rect 6176 75044 6180 75100
rect 6116 75040 6180 75044
rect 6196 75100 6260 75104
rect 6196 75044 6200 75100
rect 6200 75044 6256 75100
rect 6256 75044 6260 75100
rect 6196 75040 6260 75044
rect 86548 75100 86612 75104
rect 86548 75044 86552 75100
rect 86552 75044 86608 75100
rect 86608 75044 86612 75100
rect 86548 75040 86612 75044
rect 86628 75100 86692 75104
rect 86628 75044 86632 75100
rect 86632 75044 86688 75100
rect 86688 75044 86692 75100
rect 86628 75040 86692 75044
rect 86708 75100 86772 75104
rect 86708 75044 86712 75100
rect 86712 75044 86768 75100
rect 86768 75044 86772 75100
rect 86708 75040 86772 75044
rect 86788 75100 86852 75104
rect 86788 75044 86792 75100
rect 86792 75044 86848 75100
rect 86848 75044 86852 75100
rect 86788 75040 86852 75044
rect 6692 74556 6756 74560
rect 6692 74500 6696 74556
rect 6696 74500 6752 74556
rect 6752 74500 6756 74556
rect 6692 74496 6756 74500
rect 6772 74556 6836 74560
rect 6772 74500 6776 74556
rect 6776 74500 6832 74556
rect 6832 74500 6836 74556
rect 6772 74496 6836 74500
rect 6852 74556 6916 74560
rect 6852 74500 6856 74556
rect 6856 74500 6912 74556
rect 6912 74500 6916 74556
rect 6852 74496 6916 74500
rect 6932 74556 6996 74560
rect 6932 74500 6936 74556
rect 6936 74500 6992 74556
rect 6992 74500 6996 74556
rect 6932 74496 6996 74500
rect 87284 74556 87348 74560
rect 87284 74500 87288 74556
rect 87288 74500 87344 74556
rect 87344 74500 87348 74556
rect 87284 74496 87348 74500
rect 87364 74556 87428 74560
rect 87364 74500 87368 74556
rect 87368 74500 87424 74556
rect 87424 74500 87428 74556
rect 87364 74496 87428 74500
rect 87444 74556 87508 74560
rect 87444 74500 87448 74556
rect 87448 74500 87504 74556
rect 87504 74500 87508 74556
rect 87444 74496 87508 74500
rect 87524 74556 87588 74560
rect 87524 74500 87528 74556
rect 87528 74500 87584 74556
rect 87584 74500 87588 74556
rect 87524 74496 87588 74500
rect 5956 74012 6020 74016
rect 5956 73956 5960 74012
rect 5960 73956 6016 74012
rect 6016 73956 6020 74012
rect 5956 73952 6020 73956
rect 6036 74012 6100 74016
rect 6036 73956 6040 74012
rect 6040 73956 6096 74012
rect 6096 73956 6100 74012
rect 6036 73952 6100 73956
rect 6116 74012 6180 74016
rect 6116 73956 6120 74012
rect 6120 73956 6176 74012
rect 6176 73956 6180 74012
rect 6116 73952 6180 73956
rect 6196 74012 6260 74016
rect 6196 73956 6200 74012
rect 6200 73956 6256 74012
rect 6256 73956 6260 74012
rect 6196 73952 6260 73956
rect 86548 74012 86612 74016
rect 86548 73956 86552 74012
rect 86552 73956 86608 74012
rect 86608 73956 86612 74012
rect 86548 73952 86612 73956
rect 86628 74012 86692 74016
rect 86628 73956 86632 74012
rect 86632 73956 86688 74012
rect 86688 73956 86692 74012
rect 86628 73952 86692 73956
rect 86708 74012 86772 74016
rect 86708 73956 86712 74012
rect 86712 73956 86768 74012
rect 86768 73956 86772 74012
rect 86708 73952 86772 73956
rect 86788 74012 86852 74016
rect 86788 73956 86792 74012
rect 86792 73956 86848 74012
rect 86848 73956 86852 74012
rect 86788 73952 86852 73956
rect 6692 73468 6756 73472
rect 6692 73412 6696 73468
rect 6696 73412 6752 73468
rect 6752 73412 6756 73468
rect 6692 73408 6756 73412
rect 6772 73468 6836 73472
rect 6772 73412 6776 73468
rect 6776 73412 6832 73468
rect 6832 73412 6836 73468
rect 6772 73408 6836 73412
rect 6852 73468 6916 73472
rect 6852 73412 6856 73468
rect 6856 73412 6912 73468
rect 6912 73412 6916 73468
rect 6852 73408 6916 73412
rect 6932 73468 6996 73472
rect 6932 73412 6936 73468
rect 6936 73412 6992 73468
rect 6992 73412 6996 73468
rect 6932 73408 6996 73412
rect 87284 73468 87348 73472
rect 87284 73412 87288 73468
rect 87288 73412 87344 73468
rect 87344 73412 87348 73468
rect 87284 73408 87348 73412
rect 87364 73468 87428 73472
rect 87364 73412 87368 73468
rect 87368 73412 87424 73468
rect 87424 73412 87428 73468
rect 87364 73408 87428 73412
rect 87444 73468 87508 73472
rect 87444 73412 87448 73468
rect 87448 73412 87504 73468
rect 87504 73412 87508 73468
rect 87444 73408 87508 73412
rect 87524 73468 87588 73472
rect 87524 73412 87528 73468
rect 87528 73412 87584 73468
rect 87584 73412 87588 73468
rect 87524 73408 87588 73412
rect 5956 72924 6020 72928
rect 5956 72868 5960 72924
rect 5960 72868 6016 72924
rect 6016 72868 6020 72924
rect 5956 72864 6020 72868
rect 6036 72924 6100 72928
rect 6036 72868 6040 72924
rect 6040 72868 6096 72924
rect 6096 72868 6100 72924
rect 6036 72864 6100 72868
rect 6116 72924 6180 72928
rect 6116 72868 6120 72924
rect 6120 72868 6176 72924
rect 6176 72868 6180 72924
rect 6116 72864 6180 72868
rect 6196 72924 6260 72928
rect 6196 72868 6200 72924
rect 6200 72868 6256 72924
rect 6256 72868 6260 72924
rect 6196 72864 6260 72868
rect 86548 72924 86612 72928
rect 86548 72868 86552 72924
rect 86552 72868 86608 72924
rect 86608 72868 86612 72924
rect 86548 72864 86612 72868
rect 86628 72924 86692 72928
rect 86628 72868 86632 72924
rect 86632 72868 86688 72924
rect 86688 72868 86692 72924
rect 86628 72864 86692 72868
rect 86708 72924 86772 72928
rect 86708 72868 86712 72924
rect 86712 72868 86768 72924
rect 86768 72868 86772 72924
rect 86708 72864 86772 72868
rect 86788 72924 86852 72928
rect 86788 72868 86792 72924
rect 86792 72868 86848 72924
rect 86848 72868 86852 72924
rect 86788 72864 86852 72868
rect 6692 72380 6756 72384
rect 6692 72324 6696 72380
rect 6696 72324 6752 72380
rect 6752 72324 6756 72380
rect 6692 72320 6756 72324
rect 6772 72380 6836 72384
rect 6772 72324 6776 72380
rect 6776 72324 6832 72380
rect 6832 72324 6836 72380
rect 6772 72320 6836 72324
rect 6852 72380 6916 72384
rect 6852 72324 6856 72380
rect 6856 72324 6912 72380
rect 6912 72324 6916 72380
rect 6852 72320 6916 72324
rect 6932 72380 6996 72384
rect 6932 72324 6936 72380
rect 6936 72324 6992 72380
rect 6992 72324 6996 72380
rect 6932 72320 6996 72324
rect 87284 72380 87348 72384
rect 87284 72324 87288 72380
rect 87288 72324 87344 72380
rect 87344 72324 87348 72380
rect 87284 72320 87348 72324
rect 87364 72380 87428 72384
rect 87364 72324 87368 72380
rect 87368 72324 87424 72380
rect 87424 72324 87428 72380
rect 87364 72320 87428 72324
rect 87444 72380 87508 72384
rect 87444 72324 87448 72380
rect 87448 72324 87504 72380
rect 87504 72324 87508 72380
rect 87444 72320 87508 72324
rect 87524 72380 87588 72384
rect 87524 72324 87528 72380
rect 87528 72324 87584 72380
rect 87584 72324 87588 72380
rect 87524 72320 87588 72324
rect 5956 71836 6020 71840
rect 5956 71780 5960 71836
rect 5960 71780 6016 71836
rect 6016 71780 6020 71836
rect 5956 71776 6020 71780
rect 6036 71836 6100 71840
rect 6036 71780 6040 71836
rect 6040 71780 6096 71836
rect 6096 71780 6100 71836
rect 6036 71776 6100 71780
rect 6116 71836 6180 71840
rect 6116 71780 6120 71836
rect 6120 71780 6176 71836
rect 6176 71780 6180 71836
rect 6116 71776 6180 71780
rect 6196 71836 6260 71840
rect 6196 71780 6200 71836
rect 6200 71780 6256 71836
rect 6256 71780 6260 71836
rect 6196 71776 6260 71780
rect 86548 71836 86612 71840
rect 86548 71780 86552 71836
rect 86552 71780 86608 71836
rect 86608 71780 86612 71836
rect 86548 71776 86612 71780
rect 86628 71836 86692 71840
rect 86628 71780 86632 71836
rect 86632 71780 86688 71836
rect 86688 71780 86692 71836
rect 86628 71776 86692 71780
rect 86708 71836 86772 71840
rect 86708 71780 86712 71836
rect 86712 71780 86768 71836
rect 86768 71780 86772 71836
rect 86708 71776 86772 71780
rect 86788 71836 86852 71840
rect 86788 71780 86792 71836
rect 86792 71780 86848 71836
rect 86848 71780 86852 71836
rect 86788 71776 86852 71780
rect 6692 71292 6756 71296
rect 6692 71236 6696 71292
rect 6696 71236 6752 71292
rect 6752 71236 6756 71292
rect 6692 71232 6756 71236
rect 6772 71292 6836 71296
rect 6772 71236 6776 71292
rect 6776 71236 6832 71292
rect 6832 71236 6836 71292
rect 6772 71232 6836 71236
rect 6852 71292 6916 71296
rect 6852 71236 6856 71292
rect 6856 71236 6912 71292
rect 6912 71236 6916 71292
rect 6852 71232 6916 71236
rect 6932 71292 6996 71296
rect 6932 71236 6936 71292
rect 6936 71236 6992 71292
rect 6992 71236 6996 71292
rect 6932 71232 6996 71236
rect 87284 71292 87348 71296
rect 87284 71236 87288 71292
rect 87288 71236 87344 71292
rect 87344 71236 87348 71292
rect 87284 71232 87348 71236
rect 87364 71292 87428 71296
rect 87364 71236 87368 71292
rect 87368 71236 87424 71292
rect 87424 71236 87428 71292
rect 87364 71232 87428 71236
rect 87444 71292 87508 71296
rect 87444 71236 87448 71292
rect 87448 71236 87504 71292
rect 87504 71236 87508 71292
rect 87444 71232 87508 71236
rect 87524 71292 87588 71296
rect 87524 71236 87528 71292
rect 87528 71236 87584 71292
rect 87584 71236 87588 71292
rect 87524 71232 87588 71236
rect 5956 70748 6020 70752
rect 5956 70692 5960 70748
rect 5960 70692 6016 70748
rect 6016 70692 6020 70748
rect 5956 70688 6020 70692
rect 6036 70748 6100 70752
rect 6036 70692 6040 70748
rect 6040 70692 6096 70748
rect 6096 70692 6100 70748
rect 6036 70688 6100 70692
rect 6116 70748 6180 70752
rect 6116 70692 6120 70748
rect 6120 70692 6176 70748
rect 6176 70692 6180 70748
rect 6116 70688 6180 70692
rect 6196 70748 6260 70752
rect 6196 70692 6200 70748
rect 6200 70692 6256 70748
rect 6256 70692 6260 70748
rect 6196 70688 6260 70692
rect 86548 70748 86612 70752
rect 86548 70692 86552 70748
rect 86552 70692 86608 70748
rect 86608 70692 86612 70748
rect 86548 70688 86612 70692
rect 86628 70748 86692 70752
rect 86628 70692 86632 70748
rect 86632 70692 86688 70748
rect 86688 70692 86692 70748
rect 86628 70688 86692 70692
rect 86708 70748 86772 70752
rect 86708 70692 86712 70748
rect 86712 70692 86768 70748
rect 86768 70692 86772 70748
rect 86708 70688 86772 70692
rect 86788 70748 86852 70752
rect 86788 70692 86792 70748
rect 86792 70692 86848 70748
rect 86848 70692 86852 70748
rect 86788 70688 86852 70692
rect 6692 70204 6756 70208
rect 6692 70148 6696 70204
rect 6696 70148 6752 70204
rect 6752 70148 6756 70204
rect 6692 70144 6756 70148
rect 6772 70204 6836 70208
rect 6772 70148 6776 70204
rect 6776 70148 6832 70204
rect 6832 70148 6836 70204
rect 6772 70144 6836 70148
rect 6852 70204 6916 70208
rect 6852 70148 6856 70204
rect 6856 70148 6912 70204
rect 6912 70148 6916 70204
rect 6852 70144 6916 70148
rect 6932 70204 6996 70208
rect 6932 70148 6936 70204
rect 6936 70148 6992 70204
rect 6992 70148 6996 70204
rect 6932 70144 6996 70148
rect 87284 70204 87348 70208
rect 87284 70148 87288 70204
rect 87288 70148 87344 70204
rect 87344 70148 87348 70204
rect 87284 70144 87348 70148
rect 87364 70204 87428 70208
rect 87364 70148 87368 70204
rect 87368 70148 87424 70204
rect 87424 70148 87428 70204
rect 87364 70144 87428 70148
rect 87444 70204 87508 70208
rect 87444 70148 87448 70204
rect 87448 70148 87504 70204
rect 87504 70148 87508 70204
rect 87444 70144 87508 70148
rect 87524 70204 87588 70208
rect 87524 70148 87528 70204
rect 87528 70148 87584 70204
rect 87584 70148 87588 70204
rect 87524 70144 87588 70148
rect 5956 69660 6020 69664
rect 5956 69604 5960 69660
rect 5960 69604 6016 69660
rect 6016 69604 6020 69660
rect 5956 69600 6020 69604
rect 6036 69660 6100 69664
rect 6036 69604 6040 69660
rect 6040 69604 6096 69660
rect 6096 69604 6100 69660
rect 6036 69600 6100 69604
rect 6116 69660 6180 69664
rect 6116 69604 6120 69660
rect 6120 69604 6176 69660
rect 6176 69604 6180 69660
rect 6116 69600 6180 69604
rect 6196 69660 6260 69664
rect 6196 69604 6200 69660
rect 6200 69604 6256 69660
rect 6256 69604 6260 69660
rect 6196 69600 6260 69604
rect 86548 69660 86612 69664
rect 86548 69604 86552 69660
rect 86552 69604 86608 69660
rect 86608 69604 86612 69660
rect 86548 69600 86612 69604
rect 86628 69660 86692 69664
rect 86628 69604 86632 69660
rect 86632 69604 86688 69660
rect 86688 69604 86692 69660
rect 86628 69600 86692 69604
rect 86708 69660 86772 69664
rect 86708 69604 86712 69660
rect 86712 69604 86768 69660
rect 86768 69604 86772 69660
rect 86708 69600 86772 69604
rect 86788 69660 86852 69664
rect 86788 69604 86792 69660
rect 86792 69604 86848 69660
rect 86848 69604 86852 69660
rect 86788 69600 86852 69604
rect 6692 69116 6756 69120
rect 6692 69060 6696 69116
rect 6696 69060 6752 69116
rect 6752 69060 6756 69116
rect 6692 69056 6756 69060
rect 6772 69116 6836 69120
rect 6772 69060 6776 69116
rect 6776 69060 6832 69116
rect 6832 69060 6836 69116
rect 6772 69056 6836 69060
rect 6852 69116 6916 69120
rect 6852 69060 6856 69116
rect 6856 69060 6912 69116
rect 6912 69060 6916 69116
rect 6852 69056 6916 69060
rect 6932 69116 6996 69120
rect 6932 69060 6936 69116
rect 6936 69060 6992 69116
rect 6992 69060 6996 69116
rect 6932 69056 6996 69060
rect 87284 69116 87348 69120
rect 87284 69060 87288 69116
rect 87288 69060 87344 69116
rect 87344 69060 87348 69116
rect 87284 69056 87348 69060
rect 87364 69116 87428 69120
rect 87364 69060 87368 69116
rect 87368 69060 87424 69116
rect 87424 69060 87428 69116
rect 87364 69056 87428 69060
rect 87444 69116 87508 69120
rect 87444 69060 87448 69116
rect 87448 69060 87504 69116
rect 87504 69060 87508 69116
rect 87444 69056 87508 69060
rect 87524 69116 87588 69120
rect 87524 69060 87528 69116
rect 87528 69060 87584 69116
rect 87584 69060 87588 69116
rect 87524 69056 87588 69060
rect 5956 68572 6020 68576
rect 5956 68516 5960 68572
rect 5960 68516 6016 68572
rect 6016 68516 6020 68572
rect 5956 68512 6020 68516
rect 6036 68572 6100 68576
rect 6036 68516 6040 68572
rect 6040 68516 6096 68572
rect 6096 68516 6100 68572
rect 6036 68512 6100 68516
rect 6116 68572 6180 68576
rect 6116 68516 6120 68572
rect 6120 68516 6176 68572
rect 6176 68516 6180 68572
rect 6116 68512 6180 68516
rect 6196 68572 6260 68576
rect 6196 68516 6200 68572
rect 6200 68516 6256 68572
rect 6256 68516 6260 68572
rect 6196 68512 6260 68516
rect 86548 68572 86612 68576
rect 86548 68516 86552 68572
rect 86552 68516 86608 68572
rect 86608 68516 86612 68572
rect 86548 68512 86612 68516
rect 86628 68572 86692 68576
rect 86628 68516 86632 68572
rect 86632 68516 86688 68572
rect 86688 68516 86692 68572
rect 86628 68512 86692 68516
rect 86708 68572 86772 68576
rect 86708 68516 86712 68572
rect 86712 68516 86768 68572
rect 86768 68516 86772 68572
rect 86708 68512 86772 68516
rect 86788 68572 86852 68576
rect 86788 68516 86792 68572
rect 86792 68516 86848 68572
rect 86848 68516 86852 68572
rect 86788 68512 86852 68516
rect 6692 68028 6756 68032
rect 6692 67972 6696 68028
rect 6696 67972 6752 68028
rect 6752 67972 6756 68028
rect 6692 67968 6756 67972
rect 6772 68028 6836 68032
rect 6772 67972 6776 68028
rect 6776 67972 6832 68028
rect 6832 67972 6836 68028
rect 6772 67968 6836 67972
rect 6852 68028 6916 68032
rect 6852 67972 6856 68028
rect 6856 67972 6912 68028
rect 6912 67972 6916 68028
rect 6852 67968 6916 67972
rect 6932 68028 6996 68032
rect 6932 67972 6936 68028
rect 6936 67972 6992 68028
rect 6992 67972 6996 68028
rect 6932 67968 6996 67972
rect 87284 68028 87348 68032
rect 87284 67972 87288 68028
rect 87288 67972 87344 68028
rect 87344 67972 87348 68028
rect 87284 67968 87348 67972
rect 87364 68028 87428 68032
rect 87364 67972 87368 68028
rect 87368 67972 87424 68028
rect 87424 67972 87428 68028
rect 87364 67968 87428 67972
rect 87444 68028 87508 68032
rect 87444 67972 87448 68028
rect 87448 67972 87504 68028
rect 87504 67972 87508 68028
rect 87444 67968 87508 67972
rect 87524 68028 87588 68032
rect 87524 67972 87528 68028
rect 87528 67972 87584 68028
rect 87584 67972 87588 68028
rect 87524 67968 87588 67972
rect 5956 67484 6020 67488
rect 5956 67428 5960 67484
rect 5960 67428 6016 67484
rect 6016 67428 6020 67484
rect 5956 67424 6020 67428
rect 6036 67484 6100 67488
rect 6036 67428 6040 67484
rect 6040 67428 6096 67484
rect 6096 67428 6100 67484
rect 6036 67424 6100 67428
rect 6116 67484 6180 67488
rect 6116 67428 6120 67484
rect 6120 67428 6176 67484
rect 6176 67428 6180 67484
rect 6116 67424 6180 67428
rect 6196 67484 6260 67488
rect 6196 67428 6200 67484
rect 6200 67428 6256 67484
rect 6256 67428 6260 67484
rect 6196 67424 6260 67428
rect 86548 67484 86612 67488
rect 86548 67428 86552 67484
rect 86552 67428 86608 67484
rect 86608 67428 86612 67484
rect 86548 67424 86612 67428
rect 86628 67484 86692 67488
rect 86628 67428 86632 67484
rect 86632 67428 86688 67484
rect 86688 67428 86692 67484
rect 86628 67424 86692 67428
rect 86708 67484 86772 67488
rect 86708 67428 86712 67484
rect 86712 67428 86768 67484
rect 86768 67428 86772 67484
rect 86708 67424 86772 67428
rect 86788 67484 86852 67488
rect 86788 67428 86792 67484
rect 86792 67428 86848 67484
rect 86848 67428 86852 67484
rect 86788 67424 86852 67428
rect 6692 66940 6756 66944
rect 6692 66884 6696 66940
rect 6696 66884 6752 66940
rect 6752 66884 6756 66940
rect 6692 66880 6756 66884
rect 6772 66940 6836 66944
rect 6772 66884 6776 66940
rect 6776 66884 6832 66940
rect 6832 66884 6836 66940
rect 6772 66880 6836 66884
rect 6852 66940 6916 66944
rect 6852 66884 6856 66940
rect 6856 66884 6912 66940
rect 6912 66884 6916 66940
rect 6852 66880 6916 66884
rect 6932 66940 6996 66944
rect 6932 66884 6936 66940
rect 6936 66884 6992 66940
rect 6992 66884 6996 66940
rect 6932 66880 6996 66884
rect 87284 66940 87348 66944
rect 87284 66884 87288 66940
rect 87288 66884 87344 66940
rect 87344 66884 87348 66940
rect 87284 66880 87348 66884
rect 87364 66940 87428 66944
rect 87364 66884 87368 66940
rect 87368 66884 87424 66940
rect 87424 66884 87428 66940
rect 87364 66880 87428 66884
rect 87444 66940 87508 66944
rect 87444 66884 87448 66940
rect 87448 66884 87504 66940
rect 87504 66884 87508 66940
rect 87444 66880 87508 66884
rect 87524 66940 87588 66944
rect 87524 66884 87528 66940
rect 87528 66884 87584 66940
rect 87584 66884 87588 66940
rect 87524 66880 87588 66884
rect 5956 66396 6020 66400
rect 5956 66340 5960 66396
rect 5960 66340 6016 66396
rect 6016 66340 6020 66396
rect 5956 66336 6020 66340
rect 6036 66396 6100 66400
rect 6036 66340 6040 66396
rect 6040 66340 6096 66396
rect 6096 66340 6100 66396
rect 6036 66336 6100 66340
rect 6116 66396 6180 66400
rect 6116 66340 6120 66396
rect 6120 66340 6176 66396
rect 6176 66340 6180 66396
rect 6116 66336 6180 66340
rect 6196 66396 6260 66400
rect 6196 66340 6200 66396
rect 6200 66340 6256 66396
rect 6256 66340 6260 66396
rect 6196 66336 6260 66340
rect 86548 66396 86612 66400
rect 86548 66340 86552 66396
rect 86552 66340 86608 66396
rect 86608 66340 86612 66396
rect 86548 66336 86612 66340
rect 86628 66396 86692 66400
rect 86628 66340 86632 66396
rect 86632 66340 86688 66396
rect 86688 66340 86692 66396
rect 86628 66336 86692 66340
rect 86708 66396 86772 66400
rect 86708 66340 86712 66396
rect 86712 66340 86768 66396
rect 86768 66340 86772 66396
rect 86708 66336 86772 66340
rect 86788 66396 86852 66400
rect 86788 66340 86792 66396
rect 86792 66340 86848 66396
rect 86848 66340 86852 66396
rect 86788 66336 86852 66340
rect 6692 65852 6756 65856
rect 6692 65796 6696 65852
rect 6696 65796 6752 65852
rect 6752 65796 6756 65852
rect 6692 65792 6756 65796
rect 6772 65852 6836 65856
rect 6772 65796 6776 65852
rect 6776 65796 6832 65852
rect 6832 65796 6836 65852
rect 6772 65792 6836 65796
rect 6852 65852 6916 65856
rect 6852 65796 6856 65852
rect 6856 65796 6912 65852
rect 6912 65796 6916 65852
rect 6852 65792 6916 65796
rect 6932 65852 6996 65856
rect 6932 65796 6936 65852
rect 6936 65796 6992 65852
rect 6992 65796 6996 65852
rect 6932 65792 6996 65796
rect 87284 65852 87348 65856
rect 87284 65796 87288 65852
rect 87288 65796 87344 65852
rect 87344 65796 87348 65852
rect 87284 65792 87348 65796
rect 87364 65852 87428 65856
rect 87364 65796 87368 65852
rect 87368 65796 87424 65852
rect 87424 65796 87428 65852
rect 87364 65792 87428 65796
rect 87444 65852 87508 65856
rect 87444 65796 87448 65852
rect 87448 65796 87504 65852
rect 87504 65796 87508 65852
rect 87444 65792 87508 65796
rect 87524 65852 87588 65856
rect 87524 65796 87528 65852
rect 87528 65796 87584 65852
rect 87584 65796 87588 65852
rect 87524 65792 87588 65796
rect 5956 65308 6020 65312
rect 5956 65252 5960 65308
rect 5960 65252 6016 65308
rect 6016 65252 6020 65308
rect 5956 65248 6020 65252
rect 6036 65308 6100 65312
rect 6036 65252 6040 65308
rect 6040 65252 6096 65308
rect 6096 65252 6100 65308
rect 6036 65248 6100 65252
rect 6116 65308 6180 65312
rect 6116 65252 6120 65308
rect 6120 65252 6176 65308
rect 6176 65252 6180 65308
rect 6116 65248 6180 65252
rect 6196 65308 6260 65312
rect 6196 65252 6200 65308
rect 6200 65252 6256 65308
rect 6256 65252 6260 65308
rect 6196 65248 6260 65252
rect 86548 65308 86612 65312
rect 86548 65252 86552 65308
rect 86552 65252 86608 65308
rect 86608 65252 86612 65308
rect 86548 65248 86612 65252
rect 86628 65308 86692 65312
rect 86628 65252 86632 65308
rect 86632 65252 86688 65308
rect 86688 65252 86692 65308
rect 86628 65248 86692 65252
rect 86708 65308 86772 65312
rect 86708 65252 86712 65308
rect 86712 65252 86768 65308
rect 86768 65252 86772 65308
rect 86708 65248 86772 65252
rect 86788 65308 86852 65312
rect 86788 65252 86792 65308
rect 86792 65252 86848 65308
rect 86848 65252 86852 65308
rect 86788 65248 86852 65252
rect 6692 64764 6756 64768
rect 6692 64708 6696 64764
rect 6696 64708 6752 64764
rect 6752 64708 6756 64764
rect 6692 64704 6756 64708
rect 6772 64764 6836 64768
rect 6772 64708 6776 64764
rect 6776 64708 6832 64764
rect 6832 64708 6836 64764
rect 6772 64704 6836 64708
rect 6852 64764 6916 64768
rect 6852 64708 6856 64764
rect 6856 64708 6912 64764
rect 6912 64708 6916 64764
rect 6852 64704 6916 64708
rect 6932 64764 6996 64768
rect 6932 64708 6936 64764
rect 6936 64708 6992 64764
rect 6992 64708 6996 64764
rect 6932 64704 6996 64708
rect 87284 64764 87348 64768
rect 87284 64708 87288 64764
rect 87288 64708 87344 64764
rect 87344 64708 87348 64764
rect 87284 64704 87348 64708
rect 87364 64764 87428 64768
rect 87364 64708 87368 64764
rect 87368 64708 87424 64764
rect 87424 64708 87428 64764
rect 87364 64704 87428 64708
rect 87444 64764 87508 64768
rect 87444 64708 87448 64764
rect 87448 64708 87504 64764
rect 87504 64708 87508 64764
rect 87444 64704 87508 64708
rect 87524 64764 87588 64768
rect 87524 64708 87528 64764
rect 87528 64708 87584 64764
rect 87584 64708 87588 64764
rect 87524 64704 87588 64708
rect 5956 64220 6020 64224
rect 5956 64164 5960 64220
rect 5960 64164 6016 64220
rect 6016 64164 6020 64220
rect 5956 64160 6020 64164
rect 6036 64220 6100 64224
rect 6036 64164 6040 64220
rect 6040 64164 6096 64220
rect 6096 64164 6100 64220
rect 6036 64160 6100 64164
rect 6116 64220 6180 64224
rect 6116 64164 6120 64220
rect 6120 64164 6176 64220
rect 6176 64164 6180 64220
rect 6116 64160 6180 64164
rect 6196 64220 6260 64224
rect 6196 64164 6200 64220
rect 6200 64164 6256 64220
rect 6256 64164 6260 64220
rect 6196 64160 6260 64164
rect 86548 64220 86612 64224
rect 86548 64164 86552 64220
rect 86552 64164 86608 64220
rect 86608 64164 86612 64220
rect 86548 64160 86612 64164
rect 86628 64220 86692 64224
rect 86628 64164 86632 64220
rect 86632 64164 86688 64220
rect 86688 64164 86692 64220
rect 86628 64160 86692 64164
rect 86708 64220 86772 64224
rect 86708 64164 86712 64220
rect 86712 64164 86768 64220
rect 86768 64164 86772 64220
rect 86708 64160 86772 64164
rect 86788 64220 86852 64224
rect 86788 64164 86792 64220
rect 86792 64164 86848 64220
rect 86848 64164 86852 64220
rect 86788 64160 86852 64164
rect 6692 63676 6756 63680
rect 6692 63620 6696 63676
rect 6696 63620 6752 63676
rect 6752 63620 6756 63676
rect 6692 63616 6756 63620
rect 6772 63676 6836 63680
rect 6772 63620 6776 63676
rect 6776 63620 6832 63676
rect 6832 63620 6836 63676
rect 6772 63616 6836 63620
rect 6852 63676 6916 63680
rect 6852 63620 6856 63676
rect 6856 63620 6912 63676
rect 6912 63620 6916 63676
rect 6852 63616 6916 63620
rect 6932 63676 6996 63680
rect 6932 63620 6936 63676
rect 6936 63620 6992 63676
rect 6992 63620 6996 63676
rect 6932 63616 6996 63620
rect 87284 63676 87348 63680
rect 87284 63620 87288 63676
rect 87288 63620 87344 63676
rect 87344 63620 87348 63676
rect 87284 63616 87348 63620
rect 87364 63676 87428 63680
rect 87364 63620 87368 63676
rect 87368 63620 87424 63676
rect 87424 63620 87428 63676
rect 87364 63616 87428 63620
rect 87444 63676 87508 63680
rect 87444 63620 87448 63676
rect 87448 63620 87504 63676
rect 87504 63620 87508 63676
rect 87444 63616 87508 63620
rect 87524 63676 87588 63680
rect 87524 63620 87528 63676
rect 87528 63620 87584 63676
rect 87584 63620 87588 63676
rect 87524 63616 87588 63620
rect 5956 63132 6020 63136
rect 5956 63076 5960 63132
rect 5960 63076 6016 63132
rect 6016 63076 6020 63132
rect 5956 63072 6020 63076
rect 6036 63132 6100 63136
rect 6036 63076 6040 63132
rect 6040 63076 6096 63132
rect 6096 63076 6100 63132
rect 6036 63072 6100 63076
rect 6116 63132 6180 63136
rect 6116 63076 6120 63132
rect 6120 63076 6176 63132
rect 6176 63076 6180 63132
rect 6116 63072 6180 63076
rect 6196 63132 6260 63136
rect 6196 63076 6200 63132
rect 6200 63076 6256 63132
rect 6256 63076 6260 63132
rect 6196 63072 6260 63076
rect 86548 63132 86612 63136
rect 86548 63076 86552 63132
rect 86552 63076 86608 63132
rect 86608 63076 86612 63132
rect 86548 63072 86612 63076
rect 86628 63132 86692 63136
rect 86628 63076 86632 63132
rect 86632 63076 86688 63132
rect 86688 63076 86692 63132
rect 86628 63072 86692 63076
rect 86708 63132 86772 63136
rect 86708 63076 86712 63132
rect 86712 63076 86768 63132
rect 86768 63076 86772 63132
rect 86708 63072 86772 63076
rect 86788 63132 86852 63136
rect 86788 63076 86792 63132
rect 86792 63076 86848 63132
rect 86848 63076 86852 63132
rect 86788 63072 86852 63076
rect 6692 62588 6756 62592
rect 6692 62532 6696 62588
rect 6696 62532 6752 62588
rect 6752 62532 6756 62588
rect 6692 62528 6756 62532
rect 6772 62588 6836 62592
rect 6772 62532 6776 62588
rect 6776 62532 6832 62588
rect 6832 62532 6836 62588
rect 6772 62528 6836 62532
rect 6852 62588 6916 62592
rect 6852 62532 6856 62588
rect 6856 62532 6912 62588
rect 6912 62532 6916 62588
rect 6852 62528 6916 62532
rect 6932 62588 6996 62592
rect 6932 62532 6936 62588
rect 6936 62532 6992 62588
rect 6992 62532 6996 62588
rect 6932 62528 6996 62532
rect 87284 62588 87348 62592
rect 87284 62532 87288 62588
rect 87288 62532 87344 62588
rect 87344 62532 87348 62588
rect 87284 62528 87348 62532
rect 87364 62588 87428 62592
rect 87364 62532 87368 62588
rect 87368 62532 87424 62588
rect 87424 62532 87428 62588
rect 87364 62528 87428 62532
rect 87444 62588 87508 62592
rect 87444 62532 87448 62588
rect 87448 62532 87504 62588
rect 87504 62532 87508 62588
rect 87444 62528 87508 62532
rect 87524 62588 87588 62592
rect 87524 62532 87528 62588
rect 87528 62532 87584 62588
rect 87584 62532 87588 62588
rect 87524 62528 87588 62532
rect 5956 62044 6020 62048
rect 5956 61988 5960 62044
rect 5960 61988 6016 62044
rect 6016 61988 6020 62044
rect 5956 61984 6020 61988
rect 6036 62044 6100 62048
rect 6036 61988 6040 62044
rect 6040 61988 6096 62044
rect 6096 61988 6100 62044
rect 6036 61984 6100 61988
rect 6116 62044 6180 62048
rect 6116 61988 6120 62044
rect 6120 61988 6176 62044
rect 6176 61988 6180 62044
rect 6116 61984 6180 61988
rect 6196 62044 6260 62048
rect 6196 61988 6200 62044
rect 6200 61988 6256 62044
rect 6256 61988 6260 62044
rect 6196 61984 6260 61988
rect 86548 62044 86612 62048
rect 86548 61988 86552 62044
rect 86552 61988 86608 62044
rect 86608 61988 86612 62044
rect 86548 61984 86612 61988
rect 86628 62044 86692 62048
rect 86628 61988 86632 62044
rect 86632 61988 86688 62044
rect 86688 61988 86692 62044
rect 86628 61984 86692 61988
rect 86708 62044 86772 62048
rect 86708 61988 86712 62044
rect 86712 61988 86768 62044
rect 86768 61988 86772 62044
rect 86708 61984 86772 61988
rect 86788 62044 86852 62048
rect 86788 61988 86792 62044
rect 86792 61988 86848 62044
rect 86848 61988 86852 62044
rect 86788 61984 86852 61988
rect 6692 61500 6756 61504
rect 6692 61444 6696 61500
rect 6696 61444 6752 61500
rect 6752 61444 6756 61500
rect 6692 61440 6756 61444
rect 6772 61500 6836 61504
rect 6772 61444 6776 61500
rect 6776 61444 6832 61500
rect 6832 61444 6836 61500
rect 6772 61440 6836 61444
rect 6852 61500 6916 61504
rect 6852 61444 6856 61500
rect 6856 61444 6912 61500
rect 6912 61444 6916 61500
rect 6852 61440 6916 61444
rect 6932 61500 6996 61504
rect 6932 61444 6936 61500
rect 6936 61444 6992 61500
rect 6992 61444 6996 61500
rect 6932 61440 6996 61444
rect 87284 61500 87348 61504
rect 87284 61444 87288 61500
rect 87288 61444 87344 61500
rect 87344 61444 87348 61500
rect 87284 61440 87348 61444
rect 87364 61500 87428 61504
rect 87364 61444 87368 61500
rect 87368 61444 87424 61500
rect 87424 61444 87428 61500
rect 87364 61440 87428 61444
rect 87444 61500 87508 61504
rect 87444 61444 87448 61500
rect 87448 61444 87504 61500
rect 87504 61444 87508 61500
rect 87444 61440 87508 61444
rect 87524 61500 87588 61504
rect 87524 61444 87528 61500
rect 87528 61444 87584 61500
rect 87584 61444 87588 61500
rect 87524 61440 87588 61444
rect 5956 60956 6020 60960
rect 5956 60900 5960 60956
rect 5960 60900 6016 60956
rect 6016 60900 6020 60956
rect 5956 60896 6020 60900
rect 6036 60956 6100 60960
rect 6036 60900 6040 60956
rect 6040 60900 6096 60956
rect 6096 60900 6100 60956
rect 6036 60896 6100 60900
rect 6116 60956 6180 60960
rect 6116 60900 6120 60956
rect 6120 60900 6176 60956
rect 6176 60900 6180 60956
rect 6116 60896 6180 60900
rect 6196 60956 6260 60960
rect 6196 60900 6200 60956
rect 6200 60900 6256 60956
rect 6256 60900 6260 60956
rect 6196 60896 6260 60900
rect 86548 60956 86612 60960
rect 86548 60900 86552 60956
rect 86552 60900 86608 60956
rect 86608 60900 86612 60956
rect 86548 60896 86612 60900
rect 86628 60956 86692 60960
rect 86628 60900 86632 60956
rect 86632 60900 86688 60956
rect 86688 60900 86692 60956
rect 86628 60896 86692 60900
rect 86708 60956 86772 60960
rect 86708 60900 86712 60956
rect 86712 60900 86768 60956
rect 86768 60900 86772 60956
rect 86708 60896 86772 60900
rect 86788 60956 86852 60960
rect 86788 60900 86792 60956
rect 86792 60900 86848 60956
rect 86848 60900 86852 60956
rect 86788 60896 86852 60900
rect 6692 60412 6756 60416
rect 6692 60356 6696 60412
rect 6696 60356 6752 60412
rect 6752 60356 6756 60412
rect 6692 60352 6756 60356
rect 6772 60412 6836 60416
rect 6772 60356 6776 60412
rect 6776 60356 6832 60412
rect 6832 60356 6836 60412
rect 6772 60352 6836 60356
rect 6852 60412 6916 60416
rect 6852 60356 6856 60412
rect 6856 60356 6912 60412
rect 6912 60356 6916 60412
rect 6852 60352 6916 60356
rect 6932 60412 6996 60416
rect 6932 60356 6936 60412
rect 6936 60356 6992 60412
rect 6992 60356 6996 60412
rect 6932 60352 6996 60356
rect 87284 60412 87348 60416
rect 87284 60356 87288 60412
rect 87288 60356 87344 60412
rect 87344 60356 87348 60412
rect 87284 60352 87348 60356
rect 87364 60412 87428 60416
rect 87364 60356 87368 60412
rect 87368 60356 87424 60412
rect 87424 60356 87428 60412
rect 87364 60352 87428 60356
rect 87444 60412 87508 60416
rect 87444 60356 87448 60412
rect 87448 60356 87504 60412
rect 87504 60356 87508 60412
rect 87444 60352 87508 60356
rect 87524 60412 87588 60416
rect 87524 60356 87528 60412
rect 87528 60356 87584 60412
rect 87584 60356 87588 60412
rect 87524 60352 87588 60356
rect 5956 59868 6020 59872
rect 5956 59812 5960 59868
rect 5960 59812 6016 59868
rect 6016 59812 6020 59868
rect 5956 59808 6020 59812
rect 6036 59868 6100 59872
rect 6036 59812 6040 59868
rect 6040 59812 6096 59868
rect 6096 59812 6100 59868
rect 6036 59808 6100 59812
rect 6116 59868 6180 59872
rect 6116 59812 6120 59868
rect 6120 59812 6176 59868
rect 6176 59812 6180 59868
rect 6116 59808 6180 59812
rect 6196 59868 6260 59872
rect 6196 59812 6200 59868
rect 6200 59812 6256 59868
rect 6256 59812 6260 59868
rect 6196 59808 6260 59812
rect 86548 59868 86612 59872
rect 86548 59812 86552 59868
rect 86552 59812 86608 59868
rect 86608 59812 86612 59868
rect 86548 59808 86612 59812
rect 86628 59868 86692 59872
rect 86628 59812 86632 59868
rect 86632 59812 86688 59868
rect 86688 59812 86692 59868
rect 86628 59808 86692 59812
rect 86708 59868 86772 59872
rect 86708 59812 86712 59868
rect 86712 59812 86768 59868
rect 86768 59812 86772 59868
rect 86708 59808 86772 59812
rect 86788 59868 86852 59872
rect 86788 59812 86792 59868
rect 86792 59812 86848 59868
rect 86848 59812 86852 59868
rect 86788 59808 86852 59812
rect 6692 59324 6756 59328
rect 6692 59268 6696 59324
rect 6696 59268 6752 59324
rect 6752 59268 6756 59324
rect 6692 59264 6756 59268
rect 6772 59324 6836 59328
rect 6772 59268 6776 59324
rect 6776 59268 6832 59324
rect 6832 59268 6836 59324
rect 6772 59264 6836 59268
rect 6852 59324 6916 59328
rect 6852 59268 6856 59324
rect 6856 59268 6912 59324
rect 6912 59268 6916 59324
rect 6852 59264 6916 59268
rect 6932 59324 6996 59328
rect 6932 59268 6936 59324
rect 6936 59268 6992 59324
rect 6992 59268 6996 59324
rect 6932 59264 6996 59268
rect 87284 59324 87348 59328
rect 87284 59268 87288 59324
rect 87288 59268 87344 59324
rect 87344 59268 87348 59324
rect 87284 59264 87348 59268
rect 87364 59324 87428 59328
rect 87364 59268 87368 59324
rect 87368 59268 87424 59324
rect 87424 59268 87428 59324
rect 87364 59264 87428 59268
rect 87444 59324 87508 59328
rect 87444 59268 87448 59324
rect 87448 59268 87504 59324
rect 87504 59268 87508 59324
rect 87444 59264 87508 59268
rect 87524 59324 87588 59328
rect 87524 59268 87528 59324
rect 87528 59268 87584 59324
rect 87584 59268 87588 59324
rect 87524 59264 87588 59268
rect 5956 58780 6020 58784
rect 5956 58724 5960 58780
rect 5960 58724 6016 58780
rect 6016 58724 6020 58780
rect 5956 58720 6020 58724
rect 6036 58780 6100 58784
rect 6036 58724 6040 58780
rect 6040 58724 6096 58780
rect 6096 58724 6100 58780
rect 6036 58720 6100 58724
rect 6116 58780 6180 58784
rect 6116 58724 6120 58780
rect 6120 58724 6176 58780
rect 6176 58724 6180 58780
rect 6116 58720 6180 58724
rect 6196 58780 6260 58784
rect 6196 58724 6200 58780
rect 6200 58724 6256 58780
rect 6256 58724 6260 58780
rect 6196 58720 6260 58724
rect 86548 58780 86612 58784
rect 86548 58724 86552 58780
rect 86552 58724 86608 58780
rect 86608 58724 86612 58780
rect 86548 58720 86612 58724
rect 86628 58780 86692 58784
rect 86628 58724 86632 58780
rect 86632 58724 86688 58780
rect 86688 58724 86692 58780
rect 86628 58720 86692 58724
rect 86708 58780 86772 58784
rect 86708 58724 86712 58780
rect 86712 58724 86768 58780
rect 86768 58724 86772 58780
rect 86708 58720 86772 58724
rect 86788 58780 86852 58784
rect 86788 58724 86792 58780
rect 86792 58724 86848 58780
rect 86848 58724 86852 58780
rect 86788 58720 86852 58724
rect 6692 58236 6756 58240
rect 6692 58180 6696 58236
rect 6696 58180 6752 58236
rect 6752 58180 6756 58236
rect 6692 58176 6756 58180
rect 6772 58236 6836 58240
rect 6772 58180 6776 58236
rect 6776 58180 6832 58236
rect 6832 58180 6836 58236
rect 6772 58176 6836 58180
rect 6852 58236 6916 58240
rect 6852 58180 6856 58236
rect 6856 58180 6912 58236
rect 6912 58180 6916 58236
rect 6852 58176 6916 58180
rect 6932 58236 6996 58240
rect 6932 58180 6936 58236
rect 6936 58180 6992 58236
rect 6992 58180 6996 58236
rect 6932 58176 6996 58180
rect 87284 58236 87348 58240
rect 87284 58180 87288 58236
rect 87288 58180 87344 58236
rect 87344 58180 87348 58236
rect 87284 58176 87348 58180
rect 87364 58236 87428 58240
rect 87364 58180 87368 58236
rect 87368 58180 87424 58236
rect 87424 58180 87428 58236
rect 87364 58176 87428 58180
rect 87444 58236 87508 58240
rect 87444 58180 87448 58236
rect 87448 58180 87504 58236
rect 87504 58180 87508 58236
rect 87444 58176 87508 58180
rect 87524 58236 87588 58240
rect 87524 58180 87528 58236
rect 87528 58180 87584 58236
rect 87584 58180 87588 58236
rect 87524 58176 87588 58180
rect 5956 57692 6020 57696
rect 5956 57636 5960 57692
rect 5960 57636 6016 57692
rect 6016 57636 6020 57692
rect 5956 57632 6020 57636
rect 6036 57692 6100 57696
rect 6036 57636 6040 57692
rect 6040 57636 6096 57692
rect 6096 57636 6100 57692
rect 6036 57632 6100 57636
rect 6116 57692 6180 57696
rect 6116 57636 6120 57692
rect 6120 57636 6176 57692
rect 6176 57636 6180 57692
rect 6116 57632 6180 57636
rect 6196 57692 6260 57696
rect 6196 57636 6200 57692
rect 6200 57636 6256 57692
rect 6256 57636 6260 57692
rect 6196 57632 6260 57636
rect 86548 57692 86612 57696
rect 86548 57636 86552 57692
rect 86552 57636 86608 57692
rect 86608 57636 86612 57692
rect 86548 57632 86612 57636
rect 86628 57692 86692 57696
rect 86628 57636 86632 57692
rect 86632 57636 86688 57692
rect 86688 57636 86692 57692
rect 86628 57632 86692 57636
rect 86708 57692 86772 57696
rect 86708 57636 86712 57692
rect 86712 57636 86768 57692
rect 86768 57636 86772 57692
rect 86708 57632 86772 57636
rect 86788 57692 86852 57696
rect 86788 57636 86792 57692
rect 86792 57636 86848 57692
rect 86848 57636 86852 57692
rect 86788 57632 86852 57636
rect 6692 57148 6756 57152
rect 6692 57092 6696 57148
rect 6696 57092 6752 57148
rect 6752 57092 6756 57148
rect 6692 57088 6756 57092
rect 6772 57148 6836 57152
rect 6772 57092 6776 57148
rect 6776 57092 6832 57148
rect 6832 57092 6836 57148
rect 6772 57088 6836 57092
rect 6852 57148 6916 57152
rect 6852 57092 6856 57148
rect 6856 57092 6912 57148
rect 6912 57092 6916 57148
rect 6852 57088 6916 57092
rect 6932 57148 6996 57152
rect 6932 57092 6936 57148
rect 6936 57092 6992 57148
rect 6992 57092 6996 57148
rect 6932 57088 6996 57092
rect 87284 57148 87348 57152
rect 87284 57092 87288 57148
rect 87288 57092 87344 57148
rect 87344 57092 87348 57148
rect 87284 57088 87348 57092
rect 87364 57148 87428 57152
rect 87364 57092 87368 57148
rect 87368 57092 87424 57148
rect 87424 57092 87428 57148
rect 87364 57088 87428 57092
rect 87444 57148 87508 57152
rect 87444 57092 87448 57148
rect 87448 57092 87504 57148
rect 87504 57092 87508 57148
rect 87444 57088 87508 57092
rect 87524 57148 87588 57152
rect 87524 57092 87528 57148
rect 87528 57092 87584 57148
rect 87584 57092 87588 57148
rect 87524 57088 87588 57092
rect 5956 56604 6020 56608
rect 5956 56548 5960 56604
rect 5960 56548 6016 56604
rect 6016 56548 6020 56604
rect 5956 56544 6020 56548
rect 6036 56604 6100 56608
rect 6036 56548 6040 56604
rect 6040 56548 6096 56604
rect 6096 56548 6100 56604
rect 6036 56544 6100 56548
rect 6116 56604 6180 56608
rect 6116 56548 6120 56604
rect 6120 56548 6176 56604
rect 6176 56548 6180 56604
rect 6116 56544 6180 56548
rect 6196 56604 6260 56608
rect 6196 56548 6200 56604
rect 6200 56548 6256 56604
rect 6256 56548 6260 56604
rect 6196 56544 6260 56548
rect 86548 56604 86612 56608
rect 86548 56548 86552 56604
rect 86552 56548 86608 56604
rect 86608 56548 86612 56604
rect 86548 56544 86612 56548
rect 86628 56604 86692 56608
rect 86628 56548 86632 56604
rect 86632 56548 86688 56604
rect 86688 56548 86692 56604
rect 86628 56544 86692 56548
rect 86708 56604 86772 56608
rect 86708 56548 86712 56604
rect 86712 56548 86768 56604
rect 86768 56548 86772 56604
rect 86708 56544 86772 56548
rect 86788 56604 86852 56608
rect 86788 56548 86792 56604
rect 86792 56548 86848 56604
rect 86848 56548 86852 56604
rect 86788 56544 86852 56548
rect 6692 56060 6756 56064
rect 6692 56004 6696 56060
rect 6696 56004 6752 56060
rect 6752 56004 6756 56060
rect 6692 56000 6756 56004
rect 6772 56060 6836 56064
rect 6772 56004 6776 56060
rect 6776 56004 6832 56060
rect 6832 56004 6836 56060
rect 6772 56000 6836 56004
rect 6852 56060 6916 56064
rect 6852 56004 6856 56060
rect 6856 56004 6912 56060
rect 6912 56004 6916 56060
rect 6852 56000 6916 56004
rect 6932 56060 6996 56064
rect 6932 56004 6936 56060
rect 6936 56004 6992 56060
rect 6992 56004 6996 56060
rect 6932 56000 6996 56004
rect 87284 56060 87348 56064
rect 87284 56004 87288 56060
rect 87288 56004 87344 56060
rect 87344 56004 87348 56060
rect 87284 56000 87348 56004
rect 87364 56060 87428 56064
rect 87364 56004 87368 56060
rect 87368 56004 87424 56060
rect 87424 56004 87428 56060
rect 87364 56000 87428 56004
rect 87444 56060 87508 56064
rect 87444 56004 87448 56060
rect 87448 56004 87504 56060
rect 87504 56004 87508 56060
rect 87444 56000 87508 56004
rect 87524 56060 87588 56064
rect 87524 56004 87528 56060
rect 87528 56004 87584 56060
rect 87584 56004 87588 56060
rect 87524 56000 87588 56004
rect 5956 55516 6020 55520
rect 5956 55460 5960 55516
rect 5960 55460 6016 55516
rect 6016 55460 6020 55516
rect 5956 55456 6020 55460
rect 6036 55516 6100 55520
rect 6036 55460 6040 55516
rect 6040 55460 6096 55516
rect 6096 55460 6100 55516
rect 6036 55456 6100 55460
rect 6116 55516 6180 55520
rect 6116 55460 6120 55516
rect 6120 55460 6176 55516
rect 6176 55460 6180 55516
rect 6116 55456 6180 55460
rect 6196 55516 6260 55520
rect 6196 55460 6200 55516
rect 6200 55460 6256 55516
rect 6256 55460 6260 55516
rect 6196 55456 6260 55460
rect 86548 55516 86612 55520
rect 86548 55460 86552 55516
rect 86552 55460 86608 55516
rect 86608 55460 86612 55516
rect 86548 55456 86612 55460
rect 86628 55516 86692 55520
rect 86628 55460 86632 55516
rect 86632 55460 86688 55516
rect 86688 55460 86692 55516
rect 86628 55456 86692 55460
rect 86708 55516 86772 55520
rect 86708 55460 86712 55516
rect 86712 55460 86768 55516
rect 86768 55460 86772 55516
rect 86708 55456 86772 55460
rect 86788 55516 86852 55520
rect 86788 55460 86792 55516
rect 86792 55460 86848 55516
rect 86848 55460 86852 55516
rect 86788 55456 86852 55460
rect 6692 54972 6756 54976
rect 6692 54916 6696 54972
rect 6696 54916 6752 54972
rect 6752 54916 6756 54972
rect 6692 54912 6756 54916
rect 6772 54972 6836 54976
rect 6772 54916 6776 54972
rect 6776 54916 6832 54972
rect 6832 54916 6836 54972
rect 6772 54912 6836 54916
rect 6852 54972 6916 54976
rect 6852 54916 6856 54972
rect 6856 54916 6912 54972
rect 6912 54916 6916 54972
rect 6852 54912 6916 54916
rect 6932 54972 6996 54976
rect 6932 54916 6936 54972
rect 6936 54916 6992 54972
rect 6992 54916 6996 54972
rect 6932 54912 6996 54916
rect 87284 54972 87348 54976
rect 87284 54916 87288 54972
rect 87288 54916 87344 54972
rect 87344 54916 87348 54972
rect 87284 54912 87348 54916
rect 87364 54972 87428 54976
rect 87364 54916 87368 54972
rect 87368 54916 87424 54972
rect 87424 54916 87428 54972
rect 87364 54912 87428 54916
rect 87444 54972 87508 54976
rect 87444 54916 87448 54972
rect 87448 54916 87504 54972
rect 87504 54916 87508 54972
rect 87444 54912 87508 54916
rect 87524 54972 87588 54976
rect 87524 54916 87528 54972
rect 87528 54916 87584 54972
rect 87584 54916 87588 54972
rect 87524 54912 87588 54916
rect 5956 54428 6020 54432
rect 5956 54372 5960 54428
rect 5960 54372 6016 54428
rect 6016 54372 6020 54428
rect 5956 54368 6020 54372
rect 6036 54428 6100 54432
rect 6036 54372 6040 54428
rect 6040 54372 6096 54428
rect 6096 54372 6100 54428
rect 6036 54368 6100 54372
rect 6116 54428 6180 54432
rect 6116 54372 6120 54428
rect 6120 54372 6176 54428
rect 6176 54372 6180 54428
rect 6116 54368 6180 54372
rect 6196 54428 6260 54432
rect 6196 54372 6200 54428
rect 6200 54372 6256 54428
rect 6256 54372 6260 54428
rect 6196 54368 6260 54372
rect 86548 54428 86612 54432
rect 86548 54372 86552 54428
rect 86552 54372 86608 54428
rect 86608 54372 86612 54428
rect 86548 54368 86612 54372
rect 86628 54428 86692 54432
rect 86628 54372 86632 54428
rect 86632 54372 86688 54428
rect 86688 54372 86692 54428
rect 86628 54368 86692 54372
rect 86708 54428 86772 54432
rect 86708 54372 86712 54428
rect 86712 54372 86768 54428
rect 86768 54372 86772 54428
rect 86708 54368 86772 54372
rect 86788 54428 86852 54432
rect 86788 54372 86792 54428
rect 86792 54372 86848 54428
rect 86848 54372 86852 54428
rect 86788 54368 86852 54372
rect 6692 53884 6756 53888
rect 6692 53828 6696 53884
rect 6696 53828 6752 53884
rect 6752 53828 6756 53884
rect 6692 53824 6756 53828
rect 6772 53884 6836 53888
rect 6772 53828 6776 53884
rect 6776 53828 6832 53884
rect 6832 53828 6836 53884
rect 6772 53824 6836 53828
rect 6852 53884 6916 53888
rect 6852 53828 6856 53884
rect 6856 53828 6912 53884
rect 6912 53828 6916 53884
rect 6852 53824 6916 53828
rect 6932 53884 6996 53888
rect 6932 53828 6936 53884
rect 6936 53828 6992 53884
rect 6992 53828 6996 53884
rect 6932 53824 6996 53828
rect 87284 53884 87348 53888
rect 87284 53828 87288 53884
rect 87288 53828 87344 53884
rect 87344 53828 87348 53884
rect 87284 53824 87348 53828
rect 87364 53884 87428 53888
rect 87364 53828 87368 53884
rect 87368 53828 87424 53884
rect 87424 53828 87428 53884
rect 87364 53824 87428 53828
rect 87444 53884 87508 53888
rect 87444 53828 87448 53884
rect 87448 53828 87504 53884
rect 87504 53828 87508 53884
rect 87444 53824 87508 53828
rect 87524 53884 87588 53888
rect 87524 53828 87528 53884
rect 87528 53828 87584 53884
rect 87584 53828 87588 53884
rect 87524 53824 87588 53828
rect 5956 53340 6020 53344
rect 5956 53284 5960 53340
rect 5960 53284 6016 53340
rect 6016 53284 6020 53340
rect 5956 53280 6020 53284
rect 6036 53340 6100 53344
rect 6036 53284 6040 53340
rect 6040 53284 6096 53340
rect 6096 53284 6100 53340
rect 6036 53280 6100 53284
rect 6116 53340 6180 53344
rect 6116 53284 6120 53340
rect 6120 53284 6176 53340
rect 6176 53284 6180 53340
rect 6116 53280 6180 53284
rect 6196 53340 6260 53344
rect 6196 53284 6200 53340
rect 6200 53284 6256 53340
rect 6256 53284 6260 53340
rect 6196 53280 6260 53284
rect 86548 53340 86612 53344
rect 86548 53284 86552 53340
rect 86552 53284 86608 53340
rect 86608 53284 86612 53340
rect 86548 53280 86612 53284
rect 86628 53340 86692 53344
rect 86628 53284 86632 53340
rect 86632 53284 86688 53340
rect 86688 53284 86692 53340
rect 86628 53280 86692 53284
rect 86708 53340 86772 53344
rect 86708 53284 86712 53340
rect 86712 53284 86768 53340
rect 86768 53284 86772 53340
rect 86708 53280 86772 53284
rect 86788 53340 86852 53344
rect 86788 53284 86792 53340
rect 86792 53284 86848 53340
rect 86848 53284 86852 53340
rect 86788 53280 86852 53284
rect 6692 52796 6756 52800
rect 6692 52740 6696 52796
rect 6696 52740 6752 52796
rect 6752 52740 6756 52796
rect 6692 52736 6756 52740
rect 6772 52796 6836 52800
rect 6772 52740 6776 52796
rect 6776 52740 6832 52796
rect 6832 52740 6836 52796
rect 6772 52736 6836 52740
rect 6852 52796 6916 52800
rect 6852 52740 6856 52796
rect 6856 52740 6912 52796
rect 6912 52740 6916 52796
rect 6852 52736 6916 52740
rect 6932 52796 6996 52800
rect 6932 52740 6936 52796
rect 6936 52740 6992 52796
rect 6992 52740 6996 52796
rect 6932 52736 6996 52740
rect 87284 52796 87348 52800
rect 87284 52740 87288 52796
rect 87288 52740 87344 52796
rect 87344 52740 87348 52796
rect 87284 52736 87348 52740
rect 87364 52796 87428 52800
rect 87364 52740 87368 52796
rect 87368 52740 87424 52796
rect 87424 52740 87428 52796
rect 87364 52736 87428 52740
rect 87444 52796 87508 52800
rect 87444 52740 87448 52796
rect 87448 52740 87504 52796
rect 87504 52740 87508 52796
rect 87444 52736 87508 52740
rect 87524 52796 87588 52800
rect 87524 52740 87528 52796
rect 87528 52740 87584 52796
rect 87584 52740 87588 52796
rect 87524 52736 87588 52740
rect 5956 52252 6020 52256
rect 5956 52196 5960 52252
rect 5960 52196 6016 52252
rect 6016 52196 6020 52252
rect 5956 52192 6020 52196
rect 6036 52252 6100 52256
rect 6036 52196 6040 52252
rect 6040 52196 6096 52252
rect 6096 52196 6100 52252
rect 6036 52192 6100 52196
rect 6116 52252 6180 52256
rect 6116 52196 6120 52252
rect 6120 52196 6176 52252
rect 6176 52196 6180 52252
rect 6116 52192 6180 52196
rect 6196 52252 6260 52256
rect 6196 52196 6200 52252
rect 6200 52196 6256 52252
rect 6256 52196 6260 52252
rect 6196 52192 6260 52196
rect 86548 52252 86612 52256
rect 86548 52196 86552 52252
rect 86552 52196 86608 52252
rect 86608 52196 86612 52252
rect 86548 52192 86612 52196
rect 86628 52252 86692 52256
rect 86628 52196 86632 52252
rect 86632 52196 86688 52252
rect 86688 52196 86692 52252
rect 86628 52192 86692 52196
rect 86708 52252 86772 52256
rect 86708 52196 86712 52252
rect 86712 52196 86768 52252
rect 86768 52196 86772 52252
rect 86708 52192 86772 52196
rect 86788 52252 86852 52256
rect 86788 52196 86792 52252
rect 86792 52196 86848 52252
rect 86848 52196 86852 52252
rect 86788 52192 86852 52196
rect 6692 51708 6756 51712
rect 6692 51652 6696 51708
rect 6696 51652 6752 51708
rect 6752 51652 6756 51708
rect 6692 51648 6756 51652
rect 6772 51708 6836 51712
rect 6772 51652 6776 51708
rect 6776 51652 6832 51708
rect 6832 51652 6836 51708
rect 6772 51648 6836 51652
rect 6852 51708 6916 51712
rect 6852 51652 6856 51708
rect 6856 51652 6912 51708
rect 6912 51652 6916 51708
rect 6852 51648 6916 51652
rect 6932 51708 6996 51712
rect 6932 51652 6936 51708
rect 6936 51652 6992 51708
rect 6992 51652 6996 51708
rect 6932 51648 6996 51652
rect 87284 51708 87348 51712
rect 87284 51652 87288 51708
rect 87288 51652 87344 51708
rect 87344 51652 87348 51708
rect 87284 51648 87348 51652
rect 87364 51708 87428 51712
rect 87364 51652 87368 51708
rect 87368 51652 87424 51708
rect 87424 51652 87428 51708
rect 87364 51648 87428 51652
rect 87444 51708 87508 51712
rect 87444 51652 87448 51708
rect 87448 51652 87504 51708
rect 87504 51652 87508 51708
rect 87444 51648 87508 51652
rect 87524 51708 87588 51712
rect 87524 51652 87528 51708
rect 87528 51652 87584 51708
rect 87584 51652 87588 51708
rect 87524 51648 87588 51652
rect 5956 51164 6020 51168
rect 5956 51108 5960 51164
rect 5960 51108 6016 51164
rect 6016 51108 6020 51164
rect 5956 51104 6020 51108
rect 6036 51164 6100 51168
rect 6036 51108 6040 51164
rect 6040 51108 6096 51164
rect 6096 51108 6100 51164
rect 6036 51104 6100 51108
rect 6116 51164 6180 51168
rect 6116 51108 6120 51164
rect 6120 51108 6176 51164
rect 6176 51108 6180 51164
rect 6116 51104 6180 51108
rect 6196 51164 6260 51168
rect 6196 51108 6200 51164
rect 6200 51108 6256 51164
rect 6256 51108 6260 51164
rect 6196 51104 6260 51108
rect 86548 51164 86612 51168
rect 86548 51108 86552 51164
rect 86552 51108 86608 51164
rect 86608 51108 86612 51164
rect 86548 51104 86612 51108
rect 86628 51164 86692 51168
rect 86628 51108 86632 51164
rect 86632 51108 86688 51164
rect 86688 51108 86692 51164
rect 86628 51104 86692 51108
rect 86708 51164 86772 51168
rect 86708 51108 86712 51164
rect 86712 51108 86768 51164
rect 86768 51108 86772 51164
rect 86708 51104 86772 51108
rect 86788 51164 86852 51168
rect 86788 51108 86792 51164
rect 86792 51108 86848 51164
rect 86848 51108 86852 51164
rect 86788 51104 86852 51108
rect 6692 50620 6756 50624
rect 6692 50564 6696 50620
rect 6696 50564 6752 50620
rect 6752 50564 6756 50620
rect 6692 50560 6756 50564
rect 6772 50620 6836 50624
rect 6772 50564 6776 50620
rect 6776 50564 6832 50620
rect 6832 50564 6836 50620
rect 6772 50560 6836 50564
rect 6852 50620 6916 50624
rect 6852 50564 6856 50620
rect 6856 50564 6912 50620
rect 6912 50564 6916 50620
rect 6852 50560 6916 50564
rect 6932 50620 6996 50624
rect 6932 50564 6936 50620
rect 6936 50564 6992 50620
rect 6992 50564 6996 50620
rect 6932 50560 6996 50564
rect 87284 50620 87348 50624
rect 87284 50564 87288 50620
rect 87288 50564 87344 50620
rect 87344 50564 87348 50620
rect 87284 50560 87348 50564
rect 87364 50620 87428 50624
rect 87364 50564 87368 50620
rect 87368 50564 87424 50620
rect 87424 50564 87428 50620
rect 87364 50560 87428 50564
rect 87444 50620 87508 50624
rect 87444 50564 87448 50620
rect 87448 50564 87504 50620
rect 87504 50564 87508 50620
rect 87444 50560 87508 50564
rect 87524 50620 87588 50624
rect 87524 50564 87528 50620
rect 87528 50564 87584 50620
rect 87584 50564 87588 50620
rect 87524 50560 87588 50564
rect 5956 50076 6020 50080
rect 5956 50020 5960 50076
rect 5960 50020 6016 50076
rect 6016 50020 6020 50076
rect 5956 50016 6020 50020
rect 6036 50076 6100 50080
rect 6036 50020 6040 50076
rect 6040 50020 6096 50076
rect 6096 50020 6100 50076
rect 6036 50016 6100 50020
rect 6116 50076 6180 50080
rect 6116 50020 6120 50076
rect 6120 50020 6176 50076
rect 6176 50020 6180 50076
rect 6116 50016 6180 50020
rect 6196 50076 6260 50080
rect 6196 50020 6200 50076
rect 6200 50020 6256 50076
rect 6256 50020 6260 50076
rect 6196 50016 6260 50020
rect 86548 50076 86612 50080
rect 86548 50020 86552 50076
rect 86552 50020 86608 50076
rect 86608 50020 86612 50076
rect 86548 50016 86612 50020
rect 86628 50076 86692 50080
rect 86628 50020 86632 50076
rect 86632 50020 86688 50076
rect 86688 50020 86692 50076
rect 86628 50016 86692 50020
rect 86708 50076 86772 50080
rect 86708 50020 86712 50076
rect 86712 50020 86768 50076
rect 86768 50020 86772 50076
rect 86708 50016 86772 50020
rect 86788 50076 86852 50080
rect 86788 50020 86792 50076
rect 86792 50020 86848 50076
rect 86848 50020 86852 50076
rect 86788 50016 86852 50020
rect 6692 49532 6756 49536
rect 6692 49476 6696 49532
rect 6696 49476 6752 49532
rect 6752 49476 6756 49532
rect 6692 49472 6756 49476
rect 6772 49532 6836 49536
rect 6772 49476 6776 49532
rect 6776 49476 6832 49532
rect 6832 49476 6836 49532
rect 6772 49472 6836 49476
rect 6852 49532 6916 49536
rect 6852 49476 6856 49532
rect 6856 49476 6912 49532
rect 6912 49476 6916 49532
rect 6852 49472 6916 49476
rect 6932 49532 6996 49536
rect 6932 49476 6936 49532
rect 6936 49476 6992 49532
rect 6992 49476 6996 49532
rect 6932 49472 6996 49476
rect 87284 49532 87348 49536
rect 87284 49476 87288 49532
rect 87288 49476 87344 49532
rect 87344 49476 87348 49532
rect 87284 49472 87348 49476
rect 87364 49532 87428 49536
rect 87364 49476 87368 49532
rect 87368 49476 87424 49532
rect 87424 49476 87428 49532
rect 87364 49472 87428 49476
rect 87444 49532 87508 49536
rect 87444 49476 87448 49532
rect 87448 49476 87504 49532
rect 87504 49476 87508 49532
rect 87444 49472 87508 49476
rect 87524 49532 87588 49536
rect 87524 49476 87528 49532
rect 87528 49476 87584 49532
rect 87584 49476 87588 49532
rect 87524 49472 87588 49476
rect 5956 48988 6020 48992
rect 5956 48932 5960 48988
rect 5960 48932 6016 48988
rect 6016 48932 6020 48988
rect 5956 48928 6020 48932
rect 6036 48988 6100 48992
rect 6036 48932 6040 48988
rect 6040 48932 6096 48988
rect 6096 48932 6100 48988
rect 6036 48928 6100 48932
rect 6116 48988 6180 48992
rect 6116 48932 6120 48988
rect 6120 48932 6176 48988
rect 6176 48932 6180 48988
rect 6116 48928 6180 48932
rect 6196 48988 6260 48992
rect 6196 48932 6200 48988
rect 6200 48932 6256 48988
rect 6256 48932 6260 48988
rect 6196 48928 6260 48932
rect 86548 48988 86612 48992
rect 86548 48932 86552 48988
rect 86552 48932 86608 48988
rect 86608 48932 86612 48988
rect 86548 48928 86612 48932
rect 86628 48988 86692 48992
rect 86628 48932 86632 48988
rect 86632 48932 86688 48988
rect 86688 48932 86692 48988
rect 86628 48928 86692 48932
rect 86708 48988 86772 48992
rect 86708 48932 86712 48988
rect 86712 48932 86768 48988
rect 86768 48932 86772 48988
rect 86708 48928 86772 48932
rect 86788 48988 86852 48992
rect 86788 48932 86792 48988
rect 86792 48932 86848 48988
rect 86848 48932 86852 48988
rect 86788 48928 86852 48932
rect 6692 48444 6756 48448
rect 6692 48388 6696 48444
rect 6696 48388 6752 48444
rect 6752 48388 6756 48444
rect 6692 48384 6756 48388
rect 6772 48444 6836 48448
rect 6772 48388 6776 48444
rect 6776 48388 6832 48444
rect 6832 48388 6836 48444
rect 6772 48384 6836 48388
rect 6852 48444 6916 48448
rect 6852 48388 6856 48444
rect 6856 48388 6912 48444
rect 6912 48388 6916 48444
rect 6852 48384 6916 48388
rect 6932 48444 6996 48448
rect 6932 48388 6936 48444
rect 6936 48388 6992 48444
rect 6992 48388 6996 48444
rect 6932 48384 6996 48388
rect 87284 48444 87348 48448
rect 87284 48388 87288 48444
rect 87288 48388 87344 48444
rect 87344 48388 87348 48444
rect 87284 48384 87348 48388
rect 87364 48444 87428 48448
rect 87364 48388 87368 48444
rect 87368 48388 87424 48444
rect 87424 48388 87428 48444
rect 87364 48384 87428 48388
rect 87444 48444 87508 48448
rect 87444 48388 87448 48444
rect 87448 48388 87504 48444
rect 87504 48388 87508 48444
rect 87444 48384 87508 48388
rect 87524 48444 87588 48448
rect 87524 48388 87528 48444
rect 87528 48388 87584 48444
rect 87584 48388 87588 48444
rect 87524 48384 87588 48388
rect 5956 47900 6020 47904
rect 5956 47844 5960 47900
rect 5960 47844 6016 47900
rect 6016 47844 6020 47900
rect 5956 47840 6020 47844
rect 6036 47900 6100 47904
rect 6036 47844 6040 47900
rect 6040 47844 6096 47900
rect 6096 47844 6100 47900
rect 6036 47840 6100 47844
rect 6116 47900 6180 47904
rect 6116 47844 6120 47900
rect 6120 47844 6176 47900
rect 6176 47844 6180 47900
rect 6116 47840 6180 47844
rect 6196 47900 6260 47904
rect 6196 47844 6200 47900
rect 6200 47844 6256 47900
rect 6256 47844 6260 47900
rect 6196 47840 6260 47844
rect 86548 47900 86612 47904
rect 86548 47844 86552 47900
rect 86552 47844 86608 47900
rect 86608 47844 86612 47900
rect 86548 47840 86612 47844
rect 86628 47900 86692 47904
rect 86628 47844 86632 47900
rect 86632 47844 86688 47900
rect 86688 47844 86692 47900
rect 86628 47840 86692 47844
rect 86708 47900 86772 47904
rect 86708 47844 86712 47900
rect 86712 47844 86768 47900
rect 86768 47844 86772 47900
rect 86708 47840 86772 47844
rect 86788 47900 86852 47904
rect 86788 47844 86792 47900
rect 86792 47844 86848 47900
rect 86848 47844 86852 47900
rect 86788 47840 86852 47844
rect 6692 47356 6756 47360
rect 6692 47300 6696 47356
rect 6696 47300 6752 47356
rect 6752 47300 6756 47356
rect 6692 47296 6756 47300
rect 6772 47356 6836 47360
rect 6772 47300 6776 47356
rect 6776 47300 6832 47356
rect 6832 47300 6836 47356
rect 6772 47296 6836 47300
rect 6852 47356 6916 47360
rect 6852 47300 6856 47356
rect 6856 47300 6912 47356
rect 6912 47300 6916 47356
rect 6852 47296 6916 47300
rect 6932 47356 6996 47360
rect 6932 47300 6936 47356
rect 6936 47300 6992 47356
rect 6992 47300 6996 47356
rect 6932 47296 6996 47300
rect 87284 47356 87348 47360
rect 87284 47300 87288 47356
rect 87288 47300 87344 47356
rect 87344 47300 87348 47356
rect 87284 47296 87348 47300
rect 87364 47356 87428 47360
rect 87364 47300 87368 47356
rect 87368 47300 87424 47356
rect 87424 47300 87428 47356
rect 87364 47296 87428 47300
rect 87444 47356 87508 47360
rect 87444 47300 87448 47356
rect 87448 47300 87504 47356
rect 87504 47300 87508 47356
rect 87444 47296 87508 47300
rect 87524 47356 87588 47360
rect 87524 47300 87528 47356
rect 87528 47300 87584 47356
rect 87584 47300 87588 47356
rect 87524 47296 87588 47300
rect 5956 46812 6020 46816
rect 5956 46756 5960 46812
rect 5960 46756 6016 46812
rect 6016 46756 6020 46812
rect 5956 46752 6020 46756
rect 6036 46812 6100 46816
rect 6036 46756 6040 46812
rect 6040 46756 6096 46812
rect 6096 46756 6100 46812
rect 6036 46752 6100 46756
rect 6116 46812 6180 46816
rect 6116 46756 6120 46812
rect 6120 46756 6176 46812
rect 6176 46756 6180 46812
rect 6116 46752 6180 46756
rect 6196 46812 6260 46816
rect 6196 46756 6200 46812
rect 6200 46756 6256 46812
rect 6256 46756 6260 46812
rect 6196 46752 6260 46756
rect 86548 46812 86612 46816
rect 86548 46756 86552 46812
rect 86552 46756 86608 46812
rect 86608 46756 86612 46812
rect 86548 46752 86612 46756
rect 86628 46812 86692 46816
rect 86628 46756 86632 46812
rect 86632 46756 86688 46812
rect 86688 46756 86692 46812
rect 86628 46752 86692 46756
rect 86708 46812 86772 46816
rect 86708 46756 86712 46812
rect 86712 46756 86768 46812
rect 86768 46756 86772 46812
rect 86708 46752 86772 46756
rect 86788 46812 86852 46816
rect 86788 46756 86792 46812
rect 86792 46756 86848 46812
rect 86848 46756 86852 46812
rect 86788 46752 86852 46756
rect 6692 46268 6756 46272
rect 6692 46212 6696 46268
rect 6696 46212 6752 46268
rect 6752 46212 6756 46268
rect 6692 46208 6756 46212
rect 6772 46268 6836 46272
rect 6772 46212 6776 46268
rect 6776 46212 6832 46268
rect 6832 46212 6836 46268
rect 6772 46208 6836 46212
rect 6852 46268 6916 46272
rect 6852 46212 6856 46268
rect 6856 46212 6912 46268
rect 6912 46212 6916 46268
rect 6852 46208 6916 46212
rect 6932 46268 6996 46272
rect 6932 46212 6936 46268
rect 6936 46212 6992 46268
rect 6992 46212 6996 46268
rect 6932 46208 6996 46212
rect 87284 46268 87348 46272
rect 87284 46212 87288 46268
rect 87288 46212 87344 46268
rect 87344 46212 87348 46268
rect 87284 46208 87348 46212
rect 87364 46268 87428 46272
rect 87364 46212 87368 46268
rect 87368 46212 87424 46268
rect 87424 46212 87428 46268
rect 87364 46208 87428 46212
rect 87444 46268 87508 46272
rect 87444 46212 87448 46268
rect 87448 46212 87504 46268
rect 87504 46212 87508 46268
rect 87444 46208 87508 46212
rect 87524 46268 87588 46272
rect 87524 46212 87528 46268
rect 87528 46212 87584 46268
rect 87584 46212 87588 46268
rect 87524 46208 87588 46212
rect 5956 45724 6020 45728
rect 5956 45668 5960 45724
rect 5960 45668 6016 45724
rect 6016 45668 6020 45724
rect 5956 45664 6020 45668
rect 6036 45724 6100 45728
rect 6036 45668 6040 45724
rect 6040 45668 6096 45724
rect 6096 45668 6100 45724
rect 6036 45664 6100 45668
rect 6116 45724 6180 45728
rect 6116 45668 6120 45724
rect 6120 45668 6176 45724
rect 6176 45668 6180 45724
rect 6116 45664 6180 45668
rect 6196 45724 6260 45728
rect 6196 45668 6200 45724
rect 6200 45668 6256 45724
rect 6256 45668 6260 45724
rect 6196 45664 6260 45668
rect 86548 45724 86612 45728
rect 86548 45668 86552 45724
rect 86552 45668 86608 45724
rect 86608 45668 86612 45724
rect 86548 45664 86612 45668
rect 86628 45724 86692 45728
rect 86628 45668 86632 45724
rect 86632 45668 86688 45724
rect 86688 45668 86692 45724
rect 86628 45664 86692 45668
rect 86708 45724 86772 45728
rect 86708 45668 86712 45724
rect 86712 45668 86768 45724
rect 86768 45668 86772 45724
rect 86708 45664 86772 45668
rect 86788 45724 86852 45728
rect 86788 45668 86792 45724
rect 86792 45668 86848 45724
rect 86848 45668 86852 45724
rect 86788 45664 86852 45668
rect 6692 45180 6756 45184
rect 6692 45124 6696 45180
rect 6696 45124 6752 45180
rect 6752 45124 6756 45180
rect 6692 45120 6756 45124
rect 6772 45180 6836 45184
rect 6772 45124 6776 45180
rect 6776 45124 6832 45180
rect 6832 45124 6836 45180
rect 6772 45120 6836 45124
rect 6852 45180 6916 45184
rect 6852 45124 6856 45180
rect 6856 45124 6912 45180
rect 6912 45124 6916 45180
rect 6852 45120 6916 45124
rect 6932 45180 6996 45184
rect 6932 45124 6936 45180
rect 6936 45124 6992 45180
rect 6992 45124 6996 45180
rect 6932 45120 6996 45124
rect 87284 45180 87348 45184
rect 87284 45124 87288 45180
rect 87288 45124 87344 45180
rect 87344 45124 87348 45180
rect 87284 45120 87348 45124
rect 87364 45180 87428 45184
rect 87364 45124 87368 45180
rect 87368 45124 87424 45180
rect 87424 45124 87428 45180
rect 87364 45120 87428 45124
rect 87444 45180 87508 45184
rect 87444 45124 87448 45180
rect 87448 45124 87504 45180
rect 87504 45124 87508 45180
rect 87444 45120 87508 45124
rect 87524 45180 87588 45184
rect 87524 45124 87528 45180
rect 87528 45124 87584 45180
rect 87584 45124 87588 45180
rect 87524 45120 87588 45124
rect 5956 44636 6020 44640
rect 5956 44580 5960 44636
rect 5960 44580 6016 44636
rect 6016 44580 6020 44636
rect 5956 44576 6020 44580
rect 6036 44636 6100 44640
rect 6036 44580 6040 44636
rect 6040 44580 6096 44636
rect 6096 44580 6100 44636
rect 6036 44576 6100 44580
rect 6116 44636 6180 44640
rect 6116 44580 6120 44636
rect 6120 44580 6176 44636
rect 6176 44580 6180 44636
rect 6116 44576 6180 44580
rect 6196 44636 6260 44640
rect 6196 44580 6200 44636
rect 6200 44580 6256 44636
rect 6256 44580 6260 44636
rect 6196 44576 6260 44580
rect 86548 44636 86612 44640
rect 86548 44580 86552 44636
rect 86552 44580 86608 44636
rect 86608 44580 86612 44636
rect 86548 44576 86612 44580
rect 86628 44636 86692 44640
rect 86628 44580 86632 44636
rect 86632 44580 86688 44636
rect 86688 44580 86692 44636
rect 86628 44576 86692 44580
rect 86708 44636 86772 44640
rect 86708 44580 86712 44636
rect 86712 44580 86768 44636
rect 86768 44580 86772 44636
rect 86708 44576 86772 44580
rect 86788 44636 86852 44640
rect 86788 44580 86792 44636
rect 86792 44580 86848 44636
rect 86848 44580 86852 44636
rect 86788 44576 86852 44580
rect 6692 44092 6756 44096
rect 6692 44036 6696 44092
rect 6696 44036 6752 44092
rect 6752 44036 6756 44092
rect 6692 44032 6756 44036
rect 6772 44092 6836 44096
rect 6772 44036 6776 44092
rect 6776 44036 6832 44092
rect 6832 44036 6836 44092
rect 6772 44032 6836 44036
rect 6852 44092 6916 44096
rect 6852 44036 6856 44092
rect 6856 44036 6912 44092
rect 6912 44036 6916 44092
rect 6852 44032 6916 44036
rect 6932 44092 6996 44096
rect 6932 44036 6936 44092
rect 6936 44036 6992 44092
rect 6992 44036 6996 44092
rect 6932 44032 6996 44036
rect 87284 44092 87348 44096
rect 87284 44036 87288 44092
rect 87288 44036 87344 44092
rect 87344 44036 87348 44092
rect 87284 44032 87348 44036
rect 87364 44092 87428 44096
rect 87364 44036 87368 44092
rect 87368 44036 87424 44092
rect 87424 44036 87428 44092
rect 87364 44032 87428 44036
rect 87444 44092 87508 44096
rect 87444 44036 87448 44092
rect 87448 44036 87504 44092
rect 87504 44036 87508 44092
rect 87444 44032 87508 44036
rect 87524 44092 87588 44096
rect 87524 44036 87528 44092
rect 87528 44036 87584 44092
rect 87584 44036 87588 44092
rect 87524 44032 87588 44036
rect 5956 43548 6020 43552
rect 5956 43492 5960 43548
rect 5960 43492 6016 43548
rect 6016 43492 6020 43548
rect 5956 43488 6020 43492
rect 6036 43548 6100 43552
rect 6036 43492 6040 43548
rect 6040 43492 6096 43548
rect 6096 43492 6100 43548
rect 6036 43488 6100 43492
rect 6116 43548 6180 43552
rect 6116 43492 6120 43548
rect 6120 43492 6176 43548
rect 6176 43492 6180 43548
rect 6116 43488 6180 43492
rect 6196 43548 6260 43552
rect 6196 43492 6200 43548
rect 6200 43492 6256 43548
rect 6256 43492 6260 43548
rect 6196 43488 6260 43492
rect 86548 43548 86612 43552
rect 86548 43492 86552 43548
rect 86552 43492 86608 43548
rect 86608 43492 86612 43548
rect 86548 43488 86612 43492
rect 86628 43548 86692 43552
rect 86628 43492 86632 43548
rect 86632 43492 86688 43548
rect 86688 43492 86692 43548
rect 86628 43488 86692 43492
rect 86708 43548 86772 43552
rect 86708 43492 86712 43548
rect 86712 43492 86768 43548
rect 86768 43492 86772 43548
rect 86708 43488 86772 43492
rect 86788 43548 86852 43552
rect 86788 43492 86792 43548
rect 86792 43492 86848 43548
rect 86848 43492 86852 43548
rect 86788 43488 86852 43492
rect 6692 43004 6756 43008
rect 6692 42948 6696 43004
rect 6696 42948 6752 43004
rect 6752 42948 6756 43004
rect 6692 42944 6756 42948
rect 6772 43004 6836 43008
rect 6772 42948 6776 43004
rect 6776 42948 6832 43004
rect 6832 42948 6836 43004
rect 6772 42944 6836 42948
rect 6852 43004 6916 43008
rect 6852 42948 6856 43004
rect 6856 42948 6912 43004
rect 6912 42948 6916 43004
rect 6852 42944 6916 42948
rect 6932 43004 6996 43008
rect 6932 42948 6936 43004
rect 6936 42948 6992 43004
rect 6992 42948 6996 43004
rect 6932 42944 6996 42948
rect 87284 43004 87348 43008
rect 87284 42948 87288 43004
rect 87288 42948 87344 43004
rect 87344 42948 87348 43004
rect 87284 42944 87348 42948
rect 87364 43004 87428 43008
rect 87364 42948 87368 43004
rect 87368 42948 87424 43004
rect 87424 42948 87428 43004
rect 87364 42944 87428 42948
rect 87444 43004 87508 43008
rect 87444 42948 87448 43004
rect 87448 42948 87504 43004
rect 87504 42948 87508 43004
rect 87444 42944 87508 42948
rect 87524 43004 87588 43008
rect 87524 42948 87528 43004
rect 87528 42948 87584 43004
rect 87584 42948 87588 43004
rect 87524 42944 87588 42948
rect 5956 42460 6020 42464
rect 5956 42404 5960 42460
rect 5960 42404 6016 42460
rect 6016 42404 6020 42460
rect 5956 42400 6020 42404
rect 6036 42460 6100 42464
rect 6036 42404 6040 42460
rect 6040 42404 6096 42460
rect 6096 42404 6100 42460
rect 6036 42400 6100 42404
rect 6116 42460 6180 42464
rect 6116 42404 6120 42460
rect 6120 42404 6176 42460
rect 6176 42404 6180 42460
rect 6116 42400 6180 42404
rect 6196 42460 6260 42464
rect 6196 42404 6200 42460
rect 6200 42404 6256 42460
rect 6256 42404 6260 42460
rect 6196 42400 6260 42404
rect 86548 42460 86612 42464
rect 86548 42404 86552 42460
rect 86552 42404 86608 42460
rect 86608 42404 86612 42460
rect 86548 42400 86612 42404
rect 86628 42460 86692 42464
rect 86628 42404 86632 42460
rect 86632 42404 86688 42460
rect 86688 42404 86692 42460
rect 86628 42400 86692 42404
rect 86708 42460 86772 42464
rect 86708 42404 86712 42460
rect 86712 42404 86768 42460
rect 86768 42404 86772 42460
rect 86708 42400 86772 42404
rect 86788 42460 86852 42464
rect 86788 42404 86792 42460
rect 86792 42404 86848 42460
rect 86848 42404 86852 42460
rect 86788 42400 86852 42404
rect 6692 41916 6756 41920
rect 6692 41860 6696 41916
rect 6696 41860 6752 41916
rect 6752 41860 6756 41916
rect 6692 41856 6756 41860
rect 6772 41916 6836 41920
rect 6772 41860 6776 41916
rect 6776 41860 6832 41916
rect 6832 41860 6836 41916
rect 6772 41856 6836 41860
rect 6852 41916 6916 41920
rect 6852 41860 6856 41916
rect 6856 41860 6912 41916
rect 6912 41860 6916 41916
rect 6852 41856 6916 41860
rect 6932 41916 6996 41920
rect 6932 41860 6936 41916
rect 6936 41860 6992 41916
rect 6992 41860 6996 41916
rect 6932 41856 6996 41860
rect 87284 41916 87348 41920
rect 87284 41860 87288 41916
rect 87288 41860 87344 41916
rect 87344 41860 87348 41916
rect 87284 41856 87348 41860
rect 87364 41916 87428 41920
rect 87364 41860 87368 41916
rect 87368 41860 87424 41916
rect 87424 41860 87428 41916
rect 87364 41856 87428 41860
rect 87444 41916 87508 41920
rect 87444 41860 87448 41916
rect 87448 41860 87504 41916
rect 87504 41860 87508 41916
rect 87444 41856 87508 41860
rect 87524 41916 87588 41920
rect 87524 41860 87528 41916
rect 87528 41860 87584 41916
rect 87584 41860 87588 41916
rect 87524 41856 87588 41860
rect 5956 41372 6020 41376
rect 5956 41316 5960 41372
rect 5960 41316 6016 41372
rect 6016 41316 6020 41372
rect 5956 41312 6020 41316
rect 6036 41372 6100 41376
rect 6036 41316 6040 41372
rect 6040 41316 6096 41372
rect 6096 41316 6100 41372
rect 6036 41312 6100 41316
rect 6116 41372 6180 41376
rect 6116 41316 6120 41372
rect 6120 41316 6176 41372
rect 6176 41316 6180 41372
rect 6116 41312 6180 41316
rect 6196 41372 6260 41376
rect 6196 41316 6200 41372
rect 6200 41316 6256 41372
rect 6256 41316 6260 41372
rect 6196 41312 6260 41316
rect 86548 41372 86612 41376
rect 86548 41316 86552 41372
rect 86552 41316 86608 41372
rect 86608 41316 86612 41372
rect 86548 41312 86612 41316
rect 86628 41372 86692 41376
rect 86628 41316 86632 41372
rect 86632 41316 86688 41372
rect 86688 41316 86692 41372
rect 86628 41312 86692 41316
rect 86708 41372 86772 41376
rect 86708 41316 86712 41372
rect 86712 41316 86768 41372
rect 86768 41316 86772 41372
rect 86708 41312 86772 41316
rect 86788 41372 86852 41376
rect 86788 41316 86792 41372
rect 86792 41316 86848 41372
rect 86848 41316 86852 41372
rect 86788 41312 86852 41316
rect 6692 40828 6756 40832
rect 6692 40772 6696 40828
rect 6696 40772 6752 40828
rect 6752 40772 6756 40828
rect 6692 40768 6756 40772
rect 6772 40828 6836 40832
rect 6772 40772 6776 40828
rect 6776 40772 6832 40828
rect 6832 40772 6836 40828
rect 6772 40768 6836 40772
rect 6852 40828 6916 40832
rect 6852 40772 6856 40828
rect 6856 40772 6912 40828
rect 6912 40772 6916 40828
rect 6852 40768 6916 40772
rect 6932 40828 6996 40832
rect 6932 40772 6936 40828
rect 6936 40772 6992 40828
rect 6992 40772 6996 40828
rect 6932 40768 6996 40772
rect 87284 40828 87348 40832
rect 87284 40772 87288 40828
rect 87288 40772 87344 40828
rect 87344 40772 87348 40828
rect 87284 40768 87348 40772
rect 87364 40828 87428 40832
rect 87364 40772 87368 40828
rect 87368 40772 87424 40828
rect 87424 40772 87428 40828
rect 87364 40768 87428 40772
rect 87444 40828 87508 40832
rect 87444 40772 87448 40828
rect 87448 40772 87504 40828
rect 87504 40772 87508 40828
rect 87444 40768 87508 40772
rect 87524 40828 87588 40832
rect 87524 40772 87528 40828
rect 87528 40772 87584 40828
rect 87584 40772 87588 40828
rect 87524 40768 87588 40772
rect 5956 40284 6020 40288
rect 5956 40228 5960 40284
rect 5960 40228 6016 40284
rect 6016 40228 6020 40284
rect 5956 40224 6020 40228
rect 6036 40284 6100 40288
rect 6036 40228 6040 40284
rect 6040 40228 6096 40284
rect 6096 40228 6100 40284
rect 6036 40224 6100 40228
rect 6116 40284 6180 40288
rect 6116 40228 6120 40284
rect 6120 40228 6176 40284
rect 6176 40228 6180 40284
rect 6116 40224 6180 40228
rect 6196 40284 6260 40288
rect 6196 40228 6200 40284
rect 6200 40228 6256 40284
rect 6256 40228 6260 40284
rect 6196 40224 6260 40228
rect 86548 40284 86612 40288
rect 86548 40228 86552 40284
rect 86552 40228 86608 40284
rect 86608 40228 86612 40284
rect 86548 40224 86612 40228
rect 86628 40284 86692 40288
rect 86628 40228 86632 40284
rect 86632 40228 86688 40284
rect 86688 40228 86692 40284
rect 86628 40224 86692 40228
rect 86708 40284 86772 40288
rect 86708 40228 86712 40284
rect 86712 40228 86768 40284
rect 86768 40228 86772 40284
rect 86708 40224 86772 40228
rect 86788 40284 86852 40288
rect 86788 40228 86792 40284
rect 86792 40228 86848 40284
rect 86848 40228 86852 40284
rect 86788 40224 86852 40228
rect 6692 39740 6756 39744
rect 6692 39684 6696 39740
rect 6696 39684 6752 39740
rect 6752 39684 6756 39740
rect 6692 39680 6756 39684
rect 6772 39740 6836 39744
rect 6772 39684 6776 39740
rect 6776 39684 6832 39740
rect 6832 39684 6836 39740
rect 6772 39680 6836 39684
rect 6852 39740 6916 39744
rect 6852 39684 6856 39740
rect 6856 39684 6912 39740
rect 6912 39684 6916 39740
rect 6852 39680 6916 39684
rect 6932 39740 6996 39744
rect 6932 39684 6936 39740
rect 6936 39684 6992 39740
rect 6992 39684 6996 39740
rect 6932 39680 6996 39684
rect 87284 39740 87348 39744
rect 87284 39684 87288 39740
rect 87288 39684 87344 39740
rect 87344 39684 87348 39740
rect 87284 39680 87348 39684
rect 87364 39740 87428 39744
rect 87364 39684 87368 39740
rect 87368 39684 87424 39740
rect 87424 39684 87428 39740
rect 87364 39680 87428 39684
rect 87444 39740 87508 39744
rect 87444 39684 87448 39740
rect 87448 39684 87504 39740
rect 87504 39684 87508 39740
rect 87444 39680 87508 39684
rect 87524 39740 87588 39744
rect 87524 39684 87528 39740
rect 87528 39684 87584 39740
rect 87584 39684 87588 39740
rect 87524 39680 87588 39684
rect 5956 39196 6020 39200
rect 5956 39140 5960 39196
rect 5960 39140 6016 39196
rect 6016 39140 6020 39196
rect 5956 39136 6020 39140
rect 6036 39196 6100 39200
rect 6036 39140 6040 39196
rect 6040 39140 6096 39196
rect 6096 39140 6100 39196
rect 6036 39136 6100 39140
rect 6116 39196 6180 39200
rect 6116 39140 6120 39196
rect 6120 39140 6176 39196
rect 6176 39140 6180 39196
rect 6116 39136 6180 39140
rect 6196 39196 6260 39200
rect 6196 39140 6200 39196
rect 6200 39140 6256 39196
rect 6256 39140 6260 39196
rect 6196 39136 6260 39140
rect 86548 39196 86612 39200
rect 86548 39140 86552 39196
rect 86552 39140 86608 39196
rect 86608 39140 86612 39196
rect 86548 39136 86612 39140
rect 86628 39196 86692 39200
rect 86628 39140 86632 39196
rect 86632 39140 86688 39196
rect 86688 39140 86692 39196
rect 86628 39136 86692 39140
rect 86708 39196 86772 39200
rect 86708 39140 86712 39196
rect 86712 39140 86768 39196
rect 86768 39140 86772 39196
rect 86708 39136 86772 39140
rect 86788 39196 86852 39200
rect 86788 39140 86792 39196
rect 86792 39140 86848 39196
rect 86848 39140 86852 39196
rect 86788 39136 86852 39140
rect 6692 38652 6756 38656
rect 6692 38596 6696 38652
rect 6696 38596 6752 38652
rect 6752 38596 6756 38652
rect 6692 38592 6756 38596
rect 6772 38652 6836 38656
rect 6772 38596 6776 38652
rect 6776 38596 6832 38652
rect 6832 38596 6836 38652
rect 6772 38592 6836 38596
rect 6852 38652 6916 38656
rect 6852 38596 6856 38652
rect 6856 38596 6912 38652
rect 6912 38596 6916 38652
rect 6852 38592 6916 38596
rect 6932 38652 6996 38656
rect 6932 38596 6936 38652
rect 6936 38596 6992 38652
rect 6992 38596 6996 38652
rect 6932 38592 6996 38596
rect 87284 38652 87348 38656
rect 87284 38596 87288 38652
rect 87288 38596 87344 38652
rect 87344 38596 87348 38652
rect 87284 38592 87348 38596
rect 87364 38652 87428 38656
rect 87364 38596 87368 38652
rect 87368 38596 87424 38652
rect 87424 38596 87428 38652
rect 87364 38592 87428 38596
rect 87444 38652 87508 38656
rect 87444 38596 87448 38652
rect 87448 38596 87504 38652
rect 87504 38596 87508 38652
rect 87444 38592 87508 38596
rect 87524 38652 87588 38656
rect 87524 38596 87528 38652
rect 87528 38596 87584 38652
rect 87584 38596 87588 38652
rect 87524 38592 87588 38596
rect 5956 38108 6020 38112
rect 5956 38052 5960 38108
rect 5960 38052 6016 38108
rect 6016 38052 6020 38108
rect 5956 38048 6020 38052
rect 6036 38108 6100 38112
rect 6036 38052 6040 38108
rect 6040 38052 6096 38108
rect 6096 38052 6100 38108
rect 6036 38048 6100 38052
rect 6116 38108 6180 38112
rect 6116 38052 6120 38108
rect 6120 38052 6176 38108
rect 6176 38052 6180 38108
rect 6116 38048 6180 38052
rect 6196 38108 6260 38112
rect 6196 38052 6200 38108
rect 6200 38052 6256 38108
rect 6256 38052 6260 38108
rect 6196 38048 6260 38052
rect 86548 38108 86612 38112
rect 86548 38052 86552 38108
rect 86552 38052 86608 38108
rect 86608 38052 86612 38108
rect 86548 38048 86612 38052
rect 86628 38108 86692 38112
rect 86628 38052 86632 38108
rect 86632 38052 86688 38108
rect 86688 38052 86692 38108
rect 86628 38048 86692 38052
rect 86708 38108 86772 38112
rect 86708 38052 86712 38108
rect 86712 38052 86768 38108
rect 86768 38052 86772 38108
rect 86708 38048 86772 38052
rect 86788 38108 86852 38112
rect 86788 38052 86792 38108
rect 86792 38052 86848 38108
rect 86848 38052 86852 38108
rect 86788 38048 86852 38052
rect 6692 37564 6756 37568
rect 6692 37508 6696 37564
rect 6696 37508 6752 37564
rect 6752 37508 6756 37564
rect 6692 37504 6756 37508
rect 6772 37564 6836 37568
rect 6772 37508 6776 37564
rect 6776 37508 6832 37564
rect 6832 37508 6836 37564
rect 6772 37504 6836 37508
rect 6852 37564 6916 37568
rect 6852 37508 6856 37564
rect 6856 37508 6912 37564
rect 6912 37508 6916 37564
rect 6852 37504 6916 37508
rect 6932 37564 6996 37568
rect 6932 37508 6936 37564
rect 6936 37508 6992 37564
rect 6992 37508 6996 37564
rect 6932 37504 6996 37508
rect 87284 37564 87348 37568
rect 87284 37508 87288 37564
rect 87288 37508 87344 37564
rect 87344 37508 87348 37564
rect 87284 37504 87348 37508
rect 87364 37564 87428 37568
rect 87364 37508 87368 37564
rect 87368 37508 87424 37564
rect 87424 37508 87428 37564
rect 87364 37504 87428 37508
rect 87444 37564 87508 37568
rect 87444 37508 87448 37564
rect 87448 37508 87504 37564
rect 87504 37508 87508 37564
rect 87444 37504 87508 37508
rect 87524 37564 87588 37568
rect 87524 37508 87528 37564
rect 87528 37508 87584 37564
rect 87584 37508 87588 37564
rect 87524 37504 87588 37508
rect 5956 37020 6020 37024
rect 5956 36964 5960 37020
rect 5960 36964 6016 37020
rect 6016 36964 6020 37020
rect 5956 36960 6020 36964
rect 6036 37020 6100 37024
rect 6036 36964 6040 37020
rect 6040 36964 6096 37020
rect 6096 36964 6100 37020
rect 6036 36960 6100 36964
rect 6116 37020 6180 37024
rect 6116 36964 6120 37020
rect 6120 36964 6176 37020
rect 6176 36964 6180 37020
rect 6116 36960 6180 36964
rect 6196 37020 6260 37024
rect 6196 36964 6200 37020
rect 6200 36964 6256 37020
rect 6256 36964 6260 37020
rect 6196 36960 6260 36964
rect 86548 37020 86612 37024
rect 86548 36964 86552 37020
rect 86552 36964 86608 37020
rect 86608 36964 86612 37020
rect 86548 36960 86612 36964
rect 86628 37020 86692 37024
rect 86628 36964 86632 37020
rect 86632 36964 86688 37020
rect 86688 36964 86692 37020
rect 86628 36960 86692 36964
rect 86708 37020 86772 37024
rect 86708 36964 86712 37020
rect 86712 36964 86768 37020
rect 86768 36964 86772 37020
rect 86708 36960 86772 36964
rect 86788 37020 86852 37024
rect 86788 36964 86792 37020
rect 86792 36964 86848 37020
rect 86848 36964 86852 37020
rect 86788 36960 86852 36964
rect 6692 36476 6756 36480
rect 6692 36420 6696 36476
rect 6696 36420 6752 36476
rect 6752 36420 6756 36476
rect 6692 36416 6756 36420
rect 6772 36476 6836 36480
rect 6772 36420 6776 36476
rect 6776 36420 6832 36476
rect 6832 36420 6836 36476
rect 6772 36416 6836 36420
rect 6852 36476 6916 36480
rect 6852 36420 6856 36476
rect 6856 36420 6912 36476
rect 6912 36420 6916 36476
rect 6852 36416 6916 36420
rect 6932 36476 6996 36480
rect 6932 36420 6936 36476
rect 6936 36420 6992 36476
rect 6992 36420 6996 36476
rect 6932 36416 6996 36420
rect 87284 36476 87348 36480
rect 87284 36420 87288 36476
rect 87288 36420 87344 36476
rect 87344 36420 87348 36476
rect 87284 36416 87348 36420
rect 87364 36476 87428 36480
rect 87364 36420 87368 36476
rect 87368 36420 87424 36476
rect 87424 36420 87428 36476
rect 87364 36416 87428 36420
rect 87444 36476 87508 36480
rect 87444 36420 87448 36476
rect 87448 36420 87504 36476
rect 87504 36420 87508 36476
rect 87444 36416 87508 36420
rect 87524 36476 87588 36480
rect 87524 36420 87528 36476
rect 87528 36420 87584 36476
rect 87584 36420 87588 36476
rect 87524 36416 87588 36420
rect 5956 35932 6020 35936
rect 5956 35876 5960 35932
rect 5960 35876 6016 35932
rect 6016 35876 6020 35932
rect 5956 35872 6020 35876
rect 6036 35932 6100 35936
rect 6036 35876 6040 35932
rect 6040 35876 6096 35932
rect 6096 35876 6100 35932
rect 6036 35872 6100 35876
rect 6116 35932 6180 35936
rect 6116 35876 6120 35932
rect 6120 35876 6176 35932
rect 6176 35876 6180 35932
rect 6116 35872 6180 35876
rect 6196 35932 6260 35936
rect 6196 35876 6200 35932
rect 6200 35876 6256 35932
rect 6256 35876 6260 35932
rect 6196 35872 6260 35876
rect 86548 35932 86612 35936
rect 86548 35876 86552 35932
rect 86552 35876 86608 35932
rect 86608 35876 86612 35932
rect 86548 35872 86612 35876
rect 86628 35932 86692 35936
rect 86628 35876 86632 35932
rect 86632 35876 86688 35932
rect 86688 35876 86692 35932
rect 86628 35872 86692 35876
rect 86708 35932 86772 35936
rect 86708 35876 86712 35932
rect 86712 35876 86768 35932
rect 86768 35876 86772 35932
rect 86708 35872 86772 35876
rect 86788 35932 86852 35936
rect 86788 35876 86792 35932
rect 86792 35876 86848 35932
rect 86848 35876 86852 35932
rect 86788 35872 86852 35876
rect 6692 35388 6756 35392
rect 6692 35332 6696 35388
rect 6696 35332 6752 35388
rect 6752 35332 6756 35388
rect 6692 35328 6756 35332
rect 6772 35388 6836 35392
rect 6772 35332 6776 35388
rect 6776 35332 6832 35388
rect 6832 35332 6836 35388
rect 6772 35328 6836 35332
rect 6852 35388 6916 35392
rect 6852 35332 6856 35388
rect 6856 35332 6912 35388
rect 6912 35332 6916 35388
rect 6852 35328 6916 35332
rect 6932 35388 6996 35392
rect 6932 35332 6936 35388
rect 6936 35332 6992 35388
rect 6992 35332 6996 35388
rect 6932 35328 6996 35332
rect 87284 35388 87348 35392
rect 87284 35332 87288 35388
rect 87288 35332 87344 35388
rect 87344 35332 87348 35388
rect 87284 35328 87348 35332
rect 87364 35388 87428 35392
rect 87364 35332 87368 35388
rect 87368 35332 87424 35388
rect 87424 35332 87428 35388
rect 87364 35328 87428 35332
rect 87444 35388 87508 35392
rect 87444 35332 87448 35388
rect 87448 35332 87504 35388
rect 87504 35332 87508 35388
rect 87444 35328 87508 35332
rect 87524 35388 87588 35392
rect 87524 35332 87528 35388
rect 87528 35332 87584 35388
rect 87584 35332 87588 35388
rect 87524 35328 87588 35332
rect 5956 34844 6020 34848
rect 5956 34788 5960 34844
rect 5960 34788 6016 34844
rect 6016 34788 6020 34844
rect 5956 34784 6020 34788
rect 6036 34844 6100 34848
rect 6036 34788 6040 34844
rect 6040 34788 6096 34844
rect 6096 34788 6100 34844
rect 6036 34784 6100 34788
rect 6116 34844 6180 34848
rect 6116 34788 6120 34844
rect 6120 34788 6176 34844
rect 6176 34788 6180 34844
rect 6116 34784 6180 34788
rect 6196 34844 6260 34848
rect 6196 34788 6200 34844
rect 6200 34788 6256 34844
rect 6256 34788 6260 34844
rect 6196 34784 6260 34788
rect 86548 34844 86612 34848
rect 86548 34788 86552 34844
rect 86552 34788 86608 34844
rect 86608 34788 86612 34844
rect 86548 34784 86612 34788
rect 86628 34844 86692 34848
rect 86628 34788 86632 34844
rect 86632 34788 86688 34844
rect 86688 34788 86692 34844
rect 86628 34784 86692 34788
rect 86708 34844 86772 34848
rect 86708 34788 86712 34844
rect 86712 34788 86768 34844
rect 86768 34788 86772 34844
rect 86708 34784 86772 34788
rect 86788 34844 86852 34848
rect 86788 34788 86792 34844
rect 86792 34788 86848 34844
rect 86848 34788 86852 34844
rect 86788 34784 86852 34788
rect 6692 34300 6756 34304
rect 6692 34244 6696 34300
rect 6696 34244 6752 34300
rect 6752 34244 6756 34300
rect 6692 34240 6756 34244
rect 6772 34300 6836 34304
rect 6772 34244 6776 34300
rect 6776 34244 6832 34300
rect 6832 34244 6836 34300
rect 6772 34240 6836 34244
rect 6852 34300 6916 34304
rect 6852 34244 6856 34300
rect 6856 34244 6912 34300
rect 6912 34244 6916 34300
rect 6852 34240 6916 34244
rect 6932 34300 6996 34304
rect 6932 34244 6936 34300
rect 6936 34244 6992 34300
rect 6992 34244 6996 34300
rect 6932 34240 6996 34244
rect 87284 34300 87348 34304
rect 87284 34244 87288 34300
rect 87288 34244 87344 34300
rect 87344 34244 87348 34300
rect 87284 34240 87348 34244
rect 87364 34300 87428 34304
rect 87364 34244 87368 34300
rect 87368 34244 87424 34300
rect 87424 34244 87428 34300
rect 87364 34240 87428 34244
rect 87444 34300 87508 34304
rect 87444 34244 87448 34300
rect 87448 34244 87504 34300
rect 87504 34244 87508 34300
rect 87444 34240 87508 34244
rect 87524 34300 87588 34304
rect 87524 34244 87528 34300
rect 87528 34244 87584 34300
rect 87584 34244 87588 34300
rect 87524 34240 87588 34244
rect 5956 33756 6020 33760
rect 5956 33700 5960 33756
rect 5960 33700 6016 33756
rect 6016 33700 6020 33756
rect 5956 33696 6020 33700
rect 6036 33756 6100 33760
rect 6036 33700 6040 33756
rect 6040 33700 6096 33756
rect 6096 33700 6100 33756
rect 6036 33696 6100 33700
rect 6116 33756 6180 33760
rect 6116 33700 6120 33756
rect 6120 33700 6176 33756
rect 6176 33700 6180 33756
rect 6116 33696 6180 33700
rect 6196 33756 6260 33760
rect 6196 33700 6200 33756
rect 6200 33700 6256 33756
rect 6256 33700 6260 33756
rect 6196 33696 6260 33700
rect 86548 33756 86612 33760
rect 86548 33700 86552 33756
rect 86552 33700 86608 33756
rect 86608 33700 86612 33756
rect 86548 33696 86612 33700
rect 86628 33756 86692 33760
rect 86628 33700 86632 33756
rect 86632 33700 86688 33756
rect 86688 33700 86692 33756
rect 86628 33696 86692 33700
rect 86708 33756 86772 33760
rect 86708 33700 86712 33756
rect 86712 33700 86768 33756
rect 86768 33700 86772 33756
rect 86708 33696 86772 33700
rect 86788 33756 86852 33760
rect 86788 33700 86792 33756
rect 86792 33700 86848 33756
rect 86848 33700 86852 33756
rect 86788 33696 86852 33700
rect 6692 33212 6756 33216
rect 6692 33156 6696 33212
rect 6696 33156 6752 33212
rect 6752 33156 6756 33212
rect 6692 33152 6756 33156
rect 6772 33212 6836 33216
rect 6772 33156 6776 33212
rect 6776 33156 6832 33212
rect 6832 33156 6836 33212
rect 6772 33152 6836 33156
rect 6852 33212 6916 33216
rect 6852 33156 6856 33212
rect 6856 33156 6912 33212
rect 6912 33156 6916 33212
rect 6852 33152 6916 33156
rect 6932 33212 6996 33216
rect 6932 33156 6936 33212
rect 6936 33156 6992 33212
rect 6992 33156 6996 33212
rect 6932 33152 6996 33156
rect 87284 33212 87348 33216
rect 87284 33156 87288 33212
rect 87288 33156 87344 33212
rect 87344 33156 87348 33212
rect 87284 33152 87348 33156
rect 87364 33212 87428 33216
rect 87364 33156 87368 33212
rect 87368 33156 87424 33212
rect 87424 33156 87428 33212
rect 87364 33152 87428 33156
rect 87444 33212 87508 33216
rect 87444 33156 87448 33212
rect 87448 33156 87504 33212
rect 87504 33156 87508 33212
rect 87444 33152 87508 33156
rect 87524 33212 87588 33216
rect 87524 33156 87528 33212
rect 87528 33156 87584 33212
rect 87584 33156 87588 33212
rect 87524 33152 87588 33156
rect 5956 32668 6020 32672
rect 5956 32612 5960 32668
rect 5960 32612 6016 32668
rect 6016 32612 6020 32668
rect 5956 32608 6020 32612
rect 6036 32668 6100 32672
rect 6036 32612 6040 32668
rect 6040 32612 6096 32668
rect 6096 32612 6100 32668
rect 6036 32608 6100 32612
rect 6116 32668 6180 32672
rect 6116 32612 6120 32668
rect 6120 32612 6176 32668
rect 6176 32612 6180 32668
rect 6116 32608 6180 32612
rect 6196 32668 6260 32672
rect 6196 32612 6200 32668
rect 6200 32612 6256 32668
rect 6256 32612 6260 32668
rect 6196 32608 6260 32612
rect 86548 32668 86612 32672
rect 86548 32612 86552 32668
rect 86552 32612 86608 32668
rect 86608 32612 86612 32668
rect 86548 32608 86612 32612
rect 86628 32668 86692 32672
rect 86628 32612 86632 32668
rect 86632 32612 86688 32668
rect 86688 32612 86692 32668
rect 86628 32608 86692 32612
rect 86708 32668 86772 32672
rect 86708 32612 86712 32668
rect 86712 32612 86768 32668
rect 86768 32612 86772 32668
rect 86708 32608 86772 32612
rect 86788 32668 86852 32672
rect 86788 32612 86792 32668
rect 86792 32612 86848 32668
rect 86848 32612 86852 32668
rect 86788 32608 86852 32612
rect 6692 32124 6756 32128
rect 6692 32068 6696 32124
rect 6696 32068 6752 32124
rect 6752 32068 6756 32124
rect 6692 32064 6756 32068
rect 6772 32124 6836 32128
rect 6772 32068 6776 32124
rect 6776 32068 6832 32124
rect 6832 32068 6836 32124
rect 6772 32064 6836 32068
rect 6852 32124 6916 32128
rect 6852 32068 6856 32124
rect 6856 32068 6912 32124
rect 6912 32068 6916 32124
rect 6852 32064 6916 32068
rect 6932 32124 6996 32128
rect 6932 32068 6936 32124
rect 6936 32068 6992 32124
rect 6992 32068 6996 32124
rect 6932 32064 6996 32068
rect 87284 32124 87348 32128
rect 87284 32068 87288 32124
rect 87288 32068 87344 32124
rect 87344 32068 87348 32124
rect 87284 32064 87348 32068
rect 87364 32124 87428 32128
rect 87364 32068 87368 32124
rect 87368 32068 87424 32124
rect 87424 32068 87428 32124
rect 87364 32064 87428 32068
rect 87444 32124 87508 32128
rect 87444 32068 87448 32124
rect 87448 32068 87504 32124
rect 87504 32068 87508 32124
rect 87444 32064 87508 32068
rect 87524 32124 87588 32128
rect 87524 32068 87528 32124
rect 87528 32068 87584 32124
rect 87584 32068 87588 32124
rect 87524 32064 87588 32068
rect 5956 31580 6020 31584
rect 5956 31524 5960 31580
rect 5960 31524 6016 31580
rect 6016 31524 6020 31580
rect 5956 31520 6020 31524
rect 6036 31580 6100 31584
rect 6036 31524 6040 31580
rect 6040 31524 6096 31580
rect 6096 31524 6100 31580
rect 6036 31520 6100 31524
rect 6116 31580 6180 31584
rect 6116 31524 6120 31580
rect 6120 31524 6176 31580
rect 6176 31524 6180 31580
rect 6116 31520 6180 31524
rect 6196 31580 6260 31584
rect 6196 31524 6200 31580
rect 6200 31524 6256 31580
rect 6256 31524 6260 31580
rect 6196 31520 6260 31524
rect 86548 31580 86612 31584
rect 86548 31524 86552 31580
rect 86552 31524 86608 31580
rect 86608 31524 86612 31580
rect 86548 31520 86612 31524
rect 86628 31580 86692 31584
rect 86628 31524 86632 31580
rect 86632 31524 86688 31580
rect 86688 31524 86692 31580
rect 86628 31520 86692 31524
rect 86708 31580 86772 31584
rect 86708 31524 86712 31580
rect 86712 31524 86768 31580
rect 86768 31524 86772 31580
rect 86708 31520 86772 31524
rect 86788 31580 86852 31584
rect 86788 31524 86792 31580
rect 86792 31524 86848 31580
rect 86848 31524 86852 31580
rect 86788 31520 86852 31524
rect 6692 31036 6756 31040
rect 6692 30980 6696 31036
rect 6696 30980 6752 31036
rect 6752 30980 6756 31036
rect 6692 30976 6756 30980
rect 6772 31036 6836 31040
rect 6772 30980 6776 31036
rect 6776 30980 6832 31036
rect 6832 30980 6836 31036
rect 6772 30976 6836 30980
rect 6852 31036 6916 31040
rect 6852 30980 6856 31036
rect 6856 30980 6912 31036
rect 6912 30980 6916 31036
rect 6852 30976 6916 30980
rect 6932 31036 6996 31040
rect 6932 30980 6936 31036
rect 6936 30980 6992 31036
rect 6992 30980 6996 31036
rect 6932 30976 6996 30980
rect 87284 31036 87348 31040
rect 87284 30980 87288 31036
rect 87288 30980 87344 31036
rect 87344 30980 87348 31036
rect 87284 30976 87348 30980
rect 87364 31036 87428 31040
rect 87364 30980 87368 31036
rect 87368 30980 87424 31036
rect 87424 30980 87428 31036
rect 87364 30976 87428 30980
rect 87444 31036 87508 31040
rect 87444 30980 87448 31036
rect 87448 30980 87504 31036
rect 87504 30980 87508 31036
rect 87444 30976 87508 30980
rect 87524 31036 87588 31040
rect 87524 30980 87528 31036
rect 87528 30980 87584 31036
rect 87584 30980 87588 31036
rect 87524 30976 87588 30980
rect 5956 30492 6020 30496
rect 5956 30436 5960 30492
rect 5960 30436 6016 30492
rect 6016 30436 6020 30492
rect 5956 30432 6020 30436
rect 6036 30492 6100 30496
rect 6036 30436 6040 30492
rect 6040 30436 6096 30492
rect 6096 30436 6100 30492
rect 6036 30432 6100 30436
rect 6116 30492 6180 30496
rect 6116 30436 6120 30492
rect 6120 30436 6176 30492
rect 6176 30436 6180 30492
rect 6116 30432 6180 30436
rect 6196 30492 6260 30496
rect 6196 30436 6200 30492
rect 6200 30436 6256 30492
rect 6256 30436 6260 30492
rect 6196 30432 6260 30436
rect 86548 30492 86612 30496
rect 86548 30436 86552 30492
rect 86552 30436 86608 30492
rect 86608 30436 86612 30492
rect 86548 30432 86612 30436
rect 86628 30492 86692 30496
rect 86628 30436 86632 30492
rect 86632 30436 86688 30492
rect 86688 30436 86692 30492
rect 86628 30432 86692 30436
rect 86708 30492 86772 30496
rect 86708 30436 86712 30492
rect 86712 30436 86768 30492
rect 86768 30436 86772 30492
rect 86708 30432 86772 30436
rect 86788 30492 86852 30496
rect 86788 30436 86792 30492
rect 86792 30436 86848 30492
rect 86848 30436 86852 30492
rect 86788 30432 86852 30436
rect 6692 29948 6756 29952
rect 6692 29892 6696 29948
rect 6696 29892 6752 29948
rect 6752 29892 6756 29948
rect 6692 29888 6756 29892
rect 6772 29948 6836 29952
rect 6772 29892 6776 29948
rect 6776 29892 6832 29948
rect 6832 29892 6836 29948
rect 6772 29888 6836 29892
rect 6852 29948 6916 29952
rect 6852 29892 6856 29948
rect 6856 29892 6912 29948
rect 6912 29892 6916 29948
rect 6852 29888 6916 29892
rect 6932 29948 6996 29952
rect 6932 29892 6936 29948
rect 6936 29892 6992 29948
rect 6992 29892 6996 29948
rect 6932 29888 6996 29892
rect 87284 29948 87348 29952
rect 87284 29892 87288 29948
rect 87288 29892 87344 29948
rect 87344 29892 87348 29948
rect 87284 29888 87348 29892
rect 87364 29948 87428 29952
rect 87364 29892 87368 29948
rect 87368 29892 87424 29948
rect 87424 29892 87428 29948
rect 87364 29888 87428 29892
rect 87444 29948 87508 29952
rect 87444 29892 87448 29948
rect 87448 29892 87504 29948
rect 87504 29892 87508 29948
rect 87444 29888 87508 29892
rect 87524 29948 87588 29952
rect 87524 29892 87528 29948
rect 87528 29892 87584 29948
rect 87584 29892 87588 29948
rect 87524 29888 87588 29892
rect 5956 29404 6020 29408
rect 5956 29348 5960 29404
rect 5960 29348 6016 29404
rect 6016 29348 6020 29404
rect 5956 29344 6020 29348
rect 6036 29404 6100 29408
rect 6036 29348 6040 29404
rect 6040 29348 6096 29404
rect 6096 29348 6100 29404
rect 6036 29344 6100 29348
rect 6116 29404 6180 29408
rect 6116 29348 6120 29404
rect 6120 29348 6176 29404
rect 6176 29348 6180 29404
rect 6116 29344 6180 29348
rect 6196 29404 6260 29408
rect 6196 29348 6200 29404
rect 6200 29348 6256 29404
rect 6256 29348 6260 29404
rect 6196 29344 6260 29348
rect 86548 29404 86612 29408
rect 86548 29348 86552 29404
rect 86552 29348 86608 29404
rect 86608 29348 86612 29404
rect 86548 29344 86612 29348
rect 86628 29404 86692 29408
rect 86628 29348 86632 29404
rect 86632 29348 86688 29404
rect 86688 29348 86692 29404
rect 86628 29344 86692 29348
rect 86708 29404 86772 29408
rect 86708 29348 86712 29404
rect 86712 29348 86768 29404
rect 86768 29348 86772 29404
rect 86708 29344 86772 29348
rect 86788 29404 86852 29408
rect 86788 29348 86792 29404
rect 86792 29348 86848 29404
rect 86848 29348 86852 29404
rect 86788 29344 86852 29348
rect 6692 28860 6756 28864
rect 6692 28804 6696 28860
rect 6696 28804 6752 28860
rect 6752 28804 6756 28860
rect 6692 28800 6756 28804
rect 6772 28860 6836 28864
rect 6772 28804 6776 28860
rect 6776 28804 6832 28860
rect 6832 28804 6836 28860
rect 6772 28800 6836 28804
rect 6852 28860 6916 28864
rect 6852 28804 6856 28860
rect 6856 28804 6912 28860
rect 6912 28804 6916 28860
rect 6852 28800 6916 28804
rect 6932 28860 6996 28864
rect 6932 28804 6936 28860
rect 6936 28804 6992 28860
rect 6992 28804 6996 28860
rect 6932 28800 6996 28804
rect 87284 28860 87348 28864
rect 87284 28804 87288 28860
rect 87288 28804 87344 28860
rect 87344 28804 87348 28860
rect 87284 28800 87348 28804
rect 87364 28860 87428 28864
rect 87364 28804 87368 28860
rect 87368 28804 87424 28860
rect 87424 28804 87428 28860
rect 87364 28800 87428 28804
rect 87444 28860 87508 28864
rect 87444 28804 87448 28860
rect 87448 28804 87504 28860
rect 87504 28804 87508 28860
rect 87444 28800 87508 28804
rect 87524 28860 87588 28864
rect 87524 28804 87528 28860
rect 87528 28804 87584 28860
rect 87584 28804 87588 28860
rect 87524 28800 87588 28804
rect 5956 28316 6020 28320
rect 5956 28260 5960 28316
rect 5960 28260 6016 28316
rect 6016 28260 6020 28316
rect 5956 28256 6020 28260
rect 6036 28316 6100 28320
rect 6036 28260 6040 28316
rect 6040 28260 6096 28316
rect 6096 28260 6100 28316
rect 6036 28256 6100 28260
rect 6116 28316 6180 28320
rect 6116 28260 6120 28316
rect 6120 28260 6176 28316
rect 6176 28260 6180 28316
rect 6116 28256 6180 28260
rect 6196 28316 6260 28320
rect 6196 28260 6200 28316
rect 6200 28260 6256 28316
rect 6256 28260 6260 28316
rect 6196 28256 6260 28260
rect 86548 28316 86612 28320
rect 86548 28260 86552 28316
rect 86552 28260 86608 28316
rect 86608 28260 86612 28316
rect 86548 28256 86612 28260
rect 86628 28316 86692 28320
rect 86628 28260 86632 28316
rect 86632 28260 86688 28316
rect 86688 28260 86692 28316
rect 86628 28256 86692 28260
rect 86708 28316 86772 28320
rect 86708 28260 86712 28316
rect 86712 28260 86768 28316
rect 86768 28260 86772 28316
rect 86708 28256 86772 28260
rect 86788 28316 86852 28320
rect 86788 28260 86792 28316
rect 86792 28260 86848 28316
rect 86848 28260 86852 28316
rect 86788 28256 86852 28260
rect 6692 27772 6756 27776
rect 6692 27716 6696 27772
rect 6696 27716 6752 27772
rect 6752 27716 6756 27772
rect 6692 27712 6756 27716
rect 6772 27772 6836 27776
rect 6772 27716 6776 27772
rect 6776 27716 6832 27772
rect 6832 27716 6836 27772
rect 6772 27712 6836 27716
rect 6852 27772 6916 27776
rect 6852 27716 6856 27772
rect 6856 27716 6912 27772
rect 6912 27716 6916 27772
rect 6852 27712 6916 27716
rect 6932 27772 6996 27776
rect 6932 27716 6936 27772
rect 6936 27716 6992 27772
rect 6992 27716 6996 27772
rect 6932 27712 6996 27716
rect 87284 27772 87348 27776
rect 87284 27716 87288 27772
rect 87288 27716 87344 27772
rect 87344 27716 87348 27772
rect 87284 27712 87348 27716
rect 87364 27772 87428 27776
rect 87364 27716 87368 27772
rect 87368 27716 87424 27772
rect 87424 27716 87428 27772
rect 87364 27712 87428 27716
rect 87444 27772 87508 27776
rect 87444 27716 87448 27772
rect 87448 27716 87504 27772
rect 87504 27716 87508 27772
rect 87444 27712 87508 27716
rect 87524 27772 87588 27776
rect 87524 27716 87528 27772
rect 87528 27716 87584 27772
rect 87584 27716 87588 27772
rect 87524 27712 87588 27716
rect 5956 27228 6020 27232
rect 5956 27172 5960 27228
rect 5960 27172 6016 27228
rect 6016 27172 6020 27228
rect 5956 27168 6020 27172
rect 6036 27228 6100 27232
rect 6036 27172 6040 27228
rect 6040 27172 6096 27228
rect 6096 27172 6100 27228
rect 6036 27168 6100 27172
rect 6116 27228 6180 27232
rect 6116 27172 6120 27228
rect 6120 27172 6176 27228
rect 6176 27172 6180 27228
rect 6116 27168 6180 27172
rect 6196 27228 6260 27232
rect 6196 27172 6200 27228
rect 6200 27172 6256 27228
rect 6256 27172 6260 27228
rect 6196 27168 6260 27172
rect 86548 27228 86612 27232
rect 86548 27172 86552 27228
rect 86552 27172 86608 27228
rect 86608 27172 86612 27228
rect 86548 27168 86612 27172
rect 86628 27228 86692 27232
rect 86628 27172 86632 27228
rect 86632 27172 86688 27228
rect 86688 27172 86692 27228
rect 86628 27168 86692 27172
rect 86708 27228 86772 27232
rect 86708 27172 86712 27228
rect 86712 27172 86768 27228
rect 86768 27172 86772 27228
rect 86708 27168 86772 27172
rect 86788 27228 86852 27232
rect 86788 27172 86792 27228
rect 86792 27172 86848 27228
rect 86848 27172 86852 27228
rect 86788 27168 86852 27172
rect 6692 26684 6756 26688
rect 6692 26628 6696 26684
rect 6696 26628 6752 26684
rect 6752 26628 6756 26684
rect 6692 26624 6756 26628
rect 6772 26684 6836 26688
rect 6772 26628 6776 26684
rect 6776 26628 6832 26684
rect 6832 26628 6836 26684
rect 6772 26624 6836 26628
rect 6852 26684 6916 26688
rect 6852 26628 6856 26684
rect 6856 26628 6912 26684
rect 6912 26628 6916 26684
rect 6852 26624 6916 26628
rect 6932 26684 6996 26688
rect 6932 26628 6936 26684
rect 6936 26628 6992 26684
rect 6992 26628 6996 26684
rect 6932 26624 6996 26628
rect 87284 26684 87348 26688
rect 87284 26628 87288 26684
rect 87288 26628 87344 26684
rect 87344 26628 87348 26684
rect 87284 26624 87348 26628
rect 87364 26684 87428 26688
rect 87364 26628 87368 26684
rect 87368 26628 87424 26684
rect 87424 26628 87428 26684
rect 87364 26624 87428 26628
rect 87444 26684 87508 26688
rect 87444 26628 87448 26684
rect 87448 26628 87504 26684
rect 87504 26628 87508 26684
rect 87444 26624 87508 26628
rect 87524 26684 87588 26688
rect 87524 26628 87528 26684
rect 87528 26628 87584 26684
rect 87584 26628 87588 26684
rect 87524 26624 87588 26628
rect 5956 26140 6020 26144
rect 5956 26084 5960 26140
rect 5960 26084 6016 26140
rect 6016 26084 6020 26140
rect 5956 26080 6020 26084
rect 6036 26140 6100 26144
rect 6036 26084 6040 26140
rect 6040 26084 6096 26140
rect 6096 26084 6100 26140
rect 6036 26080 6100 26084
rect 6116 26140 6180 26144
rect 6116 26084 6120 26140
rect 6120 26084 6176 26140
rect 6176 26084 6180 26140
rect 6116 26080 6180 26084
rect 6196 26140 6260 26144
rect 6196 26084 6200 26140
rect 6200 26084 6256 26140
rect 6256 26084 6260 26140
rect 6196 26080 6260 26084
rect 86548 26140 86612 26144
rect 86548 26084 86552 26140
rect 86552 26084 86608 26140
rect 86608 26084 86612 26140
rect 86548 26080 86612 26084
rect 86628 26140 86692 26144
rect 86628 26084 86632 26140
rect 86632 26084 86688 26140
rect 86688 26084 86692 26140
rect 86628 26080 86692 26084
rect 86708 26140 86772 26144
rect 86708 26084 86712 26140
rect 86712 26084 86768 26140
rect 86768 26084 86772 26140
rect 86708 26080 86772 26084
rect 86788 26140 86852 26144
rect 86788 26084 86792 26140
rect 86792 26084 86848 26140
rect 86848 26084 86852 26140
rect 86788 26080 86852 26084
rect 6692 25596 6756 25600
rect 6692 25540 6696 25596
rect 6696 25540 6752 25596
rect 6752 25540 6756 25596
rect 6692 25536 6756 25540
rect 6772 25596 6836 25600
rect 6772 25540 6776 25596
rect 6776 25540 6832 25596
rect 6832 25540 6836 25596
rect 6772 25536 6836 25540
rect 6852 25596 6916 25600
rect 6852 25540 6856 25596
rect 6856 25540 6912 25596
rect 6912 25540 6916 25596
rect 6852 25536 6916 25540
rect 6932 25596 6996 25600
rect 6932 25540 6936 25596
rect 6936 25540 6992 25596
rect 6992 25540 6996 25596
rect 6932 25536 6996 25540
rect 87284 25596 87348 25600
rect 87284 25540 87288 25596
rect 87288 25540 87344 25596
rect 87344 25540 87348 25596
rect 87284 25536 87348 25540
rect 87364 25596 87428 25600
rect 87364 25540 87368 25596
rect 87368 25540 87424 25596
rect 87424 25540 87428 25596
rect 87364 25536 87428 25540
rect 87444 25596 87508 25600
rect 87444 25540 87448 25596
rect 87448 25540 87504 25596
rect 87504 25540 87508 25596
rect 87444 25536 87508 25540
rect 87524 25596 87588 25600
rect 87524 25540 87528 25596
rect 87528 25540 87584 25596
rect 87584 25540 87588 25596
rect 87524 25536 87588 25540
rect 5956 25052 6020 25056
rect 5956 24996 5960 25052
rect 5960 24996 6016 25052
rect 6016 24996 6020 25052
rect 5956 24992 6020 24996
rect 6036 25052 6100 25056
rect 6036 24996 6040 25052
rect 6040 24996 6096 25052
rect 6096 24996 6100 25052
rect 6036 24992 6100 24996
rect 6116 25052 6180 25056
rect 6116 24996 6120 25052
rect 6120 24996 6176 25052
rect 6176 24996 6180 25052
rect 6116 24992 6180 24996
rect 6196 25052 6260 25056
rect 6196 24996 6200 25052
rect 6200 24996 6256 25052
rect 6256 24996 6260 25052
rect 6196 24992 6260 24996
rect 86548 25052 86612 25056
rect 86548 24996 86552 25052
rect 86552 24996 86608 25052
rect 86608 24996 86612 25052
rect 86548 24992 86612 24996
rect 86628 25052 86692 25056
rect 86628 24996 86632 25052
rect 86632 24996 86688 25052
rect 86688 24996 86692 25052
rect 86628 24992 86692 24996
rect 86708 25052 86772 25056
rect 86708 24996 86712 25052
rect 86712 24996 86768 25052
rect 86768 24996 86772 25052
rect 86708 24992 86772 24996
rect 86788 25052 86852 25056
rect 86788 24996 86792 25052
rect 86792 24996 86848 25052
rect 86848 24996 86852 25052
rect 86788 24992 86852 24996
rect 6692 24508 6756 24512
rect 6692 24452 6696 24508
rect 6696 24452 6752 24508
rect 6752 24452 6756 24508
rect 6692 24448 6756 24452
rect 6772 24508 6836 24512
rect 6772 24452 6776 24508
rect 6776 24452 6832 24508
rect 6832 24452 6836 24508
rect 6772 24448 6836 24452
rect 6852 24508 6916 24512
rect 6852 24452 6856 24508
rect 6856 24452 6912 24508
rect 6912 24452 6916 24508
rect 6852 24448 6916 24452
rect 6932 24508 6996 24512
rect 6932 24452 6936 24508
rect 6936 24452 6992 24508
rect 6992 24452 6996 24508
rect 6932 24448 6996 24452
rect 87284 24508 87348 24512
rect 87284 24452 87288 24508
rect 87288 24452 87344 24508
rect 87344 24452 87348 24508
rect 87284 24448 87348 24452
rect 87364 24508 87428 24512
rect 87364 24452 87368 24508
rect 87368 24452 87424 24508
rect 87424 24452 87428 24508
rect 87364 24448 87428 24452
rect 87444 24508 87508 24512
rect 87444 24452 87448 24508
rect 87448 24452 87504 24508
rect 87504 24452 87508 24508
rect 87444 24448 87508 24452
rect 87524 24508 87588 24512
rect 87524 24452 87528 24508
rect 87528 24452 87584 24508
rect 87584 24452 87588 24508
rect 87524 24448 87588 24452
rect 5956 23964 6020 23968
rect 5956 23908 5960 23964
rect 5960 23908 6016 23964
rect 6016 23908 6020 23964
rect 5956 23904 6020 23908
rect 6036 23964 6100 23968
rect 6036 23908 6040 23964
rect 6040 23908 6096 23964
rect 6096 23908 6100 23964
rect 6036 23904 6100 23908
rect 6116 23964 6180 23968
rect 6116 23908 6120 23964
rect 6120 23908 6176 23964
rect 6176 23908 6180 23964
rect 6116 23904 6180 23908
rect 6196 23964 6260 23968
rect 6196 23908 6200 23964
rect 6200 23908 6256 23964
rect 6256 23908 6260 23964
rect 6196 23904 6260 23908
rect 86548 23964 86612 23968
rect 86548 23908 86552 23964
rect 86552 23908 86608 23964
rect 86608 23908 86612 23964
rect 86548 23904 86612 23908
rect 86628 23964 86692 23968
rect 86628 23908 86632 23964
rect 86632 23908 86688 23964
rect 86688 23908 86692 23964
rect 86628 23904 86692 23908
rect 86708 23964 86772 23968
rect 86708 23908 86712 23964
rect 86712 23908 86768 23964
rect 86768 23908 86772 23964
rect 86708 23904 86772 23908
rect 86788 23964 86852 23968
rect 86788 23908 86792 23964
rect 86792 23908 86848 23964
rect 86848 23908 86852 23964
rect 86788 23904 86852 23908
rect 6692 23420 6756 23424
rect 6692 23364 6696 23420
rect 6696 23364 6752 23420
rect 6752 23364 6756 23420
rect 6692 23360 6756 23364
rect 6772 23420 6836 23424
rect 6772 23364 6776 23420
rect 6776 23364 6832 23420
rect 6832 23364 6836 23420
rect 6772 23360 6836 23364
rect 6852 23420 6916 23424
rect 6852 23364 6856 23420
rect 6856 23364 6912 23420
rect 6912 23364 6916 23420
rect 6852 23360 6916 23364
rect 6932 23420 6996 23424
rect 6932 23364 6936 23420
rect 6936 23364 6992 23420
rect 6992 23364 6996 23420
rect 6932 23360 6996 23364
rect 87284 23420 87348 23424
rect 87284 23364 87288 23420
rect 87288 23364 87344 23420
rect 87344 23364 87348 23420
rect 87284 23360 87348 23364
rect 87364 23420 87428 23424
rect 87364 23364 87368 23420
rect 87368 23364 87424 23420
rect 87424 23364 87428 23420
rect 87364 23360 87428 23364
rect 87444 23420 87508 23424
rect 87444 23364 87448 23420
rect 87448 23364 87504 23420
rect 87504 23364 87508 23420
rect 87444 23360 87508 23364
rect 87524 23420 87588 23424
rect 87524 23364 87528 23420
rect 87528 23364 87584 23420
rect 87584 23364 87588 23420
rect 87524 23360 87588 23364
rect 5956 22876 6020 22880
rect 5956 22820 5960 22876
rect 5960 22820 6016 22876
rect 6016 22820 6020 22876
rect 5956 22816 6020 22820
rect 6036 22876 6100 22880
rect 6036 22820 6040 22876
rect 6040 22820 6096 22876
rect 6096 22820 6100 22876
rect 6036 22816 6100 22820
rect 6116 22876 6180 22880
rect 6116 22820 6120 22876
rect 6120 22820 6176 22876
rect 6176 22820 6180 22876
rect 6116 22816 6180 22820
rect 6196 22876 6260 22880
rect 6196 22820 6200 22876
rect 6200 22820 6256 22876
rect 6256 22820 6260 22876
rect 6196 22816 6260 22820
rect 86548 22876 86612 22880
rect 86548 22820 86552 22876
rect 86552 22820 86608 22876
rect 86608 22820 86612 22876
rect 86548 22816 86612 22820
rect 86628 22876 86692 22880
rect 86628 22820 86632 22876
rect 86632 22820 86688 22876
rect 86688 22820 86692 22876
rect 86628 22816 86692 22820
rect 86708 22876 86772 22880
rect 86708 22820 86712 22876
rect 86712 22820 86768 22876
rect 86768 22820 86772 22876
rect 86708 22816 86772 22820
rect 86788 22876 86852 22880
rect 86788 22820 86792 22876
rect 86792 22820 86848 22876
rect 86848 22820 86852 22876
rect 86788 22816 86852 22820
rect 6692 22332 6756 22336
rect 6692 22276 6696 22332
rect 6696 22276 6752 22332
rect 6752 22276 6756 22332
rect 6692 22272 6756 22276
rect 6772 22332 6836 22336
rect 6772 22276 6776 22332
rect 6776 22276 6832 22332
rect 6832 22276 6836 22332
rect 6772 22272 6836 22276
rect 6852 22332 6916 22336
rect 6852 22276 6856 22332
rect 6856 22276 6912 22332
rect 6912 22276 6916 22332
rect 6852 22272 6916 22276
rect 6932 22332 6996 22336
rect 6932 22276 6936 22332
rect 6936 22276 6992 22332
rect 6992 22276 6996 22332
rect 6932 22272 6996 22276
rect 87284 22332 87348 22336
rect 87284 22276 87288 22332
rect 87288 22276 87344 22332
rect 87344 22276 87348 22332
rect 87284 22272 87348 22276
rect 87364 22332 87428 22336
rect 87364 22276 87368 22332
rect 87368 22276 87424 22332
rect 87424 22276 87428 22332
rect 87364 22272 87428 22276
rect 87444 22332 87508 22336
rect 87444 22276 87448 22332
rect 87448 22276 87504 22332
rect 87504 22276 87508 22332
rect 87444 22272 87508 22276
rect 87524 22332 87588 22336
rect 87524 22276 87528 22332
rect 87528 22276 87584 22332
rect 87584 22276 87588 22332
rect 87524 22272 87588 22276
rect 5956 21788 6020 21792
rect 5956 21732 5960 21788
rect 5960 21732 6016 21788
rect 6016 21732 6020 21788
rect 5956 21728 6020 21732
rect 6036 21788 6100 21792
rect 6036 21732 6040 21788
rect 6040 21732 6096 21788
rect 6096 21732 6100 21788
rect 6036 21728 6100 21732
rect 6116 21788 6180 21792
rect 6116 21732 6120 21788
rect 6120 21732 6176 21788
rect 6176 21732 6180 21788
rect 6116 21728 6180 21732
rect 6196 21788 6260 21792
rect 6196 21732 6200 21788
rect 6200 21732 6256 21788
rect 6256 21732 6260 21788
rect 6196 21728 6260 21732
rect 86548 21788 86612 21792
rect 86548 21732 86552 21788
rect 86552 21732 86608 21788
rect 86608 21732 86612 21788
rect 86548 21728 86612 21732
rect 86628 21788 86692 21792
rect 86628 21732 86632 21788
rect 86632 21732 86688 21788
rect 86688 21732 86692 21788
rect 86628 21728 86692 21732
rect 86708 21788 86772 21792
rect 86708 21732 86712 21788
rect 86712 21732 86768 21788
rect 86768 21732 86772 21788
rect 86708 21728 86772 21732
rect 86788 21788 86852 21792
rect 86788 21732 86792 21788
rect 86792 21732 86848 21788
rect 86848 21732 86852 21788
rect 86788 21728 86852 21732
rect 6692 21244 6756 21248
rect 6692 21188 6696 21244
rect 6696 21188 6752 21244
rect 6752 21188 6756 21244
rect 6692 21184 6756 21188
rect 6772 21244 6836 21248
rect 6772 21188 6776 21244
rect 6776 21188 6832 21244
rect 6832 21188 6836 21244
rect 6772 21184 6836 21188
rect 6852 21244 6916 21248
rect 6852 21188 6856 21244
rect 6856 21188 6912 21244
rect 6912 21188 6916 21244
rect 6852 21184 6916 21188
rect 6932 21244 6996 21248
rect 6932 21188 6936 21244
rect 6936 21188 6992 21244
rect 6992 21188 6996 21244
rect 6932 21184 6996 21188
rect 87284 21244 87348 21248
rect 87284 21188 87288 21244
rect 87288 21188 87344 21244
rect 87344 21188 87348 21244
rect 87284 21184 87348 21188
rect 87364 21244 87428 21248
rect 87364 21188 87368 21244
rect 87368 21188 87424 21244
rect 87424 21188 87428 21244
rect 87364 21184 87428 21188
rect 87444 21244 87508 21248
rect 87444 21188 87448 21244
rect 87448 21188 87504 21244
rect 87504 21188 87508 21244
rect 87444 21184 87508 21188
rect 87524 21244 87588 21248
rect 87524 21188 87528 21244
rect 87528 21188 87584 21244
rect 87584 21188 87588 21244
rect 87524 21184 87588 21188
rect 5956 20700 6020 20704
rect 5956 20644 5960 20700
rect 5960 20644 6016 20700
rect 6016 20644 6020 20700
rect 5956 20640 6020 20644
rect 6036 20700 6100 20704
rect 6036 20644 6040 20700
rect 6040 20644 6096 20700
rect 6096 20644 6100 20700
rect 6036 20640 6100 20644
rect 6116 20700 6180 20704
rect 6116 20644 6120 20700
rect 6120 20644 6176 20700
rect 6176 20644 6180 20700
rect 6116 20640 6180 20644
rect 6196 20700 6260 20704
rect 6196 20644 6200 20700
rect 6200 20644 6256 20700
rect 6256 20644 6260 20700
rect 6196 20640 6260 20644
rect 86548 20700 86612 20704
rect 86548 20644 86552 20700
rect 86552 20644 86608 20700
rect 86608 20644 86612 20700
rect 86548 20640 86612 20644
rect 86628 20700 86692 20704
rect 86628 20644 86632 20700
rect 86632 20644 86688 20700
rect 86688 20644 86692 20700
rect 86628 20640 86692 20644
rect 86708 20700 86772 20704
rect 86708 20644 86712 20700
rect 86712 20644 86768 20700
rect 86768 20644 86772 20700
rect 86708 20640 86772 20644
rect 86788 20700 86852 20704
rect 86788 20644 86792 20700
rect 86792 20644 86848 20700
rect 86848 20644 86852 20700
rect 86788 20640 86852 20644
rect 6692 20156 6756 20160
rect 6692 20100 6696 20156
rect 6696 20100 6752 20156
rect 6752 20100 6756 20156
rect 6692 20096 6756 20100
rect 6772 20156 6836 20160
rect 6772 20100 6776 20156
rect 6776 20100 6832 20156
rect 6832 20100 6836 20156
rect 6772 20096 6836 20100
rect 6852 20156 6916 20160
rect 6852 20100 6856 20156
rect 6856 20100 6912 20156
rect 6912 20100 6916 20156
rect 6852 20096 6916 20100
rect 6932 20156 6996 20160
rect 6932 20100 6936 20156
rect 6936 20100 6992 20156
rect 6992 20100 6996 20156
rect 6932 20096 6996 20100
rect 87284 20156 87348 20160
rect 87284 20100 87288 20156
rect 87288 20100 87344 20156
rect 87344 20100 87348 20156
rect 87284 20096 87348 20100
rect 87364 20156 87428 20160
rect 87364 20100 87368 20156
rect 87368 20100 87424 20156
rect 87424 20100 87428 20156
rect 87364 20096 87428 20100
rect 87444 20156 87508 20160
rect 87444 20100 87448 20156
rect 87448 20100 87504 20156
rect 87504 20100 87508 20156
rect 87444 20096 87508 20100
rect 87524 20156 87588 20160
rect 87524 20100 87528 20156
rect 87528 20100 87584 20156
rect 87584 20100 87588 20156
rect 87524 20096 87588 20100
rect 5956 19612 6020 19616
rect 5956 19556 5960 19612
rect 5960 19556 6016 19612
rect 6016 19556 6020 19612
rect 5956 19552 6020 19556
rect 6036 19612 6100 19616
rect 6036 19556 6040 19612
rect 6040 19556 6096 19612
rect 6096 19556 6100 19612
rect 6036 19552 6100 19556
rect 6116 19612 6180 19616
rect 6116 19556 6120 19612
rect 6120 19556 6176 19612
rect 6176 19556 6180 19612
rect 6116 19552 6180 19556
rect 6196 19612 6260 19616
rect 6196 19556 6200 19612
rect 6200 19556 6256 19612
rect 6256 19556 6260 19612
rect 6196 19552 6260 19556
rect 86548 19612 86612 19616
rect 86548 19556 86552 19612
rect 86552 19556 86608 19612
rect 86608 19556 86612 19612
rect 86548 19552 86612 19556
rect 86628 19612 86692 19616
rect 86628 19556 86632 19612
rect 86632 19556 86688 19612
rect 86688 19556 86692 19612
rect 86628 19552 86692 19556
rect 86708 19612 86772 19616
rect 86708 19556 86712 19612
rect 86712 19556 86768 19612
rect 86768 19556 86772 19612
rect 86708 19552 86772 19556
rect 86788 19612 86852 19616
rect 86788 19556 86792 19612
rect 86792 19556 86848 19612
rect 86848 19556 86852 19612
rect 86788 19552 86852 19556
rect 6692 19068 6756 19072
rect 6692 19012 6696 19068
rect 6696 19012 6752 19068
rect 6752 19012 6756 19068
rect 6692 19008 6756 19012
rect 6772 19068 6836 19072
rect 6772 19012 6776 19068
rect 6776 19012 6832 19068
rect 6832 19012 6836 19068
rect 6772 19008 6836 19012
rect 6852 19068 6916 19072
rect 6852 19012 6856 19068
rect 6856 19012 6912 19068
rect 6912 19012 6916 19068
rect 6852 19008 6916 19012
rect 6932 19068 6996 19072
rect 6932 19012 6936 19068
rect 6936 19012 6992 19068
rect 6992 19012 6996 19068
rect 6932 19008 6996 19012
rect 87284 19068 87348 19072
rect 87284 19012 87288 19068
rect 87288 19012 87344 19068
rect 87344 19012 87348 19068
rect 87284 19008 87348 19012
rect 87364 19068 87428 19072
rect 87364 19012 87368 19068
rect 87368 19012 87424 19068
rect 87424 19012 87428 19068
rect 87364 19008 87428 19012
rect 87444 19068 87508 19072
rect 87444 19012 87448 19068
rect 87448 19012 87504 19068
rect 87504 19012 87508 19068
rect 87444 19008 87508 19012
rect 87524 19068 87588 19072
rect 87524 19012 87528 19068
rect 87528 19012 87584 19068
rect 87584 19012 87588 19068
rect 87524 19008 87588 19012
rect 5956 18524 6020 18528
rect 5956 18468 5960 18524
rect 5960 18468 6016 18524
rect 6016 18468 6020 18524
rect 5956 18464 6020 18468
rect 6036 18524 6100 18528
rect 6036 18468 6040 18524
rect 6040 18468 6096 18524
rect 6096 18468 6100 18524
rect 6036 18464 6100 18468
rect 6116 18524 6180 18528
rect 6116 18468 6120 18524
rect 6120 18468 6176 18524
rect 6176 18468 6180 18524
rect 6116 18464 6180 18468
rect 6196 18524 6260 18528
rect 6196 18468 6200 18524
rect 6200 18468 6256 18524
rect 6256 18468 6260 18524
rect 6196 18464 6260 18468
rect 86548 18524 86612 18528
rect 86548 18468 86552 18524
rect 86552 18468 86608 18524
rect 86608 18468 86612 18524
rect 86548 18464 86612 18468
rect 86628 18524 86692 18528
rect 86628 18468 86632 18524
rect 86632 18468 86688 18524
rect 86688 18468 86692 18524
rect 86628 18464 86692 18468
rect 86708 18524 86772 18528
rect 86708 18468 86712 18524
rect 86712 18468 86768 18524
rect 86768 18468 86772 18524
rect 86708 18464 86772 18468
rect 86788 18524 86852 18528
rect 86788 18468 86792 18524
rect 86792 18468 86848 18524
rect 86848 18468 86852 18524
rect 86788 18464 86852 18468
rect 6692 17980 6756 17984
rect 6692 17924 6696 17980
rect 6696 17924 6752 17980
rect 6752 17924 6756 17980
rect 6692 17920 6756 17924
rect 6772 17980 6836 17984
rect 6772 17924 6776 17980
rect 6776 17924 6832 17980
rect 6832 17924 6836 17980
rect 6772 17920 6836 17924
rect 6852 17980 6916 17984
rect 6852 17924 6856 17980
rect 6856 17924 6912 17980
rect 6912 17924 6916 17980
rect 6852 17920 6916 17924
rect 6932 17980 6996 17984
rect 6932 17924 6936 17980
rect 6936 17924 6992 17980
rect 6992 17924 6996 17980
rect 6932 17920 6996 17924
rect 87284 17980 87348 17984
rect 87284 17924 87288 17980
rect 87288 17924 87344 17980
rect 87344 17924 87348 17980
rect 87284 17920 87348 17924
rect 87364 17980 87428 17984
rect 87364 17924 87368 17980
rect 87368 17924 87424 17980
rect 87424 17924 87428 17980
rect 87364 17920 87428 17924
rect 87444 17980 87508 17984
rect 87444 17924 87448 17980
rect 87448 17924 87504 17980
rect 87504 17924 87508 17980
rect 87444 17920 87508 17924
rect 87524 17980 87588 17984
rect 87524 17924 87528 17980
rect 87528 17924 87584 17980
rect 87584 17924 87588 17980
rect 87524 17920 87588 17924
rect 5956 17436 6020 17440
rect 5956 17380 5960 17436
rect 5960 17380 6016 17436
rect 6016 17380 6020 17436
rect 5956 17376 6020 17380
rect 6036 17436 6100 17440
rect 6036 17380 6040 17436
rect 6040 17380 6096 17436
rect 6096 17380 6100 17436
rect 6036 17376 6100 17380
rect 6116 17436 6180 17440
rect 6116 17380 6120 17436
rect 6120 17380 6176 17436
rect 6176 17380 6180 17436
rect 6116 17376 6180 17380
rect 6196 17436 6260 17440
rect 6196 17380 6200 17436
rect 6200 17380 6256 17436
rect 6256 17380 6260 17436
rect 6196 17376 6260 17380
rect 86548 17436 86612 17440
rect 86548 17380 86552 17436
rect 86552 17380 86608 17436
rect 86608 17380 86612 17436
rect 86548 17376 86612 17380
rect 86628 17436 86692 17440
rect 86628 17380 86632 17436
rect 86632 17380 86688 17436
rect 86688 17380 86692 17436
rect 86628 17376 86692 17380
rect 86708 17436 86772 17440
rect 86708 17380 86712 17436
rect 86712 17380 86768 17436
rect 86768 17380 86772 17436
rect 86708 17376 86772 17380
rect 86788 17436 86852 17440
rect 86788 17380 86792 17436
rect 86792 17380 86848 17436
rect 86848 17380 86852 17436
rect 86788 17376 86852 17380
rect 6692 16892 6756 16896
rect 6692 16836 6696 16892
rect 6696 16836 6752 16892
rect 6752 16836 6756 16892
rect 6692 16832 6756 16836
rect 6772 16892 6836 16896
rect 6772 16836 6776 16892
rect 6776 16836 6832 16892
rect 6832 16836 6836 16892
rect 6772 16832 6836 16836
rect 6852 16892 6916 16896
rect 6852 16836 6856 16892
rect 6856 16836 6912 16892
rect 6912 16836 6916 16892
rect 6852 16832 6916 16836
rect 6932 16892 6996 16896
rect 6932 16836 6936 16892
rect 6936 16836 6992 16892
rect 6992 16836 6996 16892
rect 6932 16832 6996 16836
rect 87284 16892 87348 16896
rect 87284 16836 87288 16892
rect 87288 16836 87344 16892
rect 87344 16836 87348 16892
rect 87284 16832 87348 16836
rect 87364 16892 87428 16896
rect 87364 16836 87368 16892
rect 87368 16836 87424 16892
rect 87424 16836 87428 16892
rect 87364 16832 87428 16836
rect 87444 16892 87508 16896
rect 87444 16836 87448 16892
rect 87448 16836 87504 16892
rect 87504 16836 87508 16892
rect 87444 16832 87508 16836
rect 87524 16892 87588 16896
rect 87524 16836 87528 16892
rect 87528 16836 87584 16892
rect 87584 16836 87588 16892
rect 87524 16832 87588 16836
rect 5956 16348 6020 16352
rect 5956 16292 5960 16348
rect 5960 16292 6016 16348
rect 6016 16292 6020 16348
rect 5956 16288 6020 16292
rect 6036 16348 6100 16352
rect 6036 16292 6040 16348
rect 6040 16292 6096 16348
rect 6096 16292 6100 16348
rect 6036 16288 6100 16292
rect 6116 16348 6180 16352
rect 6116 16292 6120 16348
rect 6120 16292 6176 16348
rect 6176 16292 6180 16348
rect 6116 16288 6180 16292
rect 6196 16348 6260 16352
rect 6196 16292 6200 16348
rect 6200 16292 6256 16348
rect 6256 16292 6260 16348
rect 6196 16288 6260 16292
rect 86548 16348 86612 16352
rect 86548 16292 86552 16348
rect 86552 16292 86608 16348
rect 86608 16292 86612 16348
rect 86548 16288 86612 16292
rect 86628 16348 86692 16352
rect 86628 16292 86632 16348
rect 86632 16292 86688 16348
rect 86688 16292 86692 16348
rect 86628 16288 86692 16292
rect 86708 16348 86772 16352
rect 86708 16292 86712 16348
rect 86712 16292 86768 16348
rect 86768 16292 86772 16348
rect 86708 16288 86772 16292
rect 86788 16348 86852 16352
rect 86788 16292 86792 16348
rect 86792 16292 86848 16348
rect 86848 16292 86852 16348
rect 86788 16288 86852 16292
rect 6692 15804 6756 15808
rect 6692 15748 6696 15804
rect 6696 15748 6752 15804
rect 6752 15748 6756 15804
rect 6692 15744 6756 15748
rect 6772 15804 6836 15808
rect 6772 15748 6776 15804
rect 6776 15748 6832 15804
rect 6832 15748 6836 15804
rect 6772 15744 6836 15748
rect 6852 15804 6916 15808
rect 6852 15748 6856 15804
rect 6856 15748 6912 15804
rect 6912 15748 6916 15804
rect 6852 15744 6916 15748
rect 6932 15804 6996 15808
rect 6932 15748 6936 15804
rect 6936 15748 6992 15804
rect 6992 15748 6996 15804
rect 6932 15744 6996 15748
rect 87284 15804 87348 15808
rect 87284 15748 87288 15804
rect 87288 15748 87344 15804
rect 87344 15748 87348 15804
rect 87284 15744 87348 15748
rect 87364 15804 87428 15808
rect 87364 15748 87368 15804
rect 87368 15748 87424 15804
rect 87424 15748 87428 15804
rect 87364 15744 87428 15748
rect 87444 15804 87508 15808
rect 87444 15748 87448 15804
rect 87448 15748 87504 15804
rect 87504 15748 87508 15804
rect 87444 15744 87508 15748
rect 87524 15804 87588 15808
rect 87524 15748 87528 15804
rect 87528 15748 87584 15804
rect 87584 15748 87588 15804
rect 87524 15744 87588 15748
rect 5956 15260 6020 15264
rect 5956 15204 5960 15260
rect 5960 15204 6016 15260
rect 6016 15204 6020 15260
rect 5956 15200 6020 15204
rect 6036 15260 6100 15264
rect 6036 15204 6040 15260
rect 6040 15204 6096 15260
rect 6096 15204 6100 15260
rect 6036 15200 6100 15204
rect 6116 15260 6180 15264
rect 6116 15204 6120 15260
rect 6120 15204 6176 15260
rect 6176 15204 6180 15260
rect 6116 15200 6180 15204
rect 6196 15260 6260 15264
rect 6196 15204 6200 15260
rect 6200 15204 6256 15260
rect 6256 15204 6260 15260
rect 6196 15200 6260 15204
rect 86548 15260 86612 15264
rect 86548 15204 86552 15260
rect 86552 15204 86608 15260
rect 86608 15204 86612 15260
rect 86548 15200 86612 15204
rect 86628 15260 86692 15264
rect 86628 15204 86632 15260
rect 86632 15204 86688 15260
rect 86688 15204 86692 15260
rect 86628 15200 86692 15204
rect 86708 15260 86772 15264
rect 86708 15204 86712 15260
rect 86712 15204 86768 15260
rect 86768 15204 86772 15260
rect 86708 15200 86772 15204
rect 86788 15260 86852 15264
rect 86788 15204 86792 15260
rect 86792 15204 86848 15260
rect 86848 15204 86852 15260
rect 86788 15200 86852 15204
rect 6692 14716 6756 14720
rect 6692 14660 6696 14716
rect 6696 14660 6752 14716
rect 6752 14660 6756 14716
rect 6692 14656 6756 14660
rect 6772 14716 6836 14720
rect 6772 14660 6776 14716
rect 6776 14660 6832 14716
rect 6832 14660 6836 14716
rect 6772 14656 6836 14660
rect 6852 14716 6916 14720
rect 6852 14660 6856 14716
rect 6856 14660 6912 14716
rect 6912 14660 6916 14716
rect 6852 14656 6916 14660
rect 6932 14716 6996 14720
rect 6932 14660 6936 14716
rect 6936 14660 6992 14716
rect 6992 14660 6996 14716
rect 6932 14656 6996 14660
rect 87284 14716 87348 14720
rect 87284 14660 87288 14716
rect 87288 14660 87344 14716
rect 87344 14660 87348 14716
rect 87284 14656 87348 14660
rect 87364 14716 87428 14720
rect 87364 14660 87368 14716
rect 87368 14660 87424 14716
rect 87424 14660 87428 14716
rect 87364 14656 87428 14660
rect 87444 14716 87508 14720
rect 87444 14660 87448 14716
rect 87448 14660 87504 14716
rect 87504 14660 87508 14716
rect 87444 14656 87508 14660
rect 87524 14716 87588 14720
rect 87524 14660 87528 14716
rect 87528 14660 87584 14716
rect 87584 14660 87588 14716
rect 87524 14656 87588 14660
rect 5956 14172 6020 14176
rect 5956 14116 5960 14172
rect 5960 14116 6016 14172
rect 6016 14116 6020 14172
rect 5956 14112 6020 14116
rect 6036 14172 6100 14176
rect 6036 14116 6040 14172
rect 6040 14116 6096 14172
rect 6096 14116 6100 14172
rect 6036 14112 6100 14116
rect 6116 14172 6180 14176
rect 6116 14116 6120 14172
rect 6120 14116 6176 14172
rect 6176 14116 6180 14172
rect 6116 14112 6180 14116
rect 6196 14172 6260 14176
rect 6196 14116 6200 14172
rect 6200 14116 6256 14172
rect 6256 14116 6260 14172
rect 6196 14112 6260 14116
rect 86548 14172 86612 14176
rect 86548 14116 86552 14172
rect 86552 14116 86608 14172
rect 86608 14116 86612 14172
rect 86548 14112 86612 14116
rect 86628 14172 86692 14176
rect 86628 14116 86632 14172
rect 86632 14116 86688 14172
rect 86688 14116 86692 14172
rect 86628 14112 86692 14116
rect 86708 14172 86772 14176
rect 86708 14116 86712 14172
rect 86712 14116 86768 14172
rect 86768 14116 86772 14172
rect 86708 14112 86772 14116
rect 86788 14172 86852 14176
rect 86788 14116 86792 14172
rect 86792 14116 86848 14172
rect 86848 14116 86852 14172
rect 86788 14112 86852 14116
rect 6692 13628 6756 13632
rect 6692 13572 6696 13628
rect 6696 13572 6752 13628
rect 6752 13572 6756 13628
rect 6692 13568 6756 13572
rect 6772 13628 6836 13632
rect 6772 13572 6776 13628
rect 6776 13572 6832 13628
rect 6832 13572 6836 13628
rect 6772 13568 6836 13572
rect 6852 13628 6916 13632
rect 6852 13572 6856 13628
rect 6856 13572 6912 13628
rect 6912 13572 6916 13628
rect 6852 13568 6916 13572
rect 6932 13628 6996 13632
rect 6932 13572 6936 13628
rect 6936 13572 6992 13628
rect 6992 13572 6996 13628
rect 6932 13568 6996 13572
rect 87284 13628 87348 13632
rect 87284 13572 87288 13628
rect 87288 13572 87344 13628
rect 87344 13572 87348 13628
rect 87284 13568 87348 13572
rect 87364 13628 87428 13632
rect 87364 13572 87368 13628
rect 87368 13572 87424 13628
rect 87424 13572 87428 13628
rect 87364 13568 87428 13572
rect 87444 13628 87508 13632
rect 87444 13572 87448 13628
rect 87448 13572 87504 13628
rect 87504 13572 87508 13628
rect 87444 13568 87508 13572
rect 87524 13628 87588 13632
rect 87524 13572 87528 13628
rect 87528 13572 87584 13628
rect 87584 13572 87588 13628
rect 87524 13568 87588 13572
rect 5956 13084 6020 13088
rect 5956 13028 5960 13084
rect 5960 13028 6016 13084
rect 6016 13028 6020 13084
rect 5956 13024 6020 13028
rect 6036 13084 6100 13088
rect 6036 13028 6040 13084
rect 6040 13028 6096 13084
rect 6096 13028 6100 13084
rect 6036 13024 6100 13028
rect 6116 13084 6180 13088
rect 6116 13028 6120 13084
rect 6120 13028 6176 13084
rect 6176 13028 6180 13084
rect 6116 13024 6180 13028
rect 6196 13084 6260 13088
rect 6196 13028 6200 13084
rect 6200 13028 6256 13084
rect 6256 13028 6260 13084
rect 6196 13024 6260 13028
rect 86548 13084 86612 13088
rect 86548 13028 86552 13084
rect 86552 13028 86608 13084
rect 86608 13028 86612 13084
rect 86548 13024 86612 13028
rect 86628 13084 86692 13088
rect 86628 13028 86632 13084
rect 86632 13028 86688 13084
rect 86688 13028 86692 13084
rect 86628 13024 86692 13028
rect 86708 13084 86772 13088
rect 86708 13028 86712 13084
rect 86712 13028 86768 13084
rect 86768 13028 86772 13084
rect 86708 13024 86772 13028
rect 86788 13084 86852 13088
rect 86788 13028 86792 13084
rect 86792 13028 86848 13084
rect 86848 13028 86852 13084
rect 86788 13024 86852 13028
rect 6692 12540 6756 12544
rect 6692 12484 6696 12540
rect 6696 12484 6752 12540
rect 6752 12484 6756 12540
rect 6692 12480 6756 12484
rect 6772 12540 6836 12544
rect 6772 12484 6776 12540
rect 6776 12484 6832 12540
rect 6832 12484 6836 12540
rect 6772 12480 6836 12484
rect 6852 12540 6916 12544
rect 6852 12484 6856 12540
rect 6856 12484 6912 12540
rect 6912 12484 6916 12540
rect 6852 12480 6916 12484
rect 6932 12540 6996 12544
rect 6932 12484 6936 12540
rect 6936 12484 6992 12540
rect 6992 12484 6996 12540
rect 6932 12480 6996 12484
rect 87284 12540 87348 12544
rect 87284 12484 87288 12540
rect 87288 12484 87344 12540
rect 87344 12484 87348 12540
rect 87284 12480 87348 12484
rect 87364 12540 87428 12544
rect 87364 12484 87368 12540
rect 87368 12484 87424 12540
rect 87424 12484 87428 12540
rect 87364 12480 87428 12484
rect 87444 12540 87508 12544
rect 87444 12484 87448 12540
rect 87448 12484 87504 12540
rect 87504 12484 87508 12540
rect 87444 12480 87508 12484
rect 87524 12540 87588 12544
rect 87524 12484 87528 12540
rect 87528 12484 87584 12540
rect 87584 12484 87588 12540
rect 87524 12480 87588 12484
rect 5956 11996 6020 12000
rect 5956 11940 5960 11996
rect 5960 11940 6016 11996
rect 6016 11940 6020 11996
rect 5956 11936 6020 11940
rect 6036 11996 6100 12000
rect 6036 11940 6040 11996
rect 6040 11940 6096 11996
rect 6096 11940 6100 11996
rect 6036 11936 6100 11940
rect 6116 11996 6180 12000
rect 6116 11940 6120 11996
rect 6120 11940 6176 11996
rect 6176 11940 6180 11996
rect 6116 11936 6180 11940
rect 6196 11996 6260 12000
rect 6196 11940 6200 11996
rect 6200 11940 6256 11996
rect 6256 11940 6260 11996
rect 6196 11936 6260 11940
rect 86548 11996 86612 12000
rect 86548 11940 86552 11996
rect 86552 11940 86608 11996
rect 86608 11940 86612 11996
rect 86548 11936 86612 11940
rect 86628 11996 86692 12000
rect 86628 11940 86632 11996
rect 86632 11940 86688 11996
rect 86688 11940 86692 11996
rect 86628 11936 86692 11940
rect 86708 11996 86772 12000
rect 86708 11940 86712 11996
rect 86712 11940 86768 11996
rect 86768 11940 86772 11996
rect 86708 11936 86772 11940
rect 86788 11996 86852 12000
rect 86788 11940 86792 11996
rect 86792 11940 86848 11996
rect 86848 11940 86852 11996
rect 86788 11936 86852 11940
rect 6692 11452 6756 11456
rect 6692 11396 6696 11452
rect 6696 11396 6752 11452
rect 6752 11396 6756 11452
rect 6692 11392 6756 11396
rect 6772 11452 6836 11456
rect 6772 11396 6776 11452
rect 6776 11396 6832 11452
rect 6832 11396 6836 11452
rect 6772 11392 6836 11396
rect 6852 11452 6916 11456
rect 6852 11396 6856 11452
rect 6856 11396 6912 11452
rect 6912 11396 6916 11452
rect 6852 11392 6916 11396
rect 6932 11452 6996 11456
rect 6932 11396 6936 11452
rect 6936 11396 6992 11452
rect 6992 11396 6996 11452
rect 6932 11392 6996 11396
rect 87284 11452 87348 11456
rect 87284 11396 87288 11452
rect 87288 11396 87344 11452
rect 87344 11396 87348 11452
rect 87284 11392 87348 11396
rect 87364 11452 87428 11456
rect 87364 11396 87368 11452
rect 87368 11396 87424 11452
rect 87424 11396 87428 11452
rect 87364 11392 87428 11396
rect 87444 11452 87508 11456
rect 87444 11396 87448 11452
rect 87448 11396 87504 11452
rect 87504 11396 87508 11452
rect 87444 11392 87508 11396
rect 87524 11452 87588 11456
rect 87524 11396 87528 11452
rect 87528 11396 87584 11452
rect 87584 11396 87588 11452
rect 87524 11392 87588 11396
rect 5956 10908 6020 10912
rect 5956 10852 5960 10908
rect 5960 10852 6016 10908
rect 6016 10852 6020 10908
rect 5956 10848 6020 10852
rect 6036 10908 6100 10912
rect 6036 10852 6040 10908
rect 6040 10852 6096 10908
rect 6096 10852 6100 10908
rect 6036 10848 6100 10852
rect 6116 10908 6180 10912
rect 6116 10852 6120 10908
rect 6120 10852 6176 10908
rect 6176 10852 6180 10908
rect 6116 10848 6180 10852
rect 6196 10908 6260 10912
rect 6196 10852 6200 10908
rect 6200 10852 6256 10908
rect 6256 10852 6260 10908
rect 6196 10848 6260 10852
rect 86548 10908 86612 10912
rect 86548 10852 86552 10908
rect 86552 10852 86608 10908
rect 86608 10852 86612 10908
rect 86548 10848 86612 10852
rect 86628 10908 86692 10912
rect 86628 10852 86632 10908
rect 86632 10852 86688 10908
rect 86688 10852 86692 10908
rect 86628 10848 86692 10852
rect 86708 10908 86772 10912
rect 86708 10852 86712 10908
rect 86712 10852 86768 10908
rect 86768 10852 86772 10908
rect 86708 10848 86772 10852
rect 86788 10908 86852 10912
rect 86788 10852 86792 10908
rect 86792 10852 86848 10908
rect 86848 10852 86852 10908
rect 86788 10848 86852 10852
rect 6692 10364 6756 10368
rect 6692 10308 6696 10364
rect 6696 10308 6752 10364
rect 6752 10308 6756 10364
rect 6692 10304 6756 10308
rect 6772 10364 6836 10368
rect 6772 10308 6776 10364
rect 6776 10308 6832 10364
rect 6832 10308 6836 10364
rect 6772 10304 6836 10308
rect 6852 10364 6916 10368
rect 6852 10308 6856 10364
rect 6856 10308 6912 10364
rect 6912 10308 6916 10364
rect 6852 10304 6916 10308
rect 6932 10364 6996 10368
rect 6932 10308 6936 10364
rect 6936 10308 6992 10364
rect 6992 10308 6996 10364
rect 6932 10304 6996 10308
rect 87284 10364 87348 10368
rect 87284 10308 87288 10364
rect 87288 10308 87344 10364
rect 87344 10308 87348 10364
rect 87284 10304 87348 10308
rect 87364 10364 87428 10368
rect 87364 10308 87368 10364
rect 87368 10308 87424 10364
rect 87424 10308 87428 10364
rect 87364 10304 87428 10308
rect 87444 10364 87508 10368
rect 87444 10308 87448 10364
rect 87448 10308 87504 10364
rect 87504 10308 87508 10364
rect 87444 10304 87508 10308
rect 87524 10364 87588 10368
rect 87524 10308 87528 10364
rect 87528 10308 87584 10364
rect 87584 10308 87588 10364
rect 87524 10304 87588 10308
rect 5956 9820 6020 9824
rect 5956 9764 5960 9820
rect 5960 9764 6016 9820
rect 6016 9764 6020 9820
rect 5956 9760 6020 9764
rect 6036 9820 6100 9824
rect 6036 9764 6040 9820
rect 6040 9764 6096 9820
rect 6096 9764 6100 9820
rect 6036 9760 6100 9764
rect 6116 9820 6180 9824
rect 6116 9764 6120 9820
rect 6120 9764 6176 9820
rect 6176 9764 6180 9820
rect 6116 9760 6180 9764
rect 6196 9820 6260 9824
rect 6196 9764 6200 9820
rect 6200 9764 6256 9820
rect 6256 9764 6260 9820
rect 6196 9760 6260 9764
rect 86548 9820 86612 9824
rect 86548 9764 86552 9820
rect 86552 9764 86608 9820
rect 86608 9764 86612 9820
rect 86548 9760 86612 9764
rect 86628 9820 86692 9824
rect 86628 9764 86632 9820
rect 86632 9764 86688 9820
rect 86688 9764 86692 9820
rect 86628 9760 86692 9764
rect 86708 9820 86772 9824
rect 86708 9764 86712 9820
rect 86712 9764 86768 9820
rect 86768 9764 86772 9820
rect 86708 9760 86772 9764
rect 86788 9820 86852 9824
rect 86788 9764 86792 9820
rect 86792 9764 86848 9820
rect 86848 9764 86852 9820
rect 86788 9760 86852 9764
rect 6692 9276 6756 9280
rect 6692 9220 6696 9276
rect 6696 9220 6752 9276
rect 6752 9220 6756 9276
rect 6692 9216 6756 9220
rect 6772 9276 6836 9280
rect 6772 9220 6776 9276
rect 6776 9220 6832 9276
rect 6832 9220 6836 9276
rect 6772 9216 6836 9220
rect 6852 9276 6916 9280
rect 6852 9220 6856 9276
rect 6856 9220 6912 9276
rect 6912 9220 6916 9276
rect 6852 9216 6916 9220
rect 6932 9276 6996 9280
rect 6932 9220 6936 9276
rect 6936 9220 6992 9276
rect 6992 9220 6996 9276
rect 6932 9216 6996 9220
rect 87284 9276 87348 9280
rect 87284 9220 87288 9276
rect 87288 9220 87344 9276
rect 87344 9220 87348 9276
rect 87284 9216 87348 9220
rect 87364 9276 87428 9280
rect 87364 9220 87368 9276
rect 87368 9220 87424 9276
rect 87424 9220 87428 9276
rect 87364 9216 87428 9220
rect 87444 9276 87508 9280
rect 87444 9220 87448 9276
rect 87448 9220 87504 9276
rect 87504 9220 87508 9276
rect 87444 9216 87508 9220
rect 87524 9276 87588 9280
rect 87524 9220 87528 9276
rect 87528 9220 87584 9276
rect 87584 9220 87588 9276
rect 87524 9216 87588 9220
rect 5956 8732 6020 8736
rect 5956 8676 5960 8732
rect 5960 8676 6016 8732
rect 6016 8676 6020 8732
rect 5956 8672 6020 8676
rect 6036 8732 6100 8736
rect 6036 8676 6040 8732
rect 6040 8676 6096 8732
rect 6096 8676 6100 8732
rect 6036 8672 6100 8676
rect 6116 8732 6180 8736
rect 6116 8676 6120 8732
rect 6120 8676 6176 8732
rect 6176 8676 6180 8732
rect 6116 8672 6180 8676
rect 6196 8732 6260 8736
rect 6196 8676 6200 8732
rect 6200 8676 6256 8732
rect 6256 8676 6260 8732
rect 6196 8672 6260 8676
rect 86548 8732 86612 8736
rect 86548 8676 86552 8732
rect 86552 8676 86608 8732
rect 86608 8676 86612 8732
rect 86548 8672 86612 8676
rect 86628 8732 86692 8736
rect 86628 8676 86632 8732
rect 86632 8676 86688 8732
rect 86688 8676 86692 8732
rect 86628 8672 86692 8676
rect 86708 8732 86772 8736
rect 86708 8676 86712 8732
rect 86712 8676 86768 8732
rect 86768 8676 86772 8732
rect 86708 8672 86772 8676
rect 86788 8732 86852 8736
rect 86788 8676 86792 8732
rect 86792 8676 86848 8732
rect 86848 8676 86852 8732
rect 86788 8672 86852 8676
rect 6692 8188 6756 8192
rect 6692 8132 6696 8188
rect 6696 8132 6752 8188
rect 6752 8132 6756 8188
rect 6692 8128 6756 8132
rect 6772 8188 6836 8192
rect 6772 8132 6776 8188
rect 6776 8132 6832 8188
rect 6832 8132 6836 8188
rect 6772 8128 6836 8132
rect 6852 8188 6916 8192
rect 6852 8132 6856 8188
rect 6856 8132 6912 8188
rect 6912 8132 6916 8188
rect 6852 8128 6916 8132
rect 6932 8188 6996 8192
rect 6932 8132 6936 8188
rect 6936 8132 6992 8188
rect 6992 8132 6996 8188
rect 6932 8128 6996 8132
rect 87284 8188 87348 8192
rect 87284 8132 87288 8188
rect 87288 8132 87344 8188
rect 87344 8132 87348 8188
rect 87284 8128 87348 8132
rect 87364 8188 87428 8192
rect 87364 8132 87368 8188
rect 87368 8132 87424 8188
rect 87424 8132 87428 8188
rect 87364 8128 87428 8132
rect 87444 8188 87508 8192
rect 87444 8132 87448 8188
rect 87448 8132 87504 8188
rect 87504 8132 87508 8188
rect 87444 8128 87508 8132
rect 87524 8188 87588 8192
rect 87524 8132 87528 8188
rect 87528 8132 87584 8188
rect 87584 8132 87588 8188
rect 87524 8128 87588 8132
rect 5956 7644 6020 7648
rect 5956 7588 5960 7644
rect 5960 7588 6016 7644
rect 6016 7588 6020 7644
rect 5956 7584 6020 7588
rect 6036 7644 6100 7648
rect 6036 7588 6040 7644
rect 6040 7588 6096 7644
rect 6096 7588 6100 7644
rect 6036 7584 6100 7588
rect 6116 7644 6180 7648
rect 6116 7588 6120 7644
rect 6120 7588 6176 7644
rect 6176 7588 6180 7644
rect 6116 7584 6180 7588
rect 6196 7644 6260 7648
rect 6196 7588 6200 7644
rect 6200 7588 6256 7644
rect 6256 7588 6260 7644
rect 6196 7584 6260 7588
rect 17724 7644 17788 7648
rect 17724 7588 17728 7644
rect 17728 7588 17784 7644
rect 17784 7588 17788 7644
rect 17724 7584 17788 7588
rect 17804 7644 17868 7648
rect 17804 7588 17808 7644
rect 17808 7588 17864 7644
rect 17864 7588 17868 7644
rect 17804 7584 17868 7588
rect 17884 7644 17948 7648
rect 17884 7588 17888 7644
rect 17888 7588 17944 7644
rect 17944 7588 17948 7644
rect 17884 7584 17948 7588
rect 17964 7644 18028 7648
rect 17964 7588 17968 7644
rect 17968 7588 18024 7644
rect 18024 7588 18028 7644
rect 17964 7584 18028 7588
rect 36124 7644 36188 7648
rect 36124 7588 36128 7644
rect 36128 7588 36184 7644
rect 36184 7588 36188 7644
rect 36124 7584 36188 7588
rect 36204 7644 36268 7648
rect 36204 7588 36208 7644
rect 36208 7588 36264 7644
rect 36264 7588 36268 7644
rect 36204 7584 36268 7588
rect 36284 7644 36348 7648
rect 36284 7588 36288 7644
rect 36288 7588 36344 7644
rect 36344 7588 36348 7644
rect 36284 7584 36348 7588
rect 36364 7644 36428 7648
rect 36364 7588 36368 7644
rect 36368 7588 36424 7644
rect 36424 7588 36428 7644
rect 36364 7584 36428 7588
rect 54524 7644 54588 7648
rect 54524 7588 54528 7644
rect 54528 7588 54584 7644
rect 54584 7588 54588 7644
rect 54524 7584 54588 7588
rect 54604 7644 54668 7648
rect 54604 7588 54608 7644
rect 54608 7588 54664 7644
rect 54664 7588 54668 7644
rect 54604 7584 54668 7588
rect 54684 7644 54748 7648
rect 54684 7588 54688 7644
rect 54688 7588 54744 7644
rect 54744 7588 54748 7644
rect 54684 7584 54748 7588
rect 54764 7644 54828 7648
rect 54764 7588 54768 7644
rect 54768 7588 54824 7644
rect 54824 7588 54828 7644
rect 54764 7584 54828 7588
rect 72924 7644 72988 7648
rect 72924 7588 72928 7644
rect 72928 7588 72984 7644
rect 72984 7588 72988 7644
rect 72924 7584 72988 7588
rect 73004 7644 73068 7648
rect 73004 7588 73008 7644
rect 73008 7588 73064 7644
rect 73064 7588 73068 7644
rect 73004 7584 73068 7588
rect 73084 7644 73148 7648
rect 73084 7588 73088 7644
rect 73088 7588 73144 7644
rect 73144 7588 73148 7644
rect 73084 7584 73148 7588
rect 73164 7644 73228 7648
rect 73164 7588 73168 7644
rect 73168 7588 73224 7644
rect 73224 7588 73228 7644
rect 73164 7584 73228 7588
rect 86548 7644 86612 7648
rect 86548 7588 86552 7644
rect 86552 7588 86608 7644
rect 86608 7588 86612 7644
rect 86548 7584 86612 7588
rect 86628 7644 86692 7648
rect 86628 7588 86632 7644
rect 86632 7588 86688 7644
rect 86688 7588 86692 7644
rect 86628 7584 86692 7588
rect 86708 7644 86772 7648
rect 86708 7588 86712 7644
rect 86712 7588 86768 7644
rect 86768 7588 86772 7644
rect 86708 7584 86772 7588
rect 86788 7644 86852 7648
rect 86788 7588 86792 7644
rect 86792 7588 86848 7644
rect 86848 7588 86852 7644
rect 86788 7584 86852 7588
rect 6692 7100 6756 7104
rect 6692 7044 6696 7100
rect 6696 7044 6752 7100
rect 6752 7044 6756 7100
rect 6692 7040 6756 7044
rect 6772 7100 6836 7104
rect 6772 7044 6776 7100
rect 6776 7044 6832 7100
rect 6832 7044 6836 7100
rect 6772 7040 6836 7044
rect 6852 7100 6916 7104
rect 6852 7044 6856 7100
rect 6856 7044 6912 7100
rect 6912 7044 6916 7100
rect 6852 7040 6916 7044
rect 6932 7100 6996 7104
rect 6932 7044 6936 7100
rect 6936 7044 6992 7100
rect 6992 7044 6996 7100
rect 6932 7040 6996 7044
rect 18384 7100 18448 7104
rect 18384 7044 18388 7100
rect 18388 7044 18444 7100
rect 18444 7044 18448 7100
rect 18384 7040 18448 7044
rect 18464 7100 18528 7104
rect 18464 7044 18468 7100
rect 18468 7044 18524 7100
rect 18524 7044 18528 7100
rect 18464 7040 18528 7044
rect 18544 7100 18608 7104
rect 18544 7044 18548 7100
rect 18548 7044 18604 7100
rect 18604 7044 18608 7100
rect 18544 7040 18608 7044
rect 18624 7100 18688 7104
rect 18624 7044 18628 7100
rect 18628 7044 18684 7100
rect 18684 7044 18688 7100
rect 18624 7040 18688 7044
rect 36784 7100 36848 7104
rect 36784 7044 36788 7100
rect 36788 7044 36844 7100
rect 36844 7044 36848 7100
rect 36784 7040 36848 7044
rect 36864 7100 36928 7104
rect 36864 7044 36868 7100
rect 36868 7044 36924 7100
rect 36924 7044 36928 7100
rect 36864 7040 36928 7044
rect 36944 7100 37008 7104
rect 36944 7044 36948 7100
rect 36948 7044 37004 7100
rect 37004 7044 37008 7100
rect 36944 7040 37008 7044
rect 37024 7100 37088 7104
rect 37024 7044 37028 7100
rect 37028 7044 37084 7100
rect 37084 7044 37088 7100
rect 37024 7040 37088 7044
rect 55184 7100 55248 7104
rect 55184 7044 55188 7100
rect 55188 7044 55244 7100
rect 55244 7044 55248 7100
rect 55184 7040 55248 7044
rect 55264 7100 55328 7104
rect 55264 7044 55268 7100
rect 55268 7044 55324 7100
rect 55324 7044 55328 7100
rect 55264 7040 55328 7044
rect 55344 7100 55408 7104
rect 55344 7044 55348 7100
rect 55348 7044 55404 7100
rect 55404 7044 55408 7100
rect 55344 7040 55408 7044
rect 55424 7100 55488 7104
rect 55424 7044 55428 7100
rect 55428 7044 55484 7100
rect 55484 7044 55488 7100
rect 55424 7040 55488 7044
rect 73584 7100 73648 7104
rect 73584 7044 73588 7100
rect 73588 7044 73644 7100
rect 73644 7044 73648 7100
rect 73584 7040 73648 7044
rect 73664 7100 73728 7104
rect 73664 7044 73668 7100
rect 73668 7044 73724 7100
rect 73724 7044 73728 7100
rect 73664 7040 73728 7044
rect 73744 7100 73808 7104
rect 73744 7044 73748 7100
rect 73748 7044 73804 7100
rect 73804 7044 73808 7100
rect 73744 7040 73808 7044
rect 73824 7100 73888 7104
rect 73824 7044 73828 7100
rect 73828 7044 73884 7100
rect 73884 7044 73888 7100
rect 73824 7040 73888 7044
rect 87284 7100 87348 7104
rect 87284 7044 87288 7100
rect 87288 7044 87344 7100
rect 87344 7044 87348 7100
rect 87284 7040 87348 7044
rect 87364 7100 87428 7104
rect 87364 7044 87368 7100
rect 87368 7044 87424 7100
rect 87424 7044 87428 7100
rect 87364 7040 87428 7044
rect 87444 7100 87508 7104
rect 87444 7044 87448 7100
rect 87448 7044 87504 7100
rect 87504 7044 87508 7100
rect 87444 7040 87508 7044
rect 87524 7100 87588 7104
rect 87524 7044 87528 7100
rect 87528 7044 87584 7100
rect 87584 7044 87588 7100
rect 87524 7040 87588 7044
rect 17724 6556 17788 6560
rect 17724 6500 17728 6556
rect 17728 6500 17784 6556
rect 17784 6500 17788 6556
rect 17724 6496 17788 6500
rect 17804 6556 17868 6560
rect 17804 6500 17808 6556
rect 17808 6500 17864 6556
rect 17864 6500 17868 6556
rect 17804 6496 17868 6500
rect 17884 6556 17948 6560
rect 17884 6500 17888 6556
rect 17888 6500 17944 6556
rect 17944 6500 17948 6556
rect 17884 6496 17948 6500
rect 17964 6556 18028 6560
rect 17964 6500 17968 6556
rect 17968 6500 18024 6556
rect 18024 6500 18028 6556
rect 17964 6496 18028 6500
rect 36124 6556 36188 6560
rect 36124 6500 36128 6556
rect 36128 6500 36184 6556
rect 36184 6500 36188 6556
rect 36124 6496 36188 6500
rect 36204 6556 36268 6560
rect 36204 6500 36208 6556
rect 36208 6500 36264 6556
rect 36264 6500 36268 6556
rect 36204 6496 36268 6500
rect 36284 6556 36348 6560
rect 36284 6500 36288 6556
rect 36288 6500 36344 6556
rect 36344 6500 36348 6556
rect 36284 6496 36348 6500
rect 36364 6556 36428 6560
rect 36364 6500 36368 6556
rect 36368 6500 36424 6556
rect 36424 6500 36428 6556
rect 36364 6496 36428 6500
rect 54524 6556 54588 6560
rect 54524 6500 54528 6556
rect 54528 6500 54584 6556
rect 54584 6500 54588 6556
rect 54524 6496 54588 6500
rect 54604 6556 54668 6560
rect 54604 6500 54608 6556
rect 54608 6500 54664 6556
rect 54664 6500 54668 6556
rect 54604 6496 54668 6500
rect 54684 6556 54748 6560
rect 54684 6500 54688 6556
rect 54688 6500 54744 6556
rect 54744 6500 54748 6556
rect 54684 6496 54748 6500
rect 54764 6556 54828 6560
rect 54764 6500 54768 6556
rect 54768 6500 54824 6556
rect 54824 6500 54828 6556
rect 54764 6496 54828 6500
rect 72924 6556 72988 6560
rect 72924 6500 72928 6556
rect 72928 6500 72984 6556
rect 72984 6500 72988 6556
rect 72924 6496 72988 6500
rect 73004 6556 73068 6560
rect 73004 6500 73008 6556
rect 73008 6500 73064 6556
rect 73064 6500 73068 6556
rect 73004 6496 73068 6500
rect 73084 6556 73148 6560
rect 73084 6500 73088 6556
rect 73088 6500 73144 6556
rect 73144 6500 73148 6556
rect 73084 6496 73148 6500
rect 73164 6556 73228 6560
rect 73164 6500 73168 6556
rect 73168 6500 73224 6556
rect 73224 6500 73228 6556
rect 73164 6496 73228 6500
rect 18384 6012 18448 6016
rect 18384 5956 18388 6012
rect 18388 5956 18444 6012
rect 18444 5956 18448 6012
rect 18384 5952 18448 5956
rect 18464 6012 18528 6016
rect 18464 5956 18468 6012
rect 18468 5956 18524 6012
rect 18524 5956 18528 6012
rect 18464 5952 18528 5956
rect 18544 6012 18608 6016
rect 18544 5956 18548 6012
rect 18548 5956 18604 6012
rect 18604 5956 18608 6012
rect 18544 5952 18608 5956
rect 18624 6012 18688 6016
rect 18624 5956 18628 6012
rect 18628 5956 18684 6012
rect 18684 5956 18688 6012
rect 18624 5952 18688 5956
rect 36784 6012 36848 6016
rect 36784 5956 36788 6012
rect 36788 5956 36844 6012
rect 36844 5956 36848 6012
rect 36784 5952 36848 5956
rect 36864 6012 36928 6016
rect 36864 5956 36868 6012
rect 36868 5956 36924 6012
rect 36924 5956 36928 6012
rect 36864 5952 36928 5956
rect 36944 6012 37008 6016
rect 36944 5956 36948 6012
rect 36948 5956 37004 6012
rect 37004 5956 37008 6012
rect 36944 5952 37008 5956
rect 37024 6012 37088 6016
rect 37024 5956 37028 6012
rect 37028 5956 37084 6012
rect 37084 5956 37088 6012
rect 37024 5952 37088 5956
rect 55184 6012 55248 6016
rect 55184 5956 55188 6012
rect 55188 5956 55244 6012
rect 55244 5956 55248 6012
rect 55184 5952 55248 5956
rect 55264 6012 55328 6016
rect 55264 5956 55268 6012
rect 55268 5956 55324 6012
rect 55324 5956 55328 6012
rect 55264 5952 55328 5956
rect 55344 6012 55408 6016
rect 55344 5956 55348 6012
rect 55348 5956 55404 6012
rect 55404 5956 55408 6012
rect 55344 5952 55408 5956
rect 55424 6012 55488 6016
rect 55424 5956 55428 6012
rect 55428 5956 55484 6012
rect 55484 5956 55488 6012
rect 55424 5952 55488 5956
rect 73584 6012 73648 6016
rect 73584 5956 73588 6012
rect 73588 5956 73644 6012
rect 73644 5956 73648 6012
rect 73584 5952 73648 5956
rect 73664 6012 73728 6016
rect 73664 5956 73668 6012
rect 73668 5956 73724 6012
rect 73724 5956 73728 6012
rect 73664 5952 73728 5956
rect 73744 6012 73808 6016
rect 73744 5956 73748 6012
rect 73748 5956 73804 6012
rect 73804 5956 73808 6012
rect 73744 5952 73808 5956
rect 73824 6012 73888 6016
rect 73824 5956 73828 6012
rect 73828 5956 73884 6012
rect 73884 5956 73888 6012
rect 73824 5952 73888 5956
rect 17724 5468 17788 5472
rect 17724 5412 17728 5468
rect 17728 5412 17784 5468
rect 17784 5412 17788 5468
rect 17724 5408 17788 5412
rect 17804 5468 17868 5472
rect 17804 5412 17808 5468
rect 17808 5412 17864 5468
rect 17864 5412 17868 5468
rect 17804 5408 17868 5412
rect 17884 5468 17948 5472
rect 17884 5412 17888 5468
rect 17888 5412 17944 5468
rect 17944 5412 17948 5468
rect 17884 5408 17948 5412
rect 17964 5468 18028 5472
rect 17964 5412 17968 5468
rect 17968 5412 18024 5468
rect 18024 5412 18028 5468
rect 17964 5408 18028 5412
rect 36124 5468 36188 5472
rect 36124 5412 36128 5468
rect 36128 5412 36184 5468
rect 36184 5412 36188 5468
rect 36124 5408 36188 5412
rect 36204 5468 36268 5472
rect 36204 5412 36208 5468
rect 36208 5412 36264 5468
rect 36264 5412 36268 5468
rect 36204 5408 36268 5412
rect 36284 5468 36348 5472
rect 36284 5412 36288 5468
rect 36288 5412 36344 5468
rect 36344 5412 36348 5468
rect 36284 5408 36348 5412
rect 36364 5468 36428 5472
rect 36364 5412 36368 5468
rect 36368 5412 36424 5468
rect 36424 5412 36428 5468
rect 36364 5408 36428 5412
rect 54524 5468 54588 5472
rect 54524 5412 54528 5468
rect 54528 5412 54584 5468
rect 54584 5412 54588 5468
rect 54524 5408 54588 5412
rect 54604 5468 54668 5472
rect 54604 5412 54608 5468
rect 54608 5412 54664 5468
rect 54664 5412 54668 5468
rect 54604 5408 54668 5412
rect 54684 5468 54748 5472
rect 54684 5412 54688 5468
rect 54688 5412 54744 5468
rect 54744 5412 54748 5468
rect 54684 5408 54748 5412
rect 54764 5468 54828 5472
rect 54764 5412 54768 5468
rect 54768 5412 54824 5468
rect 54824 5412 54828 5468
rect 54764 5408 54828 5412
rect 72924 5468 72988 5472
rect 72924 5412 72928 5468
rect 72928 5412 72984 5468
rect 72984 5412 72988 5468
rect 72924 5408 72988 5412
rect 73004 5468 73068 5472
rect 73004 5412 73008 5468
rect 73008 5412 73064 5468
rect 73064 5412 73068 5468
rect 73004 5408 73068 5412
rect 73084 5468 73148 5472
rect 73084 5412 73088 5468
rect 73088 5412 73144 5468
rect 73144 5412 73148 5468
rect 73084 5408 73148 5412
rect 73164 5468 73228 5472
rect 73164 5412 73168 5468
rect 73168 5412 73224 5468
rect 73224 5412 73228 5468
rect 73164 5408 73228 5412
rect 18384 4924 18448 4928
rect 18384 4868 18388 4924
rect 18388 4868 18444 4924
rect 18444 4868 18448 4924
rect 18384 4864 18448 4868
rect 18464 4924 18528 4928
rect 18464 4868 18468 4924
rect 18468 4868 18524 4924
rect 18524 4868 18528 4924
rect 18464 4864 18528 4868
rect 18544 4924 18608 4928
rect 18544 4868 18548 4924
rect 18548 4868 18604 4924
rect 18604 4868 18608 4924
rect 18544 4864 18608 4868
rect 18624 4924 18688 4928
rect 18624 4868 18628 4924
rect 18628 4868 18684 4924
rect 18684 4868 18688 4924
rect 18624 4864 18688 4868
rect 36784 4924 36848 4928
rect 36784 4868 36788 4924
rect 36788 4868 36844 4924
rect 36844 4868 36848 4924
rect 36784 4864 36848 4868
rect 36864 4924 36928 4928
rect 36864 4868 36868 4924
rect 36868 4868 36924 4924
rect 36924 4868 36928 4924
rect 36864 4864 36928 4868
rect 36944 4924 37008 4928
rect 36944 4868 36948 4924
rect 36948 4868 37004 4924
rect 37004 4868 37008 4924
rect 36944 4864 37008 4868
rect 37024 4924 37088 4928
rect 37024 4868 37028 4924
rect 37028 4868 37084 4924
rect 37084 4868 37088 4924
rect 37024 4864 37088 4868
rect 55184 4924 55248 4928
rect 55184 4868 55188 4924
rect 55188 4868 55244 4924
rect 55244 4868 55248 4924
rect 55184 4864 55248 4868
rect 55264 4924 55328 4928
rect 55264 4868 55268 4924
rect 55268 4868 55324 4924
rect 55324 4868 55328 4924
rect 55264 4864 55328 4868
rect 55344 4924 55408 4928
rect 55344 4868 55348 4924
rect 55348 4868 55404 4924
rect 55404 4868 55408 4924
rect 55344 4864 55408 4868
rect 55424 4924 55488 4928
rect 55424 4868 55428 4924
rect 55428 4868 55484 4924
rect 55484 4868 55488 4924
rect 55424 4864 55488 4868
rect 73584 4924 73648 4928
rect 73584 4868 73588 4924
rect 73588 4868 73644 4924
rect 73644 4868 73648 4924
rect 73584 4864 73648 4868
rect 73664 4924 73728 4928
rect 73664 4868 73668 4924
rect 73668 4868 73724 4924
rect 73724 4868 73728 4924
rect 73664 4864 73728 4868
rect 73744 4924 73808 4928
rect 73744 4868 73748 4924
rect 73748 4868 73804 4924
rect 73804 4868 73808 4924
rect 73744 4864 73808 4868
rect 73824 4924 73888 4928
rect 73824 4868 73828 4924
rect 73828 4868 73884 4924
rect 73884 4868 73888 4924
rect 73824 4864 73888 4868
<< metal4 >>
rect 2696 89722 3016 89764
rect 2696 89486 2738 89722
rect 2974 89486 3016 89722
rect 2696 73874 3016 89486
rect 2696 73638 2738 73874
rect 2974 73638 3016 73874
rect 2696 55474 3016 73638
rect 2696 55238 2738 55474
rect 2974 55238 3016 55474
rect 2696 37074 3016 55238
rect 2696 36838 2738 37074
rect 2974 36838 3016 37074
rect 2696 18674 3016 36838
rect 2696 18438 2738 18674
rect 2974 18438 3016 18674
rect 2696 2994 3016 18438
rect 3356 89062 3676 89104
rect 3356 88826 3398 89062
rect 3634 88826 3676 89062
rect 3356 73214 3676 88826
rect 17716 89062 18036 89764
rect 17716 88826 17758 89062
rect 17994 88826 18036 89062
rect 10307 87380 10373 87381
rect 10307 87316 10308 87380
rect 10372 87316 10373 87380
rect 10307 87315 10373 87316
rect 3356 72978 3398 73214
rect 3634 72978 3676 73214
rect 3356 54814 3676 72978
rect 3356 54578 3398 54814
rect 3634 54578 3676 54814
rect 3356 36414 3676 54578
rect 3356 36178 3398 36414
rect 3634 36178 3676 36414
rect 3356 18014 3676 36178
rect 3356 17778 3398 18014
rect 3634 17778 3676 18014
rect 3356 3654 3676 17778
rect 5948 84896 6268 84912
rect 5948 84832 5956 84896
rect 6020 84832 6036 84896
rect 6100 84832 6116 84896
rect 6180 84832 6196 84896
rect 6260 84832 6268 84896
rect 5948 83808 6268 84832
rect 5948 83744 5956 83808
rect 6020 83744 6036 83808
rect 6100 83744 6116 83808
rect 6180 83744 6196 83808
rect 6260 83744 6268 83808
rect 5948 82720 6268 83744
rect 5948 82656 5956 82720
rect 6020 82656 6036 82720
rect 6100 82656 6116 82720
rect 6180 82656 6196 82720
rect 6260 82656 6268 82720
rect 5948 81632 6268 82656
rect 5948 81568 5956 81632
rect 6020 81568 6036 81632
rect 6100 81568 6116 81632
rect 6180 81568 6196 81632
rect 6260 81568 6268 81632
rect 5948 80544 6268 81568
rect 5948 80480 5956 80544
rect 6020 80480 6036 80544
rect 6100 80480 6116 80544
rect 6180 80480 6196 80544
rect 6260 80480 6268 80544
rect 5948 79456 6268 80480
rect 5948 79392 5956 79456
rect 6020 79392 6036 79456
rect 6100 79392 6116 79456
rect 6180 79392 6196 79456
rect 6260 79392 6268 79456
rect 5948 78368 6268 79392
rect 5948 78304 5956 78368
rect 6020 78304 6036 78368
rect 6100 78304 6116 78368
rect 6180 78304 6196 78368
rect 6260 78304 6268 78368
rect 5948 77280 6268 78304
rect 5948 77216 5956 77280
rect 6020 77216 6036 77280
rect 6100 77216 6116 77280
rect 6180 77216 6196 77280
rect 6260 77216 6268 77280
rect 5948 76192 6268 77216
rect 5948 76128 5956 76192
rect 6020 76128 6036 76192
rect 6100 76128 6116 76192
rect 6180 76128 6196 76192
rect 6260 76128 6268 76192
rect 5948 75104 6268 76128
rect 5948 75040 5956 75104
rect 6020 75040 6036 75104
rect 6100 75040 6116 75104
rect 6180 75040 6196 75104
rect 6260 75040 6268 75104
rect 5948 74016 6268 75040
rect 5948 73952 5956 74016
rect 6020 73952 6036 74016
rect 6100 73952 6116 74016
rect 6180 73952 6196 74016
rect 6260 73952 6268 74016
rect 5948 73214 6268 73952
rect 5948 72978 5990 73214
rect 6226 72978 6268 73214
rect 5948 72928 6268 72978
rect 5948 72864 5956 72928
rect 6020 72864 6036 72928
rect 6100 72864 6116 72928
rect 6180 72864 6196 72928
rect 6260 72864 6268 72928
rect 5948 71840 6268 72864
rect 5948 71776 5956 71840
rect 6020 71776 6036 71840
rect 6100 71776 6116 71840
rect 6180 71776 6196 71840
rect 6260 71776 6268 71840
rect 5948 70752 6268 71776
rect 5948 70688 5956 70752
rect 6020 70688 6036 70752
rect 6100 70688 6116 70752
rect 6180 70688 6196 70752
rect 6260 70688 6268 70752
rect 5948 69664 6268 70688
rect 5948 69600 5956 69664
rect 6020 69600 6036 69664
rect 6100 69600 6116 69664
rect 6180 69600 6196 69664
rect 6260 69600 6268 69664
rect 5948 68576 6268 69600
rect 5948 68512 5956 68576
rect 6020 68512 6036 68576
rect 6100 68512 6116 68576
rect 6180 68512 6196 68576
rect 6260 68512 6268 68576
rect 5948 67488 6268 68512
rect 5948 67424 5956 67488
rect 6020 67424 6036 67488
rect 6100 67424 6116 67488
rect 6180 67424 6196 67488
rect 6260 67424 6268 67488
rect 5948 66400 6268 67424
rect 5948 66336 5956 66400
rect 6020 66336 6036 66400
rect 6100 66336 6116 66400
rect 6180 66336 6196 66400
rect 6260 66336 6268 66400
rect 5948 65312 6268 66336
rect 5948 65248 5956 65312
rect 6020 65248 6036 65312
rect 6100 65248 6116 65312
rect 6180 65248 6196 65312
rect 6260 65248 6268 65312
rect 5948 64224 6268 65248
rect 5948 64160 5956 64224
rect 6020 64160 6036 64224
rect 6100 64160 6116 64224
rect 6180 64160 6196 64224
rect 6260 64160 6268 64224
rect 5948 63136 6268 64160
rect 5948 63072 5956 63136
rect 6020 63072 6036 63136
rect 6100 63072 6116 63136
rect 6180 63072 6196 63136
rect 6260 63072 6268 63136
rect 5948 62048 6268 63072
rect 5948 61984 5956 62048
rect 6020 61984 6036 62048
rect 6100 61984 6116 62048
rect 6180 61984 6196 62048
rect 6260 61984 6268 62048
rect 5948 60960 6268 61984
rect 5948 60896 5956 60960
rect 6020 60896 6036 60960
rect 6100 60896 6116 60960
rect 6180 60896 6196 60960
rect 6260 60896 6268 60960
rect 5948 59872 6268 60896
rect 5948 59808 5956 59872
rect 6020 59808 6036 59872
rect 6100 59808 6116 59872
rect 6180 59808 6196 59872
rect 6260 59808 6268 59872
rect 5948 58784 6268 59808
rect 5948 58720 5956 58784
rect 6020 58720 6036 58784
rect 6100 58720 6116 58784
rect 6180 58720 6196 58784
rect 6260 58720 6268 58784
rect 5948 57696 6268 58720
rect 5948 57632 5956 57696
rect 6020 57632 6036 57696
rect 6100 57632 6116 57696
rect 6180 57632 6196 57696
rect 6260 57632 6268 57696
rect 5948 56608 6268 57632
rect 5948 56544 5956 56608
rect 6020 56544 6036 56608
rect 6100 56544 6116 56608
rect 6180 56544 6196 56608
rect 6260 56544 6268 56608
rect 5948 55520 6268 56544
rect 5948 55456 5956 55520
rect 6020 55456 6036 55520
rect 6100 55456 6116 55520
rect 6180 55456 6196 55520
rect 6260 55456 6268 55520
rect 5948 54814 6268 55456
rect 5948 54578 5990 54814
rect 6226 54578 6268 54814
rect 5948 54432 6268 54578
rect 5948 54368 5956 54432
rect 6020 54368 6036 54432
rect 6100 54368 6116 54432
rect 6180 54368 6196 54432
rect 6260 54368 6268 54432
rect 5948 53344 6268 54368
rect 5948 53280 5956 53344
rect 6020 53280 6036 53344
rect 6100 53280 6116 53344
rect 6180 53280 6196 53344
rect 6260 53280 6268 53344
rect 5948 52256 6268 53280
rect 5948 52192 5956 52256
rect 6020 52192 6036 52256
rect 6100 52192 6116 52256
rect 6180 52192 6196 52256
rect 6260 52192 6268 52256
rect 5948 51168 6268 52192
rect 5948 51104 5956 51168
rect 6020 51104 6036 51168
rect 6100 51104 6116 51168
rect 6180 51104 6196 51168
rect 6260 51104 6268 51168
rect 5948 50080 6268 51104
rect 5948 50016 5956 50080
rect 6020 50016 6036 50080
rect 6100 50016 6116 50080
rect 6180 50016 6196 50080
rect 6260 50016 6268 50080
rect 5948 48992 6268 50016
rect 5948 48928 5956 48992
rect 6020 48928 6036 48992
rect 6100 48928 6116 48992
rect 6180 48928 6196 48992
rect 6260 48928 6268 48992
rect 5948 47904 6268 48928
rect 5948 47840 5956 47904
rect 6020 47840 6036 47904
rect 6100 47840 6116 47904
rect 6180 47840 6196 47904
rect 6260 47840 6268 47904
rect 5948 46816 6268 47840
rect 5948 46752 5956 46816
rect 6020 46752 6036 46816
rect 6100 46752 6116 46816
rect 6180 46752 6196 46816
rect 6260 46752 6268 46816
rect 5948 45728 6268 46752
rect 5948 45664 5956 45728
rect 6020 45664 6036 45728
rect 6100 45664 6116 45728
rect 6180 45664 6196 45728
rect 6260 45664 6268 45728
rect 5948 44640 6268 45664
rect 5948 44576 5956 44640
rect 6020 44576 6036 44640
rect 6100 44576 6116 44640
rect 6180 44576 6196 44640
rect 6260 44576 6268 44640
rect 5948 43552 6268 44576
rect 5948 43488 5956 43552
rect 6020 43488 6036 43552
rect 6100 43488 6116 43552
rect 6180 43488 6196 43552
rect 6260 43488 6268 43552
rect 5948 42464 6268 43488
rect 5948 42400 5956 42464
rect 6020 42400 6036 42464
rect 6100 42400 6116 42464
rect 6180 42400 6196 42464
rect 6260 42400 6268 42464
rect 5948 41376 6268 42400
rect 5948 41312 5956 41376
rect 6020 41312 6036 41376
rect 6100 41312 6116 41376
rect 6180 41312 6196 41376
rect 6260 41312 6268 41376
rect 5948 40288 6268 41312
rect 5948 40224 5956 40288
rect 6020 40224 6036 40288
rect 6100 40224 6116 40288
rect 6180 40224 6196 40288
rect 6260 40224 6268 40288
rect 5948 39200 6268 40224
rect 5948 39136 5956 39200
rect 6020 39136 6036 39200
rect 6100 39136 6116 39200
rect 6180 39136 6196 39200
rect 6260 39136 6268 39200
rect 5948 38112 6268 39136
rect 5948 38048 5956 38112
rect 6020 38048 6036 38112
rect 6100 38048 6116 38112
rect 6180 38048 6196 38112
rect 6260 38048 6268 38112
rect 5948 37024 6268 38048
rect 5948 36960 5956 37024
rect 6020 36960 6036 37024
rect 6100 36960 6116 37024
rect 6180 36960 6196 37024
rect 6260 36960 6268 37024
rect 5948 36414 6268 36960
rect 5948 36178 5990 36414
rect 6226 36178 6268 36414
rect 5948 35936 6268 36178
rect 5948 35872 5956 35936
rect 6020 35872 6036 35936
rect 6100 35872 6116 35936
rect 6180 35872 6196 35936
rect 6260 35872 6268 35936
rect 5948 34848 6268 35872
rect 5948 34784 5956 34848
rect 6020 34784 6036 34848
rect 6100 34784 6116 34848
rect 6180 34784 6196 34848
rect 6260 34784 6268 34848
rect 5948 33760 6268 34784
rect 5948 33696 5956 33760
rect 6020 33696 6036 33760
rect 6100 33696 6116 33760
rect 6180 33696 6196 33760
rect 6260 33696 6268 33760
rect 5948 32672 6268 33696
rect 5948 32608 5956 32672
rect 6020 32608 6036 32672
rect 6100 32608 6116 32672
rect 6180 32608 6196 32672
rect 6260 32608 6268 32672
rect 5948 31584 6268 32608
rect 5948 31520 5956 31584
rect 6020 31520 6036 31584
rect 6100 31520 6116 31584
rect 6180 31520 6196 31584
rect 6260 31520 6268 31584
rect 5948 30496 6268 31520
rect 5948 30432 5956 30496
rect 6020 30432 6036 30496
rect 6100 30432 6116 30496
rect 6180 30432 6196 30496
rect 6260 30432 6268 30496
rect 5948 29408 6268 30432
rect 5948 29344 5956 29408
rect 6020 29344 6036 29408
rect 6100 29344 6116 29408
rect 6180 29344 6196 29408
rect 6260 29344 6268 29408
rect 5948 28320 6268 29344
rect 5948 28256 5956 28320
rect 6020 28256 6036 28320
rect 6100 28256 6116 28320
rect 6180 28256 6196 28320
rect 6260 28256 6268 28320
rect 5948 27232 6268 28256
rect 5948 27168 5956 27232
rect 6020 27168 6036 27232
rect 6100 27168 6116 27232
rect 6180 27168 6196 27232
rect 6260 27168 6268 27232
rect 5948 26144 6268 27168
rect 5948 26080 5956 26144
rect 6020 26080 6036 26144
rect 6100 26080 6116 26144
rect 6180 26080 6196 26144
rect 6260 26080 6268 26144
rect 5948 25056 6268 26080
rect 5948 24992 5956 25056
rect 6020 24992 6036 25056
rect 6100 24992 6116 25056
rect 6180 24992 6196 25056
rect 6260 24992 6268 25056
rect 5948 23968 6268 24992
rect 5948 23904 5956 23968
rect 6020 23904 6036 23968
rect 6100 23904 6116 23968
rect 6180 23904 6196 23968
rect 6260 23904 6268 23968
rect 5948 22880 6268 23904
rect 5948 22816 5956 22880
rect 6020 22816 6036 22880
rect 6100 22816 6116 22880
rect 6180 22816 6196 22880
rect 6260 22816 6268 22880
rect 5948 21792 6268 22816
rect 5948 21728 5956 21792
rect 6020 21728 6036 21792
rect 6100 21728 6116 21792
rect 6180 21728 6196 21792
rect 6260 21728 6268 21792
rect 5948 20704 6268 21728
rect 5948 20640 5956 20704
rect 6020 20640 6036 20704
rect 6100 20640 6116 20704
rect 6180 20640 6196 20704
rect 6260 20640 6268 20704
rect 5948 19616 6268 20640
rect 5948 19552 5956 19616
rect 6020 19552 6036 19616
rect 6100 19552 6116 19616
rect 6180 19552 6196 19616
rect 6260 19552 6268 19616
rect 5948 18528 6268 19552
rect 5948 18464 5956 18528
rect 6020 18464 6036 18528
rect 6100 18464 6116 18528
rect 6180 18464 6196 18528
rect 6260 18464 6268 18528
rect 5948 18014 6268 18464
rect 5948 17778 5990 18014
rect 6226 17778 6268 18014
rect 5948 17440 6268 17778
rect 5948 17376 5956 17440
rect 6020 17376 6036 17440
rect 6100 17376 6116 17440
rect 6180 17376 6196 17440
rect 6260 17376 6268 17440
rect 5948 16352 6268 17376
rect 5948 16288 5956 16352
rect 6020 16288 6036 16352
rect 6100 16288 6116 16352
rect 6180 16288 6196 16352
rect 6260 16288 6268 16352
rect 5948 15264 6268 16288
rect 5948 15200 5956 15264
rect 6020 15200 6036 15264
rect 6100 15200 6116 15264
rect 6180 15200 6196 15264
rect 6260 15200 6268 15264
rect 5948 14176 6268 15200
rect 5948 14112 5956 14176
rect 6020 14112 6036 14176
rect 6100 14112 6116 14176
rect 6180 14112 6196 14176
rect 6260 14112 6268 14176
rect 5948 13088 6268 14112
rect 5948 13024 5956 13088
rect 6020 13024 6036 13088
rect 6100 13024 6116 13088
rect 6180 13024 6196 13088
rect 6260 13024 6268 13088
rect 5948 12000 6268 13024
rect 5948 11936 5956 12000
rect 6020 11936 6036 12000
rect 6100 11936 6116 12000
rect 6180 11936 6196 12000
rect 6260 11936 6268 12000
rect 5948 10912 6268 11936
rect 5948 10848 5956 10912
rect 6020 10848 6036 10912
rect 6100 10848 6116 10912
rect 6180 10848 6196 10912
rect 6260 10848 6268 10912
rect 5948 9824 6268 10848
rect 5948 9760 5956 9824
rect 6020 9760 6036 9824
rect 6100 9760 6116 9824
rect 6180 9760 6196 9824
rect 6260 9760 6268 9824
rect 5948 8736 6268 9760
rect 5948 8672 5956 8736
rect 6020 8672 6036 8736
rect 6100 8672 6116 8736
rect 6180 8672 6196 8736
rect 6260 8672 6268 8736
rect 5948 7648 6268 8672
rect 5948 7584 5956 7648
rect 6020 7584 6036 7648
rect 6100 7584 6116 7648
rect 6180 7584 6196 7648
rect 6260 7584 6268 7648
rect 5948 7024 6268 7584
rect 6684 84352 7004 84912
rect 6684 84288 6692 84352
rect 6756 84288 6772 84352
rect 6836 84288 6852 84352
rect 6916 84288 6932 84352
rect 6996 84288 7004 84352
rect 6684 83264 7004 84288
rect 6684 83200 6692 83264
rect 6756 83200 6772 83264
rect 6836 83200 6852 83264
rect 6916 83200 6932 83264
rect 6996 83200 7004 83264
rect 6684 82176 7004 83200
rect 6684 82112 6692 82176
rect 6756 82112 6772 82176
rect 6836 82112 6852 82176
rect 6916 82112 6932 82176
rect 6996 82112 7004 82176
rect 6684 81088 7004 82112
rect 6684 81024 6692 81088
rect 6756 81024 6772 81088
rect 6836 81024 6852 81088
rect 6916 81024 6932 81088
rect 6996 81024 7004 81088
rect 10310 81057 10370 87315
rect 17716 87072 18036 88826
rect 17716 87008 17724 87072
rect 17788 87008 17804 87072
rect 17868 87008 17884 87072
rect 17948 87008 17964 87072
rect 18028 87008 18036 87072
rect 17716 85984 18036 87008
rect 17716 85920 17724 85984
rect 17788 85920 17804 85984
rect 17868 85920 17884 85984
rect 17948 85920 17964 85984
rect 18028 85920 18036 85984
rect 17716 84896 18036 85920
rect 17716 84832 17724 84896
rect 17788 84832 17804 84896
rect 17868 84832 17884 84896
rect 17948 84832 17964 84896
rect 18028 84832 18036 84896
rect 6684 80000 7004 81024
rect 10307 81056 10373 81057
rect 10307 80992 10308 81056
rect 10372 80992 10373 81056
rect 17716 81029 18036 84832
rect 18376 89722 18696 89764
rect 18376 89486 18418 89722
rect 18654 89486 18696 89722
rect 18376 87616 18696 89486
rect 18376 87552 18384 87616
rect 18448 87552 18464 87616
rect 18528 87552 18544 87616
rect 18608 87552 18624 87616
rect 18688 87552 18696 87616
rect 18376 86528 18696 87552
rect 18376 86464 18384 86528
rect 18448 86464 18464 86528
rect 18528 86464 18544 86528
rect 18608 86464 18624 86528
rect 18688 86464 18696 86528
rect 18376 85440 18696 86464
rect 18376 85376 18384 85440
rect 18448 85376 18464 85440
rect 18528 85376 18544 85440
rect 18608 85376 18624 85440
rect 18688 85376 18696 85440
rect 18376 84352 18696 85376
rect 18376 84288 18384 84352
rect 18448 84288 18464 84352
rect 18528 84288 18544 84352
rect 18608 84288 18624 84352
rect 18688 84288 18696 84352
rect 18376 81029 18696 84288
rect 36116 89062 36436 89764
rect 36116 88826 36158 89062
rect 36394 88826 36436 89062
rect 36116 87072 36436 88826
rect 36116 87008 36124 87072
rect 36188 87008 36204 87072
rect 36268 87008 36284 87072
rect 36348 87008 36364 87072
rect 36428 87008 36436 87072
rect 36116 85984 36436 87008
rect 36116 85920 36124 85984
rect 36188 85920 36204 85984
rect 36268 85920 36284 85984
rect 36348 85920 36364 85984
rect 36428 85920 36436 85984
rect 36116 84896 36436 85920
rect 36116 84832 36124 84896
rect 36188 84832 36204 84896
rect 36268 84832 36284 84896
rect 36348 84832 36364 84896
rect 36428 84832 36436 84896
rect 36116 81029 36436 84832
rect 36776 89722 37096 89764
rect 36776 89486 36818 89722
rect 37054 89486 37096 89722
rect 36776 87616 37096 89486
rect 36776 87552 36784 87616
rect 36848 87552 36864 87616
rect 36928 87552 36944 87616
rect 37008 87552 37024 87616
rect 37088 87552 37096 87616
rect 36776 86528 37096 87552
rect 36776 86464 36784 86528
rect 36848 86464 36864 86528
rect 36928 86464 36944 86528
rect 37008 86464 37024 86528
rect 37088 86464 37096 86528
rect 36776 85440 37096 86464
rect 36776 85376 36784 85440
rect 36848 85376 36864 85440
rect 36928 85376 36944 85440
rect 37008 85376 37024 85440
rect 37088 85376 37096 85440
rect 36776 84352 37096 85376
rect 36776 84288 36784 84352
rect 36848 84288 36864 84352
rect 36928 84288 36944 84352
rect 37008 84288 37024 84352
rect 37088 84288 37096 84352
rect 36776 81029 37096 84288
rect 54516 89062 54836 89764
rect 54516 88826 54558 89062
rect 54794 88826 54836 89062
rect 54516 87072 54836 88826
rect 54516 87008 54524 87072
rect 54588 87008 54604 87072
rect 54668 87008 54684 87072
rect 54748 87008 54764 87072
rect 54828 87008 54836 87072
rect 54516 85984 54836 87008
rect 54516 85920 54524 85984
rect 54588 85920 54604 85984
rect 54668 85920 54684 85984
rect 54748 85920 54764 85984
rect 54828 85920 54836 85984
rect 54516 84896 54836 85920
rect 54516 84832 54524 84896
rect 54588 84832 54604 84896
rect 54668 84832 54684 84896
rect 54748 84832 54764 84896
rect 54828 84832 54836 84896
rect 54516 81029 54836 84832
rect 55176 89722 55496 89764
rect 55176 89486 55218 89722
rect 55454 89486 55496 89722
rect 55176 87616 55496 89486
rect 55176 87552 55184 87616
rect 55248 87552 55264 87616
rect 55328 87552 55344 87616
rect 55408 87552 55424 87616
rect 55488 87552 55496 87616
rect 55176 86528 55496 87552
rect 55176 86464 55184 86528
rect 55248 86464 55264 86528
rect 55328 86464 55344 86528
rect 55408 86464 55424 86528
rect 55488 86464 55496 86528
rect 55176 85440 55496 86464
rect 55176 85376 55184 85440
rect 55248 85376 55264 85440
rect 55328 85376 55344 85440
rect 55408 85376 55424 85440
rect 55488 85376 55496 85440
rect 55176 84352 55496 85376
rect 55176 84288 55184 84352
rect 55248 84288 55264 84352
rect 55328 84288 55344 84352
rect 55408 84288 55424 84352
rect 55488 84288 55496 84352
rect 55176 81029 55496 84288
rect 72916 89062 73236 89764
rect 72916 88826 72958 89062
rect 73194 88826 73236 89062
rect 72916 87072 73236 88826
rect 72916 87008 72924 87072
rect 72988 87008 73004 87072
rect 73068 87008 73084 87072
rect 73148 87008 73164 87072
rect 73228 87008 73236 87072
rect 72916 85984 73236 87008
rect 72916 85920 72924 85984
rect 72988 85920 73004 85984
rect 73068 85920 73084 85984
rect 73148 85920 73164 85984
rect 73228 85920 73236 85984
rect 72916 84896 73236 85920
rect 72916 84832 72924 84896
rect 72988 84832 73004 84896
rect 73068 84832 73084 84896
rect 73148 84832 73164 84896
rect 73228 84832 73236 84896
rect 72916 81029 73236 84832
rect 73576 89722 73896 89764
rect 73576 89486 73618 89722
rect 73854 89486 73896 89722
rect 73576 87616 73896 89486
rect 90456 89722 90776 89764
rect 90456 89486 90498 89722
rect 90734 89486 90776 89722
rect 73576 87552 73584 87616
rect 73648 87552 73664 87616
rect 73728 87552 73744 87616
rect 73808 87552 73824 87616
rect 73888 87552 73896 87616
rect 73576 86528 73896 87552
rect 73576 86464 73584 86528
rect 73648 86464 73664 86528
rect 73728 86464 73744 86528
rect 73808 86464 73824 86528
rect 73888 86464 73896 86528
rect 73576 85440 73896 86464
rect 73576 85376 73584 85440
rect 73648 85376 73664 85440
rect 73728 85376 73744 85440
rect 73808 85376 73824 85440
rect 73888 85376 73896 85440
rect 73576 84352 73896 85376
rect 89796 89062 90116 89104
rect 89796 88826 89838 89062
rect 90074 88826 90116 89062
rect 73576 84288 73584 84352
rect 73648 84288 73664 84352
rect 73728 84288 73744 84352
rect 73808 84288 73824 84352
rect 73888 84288 73896 84352
rect 73576 81029 73896 84288
rect 86540 84896 86860 84912
rect 86540 84832 86548 84896
rect 86612 84832 86628 84896
rect 86692 84832 86708 84896
rect 86772 84832 86788 84896
rect 86852 84832 86860 84896
rect 86540 83808 86860 84832
rect 86540 83744 86548 83808
rect 86612 83744 86628 83808
rect 86692 83744 86708 83808
rect 86772 83744 86788 83808
rect 86852 83744 86860 83808
rect 86540 82720 86860 83744
rect 86540 82656 86548 82720
rect 86612 82656 86628 82720
rect 86692 82656 86708 82720
rect 86772 82656 86788 82720
rect 86852 82656 86860 82720
rect 86540 81632 86860 82656
rect 86540 81568 86548 81632
rect 86612 81568 86628 81632
rect 86692 81568 86708 81632
rect 86772 81568 86788 81632
rect 86852 81568 86860 81632
rect 10307 80991 10373 80992
rect 11144 80630 11186 80866
rect 11422 80630 11464 80866
rect 43744 80630 43786 80866
rect 44022 80630 44064 80866
rect 48544 80630 48586 80866
rect 48822 80630 48864 80866
rect 81144 80630 81186 80866
rect 81422 80630 81464 80866
rect 86540 80544 86860 81568
rect 86540 80480 86548 80544
rect 86612 80480 86628 80544
rect 86692 80480 86708 80544
rect 86772 80480 86788 80544
rect 86852 80480 86860 80544
rect 6684 79936 6692 80000
rect 6756 79936 6772 80000
rect 6836 79936 6852 80000
rect 6916 79936 6932 80000
rect 6996 79936 7004 80000
rect 10484 79970 10526 80206
rect 10762 79970 10804 80206
rect 43084 79970 43126 80206
rect 43362 79970 43404 80206
rect 47884 79970 47926 80206
rect 48162 79970 48204 80206
rect 80484 79970 80526 80206
rect 80762 79970 80804 80206
rect 6684 78912 7004 79936
rect 6684 78848 6692 78912
rect 6756 78848 6772 78912
rect 6836 78848 6852 78912
rect 6916 78848 6932 78912
rect 6996 78848 7004 78912
rect 6684 77824 7004 78848
rect 6684 77760 6692 77824
rect 6756 77760 6772 77824
rect 6836 77760 6852 77824
rect 6916 77760 6932 77824
rect 6996 77760 7004 77824
rect 6684 76736 7004 77760
rect 6684 76672 6692 76736
rect 6756 76672 6772 76736
rect 6836 76672 6852 76736
rect 6916 76672 6932 76736
rect 6996 76672 7004 76736
rect 6684 75648 7004 76672
rect 6684 75584 6692 75648
rect 6756 75584 6772 75648
rect 6836 75584 6852 75648
rect 6916 75584 6932 75648
rect 6996 75584 7004 75648
rect 6684 74560 7004 75584
rect 6684 74496 6692 74560
rect 6756 74496 6772 74560
rect 6836 74496 6852 74560
rect 6916 74496 6932 74560
rect 6996 74496 7004 74560
rect 6684 73874 7004 74496
rect 86540 79456 86860 80480
rect 86540 79392 86548 79456
rect 86612 79392 86628 79456
rect 86692 79392 86708 79456
rect 86772 79392 86788 79456
rect 86852 79392 86860 79456
rect 86540 78368 86860 79392
rect 86540 78304 86548 78368
rect 86612 78304 86628 78368
rect 86692 78304 86708 78368
rect 86772 78304 86788 78368
rect 86852 78304 86860 78368
rect 86540 77280 86860 78304
rect 86540 77216 86548 77280
rect 86612 77216 86628 77280
rect 86692 77216 86708 77280
rect 86772 77216 86788 77280
rect 86852 77216 86860 77280
rect 86540 76192 86860 77216
rect 86540 76128 86548 76192
rect 86612 76128 86628 76192
rect 86692 76128 86708 76192
rect 86772 76128 86788 76192
rect 86852 76128 86860 76192
rect 86540 75104 86860 76128
rect 86540 75040 86548 75104
rect 86612 75040 86628 75104
rect 86692 75040 86708 75104
rect 86772 75040 86788 75104
rect 86852 75040 86860 75104
rect 86540 74016 86860 75040
rect 86540 73952 86548 74016
rect 86612 73952 86628 74016
rect 86692 73952 86708 74016
rect 86772 73952 86788 74016
rect 86852 73952 86860 74016
rect 6684 73638 6726 73874
rect 6962 73638 7004 73874
rect 11144 73638 11186 73874
rect 11422 73638 11464 73874
rect 43744 73638 43786 73874
rect 44022 73638 44064 73874
rect 48544 73638 48586 73874
rect 48822 73638 48864 73874
rect 81144 73638 81186 73874
rect 81422 73638 81464 73874
rect 6684 73472 7004 73638
rect 6684 73408 6692 73472
rect 6756 73408 6772 73472
rect 6836 73408 6852 73472
rect 6916 73408 6932 73472
rect 6996 73408 7004 73472
rect 6684 72384 7004 73408
rect 86540 73214 86860 73952
rect 10484 72978 10526 73214
rect 10762 72978 10804 73214
rect 43084 72978 43126 73214
rect 43362 72978 43404 73214
rect 47884 72978 47926 73214
rect 48162 72978 48204 73214
rect 80484 72978 80526 73214
rect 80762 72978 80804 73214
rect 86540 72978 86582 73214
rect 86818 72978 86860 73214
rect 6684 72320 6692 72384
rect 6756 72320 6772 72384
rect 6836 72320 6852 72384
rect 6916 72320 6932 72384
rect 6996 72320 7004 72384
rect 6684 71296 7004 72320
rect 6684 71232 6692 71296
rect 6756 71232 6772 71296
rect 6836 71232 6852 71296
rect 6916 71232 6932 71296
rect 6996 71232 7004 71296
rect 6684 70208 7004 71232
rect 6684 70144 6692 70208
rect 6756 70144 6772 70208
rect 6836 70144 6852 70208
rect 6916 70144 6932 70208
rect 6996 70144 7004 70208
rect 6684 69120 7004 70144
rect 6684 69056 6692 69120
rect 6756 69056 6772 69120
rect 6836 69056 6852 69120
rect 6916 69056 6932 69120
rect 6996 69056 7004 69120
rect 6684 68032 7004 69056
rect 6684 67968 6692 68032
rect 6756 67968 6772 68032
rect 6836 67968 6852 68032
rect 6916 67968 6932 68032
rect 6996 67968 7004 68032
rect 6684 66944 7004 67968
rect 6684 66880 6692 66944
rect 6756 66880 6772 66944
rect 6836 66880 6852 66944
rect 6916 66880 6932 66944
rect 6996 66880 7004 66944
rect 6684 65856 7004 66880
rect 6684 65792 6692 65856
rect 6756 65792 6772 65856
rect 6836 65792 6852 65856
rect 6916 65792 6932 65856
rect 6996 65792 7004 65856
rect 6684 64768 7004 65792
rect 6684 64704 6692 64768
rect 6756 64704 6772 64768
rect 6836 64704 6852 64768
rect 6916 64704 6932 64768
rect 6996 64704 7004 64768
rect 6684 63680 7004 64704
rect 6684 63616 6692 63680
rect 6756 63616 6772 63680
rect 6836 63616 6852 63680
rect 6916 63616 6932 63680
rect 6996 63616 7004 63680
rect 6684 62592 7004 63616
rect 6684 62528 6692 62592
rect 6756 62528 6772 62592
rect 6836 62528 6852 62592
rect 6916 62528 6932 62592
rect 6996 62528 7004 62592
rect 6684 61504 7004 62528
rect 6684 61440 6692 61504
rect 6756 61440 6772 61504
rect 6836 61440 6852 61504
rect 6916 61440 6932 61504
rect 6996 61440 7004 61504
rect 6684 60416 7004 61440
rect 6684 60352 6692 60416
rect 6756 60352 6772 60416
rect 6836 60352 6852 60416
rect 6916 60352 6932 60416
rect 6996 60352 7004 60416
rect 6684 59328 7004 60352
rect 6684 59264 6692 59328
rect 6756 59264 6772 59328
rect 6836 59264 6852 59328
rect 6916 59264 6932 59328
rect 6996 59264 7004 59328
rect 6684 58240 7004 59264
rect 6684 58176 6692 58240
rect 6756 58176 6772 58240
rect 6836 58176 6852 58240
rect 6916 58176 6932 58240
rect 6996 58176 7004 58240
rect 6684 57152 7004 58176
rect 6684 57088 6692 57152
rect 6756 57088 6772 57152
rect 6836 57088 6852 57152
rect 6916 57088 6932 57152
rect 6996 57088 7004 57152
rect 6684 56064 7004 57088
rect 6684 56000 6692 56064
rect 6756 56000 6772 56064
rect 6836 56000 6852 56064
rect 6916 56000 6932 56064
rect 6996 56000 7004 56064
rect 6684 55474 7004 56000
rect 86540 72928 86860 72978
rect 86540 72864 86548 72928
rect 86612 72864 86628 72928
rect 86692 72864 86708 72928
rect 86772 72864 86788 72928
rect 86852 72864 86860 72928
rect 86540 71840 86860 72864
rect 86540 71776 86548 71840
rect 86612 71776 86628 71840
rect 86692 71776 86708 71840
rect 86772 71776 86788 71840
rect 86852 71776 86860 71840
rect 86540 70752 86860 71776
rect 86540 70688 86548 70752
rect 86612 70688 86628 70752
rect 86692 70688 86708 70752
rect 86772 70688 86788 70752
rect 86852 70688 86860 70752
rect 86540 69664 86860 70688
rect 86540 69600 86548 69664
rect 86612 69600 86628 69664
rect 86692 69600 86708 69664
rect 86772 69600 86788 69664
rect 86852 69600 86860 69664
rect 86540 68576 86860 69600
rect 86540 68512 86548 68576
rect 86612 68512 86628 68576
rect 86692 68512 86708 68576
rect 86772 68512 86788 68576
rect 86852 68512 86860 68576
rect 86540 67488 86860 68512
rect 86540 67424 86548 67488
rect 86612 67424 86628 67488
rect 86692 67424 86708 67488
rect 86772 67424 86788 67488
rect 86852 67424 86860 67488
rect 86540 66400 86860 67424
rect 86540 66336 86548 66400
rect 86612 66336 86628 66400
rect 86692 66336 86708 66400
rect 86772 66336 86788 66400
rect 86852 66336 86860 66400
rect 86540 65312 86860 66336
rect 86540 65248 86548 65312
rect 86612 65248 86628 65312
rect 86692 65248 86708 65312
rect 86772 65248 86788 65312
rect 86852 65248 86860 65312
rect 86540 64224 86860 65248
rect 86540 64160 86548 64224
rect 86612 64160 86628 64224
rect 86692 64160 86708 64224
rect 86772 64160 86788 64224
rect 86852 64160 86860 64224
rect 86540 63136 86860 64160
rect 86540 63072 86548 63136
rect 86612 63072 86628 63136
rect 86692 63072 86708 63136
rect 86772 63072 86788 63136
rect 86852 63072 86860 63136
rect 86540 62048 86860 63072
rect 86540 61984 86548 62048
rect 86612 61984 86628 62048
rect 86692 61984 86708 62048
rect 86772 61984 86788 62048
rect 86852 61984 86860 62048
rect 86540 60960 86860 61984
rect 86540 60896 86548 60960
rect 86612 60896 86628 60960
rect 86692 60896 86708 60960
rect 86772 60896 86788 60960
rect 86852 60896 86860 60960
rect 86540 59872 86860 60896
rect 86540 59808 86548 59872
rect 86612 59808 86628 59872
rect 86692 59808 86708 59872
rect 86772 59808 86788 59872
rect 86852 59808 86860 59872
rect 86540 58784 86860 59808
rect 86540 58720 86548 58784
rect 86612 58720 86628 58784
rect 86692 58720 86708 58784
rect 86772 58720 86788 58784
rect 86852 58720 86860 58784
rect 86540 57696 86860 58720
rect 86540 57632 86548 57696
rect 86612 57632 86628 57696
rect 86692 57632 86708 57696
rect 86772 57632 86788 57696
rect 86852 57632 86860 57696
rect 86540 56608 86860 57632
rect 86540 56544 86548 56608
rect 86612 56544 86628 56608
rect 86692 56544 86708 56608
rect 86772 56544 86788 56608
rect 86852 56544 86860 56608
rect 86540 55520 86860 56544
rect 6684 55238 6726 55474
rect 6962 55238 7004 55474
rect 11144 55238 11186 55474
rect 11422 55238 11464 55474
rect 43744 55238 43786 55474
rect 44022 55238 44064 55474
rect 48544 55238 48586 55474
rect 48822 55238 48864 55474
rect 81144 55238 81186 55474
rect 81422 55238 81464 55474
rect 86540 55456 86548 55520
rect 86612 55456 86628 55520
rect 86692 55456 86708 55520
rect 86772 55456 86788 55520
rect 86852 55456 86860 55520
rect 6684 54976 7004 55238
rect 6684 54912 6692 54976
rect 6756 54912 6772 54976
rect 6836 54912 6852 54976
rect 6916 54912 6932 54976
rect 6996 54912 7004 54976
rect 6684 53888 7004 54912
rect 86540 54814 86860 55456
rect 10484 54578 10526 54814
rect 10762 54578 10804 54814
rect 43084 54578 43126 54814
rect 43362 54578 43404 54814
rect 47884 54578 47926 54814
rect 48162 54578 48204 54814
rect 80484 54578 80526 54814
rect 80762 54578 80804 54814
rect 86540 54578 86582 54814
rect 86818 54578 86860 54814
rect 6684 53824 6692 53888
rect 6756 53824 6772 53888
rect 6836 53824 6852 53888
rect 6916 53824 6932 53888
rect 6996 53824 7004 53888
rect 6684 52800 7004 53824
rect 6684 52736 6692 52800
rect 6756 52736 6772 52800
rect 6836 52736 6852 52800
rect 6916 52736 6932 52800
rect 6996 52736 7004 52800
rect 6684 51712 7004 52736
rect 6684 51648 6692 51712
rect 6756 51648 6772 51712
rect 6836 51648 6852 51712
rect 6916 51648 6932 51712
rect 6996 51648 7004 51712
rect 6684 50624 7004 51648
rect 6684 50560 6692 50624
rect 6756 50560 6772 50624
rect 6836 50560 6852 50624
rect 6916 50560 6932 50624
rect 6996 50560 7004 50624
rect 6684 49536 7004 50560
rect 6684 49472 6692 49536
rect 6756 49472 6772 49536
rect 6836 49472 6852 49536
rect 6916 49472 6932 49536
rect 6996 49472 7004 49536
rect 6684 48448 7004 49472
rect 6684 48384 6692 48448
rect 6756 48384 6772 48448
rect 6836 48384 6852 48448
rect 6916 48384 6932 48448
rect 6996 48384 7004 48448
rect 6684 47360 7004 48384
rect 86540 54432 86860 54578
rect 86540 54368 86548 54432
rect 86612 54368 86628 54432
rect 86692 54368 86708 54432
rect 86772 54368 86788 54432
rect 86852 54368 86860 54432
rect 86540 53344 86860 54368
rect 86540 53280 86548 53344
rect 86612 53280 86628 53344
rect 86692 53280 86708 53344
rect 86772 53280 86788 53344
rect 86852 53280 86860 53344
rect 86540 52256 86860 53280
rect 86540 52192 86548 52256
rect 86612 52192 86628 52256
rect 86692 52192 86708 52256
rect 86772 52192 86788 52256
rect 86852 52192 86860 52256
rect 86540 51168 86860 52192
rect 86540 51104 86548 51168
rect 86612 51104 86628 51168
rect 86692 51104 86708 51168
rect 86772 51104 86788 51168
rect 86852 51104 86860 51168
rect 86540 50080 86860 51104
rect 86540 50016 86548 50080
rect 86612 50016 86628 50080
rect 86692 50016 86708 50080
rect 86772 50016 86788 50080
rect 86852 50016 86860 50080
rect 86540 48992 86860 50016
rect 86540 48928 86548 48992
rect 86612 48928 86628 48992
rect 86692 48928 86708 48992
rect 86772 48928 86788 48992
rect 86852 48928 86860 48992
rect 11144 48030 11186 48266
rect 11422 48030 11464 48266
rect 43744 48030 43786 48266
rect 44022 48030 44064 48266
rect 48544 48030 48586 48266
rect 48822 48030 48864 48266
rect 81144 48030 81186 48266
rect 81422 48030 81464 48266
rect 86540 47904 86860 48928
rect 86540 47840 86548 47904
rect 86612 47840 86628 47904
rect 86692 47840 86708 47904
rect 86772 47840 86788 47904
rect 86852 47840 86860 47904
rect 10484 47370 10526 47606
rect 10762 47370 10804 47606
rect 43084 47370 43126 47606
rect 43362 47370 43404 47606
rect 47884 47370 47926 47606
rect 48162 47370 48204 47606
rect 80484 47370 80526 47606
rect 80762 47370 80804 47606
rect 6684 47296 6692 47360
rect 6756 47296 6772 47360
rect 6836 47296 6852 47360
rect 6916 47296 6932 47360
rect 6996 47296 7004 47360
rect 6684 46272 7004 47296
rect 6684 46208 6692 46272
rect 6756 46208 6772 46272
rect 6836 46208 6852 46272
rect 6916 46208 6932 46272
rect 6996 46208 7004 46272
rect 6684 45184 7004 46208
rect 6684 45120 6692 45184
rect 6756 45120 6772 45184
rect 6836 45120 6852 45184
rect 6916 45120 6932 45184
rect 6996 45120 7004 45184
rect 6684 44096 7004 45120
rect 86540 46816 86860 47840
rect 86540 46752 86548 46816
rect 86612 46752 86628 46816
rect 86692 46752 86708 46816
rect 86772 46752 86788 46816
rect 86852 46752 86860 46816
rect 86540 45728 86860 46752
rect 86540 45664 86548 45728
rect 86612 45664 86628 45728
rect 86692 45664 86708 45728
rect 86772 45664 86788 45728
rect 86852 45664 86860 45728
rect 86540 44640 86860 45664
rect 86540 44576 86548 44640
rect 86612 44576 86628 44640
rect 86692 44576 86708 44640
rect 86772 44576 86788 44640
rect 86852 44576 86860 44640
rect 11144 44230 11186 44466
rect 11422 44230 11464 44466
rect 43744 44230 43786 44466
rect 44022 44230 44064 44466
rect 48544 44230 48586 44466
rect 48822 44230 48864 44466
rect 81144 44230 81186 44466
rect 81422 44230 81464 44466
rect 6684 44032 6692 44096
rect 6756 44032 6772 44096
rect 6836 44032 6852 44096
rect 6916 44032 6932 44096
rect 6996 44032 7004 44096
rect 6684 43008 7004 44032
rect 10484 43570 10526 43806
rect 10762 43570 10804 43806
rect 43084 43570 43126 43806
rect 43362 43570 43404 43806
rect 47884 43570 47926 43806
rect 48162 43570 48204 43806
rect 80484 43570 80526 43806
rect 80762 43570 80804 43806
rect 6684 42944 6692 43008
rect 6756 42944 6772 43008
rect 6836 42944 6852 43008
rect 6916 42944 6932 43008
rect 6996 42944 7004 43008
rect 6684 41920 7004 42944
rect 6684 41856 6692 41920
rect 6756 41856 6772 41920
rect 6836 41856 6852 41920
rect 6916 41856 6932 41920
rect 6996 41856 7004 41920
rect 6684 40832 7004 41856
rect 6684 40768 6692 40832
rect 6756 40768 6772 40832
rect 6836 40768 6852 40832
rect 6916 40768 6932 40832
rect 6996 40768 7004 40832
rect 6684 39744 7004 40768
rect 6684 39680 6692 39744
rect 6756 39680 6772 39744
rect 6836 39680 6852 39744
rect 6916 39680 6932 39744
rect 6996 39680 7004 39744
rect 6684 38656 7004 39680
rect 6684 38592 6692 38656
rect 6756 38592 6772 38656
rect 6836 38592 6852 38656
rect 6916 38592 6932 38656
rect 6996 38592 7004 38656
rect 6684 37568 7004 38592
rect 6684 37504 6692 37568
rect 6756 37504 6772 37568
rect 6836 37504 6852 37568
rect 6916 37504 6932 37568
rect 6996 37504 7004 37568
rect 6684 37074 7004 37504
rect 86540 43552 86860 44576
rect 86540 43488 86548 43552
rect 86612 43488 86628 43552
rect 86692 43488 86708 43552
rect 86772 43488 86788 43552
rect 86852 43488 86860 43552
rect 86540 42464 86860 43488
rect 86540 42400 86548 42464
rect 86612 42400 86628 42464
rect 86692 42400 86708 42464
rect 86772 42400 86788 42464
rect 86852 42400 86860 42464
rect 86540 41376 86860 42400
rect 86540 41312 86548 41376
rect 86612 41312 86628 41376
rect 86692 41312 86708 41376
rect 86772 41312 86788 41376
rect 86852 41312 86860 41376
rect 86540 40288 86860 41312
rect 86540 40224 86548 40288
rect 86612 40224 86628 40288
rect 86692 40224 86708 40288
rect 86772 40224 86788 40288
rect 86852 40224 86860 40288
rect 86540 39200 86860 40224
rect 86540 39136 86548 39200
rect 86612 39136 86628 39200
rect 86692 39136 86708 39200
rect 86772 39136 86788 39200
rect 86852 39136 86860 39200
rect 86540 38112 86860 39136
rect 86540 38048 86548 38112
rect 86612 38048 86628 38112
rect 86692 38048 86708 38112
rect 86772 38048 86788 38112
rect 86852 38048 86860 38112
rect 6684 36838 6726 37074
rect 6962 36838 7004 37074
rect 11144 36838 11186 37074
rect 11422 36838 11464 37074
rect 43744 36838 43786 37074
rect 44022 36838 44064 37074
rect 48544 36838 48586 37074
rect 48822 36838 48864 37074
rect 81144 36838 81186 37074
rect 81422 36838 81464 37074
rect 86540 37024 86860 38048
rect 86540 36960 86548 37024
rect 86612 36960 86628 37024
rect 86692 36960 86708 37024
rect 86772 36960 86788 37024
rect 86852 36960 86860 37024
rect 6684 36480 7004 36838
rect 6684 36416 6692 36480
rect 6756 36416 6772 36480
rect 6836 36416 6852 36480
rect 6916 36416 6932 36480
rect 6996 36416 7004 36480
rect 6684 35392 7004 36416
rect 86540 36414 86860 36960
rect 10484 36178 10526 36414
rect 10762 36178 10804 36414
rect 43084 36178 43126 36414
rect 43362 36178 43404 36414
rect 47884 36178 47926 36414
rect 48162 36178 48204 36414
rect 80484 36178 80526 36414
rect 80762 36178 80804 36414
rect 86540 36178 86582 36414
rect 86818 36178 86860 36414
rect 6684 35328 6692 35392
rect 6756 35328 6772 35392
rect 6836 35328 6852 35392
rect 6916 35328 6932 35392
rect 6996 35328 7004 35392
rect 6684 34304 7004 35328
rect 6684 34240 6692 34304
rect 6756 34240 6772 34304
rect 6836 34240 6852 34304
rect 6916 34240 6932 34304
rect 6996 34240 7004 34304
rect 6684 33216 7004 34240
rect 6684 33152 6692 33216
rect 6756 33152 6772 33216
rect 6836 33152 6852 33216
rect 6916 33152 6932 33216
rect 6996 33152 7004 33216
rect 6684 32128 7004 33152
rect 6684 32064 6692 32128
rect 6756 32064 6772 32128
rect 6836 32064 6852 32128
rect 6916 32064 6932 32128
rect 6996 32064 7004 32128
rect 6684 31040 7004 32064
rect 6684 30976 6692 31040
rect 6756 30976 6772 31040
rect 6836 30976 6852 31040
rect 6916 30976 6932 31040
rect 6996 30976 7004 31040
rect 6684 29952 7004 30976
rect 6684 29888 6692 29952
rect 6756 29888 6772 29952
rect 6836 29888 6852 29952
rect 6916 29888 6932 29952
rect 6996 29888 7004 29952
rect 6684 28864 7004 29888
rect 6684 28800 6692 28864
rect 6756 28800 6772 28864
rect 6836 28800 6852 28864
rect 6916 28800 6932 28864
rect 6996 28800 7004 28864
rect 6684 27776 7004 28800
rect 6684 27712 6692 27776
rect 6756 27712 6772 27776
rect 6836 27712 6852 27776
rect 6916 27712 6932 27776
rect 6996 27712 7004 27776
rect 6684 26688 7004 27712
rect 6684 26624 6692 26688
rect 6756 26624 6772 26688
rect 6836 26624 6852 26688
rect 6916 26624 6932 26688
rect 6996 26624 7004 26688
rect 6684 25600 7004 26624
rect 6684 25536 6692 25600
rect 6756 25536 6772 25600
rect 6836 25536 6852 25600
rect 6916 25536 6932 25600
rect 6996 25536 7004 25600
rect 6684 24512 7004 25536
rect 6684 24448 6692 24512
rect 6756 24448 6772 24512
rect 6836 24448 6852 24512
rect 6916 24448 6932 24512
rect 6996 24448 7004 24512
rect 6684 23424 7004 24448
rect 6684 23360 6692 23424
rect 6756 23360 6772 23424
rect 6836 23360 6852 23424
rect 6916 23360 6932 23424
rect 6996 23360 7004 23424
rect 6684 22336 7004 23360
rect 6684 22272 6692 22336
rect 6756 22272 6772 22336
rect 6836 22272 6852 22336
rect 6916 22272 6932 22336
rect 6996 22272 7004 22336
rect 6684 21248 7004 22272
rect 6684 21184 6692 21248
rect 6756 21184 6772 21248
rect 6836 21184 6852 21248
rect 6916 21184 6932 21248
rect 6996 21184 7004 21248
rect 6684 20160 7004 21184
rect 6684 20096 6692 20160
rect 6756 20096 6772 20160
rect 6836 20096 6852 20160
rect 6916 20096 6932 20160
rect 6996 20096 7004 20160
rect 6684 19072 7004 20096
rect 6684 19008 6692 19072
rect 6756 19008 6772 19072
rect 6836 19008 6852 19072
rect 6916 19008 6932 19072
rect 6996 19008 7004 19072
rect 6684 18674 7004 19008
rect 86540 35936 86860 36178
rect 86540 35872 86548 35936
rect 86612 35872 86628 35936
rect 86692 35872 86708 35936
rect 86772 35872 86788 35936
rect 86852 35872 86860 35936
rect 86540 34848 86860 35872
rect 86540 34784 86548 34848
rect 86612 34784 86628 34848
rect 86692 34784 86708 34848
rect 86772 34784 86788 34848
rect 86852 34784 86860 34848
rect 86540 33760 86860 34784
rect 86540 33696 86548 33760
rect 86612 33696 86628 33760
rect 86692 33696 86708 33760
rect 86772 33696 86788 33760
rect 86852 33696 86860 33760
rect 86540 32672 86860 33696
rect 86540 32608 86548 32672
rect 86612 32608 86628 32672
rect 86692 32608 86708 32672
rect 86772 32608 86788 32672
rect 86852 32608 86860 32672
rect 86540 31584 86860 32608
rect 86540 31520 86548 31584
rect 86612 31520 86628 31584
rect 86692 31520 86708 31584
rect 86772 31520 86788 31584
rect 86852 31520 86860 31584
rect 86540 30496 86860 31520
rect 86540 30432 86548 30496
rect 86612 30432 86628 30496
rect 86692 30432 86708 30496
rect 86772 30432 86788 30496
rect 86852 30432 86860 30496
rect 86540 29408 86860 30432
rect 86540 29344 86548 29408
rect 86612 29344 86628 29408
rect 86692 29344 86708 29408
rect 86772 29344 86788 29408
rect 86852 29344 86860 29408
rect 86540 28320 86860 29344
rect 86540 28256 86548 28320
rect 86612 28256 86628 28320
rect 86692 28256 86708 28320
rect 86772 28256 86788 28320
rect 86852 28256 86860 28320
rect 86540 27232 86860 28256
rect 86540 27168 86548 27232
rect 86612 27168 86628 27232
rect 86692 27168 86708 27232
rect 86772 27168 86788 27232
rect 86852 27168 86860 27232
rect 86540 26144 86860 27168
rect 86540 26080 86548 26144
rect 86612 26080 86628 26144
rect 86692 26080 86708 26144
rect 86772 26080 86788 26144
rect 86852 26080 86860 26144
rect 86540 25056 86860 26080
rect 86540 24992 86548 25056
rect 86612 24992 86628 25056
rect 86692 24992 86708 25056
rect 86772 24992 86788 25056
rect 86852 24992 86860 25056
rect 86540 23968 86860 24992
rect 86540 23904 86548 23968
rect 86612 23904 86628 23968
rect 86692 23904 86708 23968
rect 86772 23904 86788 23968
rect 86852 23904 86860 23968
rect 86540 22880 86860 23904
rect 86540 22816 86548 22880
rect 86612 22816 86628 22880
rect 86692 22816 86708 22880
rect 86772 22816 86788 22880
rect 86852 22816 86860 22880
rect 86540 21792 86860 22816
rect 86540 21728 86548 21792
rect 86612 21728 86628 21792
rect 86692 21728 86708 21792
rect 86772 21728 86788 21792
rect 86852 21728 86860 21792
rect 86540 20704 86860 21728
rect 86540 20640 86548 20704
rect 86612 20640 86628 20704
rect 86692 20640 86708 20704
rect 86772 20640 86788 20704
rect 86852 20640 86860 20704
rect 86540 19616 86860 20640
rect 86540 19552 86548 19616
rect 86612 19552 86628 19616
rect 86692 19552 86708 19616
rect 86772 19552 86788 19616
rect 86852 19552 86860 19616
rect 6684 18438 6726 18674
rect 6962 18438 7004 18674
rect 11144 18438 11186 18674
rect 11422 18438 11464 18674
rect 43744 18438 43786 18674
rect 44022 18438 44064 18674
rect 48544 18438 48586 18674
rect 48822 18438 48864 18674
rect 81144 18438 81186 18674
rect 81422 18438 81464 18674
rect 86540 18528 86860 19552
rect 86540 18464 86548 18528
rect 86612 18464 86628 18528
rect 86692 18464 86708 18528
rect 86772 18464 86788 18528
rect 86852 18464 86860 18528
rect 6684 17984 7004 18438
rect 86540 18014 86860 18464
rect 6684 17920 6692 17984
rect 6756 17920 6772 17984
rect 6836 17920 6852 17984
rect 6916 17920 6932 17984
rect 6996 17920 7004 17984
rect 6684 16896 7004 17920
rect 10484 17778 10526 18014
rect 10762 17778 10804 18014
rect 43084 17778 43126 18014
rect 43362 17778 43404 18014
rect 47884 17778 47926 18014
rect 48162 17778 48204 18014
rect 80484 17778 80526 18014
rect 80762 17778 80804 18014
rect 86540 17778 86582 18014
rect 86818 17778 86860 18014
rect 6684 16832 6692 16896
rect 6756 16832 6772 16896
rect 6836 16832 6852 16896
rect 6916 16832 6932 16896
rect 6996 16832 7004 16896
rect 6684 15808 7004 16832
rect 6684 15744 6692 15808
rect 6756 15744 6772 15808
rect 6836 15744 6852 15808
rect 6916 15744 6932 15808
rect 6996 15744 7004 15808
rect 6684 14720 7004 15744
rect 6684 14656 6692 14720
rect 6756 14656 6772 14720
rect 6836 14656 6852 14720
rect 6916 14656 6932 14720
rect 6996 14656 7004 14720
rect 6684 13632 7004 14656
rect 6684 13568 6692 13632
rect 6756 13568 6772 13632
rect 6836 13568 6852 13632
rect 6916 13568 6932 13632
rect 6996 13568 7004 13632
rect 6684 12544 7004 13568
rect 6684 12480 6692 12544
rect 6756 12480 6772 12544
rect 6836 12480 6852 12544
rect 6916 12480 6932 12544
rect 6996 12480 7004 12544
rect 6684 11456 7004 12480
rect 86540 17440 86860 17778
rect 86540 17376 86548 17440
rect 86612 17376 86628 17440
rect 86692 17376 86708 17440
rect 86772 17376 86788 17440
rect 86852 17376 86860 17440
rect 86540 16352 86860 17376
rect 86540 16288 86548 16352
rect 86612 16288 86628 16352
rect 86692 16288 86708 16352
rect 86772 16288 86788 16352
rect 86852 16288 86860 16352
rect 86540 15264 86860 16288
rect 86540 15200 86548 15264
rect 86612 15200 86628 15264
rect 86692 15200 86708 15264
rect 86772 15200 86788 15264
rect 86852 15200 86860 15264
rect 86540 14176 86860 15200
rect 86540 14112 86548 14176
rect 86612 14112 86628 14176
rect 86692 14112 86708 14176
rect 86772 14112 86788 14176
rect 86852 14112 86860 14176
rect 86540 13088 86860 14112
rect 86540 13024 86548 13088
rect 86612 13024 86628 13088
rect 86692 13024 86708 13088
rect 86772 13024 86788 13088
rect 86852 13024 86860 13088
rect 86540 12000 86860 13024
rect 86540 11936 86548 12000
rect 86612 11936 86628 12000
rect 86692 11936 86708 12000
rect 86772 11936 86788 12000
rect 86852 11936 86860 12000
rect 11144 11630 11186 11866
rect 11422 11630 11464 11866
rect 43744 11630 43786 11866
rect 44022 11630 44064 11866
rect 48544 11630 48586 11866
rect 48822 11630 48864 11866
rect 81144 11630 81186 11866
rect 81422 11630 81464 11866
rect 6684 11392 6692 11456
rect 6756 11392 6772 11456
rect 6836 11392 6852 11456
rect 6916 11392 6932 11456
rect 6996 11392 7004 11456
rect 6684 10368 7004 11392
rect 10484 10970 10526 11206
rect 10762 10970 10804 11206
rect 43084 10970 43126 11206
rect 43362 10970 43404 11206
rect 47884 10970 47926 11206
rect 48162 10970 48204 11206
rect 80484 10970 80526 11206
rect 80762 10970 80804 11206
rect 6684 10304 6692 10368
rect 6756 10304 6772 10368
rect 6836 10304 6852 10368
rect 6916 10304 6932 10368
rect 6996 10304 7004 10368
rect 6684 9280 7004 10304
rect 86540 10912 86860 11936
rect 86540 10848 86548 10912
rect 86612 10848 86628 10912
rect 86692 10848 86708 10912
rect 86772 10848 86788 10912
rect 86852 10848 86860 10912
rect 6684 9216 6692 9280
rect 6756 9216 6772 9280
rect 6836 9216 6852 9280
rect 6916 9216 6932 9280
rect 6996 9216 7004 9280
rect 6684 8192 7004 9216
rect 6684 8128 6692 8192
rect 6756 8128 6772 8192
rect 6836 8128 6852 8192
rect 6916 8128 6932 8192
rect 6996 8128 7004 8192
rect 6684 7104 7004 8128
rect 6684 7040 6692 7104
rect 6756 7040 6772 7104
rect 6836 7040 6852 7104
rect 6916 7040 6932 7104
rect 6996 7040 7004 7104
rect 6684 7024 7004 7040
rect 17716 7648 18036 10187
rect 17716 7584 17724 7648
rect 17788 7584 17804 7648
rect 17868 7584 17884 7648
rect 17948 7584 17964 7648
rect 18028 7584 18036 7648
rect 3356 3418 3398 3654
rect 3634 3418 3676 3654
rect 3356 3376 3676 3418
rect 17716 6560 18036 7584
rect 17716 6496 17724 6560
rect 17788 6496 17804 6560
rect 17868 6496 17884 6560
rect 17948 6496 17964 6560
rect 18028 6496 18036 6560
rect 17716 5472 18036 6496
rect 17716 5408 17724 5472
rect 17788 5408 17804 5472
rect 17868 5408 17884 5472
rect 17948 5408 17964 5472
rect 18028 5408 18036 5472
rect 17716 3654 18036 5408
rect 17716 3418 17758 3654
rect 17994 3418 18036 3654
rect 2696 2758 2738 2994
rect 2974 2758 3016 2994
rect 2696 2716 3016 2758
rect 17716 2716 18036 3418
rect 18376 7104 18696 10187
rect 18376 7040 18384 7104
rect 18448 7040 18464 7104
rect 18528 7040 18544 7104
rect 18608 7040 18624 7104
rect 18688 7040 18696 7104
rect 18376 6016 18696 7040
rect 18376 5952 18384 6016
rect 18448 5952 18464 6016
rect 18528 5952 18544 6016
rect 18608 5952 18624 6016
rect 18688 5952 18696 6016
rect 18376 4928 18696 5952
rect 18376 4864 18384 4928
rect 18448 4864 18464 4928
rect 18528 4864 18544 4928
rect 18608 4864 18624 4928
rect 18688 4864 18696 4928
rect 18376 2994 18696 4864
rect 18376 2758 18418 2994
rect 18654 2758 18696 2994
rect 18376 2716 18696 2758
rect 36116 7648 36436 10187
rect 36116 7584 36124 7648
rect 36188 7584 36204 7648
rect 36268 7584 36284 7648
rect 36348 7584 36364 7648
rect 36428 7584 36436 7648
rect 36116 6560 36436 7584
rect 36116 6496 36124 6560
rect 36188 6496 36204 6560
rect 36268 6496 36284 6560
rect 36348 6496 36364 6560
rect 36428 6496 36436 6560
rect 36116 5472 36436 6496
rect 36116 5408 36124 5472
rect 36188 5408 36204 5472
rect 36268 5408 36284 5472
rect 36348 5408 36364 5472
rect 36428 5408 36436 5472
rect 36116 3654 36436 5408
rect 36116 3418 36158 3654
rect 36394 3418 36436 3654
rect 36116 2716 36436 3418
rect 36776 7104 37096 10187
rect 36776 7040 36784 7104
rect 36848 7040 36864 7104
rect 36928 7040 36944 7104
rect 37008 7040 37024 7104
rect 37088 7040 37096 7104
rect 36776 6016 37096 7040
rect 36776 5952 36784 6016
rect 36848 5952 36864 6016
rect 36928 5952 36944 6016
rect 37008 5952 37024 6016
rect 37088 5952 37096 6016
rect 36776 4928 37096 5952
rect 36776 4864 36784 4928
rect 36848 4864 36864 4928
rect 36928 4864 36944 4928
rect 37008 4864 37024 4928
rect 37088 4864 37096 4928
rect 36776 2994 37096 4864
rect 36776 2758 36818 2994
rect 37054 2758 37096 2994
rect 36776 2716 37096 2758
rect 54516 7648 54836 10187
rect 54516 7584 54524 7648
rect 54588 7584 54604 7648
rect 54668 7584 54684 7648
rect 54748 7584 54764 7648
rect 54828 7584 54836 7648
rect 54516 6560 54836 7584
rect 54516 6496 54524 6560
rect 54588 6496 54604 6560
rect 54668 6496 54684 6560
rect 54748 6496 54764 6560
rect 54828 6496 54836 6560
rect 54516 5472 54836 6496
rect 54516 5408 54524 5472
rect 54588 5408 54604 5472
rect 54668 5408 54684 5472
rect 54748 5408 54764 5472
rect 54828 5408 54836 5472
rect 54516 3654 54836 5408
rect 54516 3418 54558 3654
rect 54794 3418 54836 3654
rect 54516 2716 54836 3418
rect 55176 7104 55496 10187
rect 55176 7040 55184 7104
rect 55248 7040 55264 7104
rect 55328 7040 55344 7104
rect 55408 7040 55424 7104
rect 55488 7040 55496 7104
rect 55176 6016 55496 7040
rect 55176 5952 55184 6016
rect 55248 5952 55264 6016
rect 55328 5952 55344 6016
rect 55408 5952 55424 6016
rect 55488 5952 55496 6016
rect 55176 4928 55496 5952
rect 55176 4864 55184 4928
rect 55248 4864 55264 4928
rect 55328 4864 55344 4928
rect 55408 4864 55424 4928
rect 55488 4864 55496 4928
rect 55176 2994 55496 4864
rect 55176 2758 55218 2994
rect 55454 2758 55496 2994
rect 55176 2716 55496 2758
rect 72916 7648 73236 10187
rect 72916 7584 72924 7648
rect 72988 7584 73004 7648
rect 73068 7584 73084 7648
rect 73148 7584 73164 7648
rect 73228 7584 73236 7648
rect 72916 6560 73236 7584
rect 72916 6496 72924 6560
rect 72988 6496 73004 6560
rect 73068 6496 73084 6560
rect 73148 6496 73164 6560
rect 73228 6496 73236 6560
rect 72916 5472 73236 6496
rect 72916 5408 72924 5472
rect 72988 5408 73004 5472
rect 73068 5408 73084 5472
rect 73148 5408 73164 5472
rect 73228 5408 73236 5472
rect 72916 3654 73236 5408
rect 72916 3418 72958 3654
rect 73194 3418 73236 3654
rect 72916 2716 73236 3418
rect 73576 7104 73896 10187
rect 73576 7040 73584 7104
rect 73648 7040 73664 7104
rect 73728 7040 73744 7104
rect 73808 7040 73824 7104
rect 73888 7040 73896 7104
rect 73576 6016 73896 7040
rect 86540 9824 86860 10848
rect 86540 9760 86548 9824
rect 86612 9760 86628 9824
rect 86692 9760 86708 9824
rect 86772 9760 86788 9824
rect 86852 9760 86860 9824
rect 86540 8736 86860 9760
rect 86540 8672 86548 8736
rect 86612 8672 86628 8736
rect 86692 8672 86708 8736
rect 86772 8672 86788 8736
rect 86852 8672 86860 8736
rect 86540 7648 86860 8672
rect 86540 7584 86548 7648
rect 86612 7584 86628 7648
rect 86692 7584 86708 7648
rect 86772 7584 86788 7648
rect 86852 7584 86860 7648
rect 86540 7024 86860 7584
rect 87276 84352 87596 84912
rect 87276 84288 87284 84352
rect 87348 84288 87364 84352
rect 87428 84288 87444 84352
rect 87508 84288 87524 84352
rect 87588 84288 87596 84352
rect 87276 83264 87596 84288
rect 87276 83200 87284 83264
rect 87348 83200 87364 83264
rect 87428 83200 87444 83264
rect 87508 83200 87524 83264
rect 87588 83200 87596 83264
rect 87276 82176 87596 83200
rect 87276 82112 87284 82176
rect 87348 82112 87364 82176
rect 87428 82112 87444 82176
rect 87508 82112 87524 82176
rect 87588 82112 87596 82176
rect 87276 81088 87596 82112
rect 87276 81024 87284 81088
rect 87348 81024 87364 81088
rect 87428 81024 87444 81088
rect 87508 81024 87524 81088
rect 87588 81024 87596 81088
rect 87276 80000 87596 81024
rect 87276 79936 87284 80000
rect 87348 79936 87364 80000
rect 87428 79936 87444 80000
rect 87508 79936 87524 80000
rect 87588 79936 87596 80000
rect 87276 78912 87596 79936
rect 87276 78848 87284 78912
rect 87348 78848 87364 78912
rect 87428 78848 87444 78912
rect 87508 78848 87524 78912
rect 87588 78848 87596 78912
rect 87276 77824 87596 78848
rect 87276 77760 87284 77824
rect 87348 77760 87364 77824
rect 87428 77760 87444 77824
rect 87508 77760 87524 77824
rect 87588 77760 87596 77824
rect 87276 76736 87596 77760
rect 87276 76672 87284 76736
rect 87348 76672 87364 76736
rect 87428 76672 87444 76736
rect 87508 76672 87524 76736
rect 87588 76672 87596 76736
rect 87276 75648 87596 76672
rect 87276 75584 87284 75648
rect 87348 75584 87364 75648
rect 87428 75584 87444 75648
rect 87508 75584 87524 75648
rect 87588 75584 87596 75648
rect 87276 74560 87596 75584
rect 87276 74496 87284 74560
rect 87348 74496 87364 74560
rect 87428 74496 87444 74560
rect 87508 74496 87524 74560
rect 87588 74496 87596 74560
rect 87276 73874 87596 74496
rect 87276 73638 87318 73874
rect 87554 73638 87596 73874
rect 87276 73472 87596 73638
rect 87276 73408 87284 73472
rect 87348 73408 87364 73472
rect 87428 73408 87444 73472
rect 87508 73408 87524 73472
rect 87588 73408 87596 73472
rect 87276 72384 87596 73408
rect 87276 72320 87284 72384
rect 87348 72320 87364 72384
rect 87428 72320 87444 72384
rect 87508 72320 87524 72384
rect 87588 72320 87596 72384
rect 87276 71296 87596 72320
rect 87276 71232 87284 71296
rect 87348 71232 87364 71296
rect 87428 71232 87444 71296
rect 87508 71232 87524 71296
rect 87588 71232 87596 71296
rect 87276 70208 87596 71232
rect 87276 70144 87284 70208
rect 87348 70144 87364 70208
rect 87428 70144 87444 70208
rect 87508 70144 87524 70208
rect 87588 70144 87596 70208
rect 87276 69120 87596 70144
rect 87276 69056 87284 69120
rect 87348 69056 87364 69120
rect 87428 69056 87444 69120
rect 87508 69056 87524 69120
rect 87588 69056 87596 69120
rect 87276 68032 87596 69056
rect 87276 67968 87284 68032
rect 87348 67968 87364 68032
rect 87428 67968 87444 68032
rect 87508 67968 87524 68032
rect 87588 67968 87596 68032
rect 87276 66944 87596 67968
rect 87276 66880 87284 66944
rect 87348 66880 87364 66944
rect 87428 66880 87444 66944
rect 87508 66880 87524 66944
rect 87588 66880 87596 66944
rect 87276 65856 87596 66880
rect 87276 65792 87284 65856
rect 87348 65792 87364 65856
rect 87428 65792 87444 65856
rect 87508 65792 87524 65856
rect 87588 65792 87596 65856
rect 87276 64768 87596 65792
rect 87276 64704 87284 64768
rect 87348 64704 87364 64768
rect 87428 64704 87444 64768
rect 87508 64704 87524 64768
rect 87588 64704 87596 64768
rect 87276 63680 87596 64704
rect 87276 63616 87284 63680
rect 87348 63616 87364 63680
rect 87428 63616 87444 63680
rect 87508 63616 87524 63680
rect 87588 63616 87596 63680
rect 87276 62592 87596 63616
rect 87276 62528 87284 62592
rect 87348 62528 87364 62592
rect 87428 62528 87444 62592
rect 87508 62528 87524 62592
rect 87588 62528 87596 62592
rect 87276 61504 87596 62528
rect 87276 61440 87284 61504
rect 87348 61440 87364 61504
rect 87428 61440 87444 61504
rect 87508 61440 87524 61504
rect 87588 61440 87596 61504
rect 87276 60416 87596 61440
rect 87276 60352 87284 60416
rect 87348 60352 87364 60416
rect 87428 60352 87444 60416
rect 87508 60352 87524 60416
rect 87588 60352 87596 60416
rect 87276 59328 87596 60352
rect 87276 59264 87284 59328
rect 87348 59264 87364 59328
rect 87428 59264 87444 59328
rect 87508 59264 87524 59328
rect 87588 59264 87596 59328
rect 87276 58240 87596 59264
rect 87276 58176 87284 58240
rect 87348 58176 87364 58240
rect 87428 58176 87444 58240
rect 87508 58176 87524 58240
rect 87588 58176 87596 58240
rect 87276 57152 87596 58176
rect 87276 57088 87284 57152
rect 87348 57088 87364 57152
rect 87428 57088 87444 57152
rect 87508 57088 87524 57152
rect 87588 57088 87596 57152
rect 87276 56064 87596 57088
rect 87276 56000 87284 56064
rect 87348 56000 87364 56064
rect 87428 56000 87444 56064
rect 87508 56000 87524 56064
rect 87588 56000 87596 56064
rect 87276 55474 87596 56000
rect 87276 55238 87318 55474
rect 87554 55238 87596 55474
rect 87276 54976 87596 55238
rect 87276 54912 87284 54976
rect 87348 54912 87364 54976
rect 87428 54912 87444 54976
rect 87508 54912 87524 54976
rect 87588 54912 87596 54976
rect 87276 53888 87596 54912
rect 87276 53824 87284 53888
rect 87348 53824 87364 53888
rect 87428 53824 87444 53888
rect 87508 53824 87524 53888
rect 87588 53824 87596 53888
rect 87276 52800 87596 53824
rect 87276 52736 87284 52800
rect 87348 52736 87364 52800
rect 87428 52736 87444 52800
rect 87508 52736 87524 52800
rect 87588 52736 87596 52800
rect 87276 51712 87596 52736
rect 87276 51648 87284 51712
rect 87348 51648 87364 51712
rect 87428 51648 87444 51712
rect 87508 51648 87524 51712
rect 87588 51648 87596 51712
rect 87276 50624 87596 51648
rect 87276 50560 87284 50624
rect 87348 50560 87364 50624
rect 87428 50560 87444 50624
rect 87508 50560 87524 50624
rect 87588 50560 87596 50624
rect 87276 49536 87596 50560
rect 87276 49472 87284 49536
rect 87348 49472 87364 49536
rect 87428 49472 87444 49536
rect 87508 49472 87524 49536
rect 87588 49472 87596 49536
rect 87276 48448 87596 49472
rect 87276 48384 87284 48448
rect 87348 48384 87364 48448
rect 87428 48384 87444 48448
rect 87508 48384 87524 48448
rect 87588 48384 87596 48448
rect 87276 47360 87596 48384
rect 87276 47296 87284 47360
rect 87348 47296 87364 47360
rect 87428 47296 87444 47360
rect 87508 47296 87524 47360
rect 87588 47296 87596 47360
rect 87276 46272 87596 47296
rect 87276 46208 87284 46272
rect 87348 46208 87364 46272
rect 87428 46208 87444 46272
rect 87508 46208 87524 46272
rect 87588 46208 87596 46272
rect 87276 45184 87596 46208
rect 87276 45120 87284 45184
rect 87348 45120 87364 45184
rect 87428 45120 87444 45184
rect 87508 45120 87524 45184
rect 87588 45120 87596 45184
rect 87276 44096 87596 45120
rect 87276 44032 87284 44096
rect 87348 44032 87364 44096
rect 87428 44032 87444 44096
rect 87508 44032 87524 44096
rect 87588 44032 87596 44096
rect 87276 43008 87596 44032
rect 87276 42944 87284 43008
rect 87348 42944 87364 43008
rect 87428 42944 87444 43008
rect 87508 42944 87524 43008
rect 87588 42944 87596 43008
rect 87276 41920 87596 42944
rect 87276 41856 87284 41920
rect 87348 41856 87364 41920
rect 87428 41856 87444 41920
rect 87508 41856 87524 41920
rect 87588 41856 87596 41920
rect 87276 40832 87596 41856
rect 87276 40768 87284 40832
rect 87348 40768 87364 40832
rect 87428 40768 87444 40832
rect 87508 40768 87524 40832
rect 87588 40768 87596 40832
rect 87276 39744 87596 40768
rect 87276 39680 87284 39744
rect 87348 39680 87364 39744
rect 87428 39680 87444 39744
rect 87508 39680 87524 39744
rect 87588 39680 87596 39744
rect 87276 38656 87596 39680
rect 87276 38592 87284 38656
rect 87348 38592 87364 38656
rect 87428 38592 87444 38656
rect 87508 38592 87524 38656
rect 87588 38592 87596 38656
rect 87276 37568 87596 38592
rect 87276 37504 87284 37568
rect 87348 37504 87364 37568
rect 87428 37504 87444 37568
rect 87508 37504 87524 37568
rect 87588 37504 87596 37568
rect 87276 37074 87596 37504
rect 87276 36838 87318 37074
rect 87554 36838 87596 37074
rect 87276 36480 87596 36838
rect 87276 36416 87284 36480
rect 87348 36416 87364 36480
rect 87428 36416 87444 36480
rect 87508 36416 87524 36480
rect 87588 36416 87596 36480
rect 87276 35392 87596 36416
rect 87276 35328 87284 35392
rect 87348 35328 87364 35392
rect 87428 35328 87444 35392
rect 87508 35328 87524 35392
rect 87588 35328 87596 35392
rect 87276 34304 87596 35328
rect 87276 34240 87284 34304
rect 87348 34240 87364 34304
rect 87428 34240 87444 34304
rect 87508 34240 87524 34304
rect 87588 34240 87596 34304
rect 87276 33216 87596 34240
rect 87276 33152 87284 33216
rect 87348 33152 87364 33216
rect 87428 33152 87444 33216
rect 87508 33152 87524 33216
rect 87588 33152 87596 33216
rect 87276 32128 87596 33152
rect 87276 32064 87284 32128
rect 87348 32064 87364 32128
rect 87428 32064 87444 32128
rect 87508 32064 87524 32128
rect 87588 32064 87596 32128
rect 87276 31040 87596 32064
rect 87276 30976 87284 31040
rect 87348 30976 87364 31040
rect 87428 30976 87444 31040
rect 87508 30976 87524 31040
rect 87588 30976 87596 31040
rect 87276 29952 87596 30976
rect 87276 29888 87284 29952
rect 87348 29888 87364 29952
rect 87428 29888 87444 29952
rect 87508 29888 87524 29952
rect 87588 29888 87596 29952
rect 87276 28864 87596 29888
rect 87276 28800 87284 28864
rect 87348 28800 87364 28864
rect 87428 28800 87444 28864
rect 87508 28800 87524 28864
rect 87588 28800 87596 28864
rect 87276 27776 87596 28800
rect 87276 27712 87284 27776
rect 87348 27712 87364 27776
rect 87428 27712 87444 27776
rect 87508 27712 87524 27776
rect 87588 27712 87596 27776
rect 87276 26688 87596 27712
rect 87276 26624 87284 26688
rect 87348 26624 87364 26688
rect 87428 26624 87444 26688
rect 87508 26624 87524 26688
rect 87588 26624 87596 26688
rect 87276 25600 87596 26624
rect 87276 25536 87284 25600
rect 87348 25536 87364 25600
rect 87428 25536 87444 25600
rect 87508 25536 87524 25600
rect 87588 25536 87596 25600
rect 87276 24512 87596 25536
rect 87276 24448 87284 24512
rect 87348 24448 87364 24512
rect 87428 24448 87444 24512
rect 87508 24448 87524 24512
rect 87588 24448 87596 24512
rect 87276 23424 87596 24448
rect 87276 23360 87284 23424
rect 87348 23360 87364 23424
rect 87428 23360 87444 23424
rect 87508 23360 87524 23424
rect 87588 23360 87596 23424
rect 87276 22336 87596 23360
rect 87276 22272 87284 22336
rect 87348 22272 87364 22336
rect 87428 22272 87444 22336
rect 87508 22272 87524 22336
rect 87588 22272 87596 22336
rect 87276 21248 87596 22272
rect 87276 21184 87284 21248
rect 87348 21184 87364 21248
rect 87428 21184 87444 21248
rect 87508 21184 87524 21248
rect 87588 21184 87596 21248
rect 87276 20160 87596 21184
rect 87276 20096 87284 20160
rect 87348 20096 87364 20160
rect 87428 20096 87444 20160
rect 87508 20096 87524 20160
rect 87588 20096 87596 20160
rect 87276 19072 87596 20096
rect 87276 19008 87284 19072
rect 87348 19008 87364 19072
rect 87428 19008 87444 19072
rect 87508 19008 87524 19072
rect 87588 19008 87596 19072
rect 87276 18674 87596 19008
rect 87276 18438 87318 18674
rect 87554 18438 87596 18674
rect 87276 17984 87596 18438
rect 87276 17920 87284 17984
rect 87348 17920 87364 17984
rect 87428 17920 87444 17984
rect 87508 17920 87524 17984
rect 87588 17920 87596 17984
rect 87276 16896 87596 17920
rect 87276 16832 87284 16896
rect 87348 16832 87364 16896
rect 87428 16832 87444 16896
rect 87508 16832 87524 16896
rect 87588 16832 87596 16896
rect 87276 15808 87596 16832
rect 87276 15744 87284 15808
rect 87348 15744 87364 15808
rect 87428 15744 87444 15808
rect 87508 15744 87524 15808
rect 87588 15744 87596 15808
rect 87276 14720 87596 15744
rect 87276 14656 87284 14720
rect 87348 14656 87364 14720
rect 87428 14656 87444 14720
rect 87508 14656 87524 14720
rect 87588 14656 87596 14720
rect 87276 13632 87596 14656
rect 87276 13568 87284 13632
rect 87348 13568 87364 13632
rect 87428 13568 87444 13632
rect 87508 13568 87524 13632
rect 87588 13568 87596 13632
rect 87276 12544 87596 13568
rect 87276 12480 87284 12544
rect 87348 12480 87364 12544
rect 87428 12480 87444 12544
rect 87508 12480 87524 12544
rect 87588 12480 87596 12544
rect 87276 11456 87596 12480
rect 87276 11392 87284 11456
rect 87348 11392 87364 11456
rect 87428 11392 87444 11456
rect 87508 11392 87524 11456
rect 87588 11392 87596 11456
rect 87276 10368 87596 11392
rect 87276 10304 87284 10368
rect 87348 10304 87364 10368
rect 87428 10304 87444 10368
rect 87508 10304 87524 10368
rect 87588 10304 87596 10368
rect 87276 9280 87596 10304
rect 87276 9216 87284 9280
rect 87348 9216 87364 9280
rect 87428 9216 87444 9280
rect 87508 9216 87524 9280
rect 87588 9216 87596 9280
rect 87276 8192 87596 9216
rect 87276 8128 87284 8192
rect 87348 8128 87364 8192
rect 87428 8128 87444 8192
rect 87508 8128 87524 8192
rect 87588 8128 87596 8192
rect 87276 7104 87596 8128
rect 87276 7040 87284 7104
rect 87348 7040 87364 7104
rect 87428 7040 87444 7104
rect 87508 7040 87524 7104
rect 87588 7040 87596 7104
rect 87276 7024 87596 7040
rect 89796 73214 90116 88826
rect 89796 72978 89838 73214
rect 90074 72978 90116 73214
rect 89796 54814 90116 72978
rect 89796 54578 89838 54814
rect 90074 54578 90116 54814
rect 89796 36414 90116 54578
rect 89796 36178 89838 36414
rect 90074 36178 90116 36414
rect 89796 18014 90116 36178
rect 89796 17778 89838 18014
rect 90074 17778 90116 18014
rect 73576 5952 73584 6016
rect 73648 5952 73664 6016
rect 73728 5952 73744 6016
rect 73808 5952 73824 6016
rect 73888 5952 73896 6016
rect 73576 4928 73896 5952
rect 73576 4864 73584 4928
rect 73648 4864 73664 4928
rect 73728 4864 73744 4928
rect 73808 4864 73824 4928
rect 73888 4864 73896 4928
rect 73576 2994 73896 4864
rect 89796 3654 90116 17778
rect 89796 3418 89838 3654
rect 90074 3418 90116 3654
rect 89796 3376 90116 3418
rect 90456 73874 90776 89486
rect 90456 73638 90498 73874
rect 90734 73638 90776 73874
rect 90456 55474 90776 73638
rect 90456 55238 90498 55474
rect 90734 55238 90776 55474
rect 90456 37074 90776 55238
rect 90456 36838 90498 37074
rect 90734 36838 90776 37074
rect 90456 18674 90776 36838
rect 90456 18438 90498 18674
rect 90734 18438 90776 18674
rect 73576 2758 73618 2994
rect 73854 2758 73896 2994
rect 73576 2716 73896 2758
rect 90456 2994 90776 18438
rect 90456 2758 90498 2994
rect 90734 2758 90776 2994
rect 90456 2716 90776 2758
<< via4 >>
rect 2738 89486 2974 89722
rect 2738 73638 2974 73874
rect 2738 55238 2974 55474
rect 2738 36838 2974 37074
rect 2738 18438 2974 18674
rect 3398 88826 3634 89062
rect 17758 88826 17994 89062
rect 3398 72978 3634 73214
rect 3398 54578 3634 54814
rect 3398 36178 3634 36414
rect 3398 17778 3634 18014
rect 5990 72978 6226 73214
rect 5990 54578 6226 54814
rect 5990 36178 6226 36414
rect 5990 17778 6226 18014
rect 18418 89486 18654 89722
rect 36158 88826 36394 89062
rect 36818 89486 37054 89722
rect 54558 88826 54794 89062
rect 55218 89486 55454 89722
rect 72958 88826 73194 89062
rect 73618 89486 73854 89722
rect 90498 89486 90734 89722
rect 89838 88826 90074 89062
rect 11186 80630 11422 80866
rect 43786 80630 44022 80866
rect 48586 80630 48822 80866
rect 81186 80630 81422 80866
rect 10526 79970 10762 80206
rect 43126 79970 43362 80206
rect 47926 79970 48162 80206
rect 80526 79970 80762 80206
rect 6726 73638 6962 73874
rect 11186 73638 11422 73874
rect 43786 73638 44022 73874
rect 48586 73638 48822 73874
rect 81186 73638 81422 73874
rect 10526 72978 10762 73214
rect 43126 72978 43362 73214
rect 47926 72978 48162 73214
rect 80526 72978 80762 73214
rect 86582 72978 86818 73214
rect 6726 55238 6962 55474
rect 11186 55238 11422 55474
rect 43786 55238 44022 55474
rect 48586 55238 48822 55474
rect 81186 55238 81422 55474
rect 10526 54578 10762 54814
rect 43126 54578 43362 54814
rect 47926 54578 48162 54814
rect 80526 54578 80762 54814
rect 86582 54578 86818 54814
rect 11186 48030 11422 48266
rect 43786 48030 44022 48266
rect 48586 48030 48822 48266
rect 81186 48030 81422 48266
rect 10526 47370 10762 47606
rect 43126 47370 43362 47606
rect 47926 47370 48162 47606
rect 80526 47370 80762 47606
rect 11186 44230 11422 44466
rect 43786 44230 44022 44466
rect 48586 44230 48822 44466
rect 81186 44230 81422 44466
rect 10526 43570 10762 43806
rect 43126 43570 43362 43806
rect 47926 43570 48162 43806
rect 80526 43570 80762 43806
rect 6726 36838 6962 37074
rect 11186 36838 11422 37074
rect 43786 36838 44022 37074
rect 48586 36838 48822 37074
rect 81186 36838 81422 37074
rect 10526 36178 10762 36414
rect 43126 36178 43362 36414
rect 47926 36178 48162 36414
rect 80526 36178 80762 36414
rect 86582 36178 86818 36414
rect 6726 18438 6962 18674
rect 11186 18438 11422 18674
rect 43786 18438 44022 18674
rect 48586 18438 48822 18674
rect 81186 18438 81422 18674
rect 10526 17778 10762 18014
rect 43126 17778 43362 18014
rect 47926 17778 48162 18014
rect 80526 17778 80762 18014
rect 86582 17778 86818 18014
rect 11186 11630 11422 11866
rect 43786 11630 44022 11866
rect 48586 11630 48822 11866
rect 81186 11630 81422 11866
rect 10526 10970 10762 11206
rect 43126 10970 43362 11206
rect 47926 10970 48162 11206
rect 80526 10970 80762 11206
rect 3398 3418 3634 3654
rect 17758 3418 17994 3654
rect 2738 2758 2974 2994
rect 18418 2758 18654 2994
rect 36158 3418 36394 3654
rect 36818 2758 37054 2994
rect 54558 3418 54794 3654
rect 55218 2758 55454 2994
rect 72958 3418 73194 3654
rect 87318 73638 87554 73874
rect 87318 55238 87554 55474
rect 87318 36838 87554 37074
rect 87318 18438 87554 18674
rect 89838 72978 90074 73214
rect 89838 54578 90074 54814
rect 89838 36178 90074 36414
rect 89838 17778 90074 18014
rect 89838 3418 90074 3654
rect 90498 73638 90734 73874
rect 90498 55238 90734 55474
rect 90498 36838 90734 37074
rect 90498 18438 90734 18674
rect 73618 2758 73854 2994
rect 90498 2758 90734 2994
<< metal5 >>
rect 2696 89722 90776 89764
rect 2696 89486 2738 89722
rect 2974 89486 18418 89722
rect 18654 89486 36818 89722
rect 37054 89486 55218 89722
rect 55454 89486 73618 89722
rect 73854 89486 90498 89722
rect 90734 89486 90776 89722
rect 2696 89444 90776 89486
rect 3356 89062 90116 89104
rect 3356 88826 3398 89062
rect 3634 88826 17758 89062
rect 17994 88826 36158 89062
rect 36394 88826 54558 89062
rect 54794 88826 72958 89062
rect 73194 88826 89838 89062
rect 90074 88826 90116 89062
rect 3356 88784 90116 88826
rect 11162 80866 11446 80908
rect 11162 80630 11186 80866
rect 11422 80630 11446 80866
rect 11162 80588 11446 80630
rect 43762 80866 44046 80908
rect 43762 80630 43786 80866
rect 44022 80630 44046 80866
rect 43762 80588 44046 80630
rect 48562 80866 48846 80908
rect 48562 80630 48586 80866
rect 48822 80630 48846 80866
rect 48562 80588 48846 80630
rect 81162 80866 81446 80908
rect 81162 80630 81186 80866
rect 81422 80630 81446 80866
rect 81162 80588 81446 80630
rect 10502 80206 10786 80248
rect 10502 79970 10526 80206
rect 10762 79970 10786 80206
rect 10502 79928 10786 79970
rect 43102 80206 43386 80248
rect 43102 79970 43126 80206
rect 43362 79970 43386 80206
rect 43102 79928 43386 79970
rect 47902 80206 48186 80248
rect 47902 79970 47926 80206
rect 48162 79970 48186 80206
rect 47902 79928 48186 79970
rect 80502 80206 80786 80248
rect 80502 79970 80526 80206
rect 80762 79970 80786 80206
rect 80502 79928 80786 79970
rect 2696 73874 90776 73916
rect 2696 73638 2738 73874
rect 2974 73638 6726 73874
rect 6962 73638 11186 73874
rect 11422 73638 43786 73874
rect 44022 73638 48586 73874
rect 48822 73638 81186 73874
rect 81422 73638 87318 73874
rect 87554 73638 90498 73874
rect 90734 73638 90776 73874
rect 2696 73596 90776 73638
rect 2696 73214 90776 73256
rect 2696 72978 3398 73214
rect 3634 72978 5990 73214
rect 6226 72978 10526 73214
rect 10762 72978 43126 73214
rect 43362 72978 47926 73214
rect 48162 72978 80526 73214
rect 80762 72978 86582 73214
rect 86818 72978 89838 73214
rect 90074 72978 90776 73214
rect 2696 72936 90776 72978
rect 2696 55474 90776 55516
rect 2696 55238 2738 55474
rect 2974 55238 6726 55474
rect 6962 55238 11186 55474
rect 11422 55238 43786 55474
rect 44022 55238 48586 55474
rect 48822 55238 81186 55474
rect 81422 55238 87318 55474
rect 87554 55238 90498 55474
rect 90734 55238 90776 55474
rect 2696 55196 90776 55238
rect 2696 54814 90776 54856
rect 2696 54578 3398 54814
rect 3634 54578 5990 54814
rect 6226 54578 10526 54814
rect 10762 54578 43126 54814
rect 43362 54578 47926 54814
rect 48162 54578 80526 54814
rect 80762 54578 86582 54814
rect 86818 54578 89838 54814
rect 90074 54578 90776 54814
rect 2696 54536 90776 54578
rect 11162 48266 11446 48308
rect 11162 48030 11186 48266
rect 11422 48030 11446 48266
rect 11162 47988 11446 48030
rect 43762 48266 44046 48308
rect 43762 48030 43786 48266
rect 44022 48030 44046 48266
rect 43762 47988 44046 48030
rect 48562 48266 48846 48308
rect 48562 48030 48586 48266
rect 48822 48030 48846 48266
rect 48562 47988 48846 48030
rect 81162 48266 81446 48308
rect 81162 48030 81186 48266
rect 81422 48030 81446 48266
rect 81162 47988 81446 48030
rect 10502 47606 10786 47648
rect 10502 47370 10526 47606
rect 10762 47370 10786 47606
rect 10502 47328 10786 47370
rect 43102 47606 43386 47648
rect 43102 47370 43126 47606
rect 43362 47370 43386 47606
rect 43102 47328 43386 47370
rect 47902 47606 48186 47648
rect 47902 47370 47926 47606
rect 48162 47370 48186 47606
rect 47902 47328 48186 47370
rect 80502 47606 80786 47648
rect 80502 47370 80526 47606
rect 80762 47370 80786 47606
rect 80502 47328 80786 47370
rect 11162 44466 11446 44508
rect 11162 44230 11186 44466
rect 11422 44230 11446 44466
rect 11162 44188 11446 44230
rect 43762 44466 44046 44508
rect 43762 44230 43786 44466
rect 44022 44230 44046 44466
rect 43762 44188 44046 44230
rect 48562 44466 48846 44508
rect 48562 44230 48586 44466
rect 48822 44230 48846 44466
rect 48562 44188 48846 44230
rect 81162 44466 81446 44508
rect 81162 44230 81186 44466
rect 81422 44230 81446 44466
rect 81162 44188 81446 44230
rect 10502 43806 10786 43848
rect 10502 43570 10526 43806
rect 10762 43570 10786 43806
rect 10502 43528 10786 43570
rect 43102 43806 43386 43848
rect 43102 43570 43126 43806
rect 43362 43570 43386 43806
rect 43102 43528 43386 43570
rect 47902 43806 48186 43848
rect 47902 43570 47926 43806
rect 48162 43570 48186 43806
rect 47902 43528 48186 43570
rect 80502 43806 80786 43848
rect 80502 43570 80526 43806
rect 80762 43570 80786 43806
rect 80502 43528 80786 43570
rect 2696 37074 90776 37116
rect 2696 36838 2738 37074
rect 2974 36838 6726 37074
rect 6962 36838 11186 37074
rect 11422 36838 43786 37074
rect 44022 36838 48586 37074
rect 48822 36838 81186 37074
rect 81422 36838 87318 37074
rect 87554 36838 90498 37074
rect 90734 36838 90776 37074
rect 2696 36796 90776 36838
rect 2696 36414 90776 36456
rect 2696 36178 3398 36414
rect 3634 36178 5990 36414
rect 6226 36178 10526 36414
rect 10762 36178 43126 36414
rect 43362 36178 47926 36414
rect 48162 36178 80526 36414
rect 80762 36178 86582 36414
rect 86818 36178 89838 36414
rect 90074 36178 90776 36414
rect 2696 36136 90776 36178
rect 2696 18674 90776 18716
rect 2696 18438 2738 18674
rect 2974 18438 6726 18674
rect 6962 18438 11186 18674
rect 11422 18438 43786 18674
rect 44022 18438 48586 18674
rect 48822 18438 81186 18674
rect 81422 18438 87318 18674
rect 87554 18438 90498 18674
rect 90734 18438 90776 18674
rect 2696 18396 90776 18438
rect 2696 18014 90776 18056
rect 2696 17778 3398 18014
rect 3634 17778 5990 18014
rect 6226 17778 10526 18014
rect 10762 17778 43126 18014
rect 43362 17778 47926 18014
rect 48162 17778 80526 18014
rect 80762 17778 86582 18014
rect 86818 17778 89838 18014
rect 90074 17778 90776 18014
rect 2696 17736 90776 17778
rect 11162 11866 11446 11908
rect 11162 11630 11186 11866
rect 11422 11630 11446 11866
rect 11162 11588 11446 11630
rect 43762 11866 44046 11908
rect 43762 11630 43786 11866
rect 44022 11630 44046 11866
rect 43762 11588 44046 11630
rect 48562 11866 48846 11908
rect 48562 11630 48586 11866
rect 48822 11630 48846 11866
rect 48562 11588 48846 11630
rect 81162 11866 81446 11908
rect 81162 11630 81186 11866
rect 81422 11630 81446 11866
rect 81162 11588 81446 11630
rect 10502 11206 10786 11248
rect 10502 10970 10526 11206
rect 10762 10970 10786 11206
rect 10502 10928 10786 10970
rect 43102 11206 43386 11248
rect 43102 10970 43126 11206
rect 43362 10970 43386 11206
rect 43102 10928 43386 10970
rect 47902 11206 48186 11248
rect 47902 10970 47926 11206
rect 48162 10970 48186 11206
rect 47902 10928 48186 10970
rect 80502 11206 80786 11248
rect 80502 10970 80526 11206
rect 80762 10970 80786 11206
rect 80502 10928 80786 10970
rect 3356 3654 90116 3696
rect 3356 3418 3398 3654
rect 3634 3418 17758 3654
rect 17994 3418 36158 3654
rect 36394 3418 54558 3654
rect 54794 3418 72958 3654
rect 73194 3418 89838 3654
rect 90074 3418 90116 3654
rect 3356 3376 90116 3418
rect 2696 2994 90776 3036
rect 2696 2758 2738 2994
rect 2974 2758 18418 2994
rect 18654 2758 36818 2994
rect 37054 2758 55218 2994
rect 55454 2758 73618 2994
rect 73854 2758 90498 2994
rect 90734 2758 90776 2994
rect 2696 2716 90776 2758
use sky130_fd_sc_hd__diode_2  ANTENNA_cell0_clk
timestamp 18001
transform 1 0 7268 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell0_config_data_out
timestamp 18001
transform -1 0 45540 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell0_config_en
timestamp 18001
transform -1 0 7268 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell0_le_clk
timestamp 18001
transform -1 0 45724 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell0_le_en
timestamp 18001
transform -1 0 45908 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell0_le_nrst
timestamp 18001
transform -1 0 46092 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell0_nrst
timestamp 18001
transform -1 0 7636 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell1_clk
timestamp 18001
transform -1 0 85744 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell1_config_data_in
timestamp 18001
transform -1 0 85928 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell1_config_data_out
timestamp 18001
transform -1 0 85744 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell1_config_en
timestamp 18001
transform -1 0 86112 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell1_le_clk
timestamp 18001
transform 1 0 85560 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell1_le_en
timestamp 18001
transform 1 0 85560 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell1_le_nrst
timestamp 18001
transform 1 0 85560 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell1_nrst
timestamp 18001
transform -1 0 86296 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell2_clk
timestamp 18001
transform -1 0 10764 0 1 84320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell2_config_data_in
timestamp 18001
transform -1 0 14076 0 1 84320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell2_config_data_out
timestamp 18001
transform -1 0 45540 0 1 84320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell2_config_en
timestamp 18001
transform 1 0 12788 0 1 84320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell2_le_clk
timestamp 18001
transform -1 0 45724 0 1 84320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell2_le_en
timestamp 18001
transform -1 0 45908 0 1 84320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell2_le_nrst
timestamp 18001
transform -1 0 46092 0 1 84320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell2_nrst
timestamp 18001
transform 1 0 11684 0 1 84320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell3_clk
timestamp 18001
transform -1 0 48208 0 1 84320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell3_config_data_in
timestamp 18001
transform -1 0 51520 0 1 84320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell3_config_en
timestamp 18001
transform 1 0 50232 0 1 84320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell3_le_clk
timestamp 18001
transform 1 0 85560 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell3_le_en
timestamp 18001
transform 1 0 85560 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell3_le_nrst
timestamp 18001
transform 1 0 85560 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cell3_nrst
timestamp 18001
transform 1 0 49128 0 1 84320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 18001
transform 1 0 31004 0 1 84320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_X
timestamp 18001
transform -1 0 31004 0 1 84320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0__f_clk_A
timestamp 18001
transform 1 0 7452 0 -1 64736
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0__f_clk_X
timestamp 18001
transform 1 0 7452 0 -1 63648
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1__f_clk_A
timestamp 18001
transform -1 0 40940 0 1 84320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1__f_clk_X
timestamp 18001
transform -1 0 43056 0 1 84320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 18001
transform -1 0 5612 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 18001
transform -1 0 37996 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_X
timestamp 18001
transform 1 0 39836 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 18001
transform -1 0 88044 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 18001
transform -1 0 88044 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 18001
transform -1 0 88044 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 18001
transform -1 0 87860 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 18001
transform -1 0 88044 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 18001
transform -1 0 87860 0 1 66912
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 18001
transform -1 0 88044 0 -1 68000
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 18001
transform -1 0 87860 0 1 69088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 18001
transform -1 0 87860 0 1 70176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 18001
transform -1 0 88044 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 18001
transform -1 0 87860 0 1 71264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 18001
transform -1 0 87860 0 1 72352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 18001
transform -1 0 88044 0 -1 73440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 18001
transform -1 0 87860 0 1 74528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 18001
transform -1 0 87860 0 1 75616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 18001
transform -1 0 88136 0 1 76704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 18001
transform -1 0 87860 0 1 77792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 18001
transform -1 0 88044 0 -1 78880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 18001
transform -1 0 87860 0 1 79968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 18001
transform -1 0 87860 0 1 81056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 18001
transform -1 0 87860 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 18001
transform -1 0 88044 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 18001
transform -1 0 88044 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 18001
transform -1 0 88044 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 18001
transform -1 0 88044 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 18001
transform -1 0 87860 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 18001
transform -1 0 87952 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 18001
transform -1 0 88320 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 18001
transform -1 0 15180 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 18001
transform -1 0 26128 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 18001
transform -1 0 27416 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 18001
transform -1 0 28612 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 18001
transform -1 0 29348 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 18001
transform -1 0 52532 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 18001
transform -1 0 54372 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 18001
transform -1 0 54924 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 18001
transform -1 0 55752 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 18001
transform -1 0 16652 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 18001
transform -1 0 57040 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 18001
transform -1 0 57684 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 18001
transform -1 0 59524 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 18001
transform -1 0 60260 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 18001
transform -1 0 62100 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 18001
transform -1 0 62652 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 18001
transform -1 0 63480 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 18001
transform -1 0 64768 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 18001
transform -1 0 65412 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 18001
transform -1 0 67252 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 18001
transform -1 0 17112 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 18001
transform -1 0 18400 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 18001
transform -1 0 19688 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 18001
transform -1 0 20884 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 18001
transform -1 0 21620 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 18001
transform -1 0 22908 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 18001
transform -1 0 23552 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 18001
transform -1 0 24840 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 18001
transform -1 0 30636 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 18001
transform -1 0 41584 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 18001
transform -1 0 42872 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 18001
transform -1 0 44068 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 18001
transform -1 0 44804 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 18001
transform -1 0 67988 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 18001
transform -1 0 69828 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 18001
transform -1 0 70380 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 18001
transform -1 0 71208 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 18001
transform -1 0 31280 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 18001
transform -1 0 72496 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 18001
transform -1 0 73140 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 18001
transform -1 0 74980 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 18001
transform -1 0 75716 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 18001
transform -1 0 77556 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 18001
transform -1 0 78108 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 18001
transform -1 0 78936 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 18001
transform -1 0 80224 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input77_A
timestamp 18001
transform -1 0 88044 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input78_A
timestamp 18001
transform -1 0 87860 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 18001
transform -1 0 32568 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 18001
transform -1 0 33856 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input81_A
timestamp 18001
transform -1 0 35144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input82_A
timestamp 18001
transform -1 0 36340 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input83_A
timestamp 18001
transform -1 0 37076 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input84_A
timestamp 18001
transform -1 0 38364 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input85_A
timestamp 18001
transform -1 0 39008 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input86_A
timestamp 18001
transform -1 0 40296 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input87_A
timestamp 18001
transform -1 0 5612 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input88_A
timestamp 18001
transform -1 0 5612 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input89_A
timestamp 18001
transform -1 0 5612 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input90_A
timestamp 18001
transform -1 0 5612 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input91_A
timestamp 18001
transform -1 0 5612 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input92_A
timestamp 18001
transform -1 0 5612 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input93_A
timestamp 18001
transform -1 0 5612 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input94_A
timestamp 18001
transform -1 0 5612 0 1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input95_A
timestamp 18001
transform -1 0 5612 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input96_A
timestamp 18001
transform -1 0 5612 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input97_A
timestamp 18001
transform -1 0 5612 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input98_A
timestamp 18001
transform -1 0 5612 0 -1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input99_A
timestamp 18001
transform -1 0 5612 0 1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input100_A
timestamp 18001
transform -1 0 5612 0 1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input101_A
timestamp 18001
transform -1 0 5612 0 1 60384
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input102_A
timestamp 18001
transform -1 0 5612 0 1 61472
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input103_A
timestamp 18001
transform -1 0 5612 0 -1 62560
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input104_A
timestamp 18001
transform -1 0 5612 0 1 63648
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input105_A
timestamp 18001
transform -1 0 5612 0 1 64736
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input106_A
timestamp 18001
transform -1 0 5612 0 1 65824
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input107_A
timestamp 18001
transform -1 0 5612 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input108_A
timestamp 18001
transform -1 0 5612 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input109_A
timestamp 18001
transform -1 0 5612 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input110_A
timestamp 18001
transform -1 0 5612 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input111_A
timestamp 18001
transform -1 0 5612 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input112_A
timestamp 18001
transform -1 0 5612 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input113_A
timestamp 18001
transform -1 0 5612 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input114_A
timestamp 18001
transform -1 0 5612 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input115_A
timestamp 18001
transform -1 0 88136 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input115_X
timestamp 18001
transform -1 0 88228 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input116_A
timestamp 18001
transform -1 0 87768 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input116_X
timestamp 18001
transform -1 0 88320 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input117_A
timestamp 18001
transform -1 0 88136 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input117_X
timestamp 18001
transform -1 0 88320 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input118_A
timestamp 18001
transform -1 0 40940 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input118_X
timestamp 18001
transform 1 0 42044 0 -1 87584
box -38 -48 222 592
use fpgacell  cell0
timestamp 0
transform 1 0 10000 0 1 10000
box 0 0 35800 35800
use fpgacell  cell1
timestamp 0
transform 1 0 47400 0 1 10000
box 0 0 35800 35800
use fpgacell  cell2
timestamp 0
transform 1 0 10000 0 1 46400
box 0 0 35800 35800
use fpgacell  cell3
timestamp 0
transform 1 0 47400 0 1 46400
box 0 0 35800 35800
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 18001
transform -1 0 30636 0 1 84320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 18001
transform -1 0 7452 0 1 63648
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 18001
transform 1 0 41032 0 1 84320
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3
timestamp 1636986456
transform 1 0 5152 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1636986456
transform 1 0 6256 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp 18001
transform 1 0 7360 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1636986456
transform 1 0 7544 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1636986456
transform 1 0 8648 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp 18001
transform 1 0 9752 0 1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1636986456
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1636986456
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 18001
transform 1 0 12328 0 1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1636986456
transform 1 0 12696 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1636986456
transform 1 0 13800 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 18001
transform 1 0 14904 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_117
timestamp 18001
transform 1 0 15640 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_123
timestamp 18001
transform 1 0 16192 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_131
timestamp 18001
transform 1 0 16928 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 18001
transform 1 0 17480 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_141
timestamp 18001
transform 1 0 17848 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_151
timestamp 18001
transform 1 0 18768 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_159
timestamp 18001
transform 1 0 19504 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 18001
transform 1 0 20056 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_173
timestamp 18001
transform 1 0 20792 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_181
timestamp 18001
transform 1 0 21528 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_186
timestamp 18001
transform 1 0 21988 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 18001
transform 1 0 22724 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_201
timestamp 18001
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_207
timestamp 18001
transform 1 0 23920 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_215
timestamp 18001
transform 1 0 24656 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 18001
transform 1 0 25208 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_225
timestamp 18001
transform 1 0 25576 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_235
timestamp 18001
transform 1 0 26496 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_243
timestamp 18001
transform 1 0 27232 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 18001
transform 1 0 27784 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_257
timestamp 18001
transform 1 0 28520 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_265
timestamp 18001
transform 1 0 29256 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_270
timestamp 18001
transform 1 0 29716 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_284
timestamp 18001
transform 1 0 31004 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_290
timestamp 18001
transform 1 0 31556 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_298
timestamp 18001
transform 1 0 32292 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_304
timestamp 18001
transform 1 0 32844 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_309
timestamp 18001
transform 1 0 33304 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_318
timestamp 18001
transform 1 0 34132 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_326
timestamp 18001
transform 1 0 34868 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_332
timestamp 18001
transform 1 0 35420 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_342
timestamp 18001
transform 1 0 36340 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_353
timestamp 18001
transform 1 0 37352 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_361
timestamp 18001
transform 1 0 38088 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_368
timestamp 18001
transform 1 0 38732 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_374
timestamp 18001
transform 1 0 39284 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_382
timestamp 18001
transform 1 0 40020 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_388
timestamp 18001
transform 1 0 40572 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_393
timestamp 18001
transform 1 0 41032 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_402
timestamp 18001
transform 1 0 41860 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_410
timestamp 18001
transform 1 0 42596 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_416
timestamp 18001
transform 1 0 43148 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_426
timestamp 18001
transform 1 0 44068 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_437
timestamp 18001
transform 1 0 45080 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_445
timestamp 18001
transform 1 0 45816 0 1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_449
timestamp 1636986456
transform 1 0 46184 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_461
timestamp 1636986456
transform 1 0 47288 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_473
timestamp 18001
transform 1 0 48392 0 1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_477
timestamp 1636986456
transform 1 0 48760 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_489
timestamp 1636986456
transform 1 0 49864 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_501
timestamp 18001
transform 1 0 50968 0 1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_505
timestamp 1636986456
transform 1 0 51336 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_517
timestamp 18001
transform 1 0 52440 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_522
timestamp 18001
transform 1 0 52900 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_530
timestamp 18001
transform 1 0 53636 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_537
timestamp 18001
transform 1 0 54280 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_543
timestamp 18001
transform 1 0 54832 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_551
timestamp 18001
transform 1 0 55568 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_557
timestamp 18001
transform 1 0 56120 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_561
timestamp 18001
transform 1 0 56488 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_571
timestamp 18001
transform 1 0 57408 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_578
timestamp 18001
transform 1 0 58052 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_586
timestamp 18001
transform 1 0 58788 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_593
timestamp 18001
transform 1 0 59432 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_601
timestamp 18001
transform 1 0 60168 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_606
timestamp 18001
transform 1 0 60628 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_614
timestamp 18001
transform 1 0 61364 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_621
timestamp 18001
transform 1 0 62008 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_627
timestamp 18001
transform 1 0 62560 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_635
timestamp 18001
transform 1 0 63296 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_641
timestamp 18001
transform 1 0 63848 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_645
timestamp 18001
transform 1 0 64216 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_655
timestamp 18001
transform 1 0 65136 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_662
timestamp 18001
transform 1 0 65780 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_670
timestamp 18001
transform 1 0 66516 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_677
timestamp 18001
transform 1 0 67160 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_683
timestamp 18001
transform 1 0 67712 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_689
timestamp 18001
transform 1 0 68264 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_697
timestamp 18001
transform 1 0 69000 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_706
timestamp 18001
transform 1 0 69828 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_712
timestamp 18001
transform 1 0 70380 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_718
timestamp 18001
transform 1 0 70932 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_724
timestamp 18001
transform 1 0 71484 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_729
timestamp 18001
transform 1 0 71944 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_738
timestamp 18001
transform 1 0 72772 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_745
timestamp 18001
transform 1 0 73416 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_753
timestamp 18001
transform 1 0 74152 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_762
timestamp 18001
transform 1 0 74980 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_773
timestamp 18001
transform 1 0 75992 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_781
timestamp 18001
transform 1 0 76728 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_790
timestamp 18001
transform 1 0 77556 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_796
timestamp 18001
transform 1 0 78108 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_802
timestamp 18001
transform 1 0 78660 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_808
timestamp 18001
transform 1 0 79212 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_813
timestamp 18001
transform 1 0 79672 0 1 4896
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_822
timestamp 1636986456
transform 1 0 80500 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_834
timestamp 18001
transform 1 0 81604 0 1 4896
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_841
timestamp 1636986456
transform 1 0 82248 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_853
timestamp 1636986456
transform 1 0 83352 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_865
timestamp 18001
transform 1 0 84456 0 1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_869
timestamp 1636986456
transform 1 0 84824 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_881
timestamp 1636986456
transform 1 0 85928 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_893
timestamp 18001
transform 1 0 87032 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_897
timestamp 18001
transform 1 0 87400 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_905
timestamp 18001
transform 1 0 88136 0 1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1636986456
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1636986456
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1636986456
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1636986456
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 18001
transform 1 0 9568 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 18001
transform 1 0 9936 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1636986456
transform 1 0 10120 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1636986456
transform 1 0 11224 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1636986456
transform 1 0 12328 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1636986456
transform 1 0 13432 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 18001
transform 1 0 14536 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 18001
transform 1 0 15088 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1636986456
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1636986456
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1636986456
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1636986456
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 18001
transform 1 0 19688 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 18001
transform 1 0 20240 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1636986456
transform 1 0 20424 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1636986456
transform 1 0 21528 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1636986456
transform 1 0 22632 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1636986456
transform 1 0 23736 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 18001
transform 1 0 24840 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 18001
transform 1 0 25392 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1636986456
transform 1 0 25576 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1636986456
transform 1 0 26680 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1636986456
transform 1 0 27784 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1636986456
transform 1 0 28888 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 18001
transform 1 0 29992 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 18001
transform 1 0 30544 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1636986456
transform 1 0 30728 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1636986456
transform 1 0 31832 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1636986456
transform 1 0 32936 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1636986456
transform 1 0 34040 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 18001
transform 1 0 35144 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 18001
transform 1 0 35696 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1636986456
transform 1 0 35880 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1636986456
transform 1 0 36984 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1636986456
transform 1 0 38088 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1636986456
transform 1 0 39192 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 18001
transform 1 0 40296 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 18001
transform 1 0 40848 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1636986456
transform 1 0 41032 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_405
timestamp 1636986456
transform 1 0 42136 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_417
timestamp 1636986456
transform 1 0 43240 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_429
timestamp 1636986456
transform 1 0 44344 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 18001
transform 1 0 45448 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 18001
transform 1 0 46000 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_449
timestamp 1636986456
transform 1 0 46184 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_461
timestamp 1636986456
transform 1 0 47288 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_473
timestamp 1636986456
transform 1 0 48392 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_485
timestamp 1636986456
transform 1 0 49496 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_497
timestamp 18001
transform 1 0 50600 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 18001
transform 1 0 51152 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_505
timestamp 1636986456
transform 1 0 51336 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_517
timestamp 1636986456
transform 1 0 52440 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_529
timestamp 1636986456
transform 1 0 53544 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_541
timestamp 1636986456
transform 1 0 54648 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_553
timestamp 18001
transform 1 0 55752 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_559
timestamp 18001
transform 1 0 56304 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_561
timestamp 1636986456
transform 1 0 56488 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_573
timestamp 1636986456
transform 1 0 57592 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_585
timestamp 1636986456
transform 1 0 58696 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_597
timestamp 1636986456
transform 1 0 59800 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_609
timestamp 18001
transform 1 0 60904 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_615
timestamp 18001
transform 1 0 61456 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_617
timestamp 1636986456
transform 1 0 61640 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_629
timestamp 1636986456
transform 1 0 62744 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_641
timestamp 1636986456
transform 1 0 63848 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_653
timestamp 1636986456
transform 1 0 64952 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_665
timestamp 18001
transform 1 0 66056 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_671
timestamp 18001
transform 1 0 66608 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_673
timestamp 1636986456
transform 1 0 66792 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_685
timestamp 1636986456
transform 1 0 67896 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_697
timestamp 1636986456
transform 1 0 69000 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_709
timestamp 1636986456
transform 1 0 70104 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_721
timestamp 18001
transform 1 0 71208 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_727
timestamp 18001
transform 1 0 71760 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_729
timestamp 1636986456
transform 1 0 71944 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_741
timestamp 1636986456
transform 1 0 73048 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_753
timestamp 1636986456
transform 1 0 74152 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_765
timestamp 1636986456
transform 1 0 75256 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_777
timestamp 18001
transform 1 0 76360 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_783
timestamp 18001
transform 1 0 76912 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_785
timestamp 1636986456
transform 1 0 77096 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_797
timestamp 1636986456
transform 1 0 78200 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_809
timestamp 1636986456
transform 1 0 79304 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_821
timestamp 1636986456
transform 1 0 80408 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_833
timestamp 18001
transform 1 0 81512 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_839
timestamp 18001
transform 1 0 82064 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_841
timestamp 1636986456
transform 1 0 82248 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_853
timestamp 1636986456
transform 1 0 83352 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_865
timestamp 1636986456
transform 1 0 84456 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_877
timestamp 1636986456
transform 1 0 85560 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_889
timestamp 18001
transform 1 0 86664 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_895
timestamp 18001
transform 1 0 87216 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_897
timestamp 18001
transform 1 0 87400 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_905
timestamp 18001
transform 1 0 88136 0 -1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1636986456
transform 1 0 5152 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1636986456
transform 1 0 6256 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 18001
transform 1 0 7360 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1636986456
transform 1 0 7544 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1636986456
transform 1 0 8648 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1636986456
transform 1 0 9752 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1636986456
transform 1 0 10856 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 18001
transform 1 0 11960 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 18001
transform 1 0 12512 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1636986456
transform 1 0 12696 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1636986456
transform 1 0 13800 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1636986456
transform 1 0 14904 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1636986456
transform 1 0 16008 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 18001
transform 1 0 17112 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 18001
transform 1 0 17664 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1636986456
transform 1 0 17848 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1636986456
transform 1 0 18952 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1636986456
transform 1 0 20056 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1636986456
transform 1 0 21160 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 18001
transform 1 0 22264 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 18001
transform 1 0 22816 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1636986456
transform 1 0 23000 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1636986456
transform 1 0 24104 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1636986456
transform 1 0 25208 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1636986456
transform 1 0 26312 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 18001
transform 1 0 27416 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 18001
transform 1 0 27968 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1636986456
transform 1 0 28152 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1636986456
transform 1 0 29256 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1636986456
transform 1 0 30360 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1636986456
transform 1 0 31464 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 18001
transform 1 0 32568 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 18001
transform 1 0 33120 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1636986456
transform 1 0 33304 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1636986456
transform 1 0 34408 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1636986456
transform 1 0 35512 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1636986456
transform 1 0 36616 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 18001
transform 1 0 37720 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 18001
transform 1 0 38272 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1636986456
transform 1 0 38456 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1636986456
transform 1 0 39560 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1636986456
transform 1 0 40664 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1636986456
transform 1 0 41768 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 18001
transform 1 0 42872 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 18001
transform 1 0 43424 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1636986456
transform 1 0 43608 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1636986456
transform 1 0 44712 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 1636986456
transform 1 0 45816 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_457
timestamp 1636986456
transform 1 0 46920 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 18001
transform 1 0 48024 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 18001
transform 1 0 48576 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_477
timestamp 1636986456
transform 1 0 48760 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_489
timestamp 1636986456
transform 1 0 49864 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_501
timestamp 1636986456
transform 1 0 50968 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_513
timestamp 1636986456
transform 1 0 52072 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_525
timestamp 18001
transform 1 0 53176 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 18001
transform 1 0 53728 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_533
timestamp 1636986456
transform 1 0 53912 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_545
timestamp 1636986456
transform 1 0 55016 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_557
timestamp 1636986456
transform 1 0 56120 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_569
timestamp 1636986456
transform 1 0 57224 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_581
timestamp 18001
transform 1 0 58328 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 18001
transform 1 0 58880 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_589
timestamp 1636986456
transform 1 0 59064 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_601
timestamp 1636986456
transform 1 0 60168 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_613
timestamp 1636986456
transform 1 0 61272 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_625
timestamp 1636986456
transform 1 0 62376 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_637
timestamp 18001
transform 1 0 63480 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_643
timestamp 18001
transform 1 0 64032 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_645
timestamp 1636986456
transform 1 0 64216 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_657
timestamp 1636986456
transform 1 0 65320 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_669
timestamp 1636986456
transform 1 0 66424 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_681
timestamp 1636986456
transform 1 0 67528 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_693
timestamp 18001
transform 1 0 68632 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_699
timestamp 18001
transform 1 0 69184 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_701
timestamp 1636986456
transform 1 0 69368 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_713
timestamp 1636986456
transform 1 0 70472 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_725
timestamp 1636986456
transform 1 0 71576 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_737
timestamp 1636986456
transform 1 0 72680 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_749
timestamp 18001
transform 1 0 73784 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_755
timestamp 18001
transform 1 0 74336 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_757
timestamp 1636986456
transform 1 0 74520 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_769
timestamp 1636986456
transform 1 0 75624 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_781
timestamp 1636986456
transform 1 0 76728 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_793
timestamp 1636986456
transform 1 0 77832 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_805
timestamp 18001
transform 1 0 78936 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_811
timestamp 18001
transform 1 0 79488 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_813
timestamp 1636986456
transform 1 0 79672 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_825
timestamp 1636986456
transform 1 0 80776 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_837
timestamp 1636986456
transform 1 0 81880 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_849
timestamp 1636986456
transform 1 0 82984 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_861
timestamp 18001
transform 1 0 84088 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_867
timestamp 18001
transform 1 0 84640 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_869
timestamp 1636986456
transform 1 0 84824 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_881
timestamp 1636986456
transform 1 0 85928 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_893
timestamp 1636986456
transform 1 0 87032 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_905
timestamp 18001
transform 1 0 88136 0 1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1636986456
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1636986456
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1636986456
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1636986456
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 18001
transform 1 0 9568 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 18001
transform 1 0 9936 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1636986456
transform 1 0 10120 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1636986456
transform 1 0 11224 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1636986456
transform 1 0 12328 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1636986456
transform 1 0 13432 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 18001
transform 1 0 14536 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 18001
transform 1 0 15088 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1636986456
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1636986456
transform 1 0 16376 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1636986456
transform 1 0 17480 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1636986456
transform 1 0 18584 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 18001
transform 1 0 19688 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 18001
transform 1 0 20240 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1636986456
transform 1 0 20424 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1636986456
transform 1 0 21528 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1636986456
transform 1 0 22632 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1636986456
transform 1 0 23736 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 18001
transform 1 0 24840 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 18001
transform 1 0 25392 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1636986456
transform 1 0 25576 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1636986456
transform 1 0 26680 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1636986456
transform 1 0 27784 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1636986456
transform 1 0 28888 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 18001
transform 1 0 29992 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 18001
transform 1 0 30544 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1636986456
transform 1 0 30728 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1636986456
transform 1 0 31832 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1636986456
transform 1 0 32936 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1636986456
transform 1 0 34040 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 18001
transform 1 0 35144 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 18001
transform 1 0 35696 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1636986456
transform 1 0 35880 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1636986456
transform 1 0 36984 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1636986456
transform 1 0 38088 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1636986456
transform 1 0 39192 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 18001
transform 1 0 40296 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 18001
transform 1 0 40848 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1636986456
transform 1 0 41032 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1636986456
transform 1 0 42136 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1636986456
transform 1 0 43240 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1636986456
transform 1 0 44344 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 18001
transform 1 0 45448 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 18001
transform 1 0 46000 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1636986456
transform 1 0 46184 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1636986456
transform 1 0 47288 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1636986456
transform 1 0 48392 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1636986456
transform 1 0 49496 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 18001
transform 1 0 50600 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 18001
transform 1 0 51152 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_505
timestamp 1636986456
transform 1 0 51336 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_517
timestamp 1636986456
transform 1 0 52440 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_529
timestamp 1636986456
transform 1 0 53544 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_541
timestamp 1636986456
transform 1 0 54648 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_553
timestamp 18001
transform 1 0 55752 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 18001
transform 1 0 56304 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_561
timestamp 1636986456
transform 1 0 56488 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_573
timestamp 1636986456
transform 1 0 57592 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_585
timestamp 1636986456
transform 1 0 58696 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_597
timestamp 1636986456
transform 1 0 59800 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_609
timestamp 18001
transform 1 0 60904 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 18001
transform 1 0 61456 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_617
timestamp 1636986456
transform 1 0 61640 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_629
timestamp 1636986456
transform 1 0 62744 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_641
timestamp 1636986456
transform 1 0 63848 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_653
timestamp 1636986456
transform 1 0 64952 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_665
timestamp 18001
transform 1 0 66056 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_671
timestamp 18001
transform 1 0 66608 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_673
timestamp 1636986456
transform 1 0 66792 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_685
timestamp 1636986456
transform 1 0 67896 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_697
timestamp 1636986456
transform 1 0 69000 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_709
timestamp 1636986456
transform 1 0 70104 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_721
timestamp 18001
transform 1 0 71208 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_727
timestamp 18001
transform 1 0 71760 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_729
timestamp 1636986456
transform 1 0 71944 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_741
timestamp 1636986456
transform 1 0 73048 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_753
timestamp 1636986456
transform 1 0 74152 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_765
timestamp 1636986456
transform 1 0 75256 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_777
timestamp 18001
transform 1 0 76360 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_783
timestamp 18001
transform 1 0 76912 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_785
timestamp 1636986456
transform 1 0 77096 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_797
timestamp 1636986456
transform 1 0 78200 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_809
timestamp 1636986456
transform 1 0 79304 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_821
timestamp 1636986456
transform 1 0 80408 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_833
timestamp 18001
transform 1 0 81512 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_839
timestamp 18001
transform 1 0 82064 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_841
timestamp 1636986456
transform 1 0 82248 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_853
timestamp 1636986456
transform 1 0 83352 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_865
timestamp 1636986456
transform 1 0 84456 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_877
timestamp 1636986456
transform 1 0 85560 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_889
timestamp 18001
transform 1 0 86664 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_895
timestamp 18001
transform 1 0 87216 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_897
timestamp 18001
transform 1 0 87400 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_905
timestamp 18001
transform 1 0 88136 0 -1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1636986456
transform 1 0 5152 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1636986456
transform 1 0 6256 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 18001
transform 1 0 7360 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1636986456
transform 1 0 7544 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1636986456
transform 1 0 8648 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_53
timestamp 18001
transform 1 0 9752 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_57
timestamp 1636986456
transform 1 0 10120 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_69
timestamp 1636986456
transform 1 0 11224 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_81
timestamp 18001
transform 1 0 12328 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1636986456
transform 1 0 12696 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1636986456
transform 1 0 13800 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_109
timestamp 18001
transform 1 0 14904 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_113
timestamp 1636986456
transform 1 0 15272 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_125
timestamp 1636986456
transform 1 0 16376 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_137
timestamp 18001
transform 1 0 17480 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1636986456
transform 1 0 17848 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1636986456
transform 1 0 18952 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_165
timestamp 18001
transform 1 0 20056 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_169
timestamp 1636986456
transform 1 0 20424 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_181
timestamp 1636986456
transform 1 0 21528 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_193
timestamp 18001
transform 1 0 22632 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1636986456
transform 1 0 23000 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1636986456
transform 1 0 24104 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_221
timestamp 18001
transform 1 0 25208 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_225
timestamp 1636986456
transform 1 0 25576 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_237
timestamp 1636986456
transform 1 0 26680 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_249
timestamp 18001
transform 1 0 27784 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1636986456
transform 1 0 28152 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1636986456
transform 1 0 29256 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_277
timestamp 18001
transform 1 0 30360 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_281
timestamp 1636986456
transform 1 0 30728 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_293
timestamp 1636986456
transform 1 0 31832 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_305
timestamp 18001
transform 1 0 32936 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1636986456
transform 1 0 33304 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1636986456
transform 1 0 34408 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_333
timestamp 18001
transform 1 0 35512 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_337
timestamp 1636986456
transform 1 0 35880 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_349
timestamp 1636986456
transform 1 0 36984 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_361
timestamp 18001
transform 1 0 38088 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1636986456
transform 1 0 38456 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1636986456
transform 1 0 39560 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_389
timestamp 18001
transform 1 0 40664 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_393
timestamp 1636986456
transform 1 0 41032 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_405
timestamp 1636986456
transform 1 0 42136 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_417
timestamp 18001
transform 1 0 43240 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1636986456
transform 1 0 43608 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_433
timestamp 18001
transform 1 0 44712 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_439
timestamp 18001
transform 1 0 45264 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_449
timestamp 1636986456
transform 1 0 46184 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_461
timestamp 1636986456
transform 1 0 47288 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_473
timestamp 18001
transform 1 0 48392 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1636986456
transform 1 0 48760 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1636986456
transform 1 0 49864 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_501
timestamp 18001
transform 1 0 50968 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_505
timestamp 1636986456
transform 1 0 51336 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_517
timestamp 1636986456
transform 1 0 52440 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_529
timestamp 18001
transform 1 0 53544 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_533
timestamp 1636986456
transform 1 0 53912 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_545
timestamp 1636986456
transform 1 0 55016 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_557
timestamp 18001
transform 1 0 56120 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_561
timestamp 1636986456
transform 1 0 56488 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_573
timestamp 1636986456
transform 1 0 57592 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_585
timestamp 18001
transform 1 0 58696 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_589
timestamp 1636986456
transform 1 0 59064 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_601
timestamp 1636986456
transform 1 0 60168 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_613
timestamp 18001
transform 1 0 61272 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_617
timestamp 1636986456
transform 1 0 61640 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_629
timestamp 1636986456
transform 1 0 62744 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_641
timestamp 18001
transform 1 0 63848 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_645
timestamp 1636986456
transform 1 0 64216 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_657
timestamp 1636986456
transform 1 0 65320 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_669
timestamp 18001
transform 1 0 66424 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_673
timestamp 1636986456
transform 1 0 66792 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_685
timestamp 1636986456
transform 1 0 67896 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_697
timestamp 18001
transform 1 0 69000 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_701
timestamp 1636986456
transform 1 0 69368 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_713
timestamp 1636986456
transform 1 0 70472 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_725
timestamp 18001
transform 1 0 71576 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_729
timestamp 1636986456
transform 1 0 71944 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_741
timestamp 1636986456
transform 1 0 73048 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_753
timestamp 18001
transform 1 0 74152 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_757
timestamp 1636986456
transform 1 0 74520 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_769
timestamp 1636986456
transform 1 0 75624 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_781
timestamp 18001
transform 1 0 76728 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_785
timestamp 1636986456
transform 1 0 77096 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_797
timestamp 1636986456
transform 1 0 78200 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_809
timestamp 18001
transform 1 0 79304 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_813
timestamp 1636986456
transform 1 0 79672 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_825
timestamp 1636986456
transform 1 0 80776 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_837
timestamp 18001
transform 1 0 81880 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_841
timestamp 1636986456
transform 1 0 82248 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_853
timestamp 1636986456
transform 1 0 83352 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_865
timestamp 18001
transform 1 0 84456 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_869
timestamp 1636986456
transform 1 0 84824 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_881
timestamp 1636986456
transform 1 0 85928 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_893
timestamp 18001
transform 1 0 87032 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_897
timestamp 18001
transform 1 0 87400 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_905
timestamp 18001
transform 1 0 88136 0 1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1636986456
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1636986456
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_27
timestamp 18001
transform 1 0 7360 0 -1 8160
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_877
timestamp 1636986456
transform 1 0 85560 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_889
timestamp 1636986456
transform 1 0 86664 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_901
timestamp 18001
transform 1 0 87768 0 -1 8160
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1636986456
transform 1 0 5152 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1636986456
transform 1 0 6256 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 18001
transform 1 0 7360 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_29
timestamp 18001
transform 1 0 7544 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_877
timestamp 1636986456
transform 1 0 85560 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_889
timestamp 1636986456
transform 1 0 86664 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_901
timestamp 18001
transform 1 0 87768 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_903
timestamp 18001
transform 1 0 87952 0 1 8160
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1636986456
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1636986456
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_27
timestamp 18001
transform 1 0 7360 0 -1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_877
timestamp 1636986456
transform 1 0 85560 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_889
timestamp 1636986456
transform 1 0 86664 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_901
timestamp 18001
transform 1 0 87768 0 -1 9248
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1636986456
transform 1 0 5152 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1636986456
transform 1 0 6256 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 18001
transform 1 0 7360 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_29
timestamp 18001
transform 1 0 7544 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_877
timestamp 1636986456
transform 1 0 85560 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_889
timestamp 1636986456
transform 1 0 86664 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_901
timestamp 18001
transform 1 0 87768 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_903
timestamp 18001
transform 1 0 87952 0 1 9248
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1636986456
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1636986456
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_27
timestamp 18001
transform 1 0 7360 0 -1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_877
timestamp 1636986456
transform 1 0 85560 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_889
timestamp 1636986456
transform 1 0 86664 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_901
timestamp 18001
transform 1 0 87768 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1636986456
transform 1 0 5152 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1636986456
transform 1 0 6256 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 18001
transform 1 0 7360 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_29
timestamp 18001
transform 1 0 7544 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_877
timestamp 1636986456
transform 1 0 85560 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_889
timestamp 18001
transform 1 0 86664 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_897
timestamp 18001
transform 1 0 87400 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_903
timestamp 18001
transform 1 0 87952 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1636986456
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1636986456
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_27
timestamp 18001
transform 1 0 7360 0 -1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_879
timestamp 1636986456
transform 1 0 85744 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_891
timestamp 1636986456
transform 1 0 86848 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_903
timestamp 18001
transform 1 0 87952 0 -1 11424
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1636986456
transform 1 0 5152 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1636986456
transform 1 0 6256 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 18001
transform 1 0 7360 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_29
timestamp 18001
transform 1 0 7544 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_877
timestamp 1636986456
transform 1 0 85560 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_889
timestamp 1636986456
transform 1 0 86664 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_901
timestamp 18001
transform 1 0 87768 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_903
timestamp 18001
transform 1 0 87952 0 1 11424
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1636986456
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1636986456
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_27
timestamp 18001
transform 1 0 7360 0 -1 12512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_879
timestamp 1636986456
transform 1 0 85744 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_891
timestamp 1636986456
transform 1 0 86848 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_903
timestamp 18001
transform 1 0 87952 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_906
timestamp 18001
transform 1 0 88228 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1636986456
transform 1 0 5152 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1636986456
transform 1 0 6256 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 18001
transform 1 0 7360 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_29
timestamp 18001
transform 1 0 7544 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_877
timestamp 1636986456
transform 1 0 85560 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_889
timestamp 18001
transform 1 0 86664 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_895
timestamp 18001
transform 1 0 87216 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1636986456
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1636986456
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_27
timestamp 18001
transform 1 0 7360 0 -1 13600
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_879
timestamp 1636986456
transform 1 0 85744 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_891
timestamp 18001
transform 1 0 86848 0 -1 13600
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1636986456
transform 1 0 5152 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1636986456
transform 1 0 6256 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 18001
transform 1 0 7360 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_29
timestamp 18001
transform 1 0 7544 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_877
timestamp 1636986456
transform 1 0 85560 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_889
timestamp 1636986456
transform 1 0 86664 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_901
timestamp 18001
transform 1 0 87768 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_903
timestamp 18001
transform 1 0 87952 0 1 13600
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1636986456
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1636986456
transform 1 0 6256 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_27
timestamp 18001
transform 1 0 7360 0 -1 14688
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_879
timestamp 1636986456
transform 1 0 85744 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_891
timestamp 1636986456
transform 1 0 86848 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_903
timestamp 18001
transform 1 0 87952 0 -1 14688
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1636986456
transform 1 0 5152 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1636986456
transform 1 0 6256 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 18001
transform 1 0 7360 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_29
timestamp 18001
transform 1 0 7544 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_877
timestamp 1636986456
transform 1 0 85560 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_889
timestamp 18001
transform 1 0 86664 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_895
timestamp 18001
transform 1 0 87216 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_8
timestamp 1636986456
transform 1 0 5612 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_20
timestamp 18001
transform 1 0 6716 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_28
timestamp 18001
transform 1 0 7452 0 -1 15776
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_877
timestamp 1636986456
transform 1 0 85560 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_889
timestamp 1636986456
transform 1 0 86664 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_901
timestamp 18001
transform 1 0 87768 0 -1 15776
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1636986456
transform 1 0 5152 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1636986456
transform 1 0 6256 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 18001
transform 1 0 7360 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_29
timestamp 18001
transform 1 0 7544 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_877
timestamp 1636986456
transform 1 0 85560 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_889
timestamp 1636986456
transform 1 0 86664 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_901
timestamp 18001
transform 1 0 87768 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_903
timestamp 18001
transform 1 0 87952 0 1 15776
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1636986456
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1636986456
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_27
timestamp 18001
transform 1 0 7360 0 -1 16864
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_877
timestamp 1636986456
transform 1 0 85560 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_889
timestamp 1636986456
transform 1 0 86664 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_901
timestamp 18001
transform 1 0 87768 0 -1 16864
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_8
timestamp 1636986456
transform 1 0 5612 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_20
timestamp 18001
transform 1 0 6716 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_29
timestamp 18001
transform 1 0 7544 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_877
timestamp 1636986456
transform 1 0 85560 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_889
timestamp 1636986456
transform 1 0 86664 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_901
timestamp 18001
transform 1 0 87768 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_8
timestamp 1636986456
transform 1 0 5612 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_20
timestamp 18001
transform 1 0 6716 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_28
timestamp 18001
transform 1 0 7452 0 -1 17952
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_877
timestamp 1636986456
transform 1 0 85560 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_889
timestamp 1636986456
transform 1 0 86664 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_901
timestamp 18001
transform 1 0 87768 0 -1 17952
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1636986456
transform 1 0 5152 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1636986456
transform 1 0 6256 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 18001
transform 1 0 7360 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_29
timestamp 18001
transform 1 0 7544 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_877
timestamp 1636986456
transform 1 0 85560 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_889
timestamp 1636986456
transform 1 0 86664 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_901
timestamp 18001
transform 1 0 87768 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_903
timestamp 18001
transform 1 0 87952 0 1 17952
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_8
timestamp 1636986456
transform 1 0 5612 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_20
timestamp 18001
transform 1 0 6716 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_28
timestamp 18001
transform 1 0 7452 0 -1 19040
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_877
timestamp 1636986456
transform 1 0 85560 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_889
timestamp 1636986456
transform 1 0 86664 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_901
timestamp 18001
transform 1 0 87768 0 -1 19040
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1636986456
transform 1 0 5152 0 1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1636986456
transform 1 0 6256 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 18001
transform 1 0 7360 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_29
timestamp 18001
transform 1 0 7544 0 1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_877
timestamp 1636986456
transform 1 0 85560 0 1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_889
timestamp 1636986456
transform 1 0 86664 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_901
timestamp 18001
transform 1 0 87768 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_903
timestamp 18001
transform 1 0 87952 0 1 19040
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_8
timestamp 1636986456
transform 1 0 5612 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_20
timestamp 18001
transform 1 0 6716 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_28
timestamp 18001
transform 1 0 7452 0 -1 20128
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_877
timestamp 1636986456
transform 1 0 85560 0 -1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_889
timestamp 1636986456
transform 1 0 86664 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_901
timestamp 18001
transform 1 0 87768 0 -1 20128
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1636986456
transform 1 0 5152 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1636986456
transform 1 0 6256 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 18001
transform 1 0 7360 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_29
timestamp 18001
transform 1 0 7544 0 1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_877
timestamp 1636986456
transform 1 0 85560 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_889
timestamp 1636986456
transform 1 0 86664 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_901
timestamp 18001
transform 1 0 87768 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_903
timestamp 18001
transform 1 0 87952 0 1 20128
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_8
timestamp 1636986456
transform 1 0 5612 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_20
timestamp 18001
transform 1 0 6716 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_28
timestamp 18001
transform 1 0 7452 0 -1 21216
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_877
timestamp 1636986456
transform 1 0 85560 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_889
timestamp 1636986456
transform 1 0 86664 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_901
timestamp 18001
transform 1 0 87768 0 -1 21216
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1636986456
transform 1 0 5152 0 1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1636986456
transform 1 0 6256 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 18001
transform 1 0 7360 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_29
timestamp 18001
transform 1 0 7544 0 1 21216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_877
timestamp 1636986456
transform 1 0 85560 0 1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_889
timestamp 1636986456
transform 1 0 86664 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_901
timestamp 18001
transform 1 0 87768 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_903
timestamp 18001
transform 1 0 87952 0 1 21216
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1636986456
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1636986456
transform 1 0 6256 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_27
timestamp 18001
transform 1 0 7360 0 -1 22304
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_877
timestamp 1636986456
transform 1 0 85560 0 -1 22304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_889
timestamp 1636986456
transform 1 0 86664 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_901
timestamp 18001
transform 1 0 87768 0 -1 22304
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_8
timestamp 1636986456
transform 1 0 5612 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_20
timestamp 18001
transform 1 0 6716 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_29
timestamp 18001
transform 1 0 7544 0 1 22304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_877
timestamp 1636986456
transform 1 0 85560 0 1 22304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_889
timestamp 1636986456
transform 1 0 86664 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_901
timestamp 18001
transform 1 0 87768 0 1 22304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_8
timestamp 1636986456
transform 1 0 5612 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_20
timestamp 18001
transform 1 0 6716 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_28
timestamp 18001
transform 1 0 7452 0 -1 23392
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_877
timestamp 1636986456
transform 1 0 85560 0 -1 23392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_889
timestamp 1636986456
transform 1 0 86664 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_901
timestamp 18001
transform 1 0 87768 0 -1 23392
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1636986456
transform 1 0 5152 0 1 23392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1636986456
transform 1 0 6256 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 18001
transform 1 0 7360 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_29
timestamp 18001
transform 1 0 7544 0 1 23392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_877
timestamp 1636986456
transform 1 0 85560 0 1 23392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_889
timestamp 1636986456
transform 1 0 86664 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_901
timestamp 18001
transform 1 0 87768 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_903
timestamp 18001
transform 1 0 87952 0 1 23392
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_8
timestamp 1636986456
transform 1 0 5612 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_20
timestamp 18001
transform 1 0 6716 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_28
timestamp 18001
transform 1 0 7452 0 -1 24480
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_877
timestamp 1636986456
transform 1 0 85560 0 -1 24480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_889
timestamp 1636986456
transform 1 0 86664 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_901
timestamp 18001
transform 1 0 87768 0 -1 24480
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1636986456
transform 1 0 5152 0 1 24480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1636986456
transform 1 0 6256 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 18001
transform 1 0 7360 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_29
timestamp 18001
transform 1 0 7544 0 1 24480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_877
timestamp 1636986456
transform 1 0 85560 0 1 24480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_889
timestamp 1636986456
transform 1 0 86664 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_901
timestamp 18001
transform 1 0 87768 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_903
timestamp 18001
transform 1 0 87952 0 1 24480
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_8
timestamp 1636986456
transform 1 0 5612 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_20
timestamp 18001
transform 1 0 6716 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_28
timestamp 18001
transform 1 0 7452 0 -1 25568
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_877
timestamp 1636986456
transform 1 0 85560 0 -1 25568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_889
timestamp 1636986456
transform 1 0 86664 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_901
timestamp 18001
transform 1 0 87768 0 -1 25568
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1636986456
transform 1 0 5152 0 1 25568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1636986456
transform 1 0 6256 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 18001
transform 1 0 7360 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_29
timestamp 18001
transform 1 0 7544 0 1 25568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_877
timestamp 1636986456
transform 1 0 85560 0 1 25568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_889
timestamp 1636986456
transform 1 0 86664 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_901
timestamp 18001
transform 1 0 87768 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_903
timestamp 18001
transform 1 0 87952 0 1 25568
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_8
timestamp 1636986456
transform 1 0 5612 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_20
timestamp 18001
transform 1 0 6716 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_28
timestamp 18001
transform 1 0 7452 0 -1 26656
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_877
timestamp 1636986456
transform 1 0 85560 0 -1 26656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_889
timestamp 1636986456
transform 1 0 86664 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_901
timestamp 18001
transform 1 0 87768 0 -1 26656
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1636986456
transform 1 0 5152 0 1 26656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1636986456
transform 1 0 6256 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 18001
transform 1 0 7360 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_29
timestamp 18001
transform 1 0 7544 0 1 26656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_877
timestamp 1636986456
transform 1 0 85560 0 1 26656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_889
timestamp 1636986456
transform 1 0 86664 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_901
timestamp 18001
transform 1 0 87768 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_903
timestamp 18001
transform 1 0 87952 0 1 26656
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1636986456
transform 1 0 5152 0 -1 27744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1636986456
transform 1 0 6256 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_27
timestamp 18001
transform 1 0 7360 0 -1 27744
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_877
timestamp 1636986456
transform 1 0 85560 0 -1 27744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_889
timestamp 1636986456
transform 1 0 86664 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_901
timestamp 18001
transform 1 0 87768 0 -1 27744
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_8
timestamp 1636986456
transform 1 0 5612 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_20
timestamp 18001
transform 1 0 6716 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_29
timestamp 18001
transform 1 0 7544 0 1 27744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_877
timestamp 1636986456
transform 1 0 85560 0 1 27744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_889
timestamp 1636986456
transform 1 0 86664 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_901
timestamp 18001
transform 1 0 87768 0 1 27744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_8
timestamp 1636986456
transform 1 0 5612 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_20
timestamp 18001
transform 1 0 6716 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_28
timestamp 18001
transform 1 0 7452 0 -1 28832
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_877
timestamp 1636986456
transform 1 0 85560 0 -1 28832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_889
timestamp 1636986456
transform 1 0 86664 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_901
timestamp 18001
transform 1 0 87768 0 -1 28832
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1636986456
transform 1 0 5152 0 1 28832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1636986456
transform 1 0 6256 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 18001
transform 1 0 7360 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_44_29
timestamp 18001
transform 1 0 7544 0 1 28832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_877
timestamp 1636986456
transform 1 0 85560 0 1 28832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_889
timestamp 1636986456
transform 1 0 86664 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_901
timestamp 18001
transform 1 0 87768 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_903
timestamp 18001
transform 1 0 87952 0 1 28832
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_8
timestamp 1636986456
transform 1 0 5612 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_20
timestamp 18001
transform 1 0 6716 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_28
timestamp 18001
transform 1 0 7452 0 -1 29920
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_877
timestamp 1636986456
transform 1 0 85560 0 -1 29920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_889
timestamp 1636986456
transform 1 0 86664 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_901
timestamp 18001
transform 1 0 87768 0 -1 29920
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1636986456
transform 1 0 5152 0 1 29920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1636986456
transform 1 0 6256 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 18001
transform 1 0 7360 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_29
timestamp 18001
transform 1 0 7544 0 1 29920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_877
timestamp 1636986456
transform 1 0 85560 0 1 29920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_889
timestamp 1636986456
transform 1 0 86664 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_901
timestamp 18001
transform 1 0 87768 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_903
timestamp 18001
transform 1 0 87952 0 1 29920
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_7
timestamp 1636986456
transform 1 0 5520 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_19
timestamp 18001
transform 1 0 6624 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_27
timestamp 18001
transform 1 0 7360 0 -1 31008
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_877
timestamp 1636986456
transform 1 0 85560 0 -1 31008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_889
timestamp 1636986456
transform 1 0 86664 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_901
timestamp 18001
transform 1 0 87768 0 -1 31008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1636986456
transform 1 0 5152 0 1 31008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1636986456
transform 1 0 6256 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 18001
transform 1 0 7360 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_29
timestamp 18001
transform 1 0 7544 0 1 31008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_877
timestamp 1636986456
transform 1 0 85560 0 1 31008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_889
timestamp 1636986456
transform 1 0 86664 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_901
timestamp 18001
transform 1 0 87768 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_903
timestamp 18001
transform 1 0 87952 0 1 31008
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_7
timestamp 1636986456
transform 1 0 5520 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_19
timestamp 18001
transform 1 0 6624 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_27
timestamp 18001
transform 1 0 7360 0 -1 32096
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_877
timestamp 1636986456
transform 1 0 85560 0 -1 32096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_889
timestamp 1636986456
transform 1 0 86664 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_901
timestamp 18001
transform 1 0 87768 0 -1 32096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1636986456
transform 1 0 5152 0 1 32096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1636986456
transform 1 0 6256 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 18001
transform 1 0 7360 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_50_29
timestamp 18001
transform 1 0 7544 0 1 32096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_877
timestamp 1636986456
transform 1 0 85560 0 1 32096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_889
timestamp 1636986456
transform 1 0 86664 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_901
timestamp 18001
transform 1 0 87768 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_903
timestamp 18001
transform 1 0 87952 0 1 32096
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1636986456
transform 1 0 5152 0 -1 33184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1636986456
transform 1 0 6256 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_27
timestamp 18001
transform 1 0 7360 0 -1 33184
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_877
timestamp 1636986456
transform 1 0 85560 0 -1 33184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_889
timestamp 1636986456
transform 1 0 86664 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_901
timestamp 18001
transform 1 0 87768 0 -1 33184
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_7
timestamp 1636986456
transform 1 0 5520 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_19
timestamp 18001
transform 1 0 6624 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 18001
transform 1 0 7360 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_52_29
timestamp 18001
transform 1 0 7544 0 1 33184
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_877
timestamp 1636986456
transform 1 0 85560 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_889
timestamp 18001
transform 1 0 86664 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_897
timestamp 18001
transform 1 0 87400 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_52_903
timestamp 18001
transform 1 0 87952 0 1 33184
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_7
timestamp 1636986456
transform 1 0 5520 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_19
timestamp 18001
transform 1 0 6624 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_27
timestamp 18001
transform 1 0 7360 0 -1 34272
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_877
timestamp 1636986456
transform 1 0 85560 0 -1 34272
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_889
timestamp 1636986456
transform 1 0 86664 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_901
timestamp 18001
transform 1 0 87768 0 -1 34272
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1636986456
transform 1 0 5152 0 1 34272
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1636986456
transform 1 0 6256 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 18001
transform 1 0 7360 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_29
timestamp 18001
transform 1 0 7544 0 1 34272
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_877
timestamp 1636986456
transform 1 0 85560 0 1 34272
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_889
timestamp 1636986456
transform 1 0 86664 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_901
timestamp 18001
transform 1 0 87768 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_903
timestamp 18001
transform 1 0 87952 0 1 34272
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_7
timestamp 1636986456
transform 1 0 5520 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_19
timestamp 18001
transform 1 0 6624 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_27
timestamp 18001
transform 1 0 7360 0 -1 35360
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_877
timestamp 1636986456
transform 1 0 85560 0 -1 35360
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_889
timestamp 1636986456
transform 1 0 86664 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_901
timestamp 18001
transform 1 0 87768 0 -1 35360
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1636986456
transform 1 0 5152 0 1 35360
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1636986456
transform 1 0 6256 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 18001
transform 1 0 7360 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_56_29
timestamp 18001
transform 1 0 7544 0 1 35360
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_877
timestamp 1636986456
transform 1 0 85560 0 1 35360
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_889
timestamp 1636986456
transform 1 0 86664 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_901
timestamp 18001
transform 1 0 87768 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_903
timestamp 18001
transform 1 0 87952 0 1 35360
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_7
timestamp 1636986456
transform 1 0 5520 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_19
timestamp 18001
transform 1 0 6624 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_27
timestamp 18001
transform 1 0 7360 0 -1 36448
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_877
timestamp 1636986456
transform 1 0 85560 0 -1 36448
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_889
timestamp 1636986456
transform 1 0 86664 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_901
timestamp 18001
transform 1 0 87768 0 -1 36448
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1636986456
transform 1 0 5152 0 1 36448
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1636986456
transform 1 0 6256 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 18001
transform 1 0 7360 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_58_29
timestamp 18001
transform 1 0 7544 0 1 36448
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_877
timestamp 1636986456
transform 1 0 85560 0 1 36448
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_889
timestamp 1636986456
transform 1 0 86664 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_901
timestamp 18001
transform 1 0 87768 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_903
timestamp 18001
transform 1 0 87952 0 1 36448
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_7
timestamp 1636986456
transform 1 0 5520 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_19
timestamp 18001
transform 1 0 6624 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_27
timestamp 18001
transform 1 0 7360 0 -1 37536
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_877
timestamp 1636986456
transform 1 0 85560 0 -1 37536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_889
timestamp 1636986456
transform 1 0 86664 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_901
timestamp 18001
transform 1 0 87768 0 -1 37536
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1636986456
transform 1 0 5152 0 1 37536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1636986456
transform 1 0 6256 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 18001
transform 1 0 7360 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_60_29
timestamp 18001
transform 1 0 7544 0 1 37536
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_877
timestamp 1636986456
transform 1 0 85560 0 1 37536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_889
timestamp 1636986456
transform 1 0 86664 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_901
timestamp 18001
transform 1 0 87768 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_903
timestamp 18001
transform 1 0 87952 0 1 37536
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1636986456
transform 1 0 5152 0 -1 38624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1636986456
transform 1 0 6256 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_27
timestamp 18001
transform 1 0 7360 0 -1 38624
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_877
timestamp 1636986456
transform 1 0 85560 0 -1 38624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_889
timestamp 1636986456
transform 1 0 86664 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_901
timestamp 18001
transform 1 0 87768 0 -1 38624
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_62_7
timestamp 1636986456
transform 1 0 5520 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_19
timestamp 18001
transform 1 0 6624 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 18001
transform 1 0 7360 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_62_29
timestamp 18001
transform 1 0 7544 0 1 38624
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_877
timestamp 1636986456
transform 1 0 85560 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_889
timestamp 18001
transform 1 0 86664 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_897
timestamp 18001
transform 1 0 87400 0 1 38624
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_7
timestamp 1636986456
transform 1 0 5520 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_19
timestamp 18001
transform 1 0 6624 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_27
timestamp 18001
transform 1 0 7360 0 -1 39712
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_877
timestamp 1636986456
transform 1 0 85560 0 -1 39712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_889
timestamp 1636986456
transform 1 0 86664 0 -1 39712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1636986456
transform 1 0 5152 0 1 39712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1636986456
transform 1 0 6256 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 18001
transform 1 0 7360 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_64_29
timestamp 18001
transform 1 0 7544 0 1 39712
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_877
timestamp 1636986456
transform 1 0 85560 0 1 39712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_889
timestamp 1636986456
transform 1 0 86664 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_901
timestamp 18001
transform 1 0 87768 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_903
timestamp 18001
transform 1 0 87952 0 1 39712
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_7
timestamp 1636986456
transform 1 0 5520 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_19
timestamp 18001
transform 1 0 6624 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_27
timestamp 18001
transform 1 0 7360 0 -1 40800
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_65_877
timestamp 1636986456
transform 1 0 85560 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_889
timestamp 18001
transform 1 0 86664 0 -1 40800
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1636986456
transform 1 0 5152 0 1 40800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 1636986456
transform 1 0 6256 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 18001
transform 1 0 7360 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_66_29
timestamp 18001
transform 1 0 7544 0 1 40800
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_877
timestamp 1636986456
transform 1 0 85560 0 1 40800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_889
timestamp 1636986456
transform 1 0 86664 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_901
timestamp 18001
transform 1 0 87768 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_903
timestamp 18001
transform 1 0 87952 0 1 40800
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_7
timestamp 1636986456
transform 1 0 5520 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_19
timestamp 18001
transform 1 0 6624 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_27
timestamp 18001
transform 1 0 7360 0 -1 41888
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_67_877
timestamp 1636986456
transform 1 0 85560 0 -1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_889
timestamp 1636986456
transform 1 0 86664 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_901
timestamp 18001
transform 1 0 87768 0 -1 41888
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1636986456
transform 1 0 5152 0 1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1636986456
transform 1 0 6256 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 18001
transform 1 0 7360 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_68_29
timestamp 18001
transform 1 0 7544 0 1 41888
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_877
timestamp 1636986456
transform 1 0 85560 0 1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_889
timestamp 1636986456
transform 1 0 86664 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_901
timestamp 18001
transform 1 0 87768 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_903
timestamp 18001
transform 1 0 87952 0 1 41888
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_69_7
timestamp 1636986456
transform 1 0 5520 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_19
timestamp 18001
transform 1 0 6624 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_69_27
timestamp 18001
transform 1 0 7360 0 -1 42976
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_69_877
timestamp 1636986456
transform 1 0 85560 0 -1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_889
timestamp 1636986456
transform 1 0 86664 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_901
timestamp 18001
transform 1 0 87768 0 -1 42976
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1636986456
transform 1 0 5152 0 1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1636986456
transform 1 0 6256 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 18001
transform 1 0 7360 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_70_29
timestamp 18001
transform 1 0 7544 0 1 42976
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_877
timestamp 1636986456
transform 1 0 85560 0 1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_889
timestamp 1636986456
transform 1 0 86664 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_901
timestamp 18001
transform 1 0 87768 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_903
timestamp 18001
transform 1 0 87952 0 1 42976
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1636986456
transform 1 0 5152 0 -1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1636986456
transform 1 0 6256 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_71_27
timestamp 18001
transform 1 0 7360 0 -1 44064
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_71_877
timestamp 1636986456
transform 1 0 85560 0 -1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_889
timestamp 1636986456
transform 1 0 86664 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_901
timestamp 18001
transform 1 0 87768 0 -1 44064
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_72_7
timestamp 1636986456
transform 1 0 5520 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_19
timestamp 18001
transform 1 0 6624 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 18001
transform 1 0 7360 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_72_29
timestamp 18001
transform 1 0 7544 0 1 44064
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_877
timestamp 1636986456
transform 1 0 85560 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_889
timestamp 18001
transform 1 0 86664 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_72_897
timestamp 18001
transform 1 0 87400 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_72_903
timestamp 18001
transform 1 0 87952 0 1 44064
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_7
timestamp 1636986456
transform 1 0 5520 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_19
timestamp 18001
transform 1 0 6624 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_27
timestamp 18001
transform 1 0 7360 0 -1 45152
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_877
timestamp 1636986456
transform 1 0 85560 0 -1 45152
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_889
timestamp 1636986456
transform 1 0 86664 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_901
timestamp 18001
transform 1 0 87768 0 -1 45152
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_8
timestamp 1636986456
transform 1 0 5612 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_20
timestamp 18001
transform 1 0 6716 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_29
timestamp 18001
transform 1 0 7544 0 1 45152
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_885
timestamp 1636986456
transform 1 0 86296 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_897
timestamp 18001
transform 1 0 87400 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_901
timestamp 18001
transform 1 0 87768 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_74_903
timestamp 18001
transform 1 0 87952 0 1 45152
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_3
timestamp 1636986456
transform 1 0 5152 0 -1 46240
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_15
timestamp 1636986456
transform 1 0 6256 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_27
timestamp 18001
transform 1 0 7360 0 -1 46240
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_75_877
timestamp 1636986456
transform 1 0 85560 0 -1 46240
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_889
timestamp 1636986456
transform 1 0 86664 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_901
timestamp 18001
transform 1 0 87768 0 -1 46240
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1636986456
transform 1 0 5152 0 1 46240
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1636986456
transform 1 0 6256 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 18001
transform 1 0 7360 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_76_29
timestamp 18001
transform 1 0 7544 0 1 46240
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_877
timestamp 1636986456
transform 1 0 85560 0 1 46240
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_889
timestamp 1636986456
transform 1 0 86664 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_901
timestamp 18001
transform 1 0 87768 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_903
timestamp 18001
transform 1 0 87952 0 1 46240
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1636986456
transform 1 0 5152 0 -1 47328
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1636986456
transform 1 0 6256 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_77_27
timestamp 18001
transform 1 0 7360 0 -1 47328
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_77_877
timestamp 1636986456
transform 1 0 85560 0 -1 47328
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_889
timestamp 1636986456
transform 1 0 86664 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_77_901
timestamp 18001
transform 1 0 87768 0 -1 47328
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1636986456
transform 1 0 5152 0 1 47328
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1636986456
transform 1 0 6256 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 18001
transform 1 0 7360 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_78_29
timestamp 18001
transform 1 0 7544 0 1 47328
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_877
timestamp 1636986456
transform 1 0 85560 0 1 47328
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_889
timestamp 1636986456
transform 1 0 86664 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_901
timestamp 18001
transform 1 0 87768 0 1 47328
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1636986456
transform 1 0 5152 0 -1 48416
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1636986456
transform 1 0 6256 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_27
timestamp 18001
transform 1 0 7360 0 -1 48416
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_79_877
timestamp 1636986456
transform 1 0 85560 0 -1 48416
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_889
timestamp 1636986456
transform 1 0 86664 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_901
timestamp 18001
transform 1 0 87768 0 -1 48416
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_3
timestamp 1636986456
transform 1 0 5152 0 1 48416
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 1636986456
transform 1 0 6256 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 18001
transform 1 0 7360 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_80_29
timestamp 18001
transform 1 0 7544 0 1 48416
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_879
timestamp 1636986456
transform 1 0 85744 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_891
timestamp 18001
transform 1 0 86848 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_899
timestamp 18001
transform 1 0 87584 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_80_903
timestamp 18001
transform 1 0 87952 0 1 48416
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1636986456
transform 1 0 5152 0 -1 49504
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1636986456
transform 1 0 6256 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_81_27
timestamp 18001
transform 1 0 7360 0 -1 49504
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_81_877
timestamp 1636986456
transform 1 0 85560 0 -1 49504
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_889
timestamp 1636986456
transform 1 0 86664 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_901
timestamp 18001
transform 1 0 87768 0 -1 49504
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_82_3
timestamp 1636986456
transform 1 0 5152 0 1 49504
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_15
timestamp 1636986456
transform 1 0 6256 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 18001
transform 1 0 7360 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_82_29
timestamp 18001
transform 1 0 7544 0 1 49504
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_879
timestamp 1636986456
transform 1 0 85744 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_891
timestamp 18001
transform 1 0 86848 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_899
timestamp 18001
transform 1 0 87584 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_903
timestamp 18001
transform 1 0 87952 0 1 49504
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_83_3
timestamp 1636986456
transform 1 0 5152 0 -1 50592
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_15
timestamp 1636986456
transform 1 0 6256 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_83_27
timestamp 18001
transform 1 0 7360 0 -1 50592
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_83_877
timestamp 1636986456
transform 1 0 85560 0 -1 50592
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_889
timestamp 1636986456
transform 1 0 86664 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_901
timestamp 18001
transform 1 0 87768 0 -1 50592
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_84_3
timestamp 1636986456
transform 1 0 5152 0 1 50592
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_15
timestamp 1636986456
transform 1 0 6256 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 18001
transform 1 0 7360 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_84_29
timestamp 18001
transform 1 0 7544 0 1 50592
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_879
timestamp 1636986456
transform 1 0 85744 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_891
timestamp 18001
transform 1 0 86848 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_84_899
timestamp 18001
transform 1 0 87584 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_84_903
timestamp 18001
transform 1 0 87952 0 1 50592
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_85_8
timestamp 1636986456
transform 1 0 5612 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_20
timestamp 18001
transform 1 0 6716 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_85_28
timestamp 18001
transform 1 0 7452 0 -1 51680
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_85_877
timestamp 1636986456
transform 1 0 85560 0 -1 51680
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_889
timestamp 1636986456
transform 1 0 86664 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_85_901
timestamp 18001
transform 1 0 87768 0 -1 51680
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_86_3
timestamp 1636986456
transform 1 0 5152 0 1 51680
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_15
timestamp 1636986456
transform 1 0 6256 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 18001
transform 1 0 7360 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_86_29
timestamp 18001
transform 1 0 7544 0 1 51680
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_877
timestamp 1636986456
transform 1 0 85560 0 1 51680
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_889
timestamp 1636986456
transform 1 0 86664 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_901
timestamp 18001
transform 1 0 87768 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_903
timestamp 18001
transform 1 0 87952 0 1 51680
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_87_3
timestamp 1636986456
transform 1 0 5152 0 -1 52768
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_15
timestamp 1636986456
transform 1 0 6256 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_87_27
timestamp 18001
transform 1 0 7360 0 -1 52768
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_87_877
timestamp 1636986456
transform 1 0 85560 0 -1 52768
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_889
timestamp 1636986456
transform 1 0 86664 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_901
timestamp 18001
transform 1 0 87768 0 -1 52768
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_88_8
timestamp 1636986456
transform 1 0 5612 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_20
timestamp 18001
transform 1 0 6716 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_88_29
timestamp 18001
transform 1 0 7544 0 1 52768
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_877
timestamp 1636986456
transform 1 0 85560 0 1 52768
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_889
timestamp 1636986456
transform 1 0 86664 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_901
timestamp 18001
transform 1 0 87768 0 1 52768
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_3
timestamp 1636986456
transform 1 0 5152 0 -1 53856
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_15
timestamp 1636986456
transform 1 0 6256 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_89_27
timestamp 18001
transform 1 0 7360 0 -1 53856
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_89_877
timestamp 1636986456
transform 1 0 85560 0 -1 53856
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_889
timestamp 1636986456
transform 1 0 86664 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_901
timestamp 18001
transform 1 0 87768 0 -1 53856
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_90_8
timestamp 1636986456
transform 1 0 5612 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_90_20
timestamp 18001
transform 1 0 6716 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_90_29
timestamp 18001
transform 1 0 7544 0 1 53856
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_877
timestamp 1636986456
transform 1 0 85560 0 1 53856
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_889
timestamp 1636986456
transform 1 0 86664 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_901
timestamp 18001
transform 1 0 87768 0 1 53856
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_3
timestamp 1636986456
transform 1 0 5152 0 -1 54944
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_15
timestamp 1636986456
transform 1 0 6256 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_91_27
timestamp 18001
transform 1 0 7360 0 -1 54944
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_91_877
timestamp 1636986456
transform 1 0 85560 0 -1 54944
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_889
timestamp 1636986456
transform 1 0 86664 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_901
timestamp 18001
transform 1 0 87768 0 -1 54944
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_92_8
timestamp 1636986456
transform 1 0 5612 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_20
timestamp 18001
transform 1 0 6716 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_92_29
timestamp 18001
transform 1 0 7544 0 1 54944
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_877
timestamp 1636986456
transform 1 0 85560 0 1 54944
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_889
timestamp 1636986456
transform 1 0 86664 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_901
timestamp 18001
transform 1 0 87768 0 1 54944
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_3
timestamp 1636986456
transform 1 0 5152 0 -1 56032
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_15
timestamp 1636986456
transform 1 0 6256 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_93_27
timestamp 18001
transform 1 0 7360 0 -1 56032
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_93_877
timestamp 1636986456
transform 1 0 85560 0 -1 56032
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_889
timestamp 1636986456
transform 1 0 86664 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_901
timestamp 18001
transform 1 0 87768 0 -1 56032
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_94_8
timestamp 1636986456
transform 1 0 5612 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_20
timestamp 18001
transform 1 0 6716 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_94_29
timestamp 18001
transform 1 0 7544 0 1 56032
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_877
timestamp 1636986456
transform 1 0 85560 0 1 56032
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_889
timestamp 1636986456
transform 1 0 86664 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_901
timestamp 18001
transform 1 0 87768 0 1 56032
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_8
timestamp 1636986456
transform 1 0 5612 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_20
timestamp 18001
transform 1 0 6716 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_95_28
timestamp 18001
transform 1 0 7452 0 -1 57120
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_95_877
timestamp 1636986456
transform 1 0 85560 0 -1 57120
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_889
timestamp 1636986456
transform 1 0 86664 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_95_901
timestamp 18001
transform 1 0 87768 0 -1 57120
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_96_3
timestamp 1636986456
transform 1 0 5152 0 1 57120
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_15
timestamp 1636986456
transform 1 0 6256 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_27
timestamp 18001
transform 1 0 7360 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_96_29
timestamp 18001
transform 1 0 7544 0 1 57120
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_877
timestamp 1636986456
transform 1 0 85560 0 1 57120
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_889
timestamp 1636986456
transform 1 0 86664 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_901
timestamp 18001
transform 1 0 87768 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_96_903
timestamp 18001
transform 1 0 87952 0 1 57120
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_97_3
timestamp 1636986456
transform 1 0 5152 0 -1 58208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_15
timestamp 1636986456
transform 1 0 6256 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_97_27
timestamp 18001
transform 1 0 7360 0 -1 58208
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_97_877
timestamp 1636986456
transform 1 0 85560 0 -1 58208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_889
timestamp 1636986456
transform 1 0 86664 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_901
timestamp 18001
transform 1 0 87768 0 -1 58208
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_98_8
timestamp 1636986456
transform 1 0 5612 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_20
timestamp 18001
transform 1 0 6716 0 1 58208
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_98_29
timestamp 18001
transform 1 0 7544 0 1 58208
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_877
timestamp 1636986456
transform 1 0 85560 0 1 58208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_889
timestamp 1636986456
transform 1 0 86664 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_901
timestamp 18001
transform 1 0 87768 0 1 58208
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_3
timestamp 1636986456
transform 1 0 5152 0 -1 59296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_15
timestamp 1636986456
transform 1 0 6256 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_99_27
timestamp 18001
transform 1 0 7360 0 -1 59296
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_99_877
timestamp 1636986456
transform 1 0 85560 0 -1 59296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_889
timestamp 1636986456
transform 1 0 86664 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_901
timestamp 18001
transform 1 0 87768 0 -1 59296
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_100_8
timestamp 1636986456
transform 1 0 5612 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_20
timestamp 18001
transform 1 0 6716 0 1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_100_29
timestamp 18001
transform 1 0 7544 0 1 59296
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_877
timestamp 1636986456
transform 1 0 85560 0 1 59296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_889
timestamp 1636986456
transform 1 0 86664 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_901
timestamp 18001
transform 1 0 87768 0 1 59296
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_3
timestamp 1636986456
transform 1 0 5152 0 -1 60384
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_15
timestamp 1636986456
transform 1 0 6256 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_27
timestamp 18001
transform 1 0 7360 0 -1 60384
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_877
timestamp 1636986456
transform 1 0 85560 0 -1 60384
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_889
timestamp 1636986456
transform 1 0 86664 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_901
timestamp 18001
transform 1 0 87768 0 -1 60384
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_102_8
timestamp 1636986456
transform 1 0 5612 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_102_20
timestamp 18001
transform 1 0 6716 0 1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_102_29
timestamp 18001
transform 1 0 7544 0 1 60384
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_877
timestamp 1636986456
transform 1 0 85560 0 1 60384
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_889
timestamp 1636986456
transform 1 0 86664 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_102_901
timestamp 18001
transform 1 0 87768 0 1 60384
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_3
timestamp 1636986456
transform 1 0 5152 0 -1 61472
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_15
timestamp 1636986456
transform 1 0 6256 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_103_27
timestamp 18001
transform 1 0 7360 0 -1 61472
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_103_877
timestamp 1636986456
transform 1 0 85560 0 -1 61472
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_889
timestamp 1636986456
transform 1 0 86664 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_901
timestamp 18001
transform 1 0 87768 0 -1 61472
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_104_8
timestamp 1636986456
transform 1 0 5612 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_104_20
timestamp 18001
transform 1 0 6716 0 1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_104_29
timestamp 18001
transform 1 0 7544 0 1 61472
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_877
timestamp 1636986456
transform 1 0 85560 0 1 61472
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_889
timestamp 1636986456
transform 1 0 86664 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_104_901
timestamp 18001
transform 1 0 87768 0 1 61472
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_8
timestamp 1636986456
transform 1 0 5612 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_105_20
timestamp 18001
transform 1 0 6716 0 -1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_105_28
timestamp 18001
transform 1 0 7452 0 -1 62560
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_105_877
timestamp 1636986456
transform 1 0 85560 0 -1 62560
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_889
timestamp 1636986456
transform 1 0 86664 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_105_901
timestamp 18001
transform 1 0 87768 0 -1 62560
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_106_3
timestamp 1636986456
transform 1 0 5152 0 1 62560
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_15
timestamp 1636986456
transform 1 0 6256 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_106_27
timestamp 18001
transform 1 0 7360 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_106_29
timestamp 18001
transform 1 0 7544 0 1 62560
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_877
timestamp 1636986456
transform 1 0 85560 0 1 62560
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_889
timestamp 1636986456
transform 1 0 86664 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_106_901
timestamp 18001
transform 1 0 87768 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_106_903
timestamp 18001
transform 1 0 87952 0 1 62560
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_107_3
timestamp 1636986456
transform 1 0 5152 0 -1 63648
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_15
timestamp 1636986456
transform 1 0 6256 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_107_27
timestamp 18001
transform 1 0 7360 0 -1 63648
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_877
timestamp 1636986456
transform 1 0 85560 0 -1 63648
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_889
timestamp 1636986456
transform 1 0 86664 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_901
timestamp 18001
transform 1 0 87768 0 -1 63648
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_29
timestamp 18001
transform 1 0 7544 0 1 63648
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_877
timestamp 1636986456
transform 1 0 85560 0 1 63648
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_889
timestamp 1636986456
transform 1 0 86664 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_108_901
timestamp 18001
transform 1 0 87768 0 1 63648
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_3
timestamp 1636986456
transform 1 0 5152 0 -1 64736
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_15
timestamp 1636986456
transform 1 0 6256 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_109_27
timestamp 18001
transform 1 0 7360 0 -1 64736
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_877
timestamp 1636986456
transform 1 0 85560 0 -1 64736
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_889
timestamp 1636986456
transform 1 0 86664 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_901
timestamp 18001
transform 1 0 87768 0 -1 64736
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_110_8
timestamp 1636986456
transform 1 0 5612 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_110_20
timestamp 18001
transform 1 0 6716 0 1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_110_29
timestamp 18001
transform 1 0 7544 0 1 64736
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_877
timestamp 1636986456
transform 1 0 85560 0 1 64736
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_889
timestamp 1636986456
transform 1 0 86664 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_110_901
timestamp 18001
transform 1 0 87768 0 1 64736
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_3
timestamp 1636986456
transform 1 0 5152 0 -1 65824
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_15
timestamp 1636986456
transform 1 0 6256 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_111_27
timestamp 18001
transform 1 0 7360 0 -1 65824
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_111_877
timestamp 1636986456
transform 1 0 85560 0 -1 65824
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_889
timestamp 1636986456
transform 1 0 86664 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_901
timestamp 18001
transform 1 0 87768 0 -1 65824
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_112_8
timestamp 1636986456
transform 1 0 5612 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_112_20
timestamp 18001
transform 1 0 6716 0 1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_112_29
timestamp 18001
transform 1 0 7544 0 1 65824
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_877
timestamp 1636986456
transform 1 0 85560 0 1 65824
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_889
timestamp 1636986456
transform 1 0 86664 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_112_901
timestamp 18001
transform 1 0 87768 0 1 65824
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_3
timestamp 1636986456
transform 1 0 5152 0 -1 66912
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_15
timestamp 1636986456
transform 1 0 6256 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_113_27
timestamp 18001
transform 1 0 7360 0 -1 66912
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_113_877
timestamp 1636986456
transform 1 0 85560 0 -1 66912
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_889
timestamp 1636986456
transform 1 0 86664 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_901
timestamp 18001
transform 1 0 87768 0 -1 66912
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_114_7
timestamp 1636986456
transform 1 0 5520 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_114_19
timestamp 18001
transform 1 0 6624 0 1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_114_27
timestamp 18001
transform 1 0 7360 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_114_29
timestamp 18001
transform 1 0 7544 0 1 66912
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_877
timestamp 1636986456
transform 1 0 85560 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_114_889
timestamp 18001
transform 1 0 86664 0 1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_114_897
timestamp 18001
transform 1 0 87400 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_114_903
timestamp 18001
transform 1 0 87952 0 1 66912
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_7
timestamp 1636986456
transform 1 0 5520 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_115_19
timestamp 18001
transform 1 0 6624 0 -1 68000
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_115_27
timestamp 18001
transform 1 0 7360 0 -1 68000
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_115_877
timestamp 1636986456
transform 1 0 85560 0 -1 68000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_889
timestamp 1636986456
transform 1 0 86664 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_115_901
timestamp 18001
transform 1 0 87768 0 -1 68000
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_3
timestamp 1636986456
transform 1 0 5152 0 1 68000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_15
timestamp 1636986456
transform 1 0 6256 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_116_27
timestamp 18001
transform 1 0 7360 0 1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_116_29
timestamp 18001
transform 1 0 7544 0 1 68000
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_877
timestamp 1636986456
transform 1 0 85560 0 1 68000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_889
timestamp 1636986456
transform 1 0 86664 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_116_901
timestamp 18001
transform 1 0 87768 0 1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_116_903
timestamp 18001
transform 1 0 87952 0 1 68000
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_117_3
timestamp 1636986456
transform 1 0 5152 0 -1 69088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_15
timestamp 1636986456
transform 1 0 6256 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_27
timestamp 18001
transform 1 0 7360 0 -1 69088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_877
timestamp 1636986456
transform 1 0 85560 0 -1 69088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_889
timestamp 1636986456
transform 1 0 86664 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_901
timestamp 18001
transform 1 0 87768 0 -1 69088
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_118_7
timestamp 1636986456
transform 1 0 5520 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_118_19
timestamp 18001
transform 1 0 6624 0 1 69088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_118_27
timestamp 18001
transform 1 0 7360 0 1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_118_29
timestamp 18001
transform 1 0 7544 0 1 69088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_877
timestamp 1636986456
transform 1 0 85560 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_118_889
timestamp 18001
transform 1 0 86664 0 1 69088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_118_897
timestamp 18001
transform 1 0 87400 0 1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_118_903
timestamp 18001
transform 1 0 87952 0 1 69088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_3
timestamp 1636986456
transform 1 0 5152 0 -1 70176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_15
timestamp 1636986456
transform 1 0 6256 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_119_27
timestamp 18001
transform 1 0 7360 0 -1 70176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_119_877
timestamp 1636986456
transform 1 0 85560 0 -1 70176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_889
timestamp 1636986456
transform 1 0 86664 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_901
timestamp 18001
transform 1 0 87768 0 -1 70176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_120_7
timestamp 1636986456
transform 1 0 5520 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_120_19
timestamp 18001
transform 1 0 6624 0 1 70176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_120_27
timestamp 18001
transform 1 0 7360 0 1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_120_29
timestamp 18001
transform 1 0 7544 0 1 70176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_877
timestamp 1636986456
transform 1 0 85560 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_120_889
timestamp 18001
transform 1 0 86664 0 1 70176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_120_897
timestamp 18001
transform 1 0 87400 0 1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_120_903
timestamp 18001
transform 1 0 87952 0 1 70176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_3
timestamp 1636986456
transform 1 0 5152 0 -1 71264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_15
timestamp 1636986456
transform 1 0 6256 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_121_27
timestamp 18001
transform 1 0 7360 0 -1 71264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_121_877
timestamp 1636986456
transform 1 0 85560 0 -1 71264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_889
timestamp 1636986456
transform 1 0 86664 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_901
timestamp 18001
transform 1 0 87768 0 -1 71264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_122_7
timestamp 1636986456
transform 1 0 5520 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_122_19
timestamp 18001
transform 1 0 6624 0 1 71264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_122_27
timestamp 18001
transform 1 0 7360 0 1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_122_29
timestamp 18001
transform 1 0 7544 0 1 71264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_877
timestamp 1636986456
transform 1 0 85560 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_122_889
timestamp 18001
transform 1 0 86664 0 1 71264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_122_897
timestamp 18001
transform 1 0 87400 0 1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_122_903
timestamp 18001
transform 1 0 87952 0 1 71264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_3
timestamp 1636986456
transform 1 0 5152 0 -1 72352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_15
timestamp 1636986456
transform 1 0 6256 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_27
timestamp 18001
transform 1 0 7360 0 -1 72352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_123_877
timestamp 1636986456
transform 1 0 85560 0 -1 72352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_889
timestamp 1636986456
transform 1 0 86664 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_901
timestamp 18001
transform 1 0 87768 0 -1 72352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_124_7
timestamp 1636986456
transform 1 0 5520 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_124_19
timestamp 18001
transform 1 0 6624 0 1 72352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_124_27
timestamp 18001
transform 1 0 7360 0 1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_124_29
timestamp 18001
transform 1 0 7544 0 1 72352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_877
timestamp 1636986456
transform 1 0 85560 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_124_889
timestamp 18001
transform 1 0 86664 0 1 72352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_124_897
timestamp 18001
transform 1 0 87400 0 1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_124_903
timestamp 18001
transform 1 0 87952 0 1 72352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_7
timestamp 1636986456
transform 1 0 5520 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_125_19
timestamp 18001
transform 1 0 6624 0 -1 73440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_125_27
timestamp 18001
transform 1 0 7360 0 -1 73440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_125_877
timestamp 1636986456
transform 1 0 85560 0 -1 73440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_889
timestamp 1636986456
transform 1 0 86664 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_125_901
timestamp 18001
transform 1 0 87768 0 -1 73440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_3
timestamp 1636986456
transform 1 0 5152 0 1 73440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_15
timestamp 1636986456
transform 1 0 6256 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_126_27
timestamp 18001
transform 1 0 7360 0 1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_126_29
timestamp 18001
transform 1 0 7544 0 1 73440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_877
timestamp 1636986456
transform 1 0 85560 0 1 73440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_889
timestamp 1636986456
transform 1 0 86664 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_126_901
timestamp 18001
transform 1 0 87768 0 1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_126_903
timestamp 18001
transform 1 0 87952 0 1 73440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_127_3
timestamp 1636986456
transform 1 0 5152 0 -1 74528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_15
timestamp 1636986456
transform 1 0 6256 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_127_27
timestamp 18001
transform 1 0 7360 0 -1 74528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_127_877
timestamp 1636986456
transform 1 0 85560 0 -1 74528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_889
timestamp 1636986456
transform 1 0 86664 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_901
timestamp 18001
transform 1 0 87768 0 -1 74528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_128_7
timestamp 1636986456
transform 1 0 5520 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_128_19
timestamp 18001
transform 1 0 6624 0 1 74528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_128_27
timestamp 18001
transform 1 0 7360 0 1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_128_29
timestamp 18001
transform 1 0 7544 0 1 74528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_877
timestamp 1636986456
transform 1 0 85560 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_128_889
timestamp 18001
transform 1 0 86664 0 1 74528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_128_897
timestamp 18001
transform 1 0 87400 0 1 74528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_129_3
timestamp 1636986456
transform 1 0 5152 0 -1 75616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_15
timestamp 1636986456
transform 1 0 6256 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_129_27
timestamp 18001
transform 1 0 7360 0 -1 75616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_129_877
timestamp 1636986456
transform 1 0 85560 0 -1 75616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_889
timestamp 1636986456
transform 1 0 86664 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_901
timestamp 18001
transform 1 0 87768 0 -1 75616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_130_7
timestamp 1636986456
transform 1 0 5520 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_130_19
timestamp 18001
transform 1 0 6624 0 1 75616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_130_27
timestamp 18001
transform 1 0 7360 0 1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_130_29
timestamp 18001
transform 1 0 7544 0 1 75616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_877
timestamp 1636986456
transform 1 0 85560 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_130_889
timestamp 18001
transform 1 0 86664 0 1 75616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_130_897
timestamp 18001
transform 1 0 87400 0 1 75616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_131_3
timestamp 1636986456
transform 1 0 5152 0 -1 76704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_15
timestamp 1636986456
transform 1 0 6256 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_131_27
timestamp 18001
transform 1 0 7360 0 -1 76704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_131_877
timestamp 1636986456
transform 1 0 85560 0 -1 76704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_889
timestamp 1636986456
transform 1 0 86664 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_901
timestamp 18001
transform 1 0 87768 0 -1 76704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_132_7
timestamp 1636986456
transform 1 0 5520 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_132_19
timestamp 18001
transform 1 0 6624 0 1 76704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_132_27
timestamp 18001
transform 1 0 7360 0 1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_132_29
timestamp 18001
transform 1 0 7544 0 1 76704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_877
timestamp 1636986456
transform 1 0 85560 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_132_889
timestamp 18001
transform 1 0 86664 0 1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_132_905
timestamp 18001
transform 1 0 88136 0 1 76704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_133_3
timestamp 1636986456
transform 1 0 5152 0 -1 77792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_15
timestamp 1636986456
transform 1 0 6256 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_133_27
timestamp 18001
transform 1 0 7360 0 -1 77792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_133_877
timestamp 1636986456
transform 1 0 85560 0 -1 77792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_889
timestamp 1636986456
transform 1 0 86664 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_901
timestamp 18001
transform 1 0 87768 0 -1 77792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_134_7
timestamp 1636986456
transform 1 0 5520 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_134_19
timestamp 18001
transform 1 0 6624 0 1 77792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_134_27
timestamp 18001
transform 1 0 7360 0 1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_134_29
timestamp 18001
transform 1 0 7544 0 1 77792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_877
timestamp 1636986456
transform 1 0 85560 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_134_889
timestamp 18001
transform 1 0 86664 0 1 77792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_134_897
timestamp 18001
transform 1 0 87400 0 1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_134_903
timestamp 18001
transform 1 0 87952 0 1 77792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_7
timestamp 1636986456
transform 1 0 5520 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_135_19
timestamp 18001
transform 1 0 6624 0 -1 78880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_135_27
timestamp 18001
transform 1 0 7360 0 -1 78880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_135_877
timestamp 1636986456
transform 1 0 85560 0 -1 78880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_889
timestamp 1636986456
transform 1 0 86664 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_135_901
timestamp 18001
transform 1 0 87768 0 -1 78880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_3
timestamp 1636986456
transform 1 0 5152 0 1 78880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_15
timestamp 1636986456
transform 1 0 6256 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_136_27
timestamp 18001
transform 1 0 7360 0 1 78880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_136_29
timestamp 18001
transform 1 0 7544 0 1 78880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_877
timestamp 1636986456
transform 1 0 85560 0 1 78880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_889
timestamp 1636986456
transform 1 0 86664 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_136_901
timestamp 18001
transform 1 0 87768 0 1 78880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_136_903
timestamp 18001
transform 1 0 87952 0 1 78880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_137_3
timestamp 1636986456
transform 1 0 5152 0 -1 79968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_15
timestamp 1636986456
transform 1 0 6256 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_137_27
timestamp 18001
transform 1 0 7360 0 -1 79968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_137_877
timestamp 1636986456
transform 1 0 85560 0 -1 79968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_889
timestamp 1636986456
transform 1 0 86664 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_901
timestamp 18001
transform 1 0 87768 0 -1 79968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_138_7
timestamp 1636986456
transform 1 0 5520 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_138_19
timestamp 18001
transform 1 0 6624 0 1 79968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_138_27
timestamp 18001
transform 1 0 7360 0 1 79968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_138_29
timestamp 18001
transform 1 0 7544 0 1 79968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_138_877
timestamp 1636986456
transform 1 0 85560 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_138_889
timestamp 18001
transform 1 0 86664 0 1 79968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_138_897
timestamp 18001
transform 1 0 87400 0 1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_138_903
timestamp 18001
transform 1 0 87952 0 1 79968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_139_3
timestamp 1636986456
transform 1 0 5152 0 -1 81056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_15
timestamp 1636986456
transform 1 0 6256 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_139_27
timestamp 18001
transform 1 0 7360 0 -1 81056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_139_877
timestamp 1636986456
transform 1 0 85560 0 -1 81056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_889
timestamp 1636986456
transform 1 0 86664 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_139_901
timestamp 18001
transform 1 0 87768 0 -1 81056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_140_3
timestamp 1636986456
transform 1 0 5152 0 1 81056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_15
timestamp 1636986456
transform 1 0 6256 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_140_27
timestamp 18001
transform 1 0 7360 0 1 81056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_140_29
timestamp 18001
transform 1 0 7544 0 1 81056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_140_877
timestamp 1636986456
transform 1 0 85560 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_140_889
timestamp 18001
transform 1 0 86664 0 1 81056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_140_897
timestamp 18001
transform 1 0 87400 0 1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_140_903
timestamp 18001
transform 1 0 87952 0 1 81056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_141_3
timestamp 1636986456
transform 1 0 5152 0 -1 82144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_15
timestamp 1636986456
transform 1 0 6256 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_141_27
timestamp 18001
transform 1 0 7360 0 -1 82144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_141_877
timestamp 1636986456
transform 1 0 85560 0 -1 82144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_889
timestamp 1636986456
transform 1 0 86664 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_141_901
timestamp 18001
transform 1 0 87768 0 -1 82144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_142_3
timestamp 1636986456
transform 1 0 5152 0 1 82144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_15
timestamp 1636986456
transform 1 0 6256 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_142_27
timestamp 18001
transform 1 0 7360 0 1 82144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_142_29
timestamp 18001
transform 1 0 7544 0 1 82144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_142_877
timestamp 1636986456
transform 1 0 85560 0 1 82144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_889
timestamp 1636986456
transform 1 0 86664 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_142_901
timestamp 18001
transform 1 0 87768 0 1 82144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_142_903
timestamp 18001
transform 1 0 87952 0 1 82144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_143_3
timestamp 1636986456
transform 1 0 5152 0 -1 83232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_15
timestamp 1636986456
transform 1 0 6256 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_143_27
timestamp 18001
transform 1 0 7360 0 -1 83232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_143_877
timestamp 1636986456
transform 1 0 85560 0 -1 83232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_889
timestamp 1636986456
transform 1 0 86664 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_143_901
timestamp 18001
transform 1 0 87768 0 -1 83232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_144_3
timestamp 1636986456
transform 1 0 5152 0 1 83232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_15
timestamp 1636986456
transform 1 0 6256 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_144_27
timestamp 18001
transform 1 0 7360 0 1 83232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_144_29
timestamp 18001
transform 1 0 7544 0 1 83232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_144_877
timestamp 1636986456
transform 1 0 85560 0 1 83232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_889
timestamp 1636986456
transform 1 0 86664 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_144_901
timestamp 18001
transform 1 0 87768 0 1 83232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_144_903
timestamp 18001
transform 1 0 87952 0 1 83232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_145_3
timestamp 1636986456
transform 1 0 5152 0 -1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_15
timestamp 1636986456
transform 1 0 6256 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_145_27
timestamp 18001
transform 1 0 7360 0 -1 84320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_145_877
timestamp 1636986456
transform 1 0 85560 0 -1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_889
timestamp 1636986456
transform 1 0 86664 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_145_901
timestamp 18001
transform 1 0 87768 0 -1 84320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_146_3
timestamp 1636986456
transform 1 0 5152 0 1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_15
timestamp 1636986456
transform 1 0 6256 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_146_27
timestamp 18001
transform 1 0 7360 0 1 84320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_146_29
timestamp 1636986456
transform 1 0 7544 0 1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_41
timestamp 1636986456
transform 1 0 8648 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_146_53
timestamp 18001
transform 1 0 9752 0 1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_146_57
timestamp 18001
transform 1 0 10120 0 1 84320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_146_61
timestamp 18001
transform 1 0 10488 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_146_64
timestamp 18001
transform 1 0 10764 0 1 84320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_146_72
timestamp 18001
transform 1 0 11500 0 1 84320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_146_76
timestamp 18001
transform 1 0 11868 0 1 84320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_146_85
timestamp 18001
transform 1 0 12696 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_146_88
timestamp 18001
transform 1 0 12972 0 1 84320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_146_96
timestamp 18001
transform 1 0 13708 0 1 84320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_146_100
timestamp 1636986456
transform 1 0 14076 0 1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_113
timestamp 1636986456
transform 1 0 15272 0 1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_125
timestamp 1636986456
transform 1 0 16376 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_146_137
timestamp 18001
transform 1 0 17480 0 1 84320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_146_141
timestamp 1636986456
transform 1 0 17848 0 1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_153
timestamp 1636986456
transform 1 0 18952 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_146_165
timestamp 18001
transform 1 0 20056 0 1 84320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_146_169
timestamp 1636986456
transform 1 0 20424 0 1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_181
timestamp 1636986456
transform 1 0 21528 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_146_193
timestamp 18001
transform 1 0 22632 0 1 84320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_146_197
timestamp 1636986456
transform 1 0 23000 0 1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_209
timestamp 1636986456
transform 1 0 24104 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_146_221
timestamp 18001
transform 1 0 25208 0 1 84320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_146_225
timestamp 1636986456
transform 1 0 25576 0 1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_237
timestamp 1636986456
transform 1 0 26680 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_146_249
timestamp 18001
transform 1 0 27784 0 1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_146_253
timestamp 18001
transform 1 0 28152 0 1 84320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_146_259
timestamp 18001
transform 1 0 28704 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_146_281
timestamp 18001
transform 1 0 30728 0 1 84320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_146_286
timestamp 1636986456
transform 1 0 31188 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_146_298
timestamp 18001
transform 1 0 32292 0 1 84320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_146_306
timestamp 18001
transform 1 0 33028 0 1 84320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_146_309
timestamp 1636986456
transform 1 0 33304 0 1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_321
timestamp 1636986456
transform 1 0 34408 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_146_333
timestamp 18001
transform 1 0 35512 0 1 84320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_146_337
timestamp 1636986456
transform 1 0 35880 0 1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_349
timestamp 1636986456
transform 1 0 36984 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_146_361
timestamp 18001
transform 1 0 38088 0 1 84320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_146_365
timestamp 1636986456
transform 1 0 38456 0 1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_377
timestamp 1636986456
transform 1 0 39560 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_146_389
timestamp 18001
transform 1 0 40664 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_146_415
timestamp 18001
transform 1 0 43056 0 1 84320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_146_419
timestamp 18001
transform 1 0 43424 0 1 84320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_146_421
timestamp 1636986456
transform 1 0 43608 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_146_433
timestamp 18001
transform 1 0 44712 0 1 84320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_146_439
timestamp 18001
transform 1 0 45264 0 1 84320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_146_449
timestamp 1636986456
transform 1 0 46184 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_146_461
timestamp 18001
transform 1 0 47288 0 1 84320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_146_471
timestamp 18001
transform 1 0 48208 0 1 84320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_146_475
timestamp 18001
transform 1 0 48576 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_146_477
timestamp 18001
transform 1 0 48760 0 1 84320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_146_483
timestamp 18001
transform 1 0 49312 0 1 84320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_146_491
timestamp 18001
transform 1 0 50048 0 1 84320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_146_495
timestamp 18001
transform 1 0 50416 0 1 84320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_146_503
timestamp 18001
transform 1 0 51152 0 1 84320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_146_507
timestamp 1636986456
transform 1 0 51520 0 1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_519
timestamp 1636986456
transform 1 0 52624 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_146_531
timestamp 18001
transform 1 0 53728 0 1 84320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_146_533
timestamp 1636986456
transform 1 0 53912 0 1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_545
timestamp 1636986456
transform 1 0 55016 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_146_557
timestamp 18001
transform 1 0 56120 0 1 84320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_146_561
timestamp 1636986456
transform 1 0 56488 0 1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_573
timestamp 1636986456
transform 1 0 57592 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_146_585
timestamp 18001
transform 1 0 58696 0 1 84320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_146_589
timestamp 1636986456
transform 1 0 59064 0 1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_601
timestamp 1636986456
transform 1 0 60168 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_146_613
timestamp 18001
transform 1 0 61272 0 1 84320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_146_617
timestamp 1636986456
transform 1 0 61640 0 1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_629
timestamp 1636986456
transform 1 0 62744 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_146_641
timestamp 18001
transform 1 0 63848 0 1 84320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_146_645
timestamp 1636986456
transform 1 0 64216 0 1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_657
timestamp 1636986456
transform 1 0 65320 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_146_669
timestamp 18001
transform 1 0 66424 0 1 84320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_146_673
timestamp 1636986456
transform 1 0 66792 0 1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_685
timestamp 1636986456
transform 1 0 67896 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_146_697
timestamp 18001
transform 1 0 69000 0 1 84320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_146_701
timestamp 1636986456
transform 1 0 69368 0 1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_713
timestamp 1636986456
transform 1 0 70472 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_146_725
timestamp 18001
transform 1 0 71576 0 1 84320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_146_729
timestamp 1636986456
transform 1 0 71944 0 1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_741
timestamp 1636986456
transform 1 0 73048 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_146_753
timestamp 18001
transform 1 0 74152 0 1 84320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_146_757
timestamp 1636986456
transform 1 0 74520 0 1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_769
timestamp 1636986456
transform 1 0 75624 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_146_781
timestamp 18001
transform 1 0 76728 0 1 84320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_146_785
timestamp 1636986456
transform 1 0 77096 0 1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_797
timestamp 1636986456
transform 1 0 78200 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_146_809
timestamp 18001
transform 1 0 79304 0 1 84320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_146_813
timestamp 1636986456
transform 1 0 79672 0 1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_825
timestamp 1636986456
transform 1 0 80776 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_146_837
timestamp 18001
transform 1 0 81880 0 1 84320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_146_841
timestamp 1636986456
transform 1 0 82248 0 1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_853
timestamp 1636986456
transform 1 0 83352 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_146_865
timestamp 18001
transform 1 0 84456 0 1 84320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_146_869
timestamp 1636986456
transform 1 0 84824 0 1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_881
timestamp 1636986456
transform 1 0 85928 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_146_893
timestamp 18001
transform 1 0 87032 0 1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_146_897
timestamp 18001
transform 1 0 87400 0 1 84320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_146_905
timestamp 18001
transform 1 0 88136 0 1 84320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_147_3
timestamp 1636986456
transform 1 0 5152 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_15
timestamp 1636986456
transform 1 0 6256 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_27
timestamp 1636986456
transform 1 0 7360 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_39
timestamp 1636986456
transform 1 0 8464 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_147_51
timestamp 18001
transform 1 0 9568 0 -1 85408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_147_55
timestamp 18001
transform 1 0 9936 0 -1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_57
timestamp 1636986456
transform 1 0 10120 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_69
timestamp 1636986456
transform 1 0 11224 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_81
timestamp 1636986456
transform 1 0 12328 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_93
timestamp 1636986456
transform 1 0 13432 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_105
timestamp 18001
transform 1 0 14536 0 -1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_111
timestamp 18001
transform 1 0 15088 0 -1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_113
timestamp 1636986456
transform 1 0 15272 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_125
timestamp 1636986456
transform 1 0 16376 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_137
timestamp 1636986456
transform 1 0 17480 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_149
timestamp 1636986456
transform 1 0 18584 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_161
timestamp 18001
transform 1 0 19688 0 -1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_167
timestamp 18001
transform 1 0 20240 0 -1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_169
timestamp 1636986456
transform 1 0 20424 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_181
timestamp 1636986456
transform 1 0 21528 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_193
timestamp 1636986456
transform 1 0 22632 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_205
timestamp 1636986456
transform 1 0 23736 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_217
timestamp 18001
transform 1 0 24840 0 -1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_223
timestamp 18001
transform 1 0 25392 0 -1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_225
timestamp 1636986456
transform 1 0 25576 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_237
timestamp 1636986456
transform 1 0 26680 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_249
timestamp 1636986456
transform 1 0 27784 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_261
timestamp 1636986456
transform 1 0 28888 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_273
timestamp 18001
transform 1 0 29992 0 -1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_279
timestamp 18001
transform 1 0 30544 0 -1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_281
timestamp 1636986456
transform 1 0 30728 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_293
timestamp 1636986456
transform 1 0 31832 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_305
timestamp 1636986456
transform 1 0 32936 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_317
timestamp 1636986456
transform 1 0 34040 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_329
timestamp 18001
transform 1 0 35144 0 -1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_335
timestamp 18001
transform 1 0 35696 0 -1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_337
timestamp 1636986456
transform 1 0 35880 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_349
timestamp 1636986456
transform 1 0 36984 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_361
timestamp 1636986456
transform 1 0 38088 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_373
timestamp 1636986456
transform 1 0 39192 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_385
timestamp 18001
transform 1 0 40296 0 -1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_391
timestamp 18001
transform 1 0 40848 0 -1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_393
timestamp 1636986456
transform 1 0 41032 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_405
timestamp 1636986456
transform 1 0 42136 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_417
timestamp 1636986456
transform 1 0 43240 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_429
timestamp 1636986456
transform 1 0 44344 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_441
timestamp 18001
transform 1 0 45448 0 -1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_447
timestamp 18001
transform 1 0 46000 0 -1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_449
timestamp 1636986456
transform 1 0 46184 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_461
timestamp 1636986456
transform 1 0 47288 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_473
timestamp 1636986456
transform 1 0 48392 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_485
timestamp 1636986456
transform 1 0 49496 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_497
timestamp 18001
transform 1 0 50600 0 -1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_503
timestamp 18001
transform 1 0 51152 0 -1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_505
timestamp 1636986456
transform 1 0 51336 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_517
timestamp 1636986456
transform 1 0 52440 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_529
timestamp 1636986456
transform 1 0 53544 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_541
timestamp 1636986456
transform 1 0 54648 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_553
timestamp 18001
transform 1 0 55752 0 -1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_559
timestamp 18001
transform 1 0 56304 0 -1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_561
timestamp 1636986456
transform 1 0 56488 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_573
timestamp 1636986456
transform 1 0 57592 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_585
timestamp 1636986456
transform 1 0 58696 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_597
timestamp 1636986456
transform 1 0 59800 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_609
timestamp 18001
transform 1 0 60904 0 -1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_615
timestamp 18001
transform 1 0 61456 0 -1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_617
timestamp 1636986456
transform 1 0 61640 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_629
timestamp 1636986456
transform 1 0 62744 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_641
timestamp 1636986456
transform 1 0 63848 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_653
timestamp 1636986456
transform 1 0 64952 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_665
timestamp 18001
transform 1 0 66056 0 -1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_671
timestamp 18001
transform 1 0 66608 0 -1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_673
timestamp 1636986456
transform 1 0 66792 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_685
timestamp 1636986456
transform 1 0 67896 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_697
timestamp 1636986456
transform 1 0 69000 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_709
timestamp 1636986456
transform 1 0 70104 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_721
timestamp 18001
transform 1 0 71208 0 -1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_727
timestamp 18001
transform 1 0 71760 0 -1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_729
timestamp 1636986456
transform 1 0 71944 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_741
timestamp 1636986456
transform 1 0 73048 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_753
timestamp 1636986456
transform 1 0 74152 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_765
timestamp 1636986456
transform 1 0 75256 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_777
timestamp 18001
transform 1 0 76360 0 -1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_783
timestamp 18001
transform 1 0 76912 0 -1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_785
timestamp 1636986456
transform 1 0 77096 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_797
timestamp 1636986456
transform 1 0 78200 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_809
timestamp 1636986456
transform 1 0 79304 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_821
timestamp 1636986456
transform 1 0 80408 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_833
timestamp 18001
transform 1 0 81512 0 -1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_839
timestamp 18001
transform 1 0 82064 0 -1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_841
timestamp 1636986456
transform 1 0 82248 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_853
timestamp 1636986456
transform 1 0 83352 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_865
timestamp 1636986456
transform 1 0 84456 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_877
timestamp 1636986456
transform 1 0 85560 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_889
timestamp 18001
transform 1 0 86664 0 -1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_895
timestamp 18001
transform 1 0 87216 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_147_897
timestamp 18001
transform 1 0 87400 0 -1 85408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_147_905
timestamp 18001
transform 1 0 88136 0 -1 85408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_148_3
timestamp 1636986456
transform 1 0 5152 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_15
timestamp 1636986456
transform 1 0 6256 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_148_27
timestamp 18001
transform 1 0 7360 0 1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_29
timestamp 1636986456
transform 1 0 7544 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_41
timestamp 1636986456
transform 1 0 8648 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_53
timestamp 1636986456
transform 1 0 9752 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_65
timestamp 1636986456
transform 1 0 10856 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_77
timestamp 18001
transform 1 0 11960 0 1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_83
timestamp 18001
transform 1 0 12512 0 1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_85
timestamp 1636986456
transform 1 0 12696 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_97
timestamp 1636986456
transform 1 0 13800 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_109
timestamp 1636986456
transform 1 0 14904 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_121
timestamp 1636986456
transform 1 0 16008 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_133
timestamp 18001
transform 1 0 17112 0 1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_139
timestamp 18001
transform 1 0 17664 0 1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_141
timestamp 1636986456
transform 1 0 17848 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_153
timestamp 1636986456
transform 1 0 18952 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_165
timestamp 1636986456
transform 1 0 20056 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_177
timestamp 1636986456
transform 1 0 21160 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_189
timestamp 18001
transform 1 0 22264 0 1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_195
timestamp 18001
transform 1 0 22816 0 1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_197
timestamp 1636986456
transform 1 0 23000 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_209
timestamp 1636986456
transform 1 0 24104 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_221
timestamp 1636986456
transform 1 0 25208 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_233
timestamp 1636986456
transform 1 0 26312 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_245
timestamp 18001
transform 1 0 27416 0 1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_251
timestamp 18001
transform 1 0 27968 0 1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_253
timestamp 1636986456
transform 1 0 28152 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_265
timestamp 1636986456
transform 1 0 29256 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_277
timestamp 1636986456
transform 1 0 30360 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_289
timestamp 1636986456
transform 1 0 31464 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_301
timestamp 18001
transform 1 0 32568 0 1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_307
timestamp 18001
transform 1 0 33120 0 1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_309
timestamp 1636986456
transform 1 0 33304 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_321
timestamp 1636986456
transform 1 0 34408 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_333
timestamp 1636986456
transform 1 0 35512 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_345
timestamp 1636986456
transform 1 0 36616 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_357
timestamp 18001
transform 1 0 37720 0 1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_363
timestamp 18001
transform 1 0 38272 0 1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_365
timestamp 1636986456
transform 1 0 38456 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_377
timestamp 1636986456
transform 1 0 39560 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_389
timestamp 1636986456
transform 1 0 40664 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_401
timestamp 1636986456
transform 1 0 41768 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_413
timestamp 18001
transform 1 0 42872 0 1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_419
timestamp 18001
transform 1 0 43424 0 1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_421
timestamp 1636986456
transform 1 0 43608 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_433
timestamp 1636986456
transform 1 0 44712 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_445
timestamp 1636986456
transform 1 0 45816 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_457
timestamp 1636986456
transform 1 0 46920 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_469
timestamp 18001
transform 1 0 48024 0 1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_475
timestamp 18001
transform 1 0 48576 0 1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_477
timestamp 1636986456
transform 1 0 48760 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_489
timestamp 1636986456
transform 1 0 49864 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_501
timestamp 1636986456
transform 1 0 50968 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_513
timestamp 1636986456
transform 1 0 52072 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_525
timestamp 18001
transform 1 0 53176 0 1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_531
timestamp 18001
transform 1 0 53728 0 1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_533
timestamp 1636986456
transform 1 0 53912 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_545
timestamp 1636986456
transform 1 0 55016 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_557
timestamp 1636986456
transform 1 0 56120 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_569
timestamp 1636986456
transform 1 0 57224 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_581
timestamp 18001
transform 1 0 58328 0 1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_587
timestamp 18001
transform 1 0 58880 0 1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_589
timestamp 1636986456
transform 1 0 59064 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_601
timestamp 1636986456
transform 1 0 60168 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_613
timestamp 1636986456
transform 1 0 61272 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_625
timestamp 1636986456
transform 1 0 62376 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_637
timestamp 18001
transform 1 0 63480 0 1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_643
timestamp 18001
transform 1 0 64032 0 1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_645
timestamp 1636986456
transform 1 0 64216 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_657
timestamp 1636986456
transform 1 0 65320 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_669
timestamp 1636986456
transform 1 0 66424 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_681
timestamp 1636986456
transform 1 0 67528 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_693
timestamp 18001
transform 1 0 68632 0 1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_699
timestamp 18001
transform 1 0 69184 0 1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_701
timestamp 1636986456
transform 1 0 69368 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_713
timestamp 1636986456
transform 1 0 70472 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_725
timestamp 1636986456
transform 1 0 71576 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_737
timestamp 1636986456
transform 1 0 72680 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_749
timestamp 18001
transform 1 0 73784 0 1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_755
timestamp 18001
transform 1 0 74336 0 1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_757
timestamp 1636986456
transform 1 0 74520 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_769
timestamp 1636986456
transform 1 0 75624 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_781
timestamp 1636986456
transform 1 0 76728 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_793
timestamp 1636986456
transform 1 0 77832 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_805
timestamp 18001
transform 1 0 78936 0 1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_811
timestamp 18001
transform 1 0 79488 0 1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_813
timestamp 1636986456
transform 1 0 79672 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_825
timestamp 1636986456
transform 1 0 80776 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_837
timestamp 1636986456
transform 1 0 81880 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_849
timestamp 1636986456
transform 1 0 82984 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_861
timestamp 18001
transform 1 0 84088 0 1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_867
timestamp 18001
transform 1 0 84640 0 1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_869
timestamp 1636986456
transform 1 0 84824 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_881
timestamp 1636986456
transform 1 0 85928 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_893
timestamp 1636986456
transform 1 0 87032 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_148_905
timestamp 18001
transform 1 0 88136 0 1 85408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_149_3
timestamp 1636986456
transform 1 0 5152 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_15
timestamp 1636986456
transform 1 0 6256 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_27
timestamp 1636986456
transform 1 0 7360 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_39
timestamp 1636986456
transform 1 0 8464 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_149_51
timestamp 18001
transform 1 0 9568 0 -1 86496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_149_55
timestamp 18001
transform 1 0 9936 0 -1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_57
timestamp 1636986456
transform 1 0 10120 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_69
timestamp 1636986456
transform 1 0 11224 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_81
timestamp 1636986456
transform 1 0 12328 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_93
timestamp 1636986456
transform 1 0 13432 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_105
timestamp 18001
transform 1 0 14536 0 -1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_111
timestamp 18001
transform 1 0 15088 0 -1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_113
timestamp 1636986456
transform 1 0 15272 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_125
timestamp 1636986456
transform 1 0 16376 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_137
timestamp 1636986456
transform 1 0 17480 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_149
timestamp 1636986456
transform 1 0 18584 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_161
timestamp 18001
transform 1 0 19688 0 -1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_167
timestamp 18001
transform 1 0 20240 0 -1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_169
timestamp 1636986456
transform 1 0 20424 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_181
timestamp 1636986456
transform 1 0 21528 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_193
timestamp 1636986456
transform 1 0 22632 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_205
timestamp 1636986456
transform 1 0 23736 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_217
timestamp 18001
transform 1 0 24840 0 -1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_223
timestamp 18001
transform 1 0 25392 0 -1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_225
timestamp 1636986456
transform 1 0 25576 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_237
timestamp 1636986456
transform 1 0 26680 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_249
timestamp 1636986456
transform 1 0 27784 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_261
timestamp 1636986456
transform 1 0 28888 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_273
timestamp 18001
transform 1 0 29992 0 -1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_279
timestamp 18001
transform 1 0 30544 0 -1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_281
timestamp 1636986456
transform 1 0 30728 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_293
timestamp 1636986456
transform 1 0 31832 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_305
timestamp 1636986456
transform 1 0 32936 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_317
timestamp 1636986456
transform 1 0 34040 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_329
timestamp 18001
transform 1 0 35144 0 -1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_335
timestamp 18001
transform 1 0 35696 0 -1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_337
timestamp 1636986456
transform 1 0 35880 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_349
timestamp 1636986456
transform 1 0 36984 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_361
timestamp 1636986456
transform 1 0 38088 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_373
timestamp 1636986456
transform 1 0 39192 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_385
timestamp 18001
transform 1 0 40296 0 -1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_391
timestamp 18001
transform 1 0 40848 0 -1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_393
timestamp 1636986456
transform 1 0 41032 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_405
timestamp 1636986456
transform 1 0 42136 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_417
timestamp 1636986456
transform 1 0 43240 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_429
timestamp 1636986456
transform 1 0 44344 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_441
timestamp 18001
transform 1 0 45448 0 -1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_447
timestamp 18001
transform 1 0 46000 0 -1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_449
timestamp 1636986456
transform 1 0 46184 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_461
timestamp 1636986456
transform 1 0 47288 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_473
timestamp 1636986456
transform 1 0 48392 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_485
timestamp 1636986456
transform 1 0 49496 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_497
timestamp 18001
transform 1 0 50600 0 -1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_503
timestamp 18001
transform 1 0 51152 0 -1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_505
timestamp 1636986456
transform 1 0 51336 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_517
timestamp 1636986456
transform 1 0 52440 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_529
timestamp 1636986456
transform 1 0 53544 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_541
timestamp 1636986456
transform 1 0 54648 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_553
timestamp 18001
transform 1 0 55752 0 -1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_559
timestamp 18001
transform 1 0 56304 0 -1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_561
timestamp 1636986456
transform 1 0 56488 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_573
timestamp 1636986456
transform 1 0 57592 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_585
timestamp 1636986456
transform 1 0 58696 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_597
timestamp 1636986456
transform 1 0 59800 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_609
timestamp 18001
transform 1 0 60904 0 -1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_615
timestamp 18001
transform 1 0 61456 0 -1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_617
timestamp 1636986456
transform 1 0 61640 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_629
timestamp 1636986456
transform 1 0 62744 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_641
timestamp 1636986456
transform 1 0 63848 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_653
timestamp 1636986456
transform 1 0 64952 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_665
timestamp 18001
transform 1 0 66056 0 -1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_671
timestamp 18001
transform 1 0 66608 0 -1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_673
timestamp 1636986456
transform 1 0 66792 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_685
timestamp 1636986456
transform 1 0 67896 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_697
timestamp 1636986456
transform 1 0 69000 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_709
timestamp 1636986456
transform 1 0 70104 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_721
timestamp 18001
transform 1 0 71208 0 -1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_727
timestamp 18001
transform 1 0 71760 0 -1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_729
timestamp 1636986456
transform 1 0 71944 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_741
timestamp 1636986456
transform 1 0 73048 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_753
timestamp 1636986456
transform 1 0 74152 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_765
timestamp 1636986456
transform 1 0 75256 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_777
timestamp 18001
transform 1 0 76360 0 -1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_783
timestamp 18001
transform 1 0 76912 0 -1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_785
timestamp 1636986456
transform 1 0 77096 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_797
timestamp 1636986456
transform 1 0 78200 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_809
timestamp 1636986456
transform 1 0 79304 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_821
timestamp 1636986456
transform 1 0 80408 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_833
timestamp 18001
transform 1 0 81512 0 -1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_839
timestamp 18001
transform 1 0 82064 0 -1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_841
timestamp 1636986456
transform 1 0 82248 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_853
timestamp 1636986456
transform 1 0 83352 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_865
timestamp 1636986456
transform 1 0 84456 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_877
timestamp 1636986456
transform 1 0 85560 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_889
timestamp 18001
transform 1 0 86664 0 -1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_895
timestamp 18001
transform 1 0 87216 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_149_897
timestamp 18001
transform 1 0 87400 0 -1 86496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_149_905
timestamp 18001
transform 1 0 88136 0 -1 86496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_150_3
timestamp 1636986456
transform 1 0 5152 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_15
timestamp 1636986456
transform 1 0 6256 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_150_27
timestamp 18001
transform 1 0 7360 0 1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_29
timestamp 1636986456
transform 1 0 7544 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_41
timestamp 1636986456
transform 1 0 8648 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_53
timestamp 1636986456
transform 1 0 9752 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_65
timestamp 1636986456
transform 1 0 10856 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_77
timestamp 18001
transform 1 0 11960 0 1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_83
timestamp 18001
transform 1 0 12512 0 1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_85
timestamp 1636986456
transform 1 0 12696 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_97
timestamp 1636986456
transform 1 0 13800 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_109
timestamp 1636986456
transform 1 0 14904 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_121
timestamp 1636986456
transform 1 0 16008 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_133
timestamp 18001
transform 1 0 17112 0 1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_139
timestamp 18001
transform 1 0 17664 0 1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_141
timestamp 1636986456
transform 1 0 17848 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_153
timestamp 1636986456
transform 1 0 18952 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_165
timestamp 1636986456
transform 1 0 20056 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_177
timestamp 1636986456
transform 1 0 21160 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_189
timestamp 18001
transform 1 0 22264 0 1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_195
timestamp 18001
transform 1 0 22816 0 1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_197
timestamp 1636986456
transform 1 0 23000 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_209
timestamp 1636986456
transform 1 0 24104 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_221
timestamp 1636986456
transform 1 0 25208 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_233
timestamp 1636986456
transform 1 0 26312 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_245
timestamp 18001
transform 1 0 27416 0 1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_251
timestamp 18001
transform 1 0 27968 0 1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_253
timestamp 1636986456
transform 1 0 28152 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_265
timestamp 1636986456
transform 1 0 29256 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_277
timestamp 1636986456
transform 1 0 30360 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_289
timestamp 1636986456
transform 1 0 31464 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_301
timestamp 18001
transform 1 0 32568 0 1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_307
timestamp 18001
transform 1 0 33120 0 1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_309
timestamp 1636986456
transform 1 0 33304 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_321
timestamp 1636986456
transform 1 0 34408 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_333
timestamp 1636986456
transform 1 0 35512 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_345
timestamp 1636986456
transform 1 0 36616 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_357
timestamp 18001
transform 1 0 37720 0 1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_363
timestamp 18001
transform 1 0 38272 0 1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_365
timestamp 1636986456
transform 1 0 38456 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_377
timestamp 1636986456
transform 1 0 39560 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_150_389
timestamp 18001
transform 1 0 40664 0 1 86496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_150_397
timestamp 18001
transform 1 0 41400 0 1 86496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_150_403
timestamp 1636986456
transform 1 0 41952 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_150_415
timestamp 18001
transform 1 0 43056 0 1 86496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_150_419
timestamp 18001
transform 1 0 43424 0 1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_421
timestamp 1636986456
transform 1 0 43608 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_433
timestamp 1636986456
transform 1 0 44712 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_445
timestamp 1636986456
transform 1 0 45816 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_457
timestamp 1636986456
transform 1 0 46920 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_469
timestamp 18001
transform 1 0 48024 0 1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_475
timestamp 18001
transform 1 0 48576 0 1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_477
timestamp 1636986456
transform 1 0 48760 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_489
timestamp 1636986456
transform 1 0 49864 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_501
timestamp 1636986456
transform 1 0 50968 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_513
timestamp 1636986456
transform 1 0 52072 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_525
timestamp 18001
transform 1 0 53176 0 1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_531
timestamp 18001
transform 1 0 53728 0 1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_533
timestamp 1636986456
transform 1 0 53912 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_545
timestamp 1636986456
transform 1 0 55016 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_557
timestamp 1636986456
transform 1 0 56120 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_569
timestamp 1636986456
transform 1 0 57224 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_581
timestamp 18001
transform 1 0 58328 0 1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_587
timestamp 18001
transform 1 0 58880 0 1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_589
timestamp 1636986456
transform 1 0 59064 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_601
timestamp 1636986456
transform 1 0 60168 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_613
timestamp 1636986456
transform 1 0 61272 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_625
timestamp 1636986456
transform 1 0 62376 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_637
timestamp 18001
transform 1 0 63480 0 1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_643
timestamp 18001
transform 1 0 64032 0 1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_645
timestamp 1636986456
transform 1 0 64216 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_657
timestamp 1636986456
transform 1 0 65320 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_669
timestamp 1636986456
transform 1 0 66424 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_681
timestamp 1636986456
transform 1 0 67528 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_693
timestamp 18001
transform 1 0 68632 0 1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_699
timestamp 18001
transform 1 0 69184 0 1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_701
timestamp 1636986456
transform 1 0 69368 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_713
timestamp 1636986456
transform 1 0 70472 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_725
timestamp 1636986456
transform 1 0 71576 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_737
timestamp 1636986456
transform 1 0 72680 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_749
timestamp 18001
transform 1 0 73784 0 1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_755
timestamp 18001
transform 1 0 74336 0 1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_757
timestamp 1636986456
transform 1 0 74520 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_769
timestamp 1636986456
transform 1 0 75624 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_781
timestamp 1636986456
transform 1 0 76728 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_793
timestamp 1636986456
transform 1 0 77832 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_805
timestamp 18001
transform 1 0 78936 0 1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_811
timestamp 18001
transform 1 0 79488 0 1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_813
timestamp 1636986456
transform 1 0 79672 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_825
timestamp 1636986456
transform 1 0 80776 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_837
timestamp 1636986456
transform 1 0 81880 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_849
timestamp 1636986456
transform 1 0 82984 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_861
timestamp 18001
transform 1 0 84088 0 1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_867
timestamp 18001
transform 1 0 84640 0 1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_869
timestamp 1636986456
transform 1 0 84824 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_881
timestamp 1636986456
transform 1 0 85928 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_893
timestamp 1636986456
transform 1 0 87032 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_150_905
timestamp 18001
transform 1 0 88136 0 1 86496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_151_3
timestamp 1636986456
transform 1 0 5152 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_15
timestamp 1636986456
transform 1 0 6256 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_151_27
timestamp 18001
transform 1 0 7360 0 -1 87584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_151_29
timestamp 1636986456
transform 1 0 7544 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_41
timestamp 1636986456
transform 1 0 8648 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_151_53
timestamp 18001
transform 1 0 9752 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_151_57
timestamp 18001
transform 1 0 10120 0 -1 87584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_151_67
timestamp 1636986456
transform 1 0 11040 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_151_79
timestamp 18001
transform 1 0 12144 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_151_83
timestamp 18001
transform 1 0 12512 0 -1 87584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_151_85
timestamp 1636986456
transform 1 0 12696 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_97
timestamp 1636986456
transform 1 0 13800 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_151_109
timestamp 18001
transform 1 0 14904 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_151_128
timestamp 18001
transform 1 0 16652 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_151_136
timestamp 18001
transform 1 0 17388 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_151_141
timestamp 18001
transform 1 0 17848 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_151_150
timestamp 18001
transform 1 0 18676 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_151_158
timestamp 18001
transform 1 0 19412 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_151_164
timestamp 18001
transform 1 0 19964 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_151_174
timestamp 18001
transform 1 0 20884 0 -1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_151_185
timestamp 18001
transform 1 0 21896 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_151_193
timestamp 18001
transform 1 0 22632 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_151_200
timestamp 18001
transform 1 0 23276 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_151_206
timestamp 18001
transform 1 0 23828 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_151_214
timestamp 18001
transform 1 0 24564 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_151_220
timestamp 18001
transform 1 0 25116 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_151_225
timestamp 18001
transform 1 0 25576 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_151_234
timestamp 18001
transform 1 0 26404 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_151_242
timestamp 18001
transform 1 0 27140 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_151_248
timestamp 18001
transform 1 0 27692 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_151_258
timestamp 18001
transform 1 0 28612 0 -1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_151_269
timestamp 18001
transform 1 0 29624 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_151_277
timestamp 18001
transform 1 0 30360 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_151_285
timestamp 18001
transform 1 0 31096 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_151_291
timestamp 18001
transform 1 0 31648 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_151_299
timestamp 18001
transform 1 0 32384 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_151_305
timestamp 18001
transform 1 0 32936 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_151_309
timestamp 18001
transform 1 0 33304 0 -1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_151_319
timestamp 18001
transform 1 0 34224 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_151_327
timestamp 18001
transform 1 0 34960 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_151_333
timestamp 18001
transform 1 0 35512 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_151_341
timestamp 18001
transform 1 0 36248 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_151_349
timestamp 18001
transform 1 0 36984 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_151_354
timestamp 18001
transform 1 0 37444 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_151_382
timestamp 18001
transform 1 0 40020 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_151_389
timestamp 18001
transform 1 0 40664 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_151_410
timestamp 18001
transform 1 0 42596 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_151_416
timestamp 18001
transform 1 0 43148 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_151_425
timestamp 18001
transform 1 0 43976 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_151_431
timestamp 18001
transform 1 0 44528 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_151_437
timestamp 18001
transform 1 0 45080 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_151_444
timestamp 18001
transform 1 0 45724 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_151_452
timestamp 18001
transform 1 0 46460 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_151_458
timestamp 18001
transform 1 0 47012 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_151_465
timestamp 18001
transform 1 0 47656 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_151_472
timestamp 18001
transform 1 0 48300 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_151_480
timestamp 18001
transform 1 0 49036 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_151_486
timestamp 18001
transform 1 0 49588 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_151_493
timestamp 18001
transform 1 0 50232 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_151_500
timestamp 18001
transform 1 0 50876 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_151_505
timestamp 18001
transform 1 0 51336 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_151_513
timestamp 18001
transform 1 0 52072 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_151_528
timestamp 18001
transform 1 0 53452 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_151_538
timestamp 18001
transform 1 0 54372 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_151_544
timestamp 18001
transform 1 0 54924 0 -1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_550
timestamp 18001
transform 1 0 55476 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_151_556
timestamp 18001
transform 1 0 56028 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_151_561
timestamp 18001
transform 1 0 56488 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_151_570
timestamp 18001
transform 1 0 57316 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_151_577
timestamp 18001
transform 1 0 57960 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_151_585
timestamp 18001
transform 1 0 58696 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_151_594
timestamp 18001
transform 1 0 59524 0 -1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_151_605
timestamp 18001
transform 1 0 60536 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_151_613
timestamp 18001
transform 1 0 61272 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_151_622
timestamp 18001
transform 1 0 62100 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_151_628
timestamp 18001
transform 1 0 62652 0 -1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_634
timestamp 18001
transform 1 0 63204 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_151_640
timestamp 18001
transform 1 0 63756 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_151_645
timestamp 18001
transform 1 0 64216 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_151_654
timestamp 18001
transform 1 0 65044 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_151_661
timestamp 18001
transform 1 0 65688 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_151_669
timestamp 18001
transform 1 0 66424 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_151_678
timestamp 18001
transform 1 0 67252 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_151_690
timestamp 18001
transform 1 0 68356 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_151_698
timestamp 18001
transform 1 0 69092 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_151_705
timestamp 18001
transform 1 0 69736 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_151_711
timestamp 18001
transform 1 0 70288 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_151_719
timestamp 18001
transform 1 0 71024 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_151_725
timestamp 18001
transform 1 0 71576 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_151_729
timestamp 18001
transform 1 0 71944 0 -1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_151_739
timestamp 18001
transform 1 0 72864 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_151_746
timestamp 18001
transform 1 0 73508 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_151_754
timestamp 18001
transform 1 0 74244 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_151_761
timestamp 18001
transform 1 0 74888 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_151_769
timestamp 18001
transform 1 0 75624 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_151_774
timestamp 18001
transform 1 0 76084 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_151_782
timestamp 18001
transform 1 0 76820 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_151_789
timestamp 18001
transform 1 0 77464 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_151_795
timestamp 18001
transform 1 0 78016 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_151_803
timestamp 18001
transform 1 0 78752 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_151_809
timestamp 18001
transform 1 0 79304 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_151_813
timestamp 18001
transform 1 0 79672 0 -1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_151_823
timestamp 18001
transform 1 0 80592 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_151_830
timestamp 18001
transform 1 0 81236 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_151_838
timestamp 18001
transform 1 0 81972 0 -1 87584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_151_845
timestamp 1636986456
transform 1 0 82616 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_151_857
timestamp 18001
transform 1 0 83720 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_151_865
timestamp 18001
transform 1 0 84456 0 -1 87584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_151_869
timestamp 1636986456
transform 1 0 84824 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_881
timestamp 1636986456
transform 1 0 85928 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_151_893
timestamp 18001
transform 1 0 87032 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_151_897
timestamp 18001
transform 1 0 87400 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_151_905
timestamp 18001
transform 1 0 88136 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  fpga_232
timestamp 18001
transform -1 0 50876 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_233
timestamp 18001
transform -1 0 50232 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_234
timestamp 18001
transform -1 0 47656 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_235
timestamp 18001
transform -1 0 43148 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_236
timestamp 18001
transform -1 0 49036 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_237
timestamp 18001
transform 1 0 88044 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_238
timestamp 18001
transform 1 0 88044 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_239
timestamp 18001
transform -1 0 45080 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_240
timestamp 18001
transform -1 0 45724 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_241
timestamp 18001
transform -1 0 47012 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_242
timestamp 18001
transform 1 0 88044 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_243
timestamp 18001
transform 1 0 88044 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_244
timestamp 18001
transform -1 0 46460 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_245
timestamp 18001
transform 1 0 88044 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_246
timestamp 18001
transform -1 0 49588 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_247
timestamp 18001
transform -1 0 48300 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 18001
transform 1 0 5152 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  input2
timestamp 18001
transform 1 0 38456 0 -1 87584
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 18001
transform -1 0 88320 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 18001
transform 1 0 88044 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 18001
transform 1 0 88044 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 18001
transform 1 0 88044 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 18001
transform 1 0 88044 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 18001
transform -1 0 88320 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 18001
transform 1 0 88044 0 -1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 18001
transform -1 0 88320 0 1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 18001
transform 1 0 88044 0 1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 18001
transform 1 0 88044 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 18001
transform 1 0 88044 0 1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 18001
transform -1 0 88320 0 1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 18001
transform -1 0 88320 0 -1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input16
timestamp 18001
transform -1 0 88320 0 1 74528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input17
timestamp 18001
transform -1 0 88320 0 1 75616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input18
timestamp 18001
transform -1 0 87860 0 1 76704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 18001
transform 1 0 88044 0 1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 18001
transform 1 0 88044 0 -1 78880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 18001
transform 1 0 88044 0 1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 18001
transform 1 0 88044 0 1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input23
timestamp 18001
transform -1 0 88320 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 18001
transform 1 0 88044 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input25
timestamp 18001
transform -1 0 88320 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input26
timestamp 18001
transform -1 0 88320 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input27
timestamp 18001
transform -1 0 88320 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input28
timestamp 18001
transform -1 0 88320 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input29
timestamp 18001
transform -1 0 88320 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input30
timestamp 18001
transform -1 0 88320 0 -1 40800
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input31
timestamp 18001
transform 1 0 15272 0 -1 87584
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 18001
transform 1 0 26128 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input33
timestamp 18001
transform -1 0 27692 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 18001
transform 1 0 28152 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input35
timestamp 18001
transform -1 0 29624 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input36
timestamp 18001
transform 1 0 52532 0 -1 87584
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input37
timestamp 18001
transform -1 0 54188 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input38
timestamp 18001
transform 1 0 54464 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input39
timestamp 18001
transform -1 0 56028 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input40
timestamp 18001
transform -1 0 16468 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input41
timestamp 18001
transform -1 0 57316 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 18001
transform -1 0 57960 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input43
timestamp 18001
transform -1 0 59340 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input44
timestamp 18001
transform -1 0 60536 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 18001
transform 1 0 61640 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input46
timestamp 18001
transform 1 0 62192 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 18001
transform 1 0 63480 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input48
timestamp 18001
transform -1 0 65044 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 18001
transform -1 0 65688 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input50
timestamp 18001
transform -1 0 67068 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input51
timestamp 18001
transform 1 0 17112 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input52
timestamp 18001
transform -1 0 18676 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input53
timestamp 18001
transform -1 0 19964 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 18001
transform 1 0 20424 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input55
timestamp 18001
transform -1 0 21896 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input56
timestamp 18001
transform -1 0 23276 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 18001
transform -1 0 23828 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input58
timestamp 18001
transform 1 0 24840 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 18001
transform 1 0 30728 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 18001
transform 1 0 41584 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 18001
transform 1 0 42872 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 18001
transform 1 0 43608 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 18001
transform 1 0 44804 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 18001
transform 1 0 67988 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input65
timestamp 18001
transform -1 0 69644 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input66
timestamp 18001
transform 1 0 69920 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input67
timestamp 18001
transform -1 0 71484 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input68
timestamp 18001
transform 1 0 31280 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input69
timestamp 18001
transform -1 0 72772 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 18001
transform -1 0 73416 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input71
timestamp 18001
transform -1 0 74796 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input72
timestamp 18001
transform -1 0 75992 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input73
timestamp 18001
transform -1 0 77372 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input74
timestamp 18001
transform 1 0 77648 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input75
timestamp 18001
transform 1 0 78936 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input76
timestamp 18001
transform 1 0 80224 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input77
timestamp 18001
transform 1 0 88044 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input78
timestamp 18001
transform 1 0 88044 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input79
timestamp 18001
transform 1 0 32568 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input80
timestamp 18001
transform -1 0 34132 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input81
timestamp 18001
transform -1 0 35420 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input82
timestamp 18001
transform 1 0 35880 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input83
timestamp 18001
transform -1 0 37352 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input84
timestamp 18001
transform -1 0 38732 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input85
timestamp 18001
transform 1 0 39008 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input86
timestamp 18001
transform 1 0 40296 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input87
timestamp 18001
transform -1 0 5428 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input88
timestamp 18001
transform -1 0 5428 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input89
timestamp 18001
transform -1 0 5428 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input90
timestamp 18001
transform -1 0 5428 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input91
timestamp 18001
transform -1 0 5428 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input92
timestamp 18001
transform -1 0 5428 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input93
timestamp 18001
transform -1 0 5428 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input94
timestamp 18001
transform -1 0 5428 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input95
timestamp 18001
transform -1 0 5428 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input96
timestamp 18001
transform -1 0 5428 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input97
timestamp 18001
transform -1 0 5428 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input98
timestamp 18001
transform -1 0 5428 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input99
timestamp 18001
transform 1 0 5152 0 1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input100
timestamp 18001
transform -1 0 5428 0 1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input101
timestamp 18001
transform 1 0 5152 0 1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input102
timestamp 18001
transform 1 0 5152 0 1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input103
timestamp 18001
transform -1 0 5428 0 -1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input104
timestamp 18001
transform -1 0 5428 0 1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input105
timestamp 18001
transform -1 0 5428 0 1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input106
timestamp 18001
transform -1 0 5428 0 1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input107
timestamp 18001
transform -1 0 5428 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input108
timestamp 18001
transform -1 0 5428 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input109
timestamp 18001
transform -1 0 5428 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input110
timestamp 18001
transform -1 0 5428 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input111
timestamp 18001
transform 1 0 5152 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input112
timestamp 18001
transform -1 0 5428 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input113
timestamp 18001
transform 1 0 5152 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input114
timestamp 18001
transform 1 0 5152 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input115
timestamp 18001
transform -1 0 87860 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input116
timestamp 18001
transform -1 0 88320 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input117
timestamp 18001
transform -1 0 87860 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  input118
timestamp 18001
transform 1 0 41032 0 -1 87584
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_2  output119
timestamp 18001
transform 1 0 87952 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output120
timestamp 18001
transform 1 0 87952 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output121
timestamp 18001
transform 1 0 87952 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output122
timestamp 18001
transform 1 0 87952 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp 18001
transform 1 0 87952 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output124
timestamp 18001
transform 1 0 87952 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output125
timestamp 18001
transform 1 0 87952 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output126
timestamp 18001
transform 1 0 87952 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output127
timestamp 18001
transform 1 0 87952 0 1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output128
timestamp 18001
transform 1 0 87952 0 1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output129
timestamp 18001
transform 1 0 87952 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output130
timestamp 18001
transform 1 0 87952 0 1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output131
timestamp 18001
transform 1 0 87952 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output132
timestamp 18001
transform 1 0 87952 0 1 58208
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output133
timestamp 18001
transform 1 0 87952 0 1 59296
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output134
timestamp 18001
transform 1 0 87952 0 1 60384
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output135
timestamp 18001
transform 1 0 87952 0 1 61472
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output136
timestamp 18001
transform 1 0 87952 0 -1 62560
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output137
timestamp 18001
transform 1 0 87952 0 1 63648
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output138
timestamp 18001
transform 1 0 87952 0 1 64736
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp 18001
transform 1 0 87952 0 1 65824
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output140
timestamp 18001
transform 1 0 87952 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output141
timestamp 18001
transform 1 0 87952 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output142
timestamp 18001
transform 1 0 87952 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output143
timestamp 18001
transform 1 0 87952 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output144
timestamp 18001
transform 1 0 87952 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output145
timestamp 18001
transform 1 0 87952 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output146
timestamp 18001
transform 1 0 87952 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output147
timestamp 18001
transform 1 0 87952 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output148
timestamp 18001
transform 1 0 30728 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output149
timestamp 18001
transform 1 0 41584 0 1 86496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output150
timestamp 18001
transform -1 0 42596 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output151
timestamp 18001
transform 1 0 43608 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output152
timestamp 18001
transform -1 0 44528 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output153
timestamp 18001
transform 1 0 67988 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output154
timestamp 18001
transform 1 0 69368 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output155
timestamp 18001
transform -1 0 70288 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output156
timestamp 18001
transform 1 0 71208 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output157
timestamp 18001
transform -1 0 31648 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output158
timestamp 18001
transform 1 0 72496 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output159
timestamp 18001
transform -1 0 73508 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output160
timestamp 18001
transform 1 0 74520 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output161
timestamp 18001
transform 1 0 75716 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output162
timestamp 18001
transform 1 0 77096 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output163
timestamp 18001
transform -1 0 78016 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output164
timestamp 18001
transform 1 0 78936 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output165
timestamp 18001
transform 1 0 80224 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output166
timestamp 18001
transform -1 0 81236 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output167
timestamp 18001
transform 1 0 82248 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output168
timestamp 18001
transform 1 0 32568 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output169
timestamp 18001
transform 1 0 33856 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output170
timestamp 18001
transform 1 0 35144 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output171
timestamp 18001
transform 1 0 35880 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output172
timestamp 18001
transform 1 0 37076 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output173
timestamp 18001
transform 1 0 37996 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output174
timestamp 18001
transform 1 0 39468 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output175
timestamp 18001
transform 1 0 40296 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output176
timestamp 18001
transform 1 0 15272 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output177
timestamp 18001
transform 1 0 26128 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output178
timestamp 18001
transform 1 0 27416 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output179
timestamp 18001
transform 1 0 28152 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output180
timestamp 18001
transform 1 0 29348 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output181
timestamp 18001
transform 1 0 52532 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output182
timestamp 18001
transform 1 0 53912 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output183
timestamp 18001
transform -1 0 54832 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output184
timestamp 18001
transform 1 0 55752 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output185
timestamp 18001
transform -1 0 16192 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output186
timestamp 18001
transform 1 0 57040 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output187
timestamp 18001
transform -1 0 58052 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output188
timestamp 18001
transform 1 0 59064 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output189
timestamp 18001
transform 1 0 60260 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output190
timestamp 18001
transform 1 0 61640 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output191
timestamp 18001
transform -1 0 62560 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output192
timestamp 18001
transform 1 0 63480 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output193
timestamp 18001
transform 1 0 64768 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output194
timestamp 18001
transform -1 0 65780 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output195
timestamp 18001
transform 1 0 66792 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output196
timestamp 18001
transform 1 0 17112 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output197
timestamp 18001
transform 1 0 18400 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output198
timestamp 18001
transform 1 0 19688 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output199
timestamp 18001
transform 1 0 20424 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output200
timestamp 18001
transform 1 0 21620 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output201
timestamp 18001
transform 1 0 23000 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output202
timestamp 18001
transform -1 0 23920 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output203
timestamp 18001
transform 1 0 24840 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output204
timestamp 18001
transform -1 0 5520 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output205
timestamp 18001
transform -1 0 5520 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output206
timestamp 18001
transform -1 0 5520 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output207
timestamp 18001
transform -1 0 5520 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output208
timestamp 18001
transform -1 0 5520 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output209
timestamp 18001
transform -1 0 5520 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output210
timestamp 18001
transform -1 0 5520 0 -1 68000
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output211
timestamp 18001
transform -1 0 5520 0 1 69088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output212
timestamp 18001
transform -1 0 5520 0 1 70176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output213
timestamp 18001
transform -1 0 5520 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output214
timestamp 18001
transform -1 0 5520 0 1 71264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output215
timestamp 18001
transform -1 0 5520 0 1 72352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output216
timestamp 18001
transform -1 0 5520 0 -1 73440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output217
timestamp 18001
transform -1 0 5520 0 1 74528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output218
timestamp 18001
transform -1 0 5520 0 1 75616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output219
timestamp 18001
transform -1 0 5520 0 1 76704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output220
timestamp 18001
transform -1 0 5520 0 1 77792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output221
timestamp 18001
transform -1 0 5520 0 -1 78880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output222
timestamp 18001
transform -1 0 5520 0 1 79968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output223
timestamp 18001
transform 1 0 10672 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output224
timestamp 18001
transform -1 0 5520 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output225
timestamp 18001
transform -1 0 5520 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output226
timestamp 18001
transform -1 0 5520 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output227
timestamp 18001
transform -1 0 5520 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output228
timestamp 18001
transform -1 0 5520 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output229
timestamp 18001
transform -1 0 5520 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output230
timestamp 18001
transform -1 0 5520 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output231
timestamp 18001
transform -1 0 5520 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_152
timestamp 18001
transform 1 0 4876 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 18001
transform -1 0 88596 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_153
timestamp 18001
transform 1 0 4876 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 18001
transform -1 0 88596 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_154
timestamp 18001
transform 1 0 4876 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 18001
transform -1 0 88596 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_155
timestamp 18001
transform 1 0 4876 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 18001
transform -1 0 88596 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_156
timestamp 18001
transform 1 0 4876 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 18001
transform -1 0 88596 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_1_Left_303
timestamp 18001
transform 1 0 4876 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_1_Right_585
timestamp 18001
transform -1 0 7912 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_3_Left_304
timestamp 18001
transform 1 0 85284 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_3_Right_11
timestamp 18001
transform -1 0 88596 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_1_Left_157
timestamp 18001
transform 1 0 4876 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_1_Right_445
timestamp 18001
transform -1 0 7912 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_3_Left_305
timestamp 18001
transform 1 0 85284 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_3_Right_12
timestamp 18001
transform -1 0 88596 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_1_Left_158
timestamp 18001
transform 1 0 4876 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_1_Right_446
timestamp 18001
transform -1 0 7912 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_3_Left_306
timestamp 18001
transform 1 0 85284 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_3_Right_13
timestamp 18001
transform -1 0 88596 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_1_Left_159
timestamp 18001
transform 1 0 4876 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_1_Right_447
timestamp 18001
transform -1 0 7912 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_3_Left_307
timestamp 18001
transform 1 0 85284 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_3_Right_14
timestamp 18001
transform -1 0 88596 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_1_Left_160
timestamp 18001
transform 1 0 4876 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_1_Right_448
timestamp 18001
transform -1 0 7912 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_3_Left_308
timestamp 18001
transform 1 0 85284 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_3_Right_15
timestamp 18001
transform -1 0 88596 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_1_Left_161
timestamp 18001
transform 1 0 4876 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_1_Right_449
timestamp 18001
transform -1 0 7912 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_3_Left_309
timestamp 18001
transform 1 0 85284 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_3_Right_16
timestamp 18001
transform -1 0 88596 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_1_Left_162
timestamp 18001
transform 1 0 4876 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_1_Right_450
timestamp 18001
transform -1 0 7912 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_3_Left_310
timestamp 18001
transform 1 0 85284 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_3_Right_17
timestamp 18001
transform -1 0 88596 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_1_Left_163
timestamp 18001
transform 1 0 4876 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_1_Right_451
timestamp 18001
transform -1 0 7912 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_3_Left_311
timestamp 18001
transform 1 0 85284 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_3_Right_18
timestamp 18001
transform -1 0 88596 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_1_Left_164
timestamp 18001
transform 1 0 4876 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_1_Right_452
timestamp 18001
transform -1 0 7912 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_3_Left_312
timestamp 18001
transform 1 0 85284 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_3_Right_19
timestamp 18001
transform -1 0 88596 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_1_Left_165
timestamp 18001
transform 1 0 4876 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_1_Right_453
timestamp 18001
transform -1 0 7912 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_3_Left_313
timestamp 18001
transform 1 0 85284 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_3_Right_20
timestamp 18001
transform -1 0 88596 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_1_Left_166
timestamp 18001
transform 1 0 4876 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_1_Right_454
timestamp 18001
transform -1 0 7912 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_3_Left_314
timestamp 18001
transform 1 0 85284 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_3_Right_21
timestamp 18001
transform -1 0 88596 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_1_Left_167
timestamp 18001
transform 1 0 4876 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_1_Right_455
timestamp 18001
transform -1 0 7912 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_3_Left_315
timestamp 18001
transform 1 0 85284 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_3_Right_22
timestamp 18001
transform -1 0 88596 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_1_Left_168
timestamp 18001
transform 1 0 4876 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_1_Right_456
timestamp 18001
transform -1 0 7912 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_3_Left_316
timestamp 18001
transform 1 0 85284 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_3_Right_23
timestamp 18001
transform -1 0 88596 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_1_Left_169
timestamp 18001
transform 1 0 4876 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_1_Right_457
timestamp 18001
transform -1 0 7912 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_3_Left_317
timestamp 18001
transform 1 0 85284 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_3_Right_24
timestamp 18001
transform -1 0 88596 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_1_Left_170
timestamp 18001
transform 1 0 4876 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_1_Right_458
timestamp 18001
transform -1 0 7912 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_3_Left_318
timestamp 18001
transform 1 0 85284 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_3_Right_25
timestamp 18001
transform -1 0 88596 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_1_Left_171
timestamp 18001
transform 1 0 4876 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_1_Right_459
timestamp 18001
transform -1 0 7912 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_3_Left_319
timestamp 18001
transform 1 0 85284 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_3_Right_26
timestamp 18001
transform -1 0 88596 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_1_Left_172
timestamp 18001
transform 1 0 4876 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_1_Right_460
timestamp 18001
transform -1 0 7912 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_3_Left_320
timestamp 18001
transform 1 0 85284 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_3_Right_27
timestamp 18001
transform -1 0 88596 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_1_Left_173
timestamp 18001
transform 1 0 4876 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_1_Right_461
timestamp 18001
transform -1 0 7912 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_3_Left_321
timestamp 18001
transform 1 0 85284 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_3_Right_28
timestamp 18001
transform -1 0 88596 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_1_Left_174
timestamp 18001
transform 1 0 4876 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_1_Right_462
timestamp 18001
transform -1 0 7912 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_3_Left_322
timestamp 18001
transform 1 0 85284 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_3_Right_29
timestamp 18001
transform -1 0 88596 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_1_Left_175
timestamp 18001
transform 1 0 4876 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_1_Right_463
timestamp 18001
transform -1 0 7912 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_3_Left_323
timestamp 18001
transform 1 0 85284 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_3_Right_30
timestamp 18001
transform -1 0 88596 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_1_Left_176
timestamp 18001
transform 1 0 4876 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_1_Right_464
timestamp 18001
transform -1 0 7912 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_3_Left_324
timestamp 18001
transform 1 0 85284 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_3_Right_31
timestamp 18001
transform -1 0 88596 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_1_Left_177
timestamp 18001
transform 1 0 4876 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_1_Right_465
timestamp 18001
transform -1 0 7912 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_3_Left_325
timestamp 18001
transform 1 0 85284 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_3_Right_32
timestamp 18001
transform -1 0 88596 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_1_Left_178
timestamp 18001
transform 1 0 4876 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_1_Right_466
timestamp 18001
transform -1 0 7912 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_3_Left_326
timestamp 18001
transform 1 0 85284 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_3_Right_33
timestamp 18001
transform -1 0 88596 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_1_Left_179
timestamp 18001
transform 1 0 4876 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_1_Right_467
timestamp 18001
transform -1 0 7912 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_3_Left_327
timestamp 18001
transform 1 0 85284 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_3_Right_34
timestamp 18001
transform -1 0 88596 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_1_Left_180
timestamp 18001
transform 1 0 4876 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_1_Right_468
timestamp 18001
transform -1 0 7912 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_3_Left_328
timestamp 18001
transform 1 0 85284 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_3_Right_35
timestamp 18001
transform -1 0 88596 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_1_Left_181
timestamp 18001
transform 1 0 4876 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_1_Right_469
timestamp 18001
transform -1 0 7912 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_3_Left_329
timestamp 18001
transform 1 0 85284 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_3_Right_36
timestamp 18001
transform -1 0 88596 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_1_Left_182
timestamp 18001
transform 1 0 4876 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_1_Right_470
timestamp 18001
transform -1 0 7912 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_3_Left_330
timestamp 18001
transform 1 0 85284 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_3_Right_37
timestamp 18001
transform -1 0 88596 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_1_Left_183
timestamp 18001
transform 1 0 4876 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_1_Right_471
timestamp 18001
transform -1 0 7912 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_3_Left_331
timestamp 18001
transform 1 0 85284 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_3_Right_38
timestamp 18001
transform -1 0 88596 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_1_Left_184
timestamp 18001
transform 1 0 4876 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_1_Right_472
timestamp 18001
transform -1 0 7912 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_3_Left_332
timestamp 18001
transform 1 0 85284 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_3_Right_39
timestamp 18001
transform -1 0 88596 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_1_Left_185
timestamp 18001
transform 1 0 4876 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_1_Right_473
timestamp 18001
transform -1 0 7912 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_3_Left_333
timestamp 18001
transform 1 0 85284 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_3_Right_40
timestamp 18001
transform -1 0 88596 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_1_Left_186
timestamp 18001
transform 1 0 4876 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_1_Right_474
timestamp 18001
transform -1 0 7912 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_3_Left_334
timestamp 18001
transform 1 0 85284 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_3_Right_41
timestamp 18001
transform -1 0 88596 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_1_Left_187
timestamp 18001
transform 1 0 4876 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_1_Right_475
timestamp 18001
transform -1 0 7912 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_3_Left_335
timestamp 18001
transform 1 0 85284 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_3_Right_42
timestamp 18001
transform -1 0 88596 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_1_Left_188
timestamp 18001
transform 1 0 4876 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_1_Right_476
timestamp 18001
transform -1 0 7912 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_3_Left_336
timestamp 18001
transform 1 0 85284 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_3_Right_43
timestamp 18001
transform -1 0 88596 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_1_Left_189
timestamp 18001
transform 1 0 4876 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_1_Right_477
timestamp 18001
transform -1 0 7912 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_3_Left_337
timestamp 18001
transform 1 0 85284 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_3_Right_44
timestamp 18001
transform -1 0 88596 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_1_Left_190
timestamp 18001
transform 1 0 4876 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_1_Right_478
timestamp 18001
transform -1 0 7912 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_3_Left_338
timestamp 18001
transform 1 0 85284 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_3_Right_45
timestamp 18001
transform -1 0 88596 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_1_Left_191
timestamp 18001
transform 1 0 4876 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_1_Right_479
timestamp 18001
transform -1 0 7912 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_3_Left_339
timestamp 18001
transform 1 0 85284 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_3_Right_46
timestamp 18001
transform -1 0 88596 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_1_Left_192
timestamp 18001
transform 1 0 4876 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_1_Right_480
timestamp 18001
transform -1 0 7912 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_3_Left_340
timestamp 18001
transform 1 0 85284 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_3_Right_47
timestamp 18001
transform -1 0 88596 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_1_Left_193
timestamp 18001
transform 1 0 4876 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_1_Right_481
timestamp 18001
transform -1 0 7912 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_3_Left_341
timestamp 18001
transform 1 0 85284 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_3_Right_48
timestamp 18001
transform -1 0 88596 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_1_Left_194
timestamp 18001
transform 1 0 4876 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_1_Right_482
timestamp 18001
transform -1 0 7912 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_3_Left_342
timestamp 18001
transform 1 0 85284 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_3_Right_49
timestamp 18001
transform -1 0 88596 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_1_Left_195
timestamp 18001
transform 1 0 4876 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_1_Right_483
timestamp 18001
transform -1 0 7912 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_3_Left_343
timestamp 18001
transform 1 0 85284 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_3_Right_50
timestamp 18001
transform -1 0 88596 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_1_Left_196
timestamp 18001
transform 1 0 4876 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_1_Right_484
timestamp 18001
transform -1 0 7912 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_3_Left_344
timestamp 18001
transform 1 0 85284 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_3_Right_51
timestamp 18001
transform -1 0 88596 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_1_Left_197
timestamp 18001
transform 1 0 4876 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_1_Right_485
timestamp 18001
transform -1 0 7912 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_3_Left_345
timestamp 18001
transform 1 0 85284 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_3_Right_52
timestamp 18001
transform -1 0 88596 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_1_Left_198
timestamp 18001
transform 1 0 4876 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_1_Right_486
timestamp 18001
transform -1 0 7912 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_3_Left_346
timestamp 18001
transform 1 0 85284 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_3_Right_53
timestamp 18001
transform -1 0 88596 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_1_Left_199
timestamp 18001
transform 1 0 4876 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_1_Right_487
timestamp 18001
transform -1 0 7912 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_3_Left_347
timestamp 18001
transform 1 0 85284 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_3_Right_54
timestamp 18001
transform -1 0 88596 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_1_Left_200
timestamp 18001
transform 1 0 4876 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_1_Right_488
timestamp 18001
transform -1 0 7912 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_3_Left_348
timestamp 18001
transform 1 0 85284 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_3_Right_55
timestamp 18001
transform -1 0 88596 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_1_Left_201
timestamp 18001
transform 1 0 4876 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_1_Right_489
timestamp 18001
transform -1 0 7912 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_3_Left_349
timestamp 18001
transform 1 0 85284 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_3_Right_56
timestamp 18001
transform -1 0 88596 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_1_Left_202
timestamp 18001
transform 1 0 4876 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_1_Right_490
timestamp 18001
transform -1 0 7912 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_3_Left_350
timestamp 18001
transform 1 0 85284 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_3_Right_57
timestamp 18001
transform -1 0 88596 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_1_Left_203
timestamp 18001
transform 1 0 4876 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_1_Right_491
timestamp 18001
transform -1 0 7912 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_3_Left_351
timestamp 18001
transform 1 0 85284 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_3_Right_58
timestamp 18001
transform -1 0 88596 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_1_Left_204
timestamp 18001
transform 1 0 4876 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_1_Right_492
timestamp 18001
transform -1 0 7912 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_3_Left_352
timestamp 18001
transform 1 0 85284 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_3_Right_59
timestamp 18001
transform -1 0 88596 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_1_Left_205
timestamp 18001
transform 1 0 4876 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_1_Right_493
timestamp 18001
transform -1 0 7912 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_3_Left_353
timestamp 18001
transform 1 0 85284 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_3_Right_60
timestamp 18001
transform -1 0 88596 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_1_Left_206
timestamp 18001
transform 1 0 4876 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_1_Right_494
timestamp 18001
transform -1 0 7912 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_3_Left_354
timestamp 18001
transform 1 0 85284 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_3_Right_61
timestamp 18001
transform -1 0 88596 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_1_Left_207
timestamp 18001
transform 1 0 4876 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_1_Right_495
timestamp 18001
transform -1 0 7912 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_3_Left_355
timestamp 18001
transform 1 0 85284 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_3_Right_62
timestamp 18001
transform -1 0 88596 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_1_Left_208
timestamp 18001
transform 1 0 4876 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_1_Right_496
timestamp 18001
transform -1 0 7912 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_3_Left_356
timestamp 18001
transform 1 0 85284 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_3_Right_63
timestamp 18001
transform -1 0 88596 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_1_Left_209
timestamp 18001
transform 1 0 4876 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_1_Right_497
timestamp 18001
transform -1 0 7912 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_3_Left_357
timestamp 18001
transform 1 0 85284 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_3_Right_64
timestamp 18001
transform -1 0 88596 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_1_Left_210
timestamp 18001
transform 1 0 4876 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_1_Right_498
timestamp 18001
transform -1 0 7912 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_3_Left_358
timestamp 18001
transform 1 0 85284 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_3_Right_65
timestamp 18001
transform -1 0 88596 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_1_Left_211
timestamp 18001
transform 1 0 4876 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_1_Right_499
timestamp 18001
transform -1 0 7912 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_3_Left_359
timestamp 18001
transform 1 0 85284 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_3_Right_66
timestamp 18001
transform -1 0 88596 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_1_Left_212
timestamp 18001
transform 1 0 4876 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_1_Right_500
timestamp 18001
transform -1 0 7912 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_3_Left_360
timestamp 18001
transform 1 0 85284 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_3_Right_67
timestamp 18001
transform -1 0 88596 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_1_Left_213
timestamp 18001
transform 1 0 4876 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_1_Right_501
timestamp 18001
transform -1 0 7912 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_3_Left_361
timestamp 18001
transform 1 0 85284 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_3_Right_68
timestamp 18001
transform -1 0 88596 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_1_Left_214
timestamp 18001
transform 1 0 4876 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_1_Right_502
timestamp 18001
transform -1 0 7912 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_3_Left_362
timestamp 18001
transform 1 0 85284 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_3_Right_69
timestamp 18001
transform -1 0 88596 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_1_Left_215
timestamp 18001
transform 1 0 4876 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_1_Right_503
timestamp 18001
transform -1 0 7912 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_3_Left_363
timestamp 18001
transform 1 0 85284 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_3_Right_70
timestamp 18001
transform -1 0 88596 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_1_Left_216
timestamp 18001
transform 1 0 4876 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_1_Right_504
timestamp 18001
transform -1 0 7912 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_3_Left_364
timestamp 18001
transform 1 0 85284 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_3_Right_71
timestamp 18001
transform -1 0 88596 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_1_Left_217
timestamp 18001
transform 1 0 4876 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_1_Right_505
timestamp 18001
transform -1 0 7912 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_3_Left_365
timestamp 18001
transform 1 0 85284 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_3_Right_72
timestamp 18001
transform -1 0 88596 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_1_Left_218
timestamp 18001
transform 1 0 4876 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_1_Right_506
timestamp 18001
transform -1 0 7912 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_3_Left_366
timestamp 18001
transform 1 0 85284 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_3_Right_73
timestamp 18001
transform -1 0 88596 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_1_Left_219
timestamp 18001
transform 1 0 4876 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_1_Right_507
timestamp 18001
transform -1 0 7912 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_3_Left_367
timestamp 18001
transform 1 0 85284 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_3_Right_74
timestamp 18001
transform -1 0 88596 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_1_Left_220
timestamp 18001
transform 1 0 4876 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_1_Right_508
timestamp 18001
transform -1 0 7912 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_3_Left_368
timestamp 18001
transform 1 0 85284 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_3_Right_75
timestamp 18001
transform -1 0 88596 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_1_Left_221
timestamp 18001
transform 1 0 4876 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_1_Right_509
timestamp 18001
transform -1 0 7912 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_3_Left_369
timestamp 18001
transform 1 0 85284 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_3_Right_76
timestamp 18001
transform -1 0 88596 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_1_Left_222
timestamp 18001
transform 1 0 4876 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_1_Right_510
timestamp 18001
transform -1 0 7912 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_3_Left_370
timestamp 18001
transform 1 0 85284 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_3_Right_77
timestamp 18001
transform -1 0 88596 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_1_Left_223
timestamp 18001
transform 1 0 4876 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_1_Right_511
timestamp 18001
transform -1 0 7912 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_5_Left_371
timestamp 18001
transform 1 0 85284 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_5_Right_78
timestamp 18001
transform -1 0 88596 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_1_Left_224
timestamp 18001
transform 1 0 4876 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_1_Right_512
timestamp 18001
transform -1 0 7912 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_5_Left_372
timestamp 18001
transform 1 0 85284 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_5_Right_79
timestamp 18001
transform -1 0 88596 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_1_Left_225
timestamp 18001
transform 1 0 4876 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_1_Right_513
timestamp 18001
transform -1 0 7912 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_5_Left_373
timestamp 18001
transform 1 0 85284 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_5_Right_80
timestamp 18001
transform -1 0 88596 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_1_Left_226
timestamp 18001
transform 1 0 4876 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_1_Right_514
timestamp 18001
transform -1 0 7912 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_5_Left_374
timestamp 18001
transform 1 0 85284 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_5_Right_81
timestamp 18001
transform -1 0 88596 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_1_Left_227
timestamp 18001
transform 1 0 4876 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_1_Right_515
timestamp 18001
transform -1 0 7912 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_5_Left_375
timestamp 18001
transform 1 0 85284 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_5_Right_82
timestamp 18001
transform -1 0 88596 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_1_Left_228
timestamp 18001
transform 1 0 4876 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_1_Right_516
timestamp 18001
transform -1 0 7912 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_5_Left_376
timestamp 18001
transform 1 0 85284 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_5_Right_83
timestamp 18001
transform -1 0 88596 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_1_Left_229
timestamp 18001
transform 1 0 4876 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_1_Right_517
timestamp 18001
transform -1 0 7912 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_5_Left_377
timestamp 18001
transform 1 0 85284 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_5_Right_84
timestamp 18001
transform -1 0 88596 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_1_Left_230
timestamp 18001
transform 1 0 4876 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_1_Right_518
timestamp 18001
transform -1 0 7912 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_3_Left_378
timestamp 18001
transform 1 0 85284 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_3_Right_85
timestamp 18001
transform -1 0 88596 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_1_Left_231
timestamp 18001
transform 1 0 4876 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_1_Right_519
timestamp 18001
transform -1 0 7912 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_3_Left_379
timestamp 18001
transform 1 0 85284 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_3_Right_86
timestamp 18001
transform -1 0 88596 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_1_Left_232
timestamp 18001
transform 1 0 4876 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_1_Right_520
timestamp 18001
transform -1 0 7912 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_3_Left_380
timestamp 18001
transform 1 0 85284 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_3_Right_87
timestamp 18001
transform -1 0 88596 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_1_Left_233
timestamp 18001
transform 1 0 4876 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_1_Right_521
timestamp 18001
transform -1 0 7912 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_3_Left_381
timestamp 18001
transform 1 0 85284 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_3_Right_88
timestamp 18001
transform -1 0 88596 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_1_Left_234
timestamp 18001
transform 1 0 4876 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_1_Right_522
timestamp 18001
transform -1 0 7912 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_3_Left_382
timestamp 18001
transform 1 0 85284 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_3_Right_89
timestamp 18001
transform -1 0 88596 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_1_Left_235
timestamp 18001
transform 1 0 4876 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_1_Right_523
timestamp 18001
transform -1 0 7912 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_3_Left_383
timestamp 18001
transform 1 0 85284 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_3_Right_90
timestamp 18001
transform -1 0 88596 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_1_Left_236
timestamp 18001
transform 1 0 4876 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_1_Right_524
timestamp 18001
transform -1 0 7912 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_3_Left_384
timestamp 18001
transform 1 0 85284 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_3_Right_91
timestamp 18001
transform -1 0 88596 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_1_Left_237
timestamp 18001
transform 1 0 4876 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_1_Right_525
timestamp 18001
transform -1 0 7912 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_3_Left_385
timestamp 18001
transform 1 0 85284 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_3_Right_92
timestamp 18001
transform -1 0 88596 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_1_Left_238
timestamp 18001
transform 1 0 4876 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_1_Right_526
timestamp 18001
transform -1 0 7912 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_3_Left_386
timestamp 18001
transform 1 0 85284 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_3_Right_93
timestamp 18001
transform -1 0 88596 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_1_Left_239
timestamp 18001
transform 1 0 4876 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_1_Right_527
timestamp 18001
transform -1 0 7912 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_3_Left_387
timestamp 18001
transform 1 0 85284 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_3_Right_94
timestamp 18001
transform -1 0 88596 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_1_Left_240
timestamp 18001
transform 1 0 4876 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_1_Right_528
timestamp 18001
transform -1 0 7912 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_3_Left_388
timestamp 18001
transform 1 0 85284 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_3_Right_95
timestamp 18001
transform -1 0 88596 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_1_Left_241
timestamp 18001
transform 1 0 4876 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_1_Right_529
timestamp 18001
transform -1 0 7912 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_3_Left_389
timestamp 18001
transform 1 0 85284 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_3_Right_96
timestamp 18001
transform -1 0 88596 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_1_Left_242
timestamp 18001
transform 1 0 4876 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_1_Right_530
timestamp 18001
transform -1 0 7912 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_3_Left_390
timestamp 18001
transform 1 0 85284 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_3_Right_97
timestamp 18001
transform -1 0 88596 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_1_Left_243
timestamp 18001
transform 1 0 4876 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_1_Right_531
timestamp 18001
transform -1 0 7912 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_3_Left_391
timestamp 18001
transform 1 0 85284 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_3_Right_98
timestamp 18001
transform -1 0 88596 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_1_Left_244
timestamp 18001
transform 1 0 4876 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_1_Right_532
timestamp 18001
transform -1 0 7912 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_3_Left_392
timestamp 18001
transform 1 0 85284 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_3_Right_99
timestamp 18001
transform -1 0 88596 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_1_Left_245
timestamp 18001
transform 1 0 4876 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_1_Right_533
timestamp 18001
transform -1 0 7912 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_3_Left_393
timestamp 18001
transform 1 0 85284 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_3_Right_100
timestamp 18001
transform -1 0 88596 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_1_Left_246
timestamp 18001
transform 1 0 4876 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_1_Right_534
timestamp 18001
transform -1 0 7912 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_3_Left_394
timestamp 18001
transform 1 0 85284 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_3_Right_101
timestamp 18001
transform -1 0 88596 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_1_Left_247
timestamp 18001
transform 1 0 4876 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_1_Right_535
timestamp 18001
transform -1 0 7912 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_3_Left_395
timestamp 18001
transform 1 0 85284 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_3_Right_102
timestamp 18001
transform -1 0 88596 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_1_Left_248
timestamp 18001
transform 1 0 4876 0 -1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_1_Right_536
timestamp 18001
transform -1 0 7912 0 -1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_3_Left_396
timestamp 18001
transform 1 0 85284 0 -1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_3_Right_103
timestamp 18001
transform -1 0 88596 0 -1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_1_Left_249
timestamp 18001
transform 1 0 4876 0 1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_1_Right_537
timestamp 18001
transform -1 0 7912 0 1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_3_Left_397
timestamp 18001
transform 1 0 85284 0 1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_3_Right_104
timestamp 18001
transform -1 0 88596 0 1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_1_Left_250
timestamp 18001
transform 1 0 4876 0 -1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_1_Right_538
timestamp 18001
transform -1 0 7912 0 -1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_3_Left_398
timestamp 18001
transform 1 0 85284 0 -1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_3_Right_105
timestamp 18001
transform -1 0 88596 0 -1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_1_Left_251
timestamp 18001
transform 1 0 4876 0 1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_1_Right_539
timestamp 18001
transform -1 0 7912 0 1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_3_Left_399
timestamp 18001
transform 1 0 85284 0 1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_3_Right_106
timestamp 18001
transform -1 0 88596 0 1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_1_Left_252
timestamp 18001
transform 1 0 4876 0 -1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_1_Right_540
timestamp 18001
transform -1 0 7912 0 -1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_3_Left_400
timestamp 18001
transform 1 0 85284 0 -1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_3_Right_107
timestamp 18001
transform -1 0 88596 0 -1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_1_Left_253
timestamp 18001
transform 1 0 4876 0 1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_1_Right_541
timestamp 18001
transform -1 0 7912 0 1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_3_Left_401
timestamp 18001
transform 1 0 85284 0 1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_3_Right_108
timestamp 18001
transform -1 0 88596 0 1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_1_Left_254
timestamp 18001
transform 1 0 4876 0 -1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_1_Right_542
timestamp 18001
transform -1 0 7912 0 -1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_3_Left_402
timestamp 18001
transform 1 0 85284 0 -1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_3_Right_109
timestamp 18001
transform -1 0 88596 0 -1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_1_Left_255
timestamp 18001
transform 1 0 4876 0 1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_1_Right_543
timestamp 18001
transform -1 0 7912 0 1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_3_Left_403
timestamp 18001
transform 1 0 85284 0 1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_3_Right_110
timestamp 18001
transform -1 0 88596 0 1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_1_Left_256
timestamp 18001
transform 1 0 4876 0 -1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_1_Right_544
timestamp 18001
transform -1 0 7912 0 -1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_3_Left_404
timestamp 18001
transform 1 0 85284 0 -1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_3_Right_111
timestamp 18001
transform -1 0 88596 0 -1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_1_Left_257
timestamp 18001
transform 1 0 4876 0 1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_1_Right_545
timestamp 18001
transform -1 0 7912 0 1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_3_Left_405
timestamp 18001
transform 1 0 85284 0 1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_3_Right_112
timestamp 18001
transform -1 0 88596 0 1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_1_Left_258
timestamp 18001
transform 1 0 4876 0 -1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_1_Right_546
timestamp 18001
transform -1 0 7912 0 -1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_3_Left_406
timestamp 18001
transform 1 0 85284 0 -1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_3_Right_113
timestamp 18001
transform -1 0 88596 0 -1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_1_Left_259
timestamp 18001
transform 1 0 4876 0 1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_1_Right_547
timestamp 18001
transform -1 0 7912 0 1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_3_Left_407
timestamp 18001
transform 1 0 85284 0 1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_3_Right_114
timestamp 18001
transform -1 0 88596 0 1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_1_Left_260
timestamp 18001
transform 1 0 4876 0 -1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_1_Right_548
timestamp 18001
transform -1 0 7912 0 -1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_3_Left_408
timestamp 18001
transform 1 0 85284 0 -1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_3_Right_115
timestamp 18001
transform -1 0 88596 0 -1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_1_Left_261
timestamp 18001
transform 1 0 4876 0 1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_1_Right_549
timestamp 18001
transform -1 0 7912 0 1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_3_Left_409
timestamp 18001
transform 1 0 85284 0 1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_3_Right_116
timestamp 18001
transform -1 0 88596 0 1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_1_Left_262
timestamp 18001
transform 1 0 4876 0 -1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_1_Right_550
timestamp 18001
transform -1 0 7912 0 -1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_3_Left_410
timestamp 18001
transform 1 0 85284 0 -1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_3_Right_117
timestamp 18001
transform -1 0 88596 0 -1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_1_Left_263
timestamp 18001
transform 1 0 4876 0 1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_1_Right_551
timestamp 18001
transform -1 0 7912 0 1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_3_Left_411
timestamp 18001
transform 1 0 85284 0 1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_3_Right_118
timestamp 18001
transform -1 0 88596 0 1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_1_Left_264
timestamp 18001
transform 1 0 4876 0 -1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_1_Right_552
timestamp 18001
transform -1 0 7912 0 -1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_3_Left_412
timestamp 18001
transform 1 0 85284 0 -1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_3_Right_119
timestamp 18001
transform -1 0 88596 0 -1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_1_Left_265
timestamp 18001
transform 1 0 4876 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_1_Right_553
timestamp 18001
transform -1 0 7912 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_3_Left_413
timestamp 18001
transform 1 0 85284 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_3_Right_120
timestamp 18001
transform -1 0 88596 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_1_Left_266
timestamp 18001
transform 1 0 4876 0 -1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_1_Right_554
timestamp 18001
transform -1 0 7912 0 -1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_3_Left_414
timestamp 18001
transform 1 0 85284 0 -1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_3_Right_121
timestamp 18001
transform -1 0 88596 0 -1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_1_Left_267
timestamp 18001
transform 1 0 4876 0 1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_1_Right_555
timestamp 18001
transform -1 0 7912 0 1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_3_Left_415
timestamp 18001
transform 1 0 85284 0 1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_3_Right_122
timestamp 18001
transform -1 0 88596 0 1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_117_1_Left_268
timestamp 18001
transform 1 0 4876 0 -1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_117_1_Right_556
timestamp 18001
transform -1 0 7912 0 -1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_117_3_Left_416
timestamp 18001
transform 1 0 85284 0 -1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_117_3_Right_123
timestamp 18001
transform -1 0 88596 0 -1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_118_1_Left_269
timestamp 18001
transform 1 0 4876 0 1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_118_1_Right_557
timestamp 18001
transform -1 0 7912 0 1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_118_3_Left_417
timestamp 18001
transform 1 0 85284 0 1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_118_3_Right_124
timestamp 18001
transform -1 0 88596 0 1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_119_1_Left_270
timestamp 18001
transform 1 0 4876 0 -1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_119_1_Right_558
timestamp 18001
transform -1 0 7912 0 -1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_119_3_Left_418
timestamp 18001
transform 1 0 85284 0 -1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_119_3_Right_125
timestamp 18001
transform -1 0 88596 0 -1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_120_1_Left_271
timestamp 18001
transform 1 0 4876 0 1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_120_1_Right_559
timestamp 18001
transform -1 0 7912 0 1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_120_3_Left_419
timestamp 18001
transform 1 0 85284 0 1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_120_3_Right_126
timestamp 18001
transform -1 0 88596 0 1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_121_1_Left_272
timestamp 18001
transform 1 0 4876 0 -1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_121_1_Right_560
timestamp 18001
transform -1 0 7912 0 -1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_121_3_Left_420
timestamp 18001
transform 1 0 85284 0 -1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_121_3_Right_127
timestamp 18001
transform -1 0 88596 0 -1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_122_1_Left_273
timestamp 18001
transform 1 0 4876 0 1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_122_1_Right_561
timestamp 18001
transform -1 0 7912 0 1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_122_3_Left_421
timestamp 18001
transform 1 0 85284 0 1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_122_3_Right_128
timestamp 18001
transform -1 0 88596 0 1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_123_1_Left_274
timestamp 18001
transform 1 0 4876 0 -1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_123_1_Right_562
timestamp 18001
transform -1 0 7912 0 -1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_123_3_Left_422
timestamp 18001
transform 1 0 85284 0 -1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_123_3_Right_129
timestamp 18001
transform -1 0 88596 0 -1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_124_1_Left_275
timestamp 18001
transform 1 0 4876 0 1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_124_1_Right_563
timestamp 18001
transform -1 0 7912 0 1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_124_3_Left_423
timestamp 18001
transform 1 0 85284 0 1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_124_3_Right_130
timestamp 18001
transform -1 0 88596 0 1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_125_1_Left_276
timestamp 18001
transform 1 0 4876 0 -1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_125_1_Right_564
timestamp 18001
transform -1 0 7912 0 -1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_125_3_Left_424
timestamp 18001
transform 1 0 85284 0 -1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_125_3_Right_131
timestamp 18001
transform -1 0 88596 0 -1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_126_1_Left_277
timestamp 18001
transform 1 0 4876 0 1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_126_1_Right_565
timestamp 18001
transform -1 0 7912 0 1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_126_3_Left_425
timestamp 18001
transform 1 0 85284 0 1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_126_3_Right_132
timestamp 18001
transform -1 0 88596 0 1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_127_1_Left_278
timestamp 18001
transform 1 0 4876 0 -1 74528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_127_1_Right_566
timestamp 18001
transform -1 0 7912 0 -1 74528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_127_3_Left_426
timestamp 18001
transform 1 0 85284 0 -1 74528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_127_3_Right_133
timestamp 18001
transform -1 0 88596 0 -1 74528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_128_1_Left_279
timestamp 18001
transform 1 0 4876 0 1 74528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_128_1_Right_567
timestamp 18001
transform -1 0 7912 0 1 74528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_128_3_Left_427
timestamp 18001
transform 1 0 85284 0 1 74528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_128_3_Right_134
timestamp 18001
transform -1 0 88596 0 1 74528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_129_1_Left_280
timestamp 18001
transform 1 0 4876 0 -1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_129_1_Right_568
timestamp 18001
transform -1 0 7912 0 -1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_129_3_Left_428
timestamp 18001
transform 1 0 85284 0 -1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_129_3_Right_135
timestamp 18001
transform -1 0 88596 0 -1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_130_1_Left_281
timestamp 18001
transform 1 0 4876 0 1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_130_1_Right_569
timestamp 18001
transform -1 0 7912 0 1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_130_3_Left_429
timestamp 18001
transform 1 0 85284 0 1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_130_3_Right_136
timestamp 18001
transform -1 0 88596 0 1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_131_1_Left_282
timestamp 18001
transform 1 0 4876 0 -1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_131_1_Right_570
timestamp 18001
transform -1 0 7912 0 -1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_131_3_Left_430
timestamp 18001
transform 1 0 85284 0 -1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_131_3_Right_137
timestamp 18001
transform -1 0 88596 0 -1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_132_1_Left_283
timestamp 18001
transform 1 0 4876 0 1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_132_1_Right_571
timestamp 18001
transform -1 0 7912 0 1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_132_3_Left_431
timestamp 18001
transform 1 0 85284 0 1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_132_3_Right_138
timestamp 18001
transform -1 0 88596 0 1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_133_1_Left_284
timestamp 18001
transform 1 0 4876 0 -1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_133_1_Right_572
timestamp 18001
transform -1 0 7912 0 -1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_133_3_Left_432
timestamp 18001
transform 1 0 85284 0 -1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_133_3_Right_139
timestamp 18001
transform -1 0 88596 0 -1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_134_1_Left_285
timestamp 18001
transform 1 0 4876 0 1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_134_1_Right_573
timestamp 18001
transform -1 0 7912 0 1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_134_3_Left_433
timestamp 18001
transform 1 0 85284 0 1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_134_3_Right_140
timestamp 18001
transform -1 0 88596 0 1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_135_1_Left_286
timestamp 18001
transform 1 0 4876 0 -1 78880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_135_1_Right_574
timestamp 18001
transform -1 0 7912 0 -1 78880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_135_3_Left_434
timestamp 18001
transform 1 0 85284 0 -1 78880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_135_3_Right_141
timestamp 18001
transform -1 0 88596 0 -1 78880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_136_1_Left_287
timestamp 18001
transform 1 0 4876 0 1 78880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_136_1_Right_575
timestamp 18001
transform -1 0 7912 0 1 78880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_136_3_Left_435
timestamp 18001
transform 1 0 85284 0 1 78880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_136_3_Right_142
timestamp 18001
transform -1 0 88596 0 1 78880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_137_1_Left_288
timestamp 18001
transform 1 0 4876 0 -1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_137_1_Right_576
timestamp 18001
transform -1 0 7912 0 -1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_137_3_Left_436
timestamp 18001
transform 1 0 85284 0 -1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_137_3_Right_143
timestamp 18001
transform -1 0 88596 0 -1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_138_1_Left_289
timestamp 18001
transform 1 0 4876 0 1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_138_1_Right_577
timestamp 18001
transform -1 0 7912 0 1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_138_3_Left_437
timestamp 18001
transform 1 0 85284 0 1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_138_3_Right_144
timestamp 18001
transform -1 0 88596 0 1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_139_1_Left_290
timestamp 18001
transform 1 0 4876 0 -1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_139_1_Right_578
timestamp 18001
transform -1 0 7912 0 -1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_139_3_Left_438
timestamp 18001
transform 1 0 85284 0 -1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_139_3_Right_145
timestamp 18001
transform -1 0 88596 0 -1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_140_1_Left_291
timestamp 18001
transform 1 0 4876 0 1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_140_1_Right_579
timestamp 18001
transform -1 0 7912 0 1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_140_3_Left_439
timestamp 18001
transform 1 0 85284 0 1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_140_3_Right_146
timestamp 18001
transform -1 0 88596 0 1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_141_1_Left_292
timestamp 18001
transform 1 0 4876 0 -1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_141_1_Right_580
timestamp 18001
transform -1 0 7912 0 -1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_141_3_Left_440
timestamp 18001
transform 1 0 85284 0 -1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_141_3_Right_147
timestamp 18001
transform -1 0 88596 0 -1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_142_1_Left_293
timestamp 18001
transform 1 0 4876 0 1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_142_1_Right_581
timestamp 18001
transform -1 0 7912 0 1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_142_3_Left_441
timestamp 18001
transform 1 0 85284 0 1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_142_3_Right_148
timestamp 18001
transform -1 0 88596 0 1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_143_1_Left_294
timestamp 18001
transform 1 0 4876 0 -1 83232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_143_1_Right_582
timestamp 18001
transform -1 0 7912 0 -1 83232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_143_3_Left_442
timestamp 18001
transform 1 0 85284 0 -1 83232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_143_3_Right_149
timestamp 18001
transform -1 0 88596 0 -1 83232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_144_1_Left_295
timestamp 18001
transform 1 0 4876 0 1 83232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_144_1_Right_583
timestamp 18001
transform -1 0 7912 0 1 83232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_144_3_Left_443
timestamp 18001
transform 1 0 85284 0 1 83232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_144_3_Right_150
timestamp 18001
transform -1 0 88596 0 1 83232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_145_1_Left_296
timestamp 18001
transform 1 0 4876 0 -1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_145_1_Right_584
timestamp 18001
transform -1 0 7912 0 -1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_145_3_Left_444
timestamp 18001
transform 1 0 85284 0 -1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_145_3_Right_151
timestamp 18001
transform -1 0 88596 0 -1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_146_Left_297
timestamp 18001
transform 1 0 4876 0 1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_146_Right_5
timestamp 18001
transform -1 0 88596 0 1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_147_Left_298
timestamp 18001
transform 1 0 4876 0 -1 85408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_147_Right_6
timestamp 18001
transform -1 0 88596 0 -1 85408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_148_Left_299
timestamp 18001
transform 1 0 4876 0 1 85408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_148_Right_7
timestamp 18001
transform -1 0 88596 0 1 85408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_149_Left_300
timestamp 18001
transform 1 0 4876 0 -1 86496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_149_Right_8
timestamp 18001
transform -1 0 88596 0 -1 86496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_150_Left_301
timestamp 18001
transform 1 0 4876 0 1 86496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_150_Right_9
timestamp 18001
transform -1 0 88596 0 1 86496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_151_Left_302
timestamp 18001
transform 1 0 4876 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_151_Right_10
timestamp 18001
transform -1 0 88596 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_586
timestamp 18001
transform 1 0 7452 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_587
timestamp 18001
transform 1 0 10028 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_588
timestamp 18001
transform 1 0 12604 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_589
timestamp 18001
transform 1 0 15180 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_590
timestamp 18001
transform 1 0 17756 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_591
timestamp 18001
transform 1 0 20332 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_592
timestamp 18001
transform 1 0 22908 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_593
timestamp 18001
transform 1 0 25484 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_594
timestamp 18001
transform 1 0 28060 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_595
timestamp 18001
transform 1 0 30636 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_596
timestamp 18001
transform 1 0 33212 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_597
timestamp 18001
transform 1 0 35788 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_598
timestamp 18001
transform 1 0 38364 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_599
timestamp 18001
transform 1 0 40940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_600
timestamp 18001
transform 1 0 43516 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_601
timestamp 18001
transform 1 0 46092 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_602
timestamp 18001
transform 1 0 48668 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_603
timestamp 18001
transform 1 0 51244 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_604
timestamp 18001
transform 1 0 53820 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_605
timestamp 18001
transform 1 0 56396 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_606
timestamp 18001
transform 1 0 58972 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_607
timestamp 18001
transform 1 0 61548 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_608
timestamp 18001
transform 1 0 64124 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_609
timestamp 18001
transform 1 0 66700 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_610
timestamp 18001
transform 1 0 69276 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_611
timestamp 18001
transform 1 0 71852 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_612
timestamp 18001
transform 1 0 74428 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_613
timestamp 18001
transform 1 0 77004 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_614
timestamp 18001
transform 1 0 79580 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_615
timestamp 18001
transform 1 0 82156 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_616
timestamp 18001
transform 1 0 84732 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_617
timestamp 18001
transform 1 0 87308 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_618
timestamp 18001
transform 1 0 10028 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_619
timestamp 18001
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_620
timestamp 18001
transform 1 0 20332 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_621
timestamp 18001
transform 1 0 25484 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_622
timestamp 18001
transform 1 0 30636 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_623
timestamp 18001
transform 1 0 35788 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_624
timestamp 18001
transform 1 0 40940 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_625
timestamp 18001
transform 1 0 46092 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_626
timestamp 18001
transform 1 0 51244 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_627
timestamp 18001
transform 1 0 56396 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_628
timestamp 18001
transform 1 0 61548 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_629
timestamp 18001
transform 1 0 66700 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_630
timestamp 18001
transform 1 0 71852 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_631
timestamp 18001
transform 1 0 77004 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_632
timestamp 18001
transform 1 0 82156 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_633
timestamp 18001
transform 1 0 87308 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_634
timestamp 18001
transform 1 0 7452 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_635
timestamp 18001
transform 1 0 12604 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_636
timestamp 18001
transform 1 0 17756 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_637
timestamp 18001
transform 1 0 22908 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_638
timestamp 18001
transform 1 0 28060 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_639
timestamp 18001
transform 1 0 33212 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_640
timestamp 18001
transform 1 0 38364 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_641
timestamp 18001
transform 1 0 43516 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_642
timestamp 18001
transform 1 0 48668 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_643
timestamp 18001
transform 1 0 53820 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_644
timestamp 18001
transform 1 0 58972 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_645
timestamp 18001
transform 1 0 64124 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_646
timestamp 18001
transform 1 0 69276 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_647
timestamp 18001
transform 1 0 74428 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_648
timestamp 18001
transform 1 0 79580 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_649
timestamp 18001
transform 1 0 84732 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_650
timestamp 18001
transform 1 0 10028 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_651
timestamp 18001
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_652
timestamp 18001
transform 1 0 20332 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_653
timestamp 18001
transform 1 0 25484 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_654
timestamp 18001
transform 1 0 30636 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_655
timestamp 18001
transform 1 0 35788 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_656
timestamp 18001
transform 1 0 40940 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_657
timestamp 18001
transform 1 0 46092 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_658
timestamp 18001
transform 1 0 51244 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_659
timestamp 18001
transform 1 0 56396 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_660
timestamp 18001
transform 1 0 61548 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_661
timestamp 18001
transform 1 0 66700 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_662
timestamp 18001
transform 1 0 71852 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_663
timestamp 18001
transform 1 0 77004 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_664
timestamp 18001
transform 1 0 82156 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_665
timestamp 18001
transform 1 0 87308 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_666
timestamp 18001
transform 1 0 7452 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_667
timestamp 18001
transform 1 0 10028 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_668
timestamp 18001
transform 1 0 12604 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_669
timestamp 18001
transform 1 0 15180 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_670
timestamp 18001
transform 1 0 17756 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_671
timestamp 18001
transform 1 0 20332 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_672
timestamp 18001
transform 1 0 22908 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_673
timestamp 18001
transform 1 0 25484 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_674
timestamp 18001
transform 1 0 28060 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_675
timestamp 18001
transform 1 0 30636 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_676
timestamp 18001
transform 1 0 33212 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_677
timestamp 18001
transform 1 0 35788 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_678
timestamp 18001
transform 1 0 38364 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_679
timestamp 18001
transform 1 0 40940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_680
timestamp 18001
transform 1 0 43516 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_681
timestamp 18001
transform 1 0 46092 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_682
timestamp 18001
transform 1 0 48668 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_683
timestamp 18001
transform 1 0 51244 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_684
timestamp 18001
transform 1 0 53820 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_685
timestamp 18001
transform 1 0 56396 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_686
timestamp 18001
transform 1 0 58972 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_687
timestamp 18001
transform 1 0 61548 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_688
timestamp 18001
transform 1 0 64124 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_689
timestamp 18001
transform 1 0 66700 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_690
timestamp 18001
transform 1 0 69276 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_691
timestamp 18001
transform 1 0 71852 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_692
timestamp 18001
transform 1 0 74428 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_693
timestamp 18001
transform 1 0 77004 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_694
timestamp 18001
transform 1 0 79580 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_695
timestamp 18001
transform 1 0 82156 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_696
timestamp 18001
transform 1 0 84732 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_697
timestamp 18001
transform 1 0 87308 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1_698
timestamp 18001
transform 1 0 7452 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_3_896
timestamp 18001
transform 1 0 87860 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1_699
timestamp 18001
transform 1 0 7452 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_3_897
timestamp 18001
transform 1 0 87860 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_1_700
timestamp 18001
transform 1 0 7452 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_3_898
timestamp 18001
transform 1 0 87860 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_1_701
timestamp 18001
transform 1 0 7452 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_3_899
timestamp 18001
transform 1 0 87860 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_1_702
timestamp 18001
transform 1 0 7452 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_3_900
timestamp 18001
transform 1 0 87860 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_1_703
timestamp 18001
transform 1 0 7452 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_3_901
timestamp 18001
transform 1 0 87860 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_1_704
timestamp 18001
transform 1 0 7452 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_3_902
timestamp 18001
transform 1 0 87860 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_1_705
timestamp 18001
transform 1 0 7452 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_3_903
timestamp 18001
transform 1 0 87860 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_1_706
timestamp 18001
transform 1 0 7452 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_3_904
timestamp 18001
transform 1 0 87860 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_1_707
timestamp 18001
transform 1 0 7452 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_3_905
timestamp 18001
transform 1 0 87860 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_1_708
timestamp 18001
transform 1 0 7452 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_3_906
timestamp 18001
transform 1 0 87860 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_1_709
timestamp 18001
transform 1 0 7452 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_3_907
timestamp 18001
transform 1 0 87860 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_1_710
timestamp 18001
transform 1 0 7452 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_3_908
timestamp 18001
transform 1 0 87860 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_1_711
timestamp 18001
transform 1 0 7452 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_3_909
timestamp 18001
transform 1 0 87860 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_1_712
timestamp 18001
transform 1 0 7452 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_3_910
timestamp 18001
transform 1 0 87860 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_1_713
timestamp 18001
transform 1 0 7452 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_3_911
timestamp 18001
transform 1 0 87860 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_1_714
timestamp 18001
transform 1 0 7452 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_3_912
timestamp 18001
transform 1 0 87860 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_1_715
timestamp 18001
transform 1 0 7452 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_3_913
timestamp 18001
transform 1 0 87860 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_1_716
timestamp 18001
transform 1 0 7452 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_3_914
timestamp 18001
transform 1 0 87860 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_1_717
timestamp 18001
transform 1 0 7452 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_3_915
timestamp 18001
transform 1 0 87860 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_1_718
timestamp 18001
transform 1 0 7452 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_3_916
timestamp 18001
transform 1 0 87860 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_1_719
timestamp 18001
transform 1 0 7452 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_3_917
timestamp 18001
transform 1 0 87860 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_1_720
timestamp 18001
transform 1 0 7452 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_3_918
timestamp 18001
transform 1 0 87860 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_1_721
timestamp 18001
transform 1 0 7452 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_3_919
timestamp 18001
transform 1 0 87860 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_1_722
timestamp 18001
transform 1 0 7452 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_3_920
timestamp 18001
transform 1 0 87860 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_1_723
timestamp 18001
transform 1 0 7452 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_3_921
timestamp 18001
transform 1 0 87860 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_1_724
timestamp 18001
transform 1 0 7452 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_3_922
timestamp 18001
transform 1 0 87860 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1_725
timestamp 18001
transform 1 0 7452 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_3_923
timestamp 18001
transform 1 0 87860 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1_726
timestamp 18001
transform 1 0 7452 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_3_924
timestamp 18001
transform 1 0 87860 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1_727
timestamp 18001
transform 1 0 7452 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_3_925
timestamp 18001
transform 1 0 87860 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_1_728
timestamp 18001
transform 1 0 7452 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_3_926
timestamp 18001
transform 1 0 87860 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_1_729
timestamp 18001
transform 1 0 7452 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_3_927
timestamp 18001
transform 1 0 87860 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_1_730
timestamp 18001
transform 1 0 7452 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_3_928
timestamp 18001
transform 1 0 87860 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1_731
timestamp 18001
transform 1 0 7452 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_5_929
timestamp 18001
transform 1 0 87860 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1_732
timestamp 18001
transform 1 0 7452 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_5_930
timestamp 18001
transform 1 0 87860 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1_733
timestamp 18001
transform 1 0 7452 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_5_931
timestamp 18001
transform 1 0 87860 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1_734
timestamp 18001
transform 1 0 7452 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_5_932
timestamp 18001
transform 1 0 87860 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1_735
timestamp 18001
transform 1 0 7452 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_3_933
timestamp 18001
transform 1 0 87860 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1_736
timestamp 18001
transform 1 0 7452 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_3_934
timestamp 18001
transform 1 0 87860 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1_737
timestamp 18001
transform 1 0 7452 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_3_935
timestamp 18001
transform 1 0 87860 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1_738
timestamp 18001
transform 1 0 7452 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_3_936
timestamp 18001
transform 1 0 87860 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1_739
timestamp 18001
transform 1 0 7452 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_3_937
timestamp 18001
transform 1 0 87860 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1_740
timestamp 18001
transform 1 0 7452 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_3_938
timestamp 18001
transform 1 0 87860 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1_741
timestamp 18001
transform 1 0 7452 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_3_939
timestamp 18001
transform 1 0 87860 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1_742
timestamp 18001
transform 1 0 7452 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_3_940
timestamp 18001
transform 1 0 87860 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1_743
timestamp 18001
transform 1 0 7452 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_3_941
timestamp 18001
transform 1 0 87860 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1_744
timestamp 18001
transform 1 0 7452 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_3_942
timestamp 18001
transform 1 0 87860 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1_745
timestamp 18001
transform 1 0 7452 0 1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_3_943
timestamp 18001
transform 1 0 87860 0 1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_1_746
timestamp 18001
transform 1 0 7452 0 1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_3_944
timestamp 18001
transform 1 0 87860 0 1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_1_747
timestamp 18001
transform 1 0 7452 0 1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_3_945
timestamp 18001
transform 1 0 87860 0 1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_1_748
timestamp 18001
transform 1 0 7452 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_3_946
timestamp 18001
transform 1 0 87860 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_1_749
timestamp 18001
transform 1 0 7452 0 1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_3_947
timestamp 18001
transform 1 0 87860 0 1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_1_750
timestamp 18001
transform 1 0 7452 0 1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_3_948
timestamp 18001
transform 1 0 87860 0 1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_1_751
timestamp 18001
transform 1 0 7452 0 1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_3_949
timestamp 18001
transform 1 0 87860 0 1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_1_752
timestamp 18001
transform 1 0 7452 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_3_950
timestamp 18001
transform 1 0 87860 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_1_753
timestamp 18001
transform 1 0 7452 0 1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_3_951
timestamp 18001
transform 1 0 87860 0 1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1_754
timestamp 18001
transform 1 0 7452 0 1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_3_952
timestamp 18001
transform 1 0 87860 0 1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1_755
timestamp 18001
transform 1 0 7452 0 1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_3_953
timestamp 18001
transform 1 0 87860 0 1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1_756
timestamp 18001
transform 1 0 7452 0 1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_3_954
timestamp 18001
transform 1 0 87860 0 1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1_757
timestamp 18001
transform 1 0 7452 0 1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_3_955
timestamp 18001
transform 1 0 87860 0 1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1_758
timestamp 18001
transform 1 0 7452 0 1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_3_956
timestamp 18001
transform 1 0 87860 0 1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1_759
timestamp 18001
transform 1 0 7452 0 1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_3_957
timestamp 18001
transform 1 0 87860 0 1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1_760
timestamp 18001
transform 1 0 7452 0 1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_3_958
timestamp 18001
transform 1 0 87860 0 1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1_761
timestamp 18001
transform 1 0 7452 0 1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_3_959
timestamp 18001
transform 1 0 87860 0 1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1_762
timestamp 18001
transform 1 0 7452 0 1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_3_960
timestamp 18001
transform 1 0 87860 0 1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1_763
timestamp 18001
transform 1 0 7452 0 1 78880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_3_961
timestamp 18001
transform 1 0 87860 0 1 78880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1_764
timestamp 18001
transform 1 0 7452 0 1 79968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_3_962
timestamp 18001
transform 1 0 87860 0 1 79968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_140_1_765
timestamp 18001
transform 1 0 7452 0 1 81056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_140_3_963
timestamp 18001
transform 1 0 87860 0 1 81056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_142_1_766
timestamp 18001
transform 1 0 7452 0 1 82144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_142_3_964
timestamp 18001
transform 1 0 87860 0 1 82144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_144_1_767
timestamp 18001
transform 1 0 7452 0 1 83232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_144_3_965
timestamp 18001
transform 1 0 87860 0 1 83232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_768
timestamp 18001
transform 1 0 7452 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_769
timestamp 18001
transform 1 0 10028 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_770
timestamp 18001
transform 1 0 12604 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_771
timestamp 18001
transform 1 0 15180 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_772
timestamp 18001
transform 1 0 17756 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_773
timestamp 18001
transform 1 0 20332 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_774
timestamp 18001
transform 1 0 22908 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_775
timestamp 18001
transform 1 0 25484 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_776
timestamp 18001
transform 1 0 28060 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_777
timestamp 18001
transform 1 0 30636 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_778
timestamp 18001
transform 1 0 33212 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_779
timestamp 18001
transform 1 0 35788 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_780
timestamp 18001
transform 1 0 38364 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_781
timestamp 18001
transform 1 0 40940 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_782
timestamp 18001
transform 1 0 43516 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_783
timestamp 18001
transform 1 0 46092 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_784
timestamp 18001
transform 1 0 48668 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_785
timestamp 18001
transform 1 0 51244 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_786
timestamp 18001
transform 1 0 53820 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_787
timestamp 18001
transform 1 0 56396 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_788
timestamp 18001
transform 1 0 58972 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_789
timestamp 18001
transform 1 0 61548 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_790
timestamp 18001
transform 1 0 64124 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_791
timestamp 18001
transform 1 0 66700 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_792
timestamp 18001
transform 1 0 69276 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_793
timestamp 18001
transform 1 0 71852 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_794
timestamp 18001
transform 1 0 74428 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_795
timestamp 18001
transform 1 0 77004 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_796
timestamp 18001
transform 1 0 79580 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_797
timestamp 18001
transform 1 0 82156 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_798
timestamp 18001
transform 1 0 84732 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_799
timestamp 18001
transform 1 0 87308 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_800
timestamp 18001
transform 1 0 10028 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_801
timestamp 18001
transform 1 0 15180 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_802
timestamp 18001
transform 1 0 20332 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_803
timestamp 18001
transform 1 0 25484 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_804
timestamp 18001
transform 1 0 30636 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_805
timestamp 18001
transform 1 0 35788 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_806
timestamp 18001
transform 1 0 40940 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_807
timestamp 18001
transform 1 0 46092 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_808
timestamp 18001
transform 1 0 51244 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_809
timestamp 18001
transform 1 0 56396 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_810
timestamp 18001
transform 1 0 61548 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_811
timestamp 18001
transform 1 0 66700 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_812
timestamp 18001
transform 1 0 71852 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_813
timestamp 18001
transform 1 0 77004 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_814
timestamp 18001
transform 1 0 82156 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_815
timestamp 18001
transform 1 0 87308 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_816
timestamp 18001
transform 1 0 7452 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_817
timestamp 18001
transform 1 0 12604 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_818
timestamp 18001
transform 1 0 17756 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_819
timestamp 18001
transform 1 0 22908 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_820
timestamp 18001
transform 1 0 28060 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_821
timestamp 18001
transform 1 0 33212 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_822
timestamp 18001
transform 1 0 38364 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_823
timestamp 18001
transform 1 0 43516 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_824
timestamp 18001
transform 1 0 48668 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_825
timestamp 18001
transform 1 0 53820 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_826
timestamp 18001
transform 1 0 58972 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_827
timestamp 18001
transform 1 0 64124 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_828
timestamp 18001
transform 1 0 69276 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_829
timestamp 18001
transform 1 0 74428 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_830
timestamp 18001
transform 1 0 79580 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_831
timestamp 18001
transform 1 0 84732 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_832
timestamp 18001
transform 1 0 10028 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_833
timestamp 18001
transform 1 0 15180 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_834
timestamp 18001
transform 1 0 20332 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_835
timestamp 18001
transform 1 0 25484 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_836
timestamp 18001
transform 1 0 30636 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_837
timestamp 18001
transform 1 0 35788 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_838
timestamp 18001
transform 1 0 40940 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_839
timestamp 18001
transform 1 0 46092 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_840
timestamp 18001
transform 1 0 51244 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_841
timestamp 18001
transform 1 0 56396 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_842
timestamp 18001
transform 1 0 61548 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_843
timestamp 18001
transform 1 0 66700 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_844
timestamp 18001
transform 1 0 71852 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_845
timestamp 18001
transform 1 0 77004 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_846
timestamp 18001
transform 1 0 82156 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_847
timestamp 18001
transform 1 0 87308 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_848
timestamp 18001
transform 1 0 7452 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_849
timestamp 18001
transform 1 0 12604 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_850
timestamp 18001
transform 1 0 17756 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_851
timestamp 18001
transform 1 0 22908 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_852
timestamp 18001
transform 1 0 28060 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_853
timestamp 18001
transform 1 0 33212 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_854
timestamp 18001
transform 1 0 38364 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_855
timestamp 18001
transform 1 0 43516 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_856
timestamp 18001
transform 1 0 48668 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_857
timestamp 18001
transform 1 0 53820 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_858
timestamp 18001
transform 1 0 58972 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_859
timestamp 18001
transform 1 0 64124 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_860
timestamp 18001
transform 1 0 69276 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_861
timestamp 18001
transform 1 0 74428 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_862
timestamp 18001
transform 1 0 79580 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_863
timestamp 18001
transform 1 0 84732 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_864
timestamp 18001
transform 1 0 7452 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_865
timestamp 18001
transform 1 0 10028 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_866
timestamp 18001
transform 1 0 12604 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_867
timestamp 18001
transform 1 0 15180 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_868
timestamp 18001
transform 1 0 17756 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_869
timestamp 18001
transform 1 0 20332 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_870
timestamp 18001
transform 1 0 22908 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_871
timestamp 18001
transform 1 0 25484 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_872
timestamp 18001
transform 1 0 28060 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_873
timestamp 18001
transform 1 0 30636 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_874
timestamp 18001
transform 1 0 33212 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_875
timestamp 18001
transform 1 0 35788 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_876
timestamp 18001
transform 1 0 38364 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_877
timestamp 18001
transform 1 0 40940 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_878
timestamp 18001
transform 1 0 43516 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_879
timestamp 18001
transform 1 0 46092 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_880
timestamp 18001
transform 1 0 48668 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_881
timestamp 18001
transform 1 0 51244 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_882
timestamp 18001
transform 1 0 53820 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_883
timestamp 18001
transform 1 0 56396 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_884
timestamp 18001
transform 1 0 58972 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_885
timestamp 18001
transform 1 0 61548 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_886
timestamp 18001
transform 1 0 64124 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_887
timestamp 18001
transform 1 0 66700 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_888
timestamp 18001
transform 1 0 69276 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_889
timestamp 18001
transform 1 0 71852 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_890
timestamp 18001
transform 1 0 74428 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_891
timestamp 18001
transform 1 0 77004 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_892
timestamp 18001
transform 1 0 79580 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_893
timestamp 18001
transform 1 0 82156 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_894
timestamp 18001
transform 1 0 84732 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_895
timestamp 18001
transform 1 0 87308 0 -1 87584
box -38 -48 130 592
<< labels >>
flabel metal2 s 39614 88000 39670 88800 0 FreeSans 224 90 0 0 clk
port 0 nsew signal input
flabel metal3 s 1600 45128 2400 45248 0 FreeSans 480 0 0 0 config_data_in
port 1 nsew signal input
flabel metal3 s 89200 47168 90000 47288 0 FreeSans 480 0 0 0 config_data_out
port 2 nsew signal output
flabel metal2 s 37682 88000 37738 88800 0 FreeSans 224 90 0 0 config_en
port 3 nsew signal input
flabel metal3 s 89200 30168 90000 30288 0 FreeSans 480 0 0 0 io_east_in[0]
port 4 nsew signal input
flabel metal3 s 89200 41048 90000 41168 0 FreeSans 480 0 0 0 io_east_in[10]
port 5 nsew signal input
flabel metal3 s 89200 42408 90000 42528 0 FreeSans 480 0 0 0 io_east_in[11]
port 6 nsew signal input
flabel metal3 s 89200 43768 90000 43888 0 FreeSans 480 0 0 0 io_east_in[12]
port 7 nsew signal input
flabel metal3 s 89200 44448 90000 44568 0 FreeSans 480 0 0 0 io_east_in[13]
port 8 nsew signal input
flabel metal2 s 1618 1600 1674 2400 0 FreeSans 224 90 0 0 io_east_in[14]
port 9 nsew signal input
flabel metal2 s 2262 1600 2318 2400 0 FreeSans 224 90 0 0 io_east_in[15]
port 10 nsew signal input
flabel metal3 s 89200 66888 90000 67008 0 FreeSans 480 0 0 0 io_east_in[16]
port 11 nsew signal input
flabel metal3 s 89200 67568 90000 67688 0 FreeSans 480 0 0 0 io_east_in[17]
port 12 nsew signal input
flabel metal3 s 89200 68928 90000 69048 0 FreeSans 480 0 0 0 io_east_in[18]
port 13 nsew signal input
flabel metal3 s 89200 70288 90000 70408 0 FreeSans 480 0 0 0 io_east_in[19]
port 14 nsew signal input
flabel metal3 s 89200 31528 90000 31648 0 FreeSans 480 0 0 0 io_east_in[1]
port 15 nsew signal input
flabel metal3 s 89200 70968 90000 71088 0 FreeSans 480 0 0 0 io_east_in[20]
port 16 nsew signal input
flabel metal3 s 89200 72328 90000 72448 0 FreeSans 480 0 0 0 io_east_in[21]
port 17 nsew signal input
flabel metal3 s 89200 73008 90000 73128 0 FreeSans 480 0 0 0 io_east_in[22]
port 18 nsew signal input
flabel metal3 s 89200 74368 90000 74488 0 FreeSans 480 0 0 0 io_east_in[23]
port 19 nsew signal input
flabel metal3 s 89200 75728 90000 75848 0 FreeSans 480 0 0 0 io_east_in[24]
port 20 nsew signal input
flabel metal3 s 89200 76408 90000 76528 0 FreeSans 480 0 0 0 io_east_in[25]
port 21 nsew signal input
flabel metal3 s 89200 77768 90000 77888 0 FreeSans 480 0 0 0 io_east_in[26]
port 22 nsew signal input
flabel metal3 s 89200 78448 90000 78568 0 FreeSans 480 0 0 0 io_east_in[27]
port 23 nsew signal input
flabel metal3 s 89200 79808 90000 79928 0 FreeSans 480 0 0 0 io_east_in[28]
port 24 nsew signal input
flabel metal3 s 89200 81168 90000 81288 0 FreeSans 480 0 0 0 io_east_in[29]
port 25 nsew signal input
flabel metal3 s 89200 32888 90000 33008 0 FreeSans 480 0 0 0 io_east_in[2]
port 26 nsew signal input
flabel metal2 s 2906 1600 2962 2400 0 FreeSans 224 90 0 0 io_east_in[30]
port 27 nsew signal input
flabel metal2 s 3550 1600 3606 2400 0 FreeSans 224 90 0 0 io_east_in[31]
port 28 nsew signal input
flabel metal3 s 89200 33568 90000 33688 0 FreeSans 480 0 0 0 io_east_in[3]
port 29 nsew signal input
flabel metal3 s 89200 34928 90000 35048 0 FreeSans 480 0 0 0 io_east_in[4]
port 30 nsew signal input
flabel metal3 s 89200 35608 90000 35728 0 FreeSans 480 0 0 0 io_east_in[5]
port 31 nsew signal input
flabel metal3 s 89200 36968 90000 37088 0 FreeSans 480 0 0 0 io_east_in[6]
port 32 nsew signal input
flabel metal3 s 89200 38328 90000 38448 0 FreeSans 480 0 0 0 io_east_in[7]
port 33 nsew signal input
flabel metal3 s 89200 39008 90000 39128 0 FreeSans 480 0 0 0 io_east_in[8]
port 34 nsew signal input
flabel metal3 s 89200 40368 90000 40488 0 FreeSans 480 0 0 0 io_east_in[9]
port 35 nsew signal input
flabel metal3 s 89200 15208 90000 15328 0 FreeSans 480 0 0 0 io_east_out[0]
port 36 nsew signal output
flabel metal3 s 89200 26088 90000 26208 0 FreeSans 480 0 0 0 io_east_out[10]
port 37 nsew signal output
flabel metal3 s 89200 27448 90000 27568 0 FreeSans 480 0 0 0 io_east_out[11]
port 38 nsew signal output
flabel metal3 s 89200 28128 90000 28248 0 FreeSans 480 0 0 0 io_east_out[12]
port 39 nsew signal output
flabel metal3 s 89200 29488 90000 29608 0 FreeSans 480 0 0 0 io_east_out[13]
port 40 nsew signal output
flabel metal2 s 50562 88000 50618 88800 0 FreeSans 224 90 0 0 io_east_out[14]
port 41 nsew signal output
flabel metal2 s 49918 88000 49974 88800 0 FreeSans 224 90 0 0 io_east_out[15]
port 42 nsew signal output
flabel metal3 s 89200 51248 90000 51368 0 FreeSans 480 0 0 0 io_east_out[16]
port 43 nsew signal output
flabel metal3 s 89200 52608 90000 52728 0 FreeSans 480 0 0 0 io_east_out[17]
port 44 nsew signal output
flabel metal3 s 89200 53968 90000 54088 0 FreeSans 480 0 0 0 io_east_out[18]
port 45 nsew signal output
flabel metal3 s 89200 54648 90000 54768 0 FreeSans 480 0 0 0 io_east_out[19]
port 46 nsew signal output
flabel metal3 s 89200 16568 90000 16688 0 FreeSans 480 0 0 0 io_east_out[1]
port 47 nsew signal output
flabel metal3 s 89200 56008 90000 56128 0 FreeSans 480 0 0 0 io_east_out[20]
port 48 nsew signal output
flabel metal3 s 89200 56688 90000 56808 0 FreeSans 480 0 0 0 io_east_out[21]
port 49 nsew signal output
flabel metal3 s 89200 58048 90000 58168 0 FreeSans 480 0 0 0 io_east_out[22]
port 50 nsew signal output
flabel metal3 s 89200 59408 90000 59528 0 FreeSans 480 0 0 0 io_east_out[23]
port 51 nsew signal output
flabel metal3 s 89200 60088 90000 60208 0 FreeSans 480 0 0 0 io_east_out[24]
port 52 nsew signal output
flabel metal3 s 89200 61448 90000 61568 0 FreeSans 480 0 0 0 io_east_out[25]
port 53 nsew signal output
flabel metal3 s 89200 62128 90000 62248 0 FreeSans 480 0 0 0 io_east_out[26]
port 54 nsew signal output
flabel metal3 s 89200 63488 90000 63608 0 FreeSans 480 0 0 0 io_east_out[27]
port 55 nsew signal output
flabel metal3 s 89200 64848 90000 64968 0 FreeSans 480 0 0 0 io_east_out[28]
port 56 nsew signal output
flabel metal3 s 89200 65528 90000 65648 0 FreeSans 480 0 0 0 io_east_out[29]
port 57 nsew signal output
flabel metal3 s 89200 17248 90000 17368 0 FreeSans 480 0 0 0 io_east_out[2]
port 58 nsew signal output
flabel metal2 s 47342 88000 47398 88800 0 FreeSans 224 90 0 0 io_east_out[30]
port 59 nsew signal output
flabel metal2 s 42834 88000 42890 88800 0 FreeSans 224 90 0 0 io_east_out[31]
port 60 nsew signal output
flabel metal3 s 89200 18608 90000 18728 0 FreeSans 480 0 0 0 io_east_out[3]
port 61 nsew signal output
flabel metal3 s 89200 19288 90000 19408 0 FreeSans 480 0 0 0 io_east_out[4]
port 62 nsew signal output
flabel metal3 s 89200 20648 90000 20768 0 FreeSans 480 0 0 0 io_east_out[5]
port 63 nsew signal output
flabel metal3 s 89200 22008 90000 22128 0 FreeSans 480 0 0 0 io_east_out[6]
port 64 nsew signal output
flabel metal3 s 89200 22688 90000 22808 0 FreeSans 480 0 0 0 io_east_out[7]
port 65 nsew signal output
flabel metal3 s 89200 24048 90000 24168 0 FreeSans 480 0 0 0 io_east_out[8]
port 66 nsew signal output
flabel metal3 s 89200 24728 90000 24848 0 FreeSans 480 0 0 0 io_east_out[9]
port 67 nsew signal output
flabel metal2 s 15142 88000 15198 88800 0 FreeSans 224 90 0 0 io_north_in[0]
port 68 nsew signal input
flabel metal2 s 26090 88000 26146 88800 0 FreeSans 224 90 0 0 io_north_in[10]
port 69 nsew signal input
flabel metal2 s 27378 88000 27434 88800 0 FreeSans 224 90 0 0 io_north_in[11]
port 70 nsew signal input
flabel metal2 s 28022 88000 28078 88800 0 FreeSans 224 90 0 0 io_north_in[12]
port 71 nsew signal input
flabel metal2 s 29310 88000 29366 88800 0 FreeSans 224 90 0 0 io_north_in[13]
port 72 nsew signal input
flabel metal2 s 4194 1600 4250 2400 0 FreeSans 224 90 0 0 io_north_in[14]
port 73 nsew signal input
flabel metal2 s 4838 1600 4894 2400 0 FreeSans 224 90 0 0 io_north_in[15]
port 74 nsew signal input
flabel metal2 s 52494 88000 52550 88800 0 FreeSans 224 90 0 0 io_north_in[16]
port 75 nsew signal input
flabel metal2 s 53782 88000 53838 88800 0 FreeSans 224 90 0 0 io_north_in[17]
port 76 nsew signal input
flabel metal2 s 54426 88000 54482 88800 0 FreeSans 224 90 0 0 io_north_in[18]
port 77 nsew signal input
flabel metal2 s 55714 88000 55770 88800 0 FreeSans 224 90 0 0 io_north_in[19]
port 78 nsew signal input
flabel metal2 s 15786 88000 15842 88800 0 FreeSans 224 90 0 0 io_north_in[1]
port 79 nsew signal input
flabel metal2 s 57002 88000 57058 88800 0 FreeSans 224 90 0 0 io_north_in[20]
port 80 nsew signal input
flabel metal2 s 57646 88000 57702 88800 0 FreeSans 224 90 0 0 io_north_in[21]
port 81 nsew signal input
flabel metal2 s 58934 88000 58990 88800 0 FreeSans 224 90 0 0 io_north_in[22]
port 82 nsew signal input
flabel metal2 s 60222 88000 60278 88800 0 FreeSans 224 90 0 0 io_north_in[23]
port 83 nsew signal input
flabel metal2 s 61510 88000 61566 88800 0 FreeSans 224 90 0 0 io_north_in[24]
port 84 nsew signal input
flabel metal2 s 62154 88000 62210 88800 0 FreeSans 224 90 0 0 io_north_in[25]
port 85 nsew signal input
flabel metal2 s 63442 88000 63498 88800 0 FreeSans 224 90 0 0 io_north_in[26]
port 86 nsew signal input
flabel metal2 s 64730 88000 64786 88800 0 FreeSans 224 90 0 0 io_north_in[27]
port 87 nsew signal input
flabel metal2 s 65374 88000 65430 88800 0 FreeSans 224 90 0 0 io_north_in[28]
port 88 nsew signal input
flabel metal2 s 66662 88000 66718 88800 0 FreeSans 224 90 0 0 io_north_in[29]
port 89 nsew signal input
flabel metal2 s 17074 88000 17130 88800 0 FreeSans 224 90 0 0 io_north_in[2]
port 90 nsew signal input
flabel metal2 s 5482 1600 5538 2400 0 FreeSans 224 90 0 0 io_north_in[30]
port 91 nsew signal input
flabel metal2 s 6126 1600 6182 2400 0 FreeSans 224 90 0 0 io_north_in[31]
port 92 nsew signal input
flabel metal2 s 18362 88000 18418 88800 0 FreeSans 224 90 0 0 io_north_in[3]
port 93 nsew signal input
flabel metal2 s 19650 88000 19706 88800 0 FreeSans 224 90 0 0 io_north_in[4]
port 94 nsew signal input
flabel metal2 s 20294 88000 20350 88800 0 FreeSans 224 90 0 0 io_north_in[5]
port 95 nsew signal input
flabel metal2 s 21582 88000 21638 88800 0 FreeSans 224 90 0 0 io_north_in[6]
port 96 nsew signal input
flabel metal2 s 22870 88000 22926 88800 0 FreeSans 224 90 0 0 io_north_in[7]
port 97 nsew signal input
flabel metal2 s 23514 88000 23570 88800 0 FreeSans 224 90 0 0 io_north_in[8]
port 98 nsew signal input
flabel metal2 s 24802 88000 24858 88800 0 FreeSans 224 90 0 0 io_north_in[9]
port 99 nsew signal input
flabel metal2 s 30598 88000 30654 88800 0 FreeSans 224 90 0 0 io_north_out[0]
port 100 nsew signal output
flabel metal2 s 41546 88000 41602 88800 0 FreeSans 224 90 0 0 io_north_out[10]
port 101 nsew signal output
flabel metal2 s 42190 88000 42246 88800 0 FreeSans 224 90 0 0 io_north_out[11]
port 102 nsew signal output
flabel metal2 s 43478 88000 43534 88800 0 FreeSans 224 90 0 0 io_north_out[12]
port 103 nsew signal output
flabel metal2 s 44122 88000 44178 88800 0 FreeSans 224 90 0 0 io_north_out[13]
port 104 nsew signal output
flabel metal2 s 48630 88000 48686 88800 0 FreeSans 224 90 0 0 io_north_out[14]
port 105 nsew signal output
flabel metal3 s 89200 47848 90000 47968 0 FreeSans 480 0 0 0 io_north_out[15]
port 106 nsew signal output
flabel metal2 s 67950 88000 68006 88800 0 FreeSans 224 90 0 0 io_north_out[16]
port 107 nsew signal output
flabel metal2 s 69238 88000 69294 88800 0 FreeSans 224 90 0 0 io_north_out[17]
port 108 nsew signal output
flabel metal2 s 69882 88000 69938 88800 0 FreeSans 224 90 0 0 io_north_out[18]
port 109 nsew signal output
flabel metal2 s 71170 88000 71226 88800 0 FreeSans 224 90 0 0 io_north_out[19]
port 110 nsew signal output
flabel metal2 s 31242 88000 31298 88800 0 FreeSans 224 90 0 0 io_north_out[1]
port 111 nsew signal output
flabel metal2 s 72458 88000 72514 88800 0 FreeSans 224 90 0 0 io_north_out[20]
port 112 nsew signal output
flabel metal2 s 73102 88000 73158 88800 0 FreeSans 224 90 0 0 io_north_out[21]
port 113 nsew signal output
flabel metal2 s 74390 88000 74446 88800 0 FreeSans 224 90 0 0 io_north_out[22]
port 114 nsew signal output
flabel metal2 s 75678 88000 75734 88800 0 FreeSans 224 90 0 0 io_north_out[23]
port 115 nsew signal output
flabel metal2 s 76966 88000 77022 88800 0 FreeSans 224 90 0 0 io_north_out[24]
port 116 nsew signal output
flabel metal2 s 77610 88000 77666 88800 0 FreeSans 224 90 0 0 io_north_out[25]
port 117 nsew signal output
flabel metal2 s 78898 88000 78954 88800 0 FreeSans 224 90 0 0 io_north_out[26]
port 118 nsew signal output
flabel metal2 s 80186 88000 80242 88800 0 FreeSans 224 90 0 0 io_north_out[27]
port 119 nsew signal output
flabel metal2 s 80830 88000 80886 88800 0 FreeSans 224 90 0 0 io_north_out[28]
port 120 nsew signal output
flabel metal2 s 82118 88000 82174 88800 0 FreeSans 224 90 0 0 io_north_out[29]
port 121 nsew signal output
flabel metal2 s 32530 88000 32586 88800 0 FreeSans 224 90 0 0 io_north_out[2]
port 122 nsew signal output
flabel metal3 s 89200 45808 90000 45928 0 FreeSans 480 0 0 0 io_north_out[30]
port 123 nsew signal output
flabel metal2 s 44766 88000 44822 88800 0 FreeSans 224 90 0 0 io_north_out[31]
port 124 nsew signal output
flabel metal2 s 33818 88000 33874 88800 0 FreeSans 224 90 0 0 io_north_out[3]
port 125 nsew signal output
flabel metal2 s 35106 88000 35162 88800 0 FreeSans 224 90 0 0 io_north_out[4]
port 126 nsew signal output
flabel metal2 s 35750 88000 35806 88800 0 FreeSans 224 90 0 0 io_north_out[5]
port 127 nsew signal output
flabel metal2 s 37038 88000 37094 88800 0 FreeSans 224 90 0 0 io_north_out[6]
port 128 nsew signal output
flabel metal2 s 38326 88000 38382 88800 0 FreeSans 224 90 0 0 io_north_out[7]
port 129 nsew signal output
flabel metal2 s 38970 88000 39026 88800 0 FreeSans 224 90 0 0 io_north_out[8]
port 130 nsew signal output
flabel metal2 s 40258 88000 40314 88800 0 FreeSans 224 90 0 0 io_north_out[9]
port 131 nsew signal output
flabel metal2 s 30598 1600 30654 2400 0 FreeSans 224 90 0 0 io_south_in[0]
port 132 nsew signal input
flabel metal2 s 41546 1600 41602 2400 0 FreeSans 224 90 0 0 io_south_in[10]
port 133 nsew signal input
flabel metal2 s 42834 1600 42890 2400 0 FreeSans 224 90 0 0 io_south_in[11]
port 134 nsew signal input
flabel metal2 s 43478 1600 43534 2400 0 FreeSans 224 90 0 0 io_south_in[12]
port 135 nsew signal input
flabel metal2 s 44766 1600 44822 2400 0 FreeSans 224 90 0 0 io_south_in[13]
port 136 nsew signal input
flabel metal2 s 6770 1600 6826 2400 0 FreeSans 224 90 0 0 io_south_in[14]
port 137 nsew signal input
flabel metal2 s 7414 1600 7470 2400 0 FreeSans 224 90 0 0 io_south_in[15]
port 138 nsew signal input
flabel metal2 s 67950 1600 68006 2400 0 FreeSans 224 90 0 0 io_south_in[16]
port 139 nsew signal input
flabel metal2 s 69238 1600 69294 2400 0 FreeSans 224 90 0 0 io_south_in[17]
port 140 nsew signal input
flabel metal2 s 69882 1600 69938 2400 0 FreeSans 224 90 0 0 io_south_in[18]
port 141 nsew signal input
flabel metal2 s 71170 1600 71226 2400 0 FreeSans 224 90 0 0 io_south_in[19]
port 142 nsew signal input
flabel metal2 s 31242 1600 31298 2400 0 FreeSans 224 90 0 0 io_south_in[1]
port 143 nsew signal input
flabel metal2 s 72458 1600 72514 2400 0 FreeSans 224 90 0 0 io_south_in[20]
port 144 nsew signal input
flabel metal2 s 73102 1600 73158 2400 0 FreeSans 224 90 0 0 io_south_in[21]
port 145 nsew signal input
flabel metal2 s 74390 1600 74446 2400 0 FreeSans 224 90 0 0 io_south_in[22]
port 146 nsew signal input
flabel metal2 s 75678 1600 75734 2400 0 FreeSans 224 90 0 0 io_south_in[23]
port 147 nsew signal input
flabel metal2 s 76966 1600 77022 2400 0 FreeSans 224 90 0 0 io_south_in[24]
port 148 nsew signal input
flabel metal2 s 77610 1600 77666 2400 0 FreeSans 224 90 0 0 io_south_in[25]
port 149 nsew signal input
flabel metal2 s 78898 1600 78954 2400 0 FreeSans 224 90 0 0 io_south_in[26]
port 150 nsew signal input
flabel metal2 s 80186 1600 80242 2400 0 FreeSans 224 90 0 0 io_south_in[27]
port 151 nsew signal input
flabel metal3 s 89200 9768 90000 9888 0 FreeSans 480 0 0 0 io_south_in[28]
port 152 nsew signal input
flabel metal3 s 89200 10448 90000 10568 0 FreeSans 480 0 0 0 io_south_in[29]
port 153 nsew signal input
flabel metal2 s 32530 1600 32586 2400 0 FreeSans 224 90 0 0 io_south_in[2]
port 154 nsew signal input
flabel metal2 s 8058 1600 8114 2400 0 FreeSans 224 90 0 0 io_south_in[30]
port 155 nsew signal input
flabel metal2 s 8702 1600 8758 2400 0 FreeSans 224 90 0 0 io_south_in[31]
port 156 nsew signal input
flabel metal2 s 33818 1600 33874 2400 0 FreeSans 224 90 0 0 io_south_in[3]
port 157 nsew signal input
flabel metal2 s 35106 1600 35162 2400 0 FreeSans 224 90 0 0 io_south_in[4]
port 158 nsew signal input
flabel metal2 s 35750 1600 35806 2400 0 FreeSans 224 90 0 0 io_south_in[5]
port 159 nsew signal input
flabel metal2 s 37038 1600 37094 2400 0 FreeSans 224 90 0 0 io_south_in[6]
port 160 nsew signal input
flabel metal2 s 38326 1600 38382 2400 0 FreeSans 224 90 0 0 io_south_in[7]
port 161 nsew signal input
flabel metal2 s 38970 1600 39026 2400 0 FreeSans 224 90 0 0 io_south_in[8]
port 162 nsew signal input
flabel metal2 s 40258 1600 40314 2400 0 FreeSans 224 90 0 0 io_south_in[9]
port 163 nsew signal input
flabel metal2 s 15142 1600 15198 2400 0 FreeSans 224 90 0 0 io_south_out[0]
port 164 nsew signal output
flabel metal2 s 26090 1600 26146 2400 0 FreeSans 224 90 0 0 io_south_out[10]
port 165 nsew signal output
flabel metal2 s 27378 1600 27434 2400 0 FreeSans 224 90 0 0 io_south_out[11]
port 166 nsew signal output
flabel metal2 s 28022 1600 28078 2400 0 FreeSans 224 90 0 0 io_south_out[12]
port 167 nsew signal output
flabel metal2 s 29310 1600 29366 2400 0 FreeSans 224 90 0 0 io_south_out[13]
port 168 nsew signal output
flabel metal2 s 45410 88000 45466 88800 0 FreeSans 224 90 0 0 io_south_out[14]
port 169 nsew signal output
flabel metal2 s 46698 88000 46754 88800 0 FreeSans 224 90 0 0 io_south_out[15]
port 170 nsew signal output
flabel metal2 s 52494 1600 52550 2400 0 FreeSans 224 90 0 0 io_south_out[16]
port 171 nsew signal output
flabel metal2 s 53782 1600 53838 2400 0 FreeSans 224 90 0 0 io_south_out[17]
port 172 nsew signal output
flabel metal2 s 54426 1600 54482 2400 0 FreeSans 224 90 0 0 io_south_out[18]
port 173 nsew signal output
flabel metal2 s 55714 1600 55770 2400 0 FreeSans 224 90 0 0 io_south_out[19]
port 174 nsew signal output
flabel metal2 s 15786 1600 15842 2400 0 FreeSans 224 90 0 0 io_south_out[1]
port 175 nsew signal output
flabel metal2 s 57002 1600 57058 2400 0 FreeSans 224 90 0 0 io_south_out[20]
port 176 nsew signal output
flabel metal2 s 57646 1600 57702 2400 0 FreeSans 224 90 0 0 io_south_out[21]
port 177 nsew signal output
flabel metal2 s 58934 1600 58990 2400 0 FreeSans 224 90 0 0 io_south_out[22]
port 178 nsew signal output
flabel metal2 s 60222 1600 60278 2400 0 FreeSans 224 90 0 0 io_south_out[23]
port 179 nsew signal output
flabel metal2 s 61510 1600 61566 2400 0 FreeSans 224 90 0 0 io_south_out[24]
port 180 nsew signal output
flabel metal2 s 62154 1600 62210 2400 0 FreeSans 224 90 0 0 io_south_out[25]
port 181 nsew signal output
flabel metal2 s 63442 1600 63498 2400 0 FreeSans 224 90 0 0 io_south_out[26]
port 182 nsew signal output
flabel metal2 s 64730 1600 64786 2400 0 FreeSans 224 90 0 0 io_south_out[27]
port 183 nsew signal output
flabel metal2 s 65374 1600 65430 2400 0 FreeSans 224 90 0 0 io_south_out[28]
port 184 nsew signal output
flabel metal2 s 66662 1600 66718 2400 0 FreeSans 224 90 0 0 io_south_out[29]
port 185 nsew signal output
flabel metal2 s 17074 1600 17130 2400 0 FreeSans 224 90 0 0 io_south_out[2]
port 186 nsew signal output
flabel metal3 s 89200 45128 90000 45248 0 FreeSans 480 0 0 0 io_south_out[30]
port 187 nsew signal output
flabel metal3 s 89200 46488 90000 46608 0 FreeSans 480 0 0 0 io_south_out[31]
port 188 nsew signal output
flabel metal2 s 18362 1600 18418 2400 0 FreeSans 224 90 0 0 io_south_out[3]
port 189 nsew signal output
flabel metal2 s 19650 1600 19706 2400 0 FreeSans 224 90 0 0 io_south_out[4]
port 190 nsew signal output
flabel metal2 s 20294 1600 20350 2400 0 FreeSans 224 90 0 0 io_south_out[5]
port 191 nsew signal output
flabel metal2 s 21582 1600 21638 2400 0 FreeSans 224 90 0 0 io_south_out[6]
port 192 nsew signal output
flabel metal2 s 22870 1600 22926 2400 0 FreeSans 224 90 0 0 io_south_out[7]
port 193 nsew signal output
flabel metal2 s 23514 1600 23570 2400 0 FreeSans 224 90 0 0 io_south_out[8]
port 194 nsew signal output
flabel metal2 s 24802 1600 24858 2400 0 FreeSans 224 90 0 0 io_south_out[9]
port 195 nsew signal output
flabel metal3 s 1600 15208 2400 15328 0 FreeSans 480 0 0 0 io_west_in[0]
port 196 nsew signal input
flabel metal3 s 1600 26088 2400 26208 0 FreeSans 480 0 0 0 io_west_in[10]
port 197 nsew signal input
flabel metal3 s 1600 27448 2400 27568 0 FreeSans 480 0 0 0 io_west_in[11]
port 198 nsew signal input
flabel metal3 s 1600 28128 2400 28248 0 FreeSans 480 0 0 0 io_west_in[12]
port 199 nsew signal input
flabel metal3 s 1600 29488 2400 29608 0 FreeSans 480 0 0 0 io_west_in[13]
port 200 nsew signal input
flabel metal2 s 9346 1600 9402 2400 0 FreeSans 224 90 0 0 io_west_in[14]
port 201 nsew signal input
flabel metal2 s 9990 1600 10046 2400 0 FreeSans 224 90 0 0 io_west_in[15]
port 202 nsew signal input
flabel metal3 s 1600 51248 2400 51368 0 FreeSans 480 0 0 0 io_west_in[16]
port 203 nsew signal input
flabel metal3 s 1600 52608 2400 52728 0 FreeSans 480 0 0 0 io_west_in[17]
port 204 nsew signal input
flabel metal3 s 1600 53968 2400 54088 0 FreeSans 480 0 0 0 io_west_in[18]
port 205 nsew signal input
flabel metal3 s 1600 54648 2400 54768 0 FreeSans 480 0 0 0 io_west_in[19]
port 206 nsew signal input
flabel metal3 s 1600 16568 2400 16688 0 FreeSans 480 0 0 0 io_west_in[1]
port 207 nsew signal input
flabel metal3 s 1600 56008 2400 56128 0 FreeSans 480 0 0 0 io_west_in[20]
port 208 nsew signal input
flabel metal3 s 1600 56688 2400 56808 0 FreeSans 480 0 0 0 io_west_in[21]
port 209 nsew signal input
flabel metal3 s 1600 58048 2400 58168 0 FreeSans 480 0 0 0 io_west_in[22]
port 210 nsew signal input
flabel metal3 s 1600 59408 2400 59528 0 FreeSans 480 0 0 0 io_west_in[23]
port 211 nsew signal input
flabel metal3 s 1600 60088 2400 60208 0 FreeSans 480 0 0 0 io_west_in[24]
port 212 nsew signal input
flabel metal3 s 1600 61448 2400 61568 0 FreeSans 480 0 0 0 io_west_in[25]
port 213 nsew signal input
flabel metal3 s 1600 62128 2400 62248 0 FreeSans 480 0 0 0 io_west_in[26]
port 214 nsew signal input
flabel metal3 s 1600 63488 2400 63608 0 FreeSans 480 0 0 0 io_west_in[27]
port 215 nsew signal input
flabel metal3 s 1600 64848 2400 64968 0 FreeSans 480 0 0 0 io_west_in[28]
port 216 nsew signal input
flabel metal3 s 1600 65528 2400 65648 0 FreeSans 480 0 0 0 io_west_in[29]
port 217 nsew signal input
flabel metal3 s 1600 17248 2400 17368 0 FreeSans 480 0 0 0 io_west_in[2]
port 218 nsew signal input
flabel metal2 s 10634 1600 10690 2400 0 FreeSans 224 90 0 0 io_west_in[30]
port 219 nsew signal input
flabel metal2 s 11278 1600 11334 2400 0 FreeSans 224 90 0 0 io_west_in[31]
port 220 nsew signal input
flabel metal3 s 1600 18608 2400 18728 0 FreeSans 480 0 0 0 io_west_in[3]
port 221 nsew signal input
flabel metal3 s 1600 19288 2400 19408 0 FreeSans 480 0 0 0 io_west_in[4]
port 222 nsew signal input
flabel metal3 s 1600 20648 2400 20768 0 FreeSans 480 0 0 0 io_west_in[5]
port 223 nsew signal input
flabel metal3 s 1600 22008 2400 22128 0 FreeSans 480 0 0 0 io_west_in[6]
port 224 nsew signal input
flabel metal3 s 1600 22688 2400 22808 0 FreeSans 480 0 0 0 io_west_in[7]
port 225 nsew signal input
flabel metal3 s 1600 24048 2400 24168 0 FreeSans 480 0 0 0 io_west_in[8]
port 226 nsew signal input
flabel metal3 s 1600 24728 2400 24848 0 FreeSans 480 0 0 0 io_west_in[9]
port 227 nsew signal input
flabel metal3 s 1600 30168 2400 30288 0 FreeSans 480 0 0 0 io_west_out[0]
port 228 nsew signal output
flabel metal3 s 1600 41048 2400 41168 0 FreeSans 480 0 0 0 io_west_out[10]
port 229 nsew signal output
flabel metal3 s 1600 42408 2400 42528 0 FreeSans 480 0 0 0 io_west_out[11]
port 230 nsew signal output
flabel metal3 s 1600 43768 2400 43888 0 FreeSans 480 0 0 0 io_west_out[12]
port 231 nsew signal output
flabel metal3 s 1600 44448 2400 44568 0 FreeSans 480 0 0 0 io_west_out[13]
port 232 nsew signal output
flabel metal2 s 46054 88000 46110 88800 0 FreeSans 224 90 0 0 io_west_out[14]
port 233 nsew signal output
flabel metal3 s 89200 48528 90000 48648 0 FreeSans 480 0 0 0 io_west_out[15]
port 234 nsew signal output
flabel metal3 s 1600 66888 2400 67008 0 FreeSans 480 0 0 0 io_west_out[16]
port 235 nsew signal output
flabel metal3 s 1600 67568 2400 67688 0 FreeSans 480 0 0 0 io_west_out[17]
port 236 nsew signal output
flabel metal3 s 1600 68928 2400 69048 0 FreeSans 480 0 0 0 io_west_out[18]
port 237 nsew signal output
flabel metal3 s 1600 70288 2400 70408 0 FreeSans 480 0 0 0 io_west_out[19]
port 238 nsew signal output
flabel metal3 s 1600 31528 2400 31648 0 FreeSans 480 0 0 0 io_west_out[1]
port 239 nsew signal output
flabel metal3 s 1600 70968 2400 71088 0 FreeSans 480 0 0 0 io_west_out[20]
port 240 nsew signal output
flabel metal3 s 1600 72328 2400 72448 0 FreeSans 480 0 0 0 io_west_out[21]
port 241 nsew signal output
flabel metal3 s 1600 73008 2400 73128 0 FreeSans 480 0 0 0 io_west_out[22]
port 242 nsew signal output
flabel metal3 s 1600 74368 2400 74488 0 FreeSans 480 0 0 0 io_west_out[23]
port 243 nsew signal output
flabel metal3 s 1600 75728 2400 75848 0 FreeSans 480 0 0 0 io_west_out[24]
port 244 nsew signal output
flabel metal3 s 1600 76408 2400 76528 0 FreeSans 480 0 0 0 io_west_out[25]
port 245 nsew signal output
flabel metal3 s 1600 77768 2400 77888 0 FreeSans 480 0 0 0 io_west_out[26]
port 246 nsew signal output
flabel metal3 s 1600 78448 2400 78568 0 FreeSans 480 0 0 0 io_west_out[27]
port 247 nsew signal output
flabel metal3 s 1600 79808 2400 79928 0 FreeSans 480 0 0 0 io_west_out[28]
port 248 nsew signal output
flabel metal2 s 10634 88000 10690 88800 0 FreeSans 224 90 0 0 io_west_out[29]
port 249 nsew signal output
flabel metal3 s 1600 32888 2400 33008 0 FreeSans 480 0 0 0 io_west_out[2]
port 250 nsew signal output
flabel metal2 s 49274 88000 49330 88800 0 FreeSans 224 90 0 0 io_west_out[30]
port 251 nsew signal output
flabel metal2 s 47986 88000 48042 88800 0 FreeSans 224 90 0 0 io_west_out[31]
port 252 nsew signal output
flabel metal3 s 1600 33568 2400 33688 0 FreeSans 480 0 0 0 io_west_out[3]
port 253 nsew signal output
flabel metal3 s 1600 34928 2400 35048 0 FreeSans 480 0 0 0 io_west_out[4]
port 254 nsew signal output
flabel metal3 s 1600 35608 2400 35728 0 FreeSans 480 0 0 0 io_west_out[5]
port 255 nsew signal output
flabel metal3 s 1600 36968 2400 37088 0 FreeSans 480 0 0 0 io_west_out[6]
port 256 nsew signal output
flabel metal3 s 1600 38328 2400 38448 0 FreeSans 480 0 0 0 io_west_out[7]
port 257 nsew signal output
flabel metal3 s 1600 39008 2400 39128 0 FreeSans 480 0 0 0 io_west_out[8]
port 258 nsew signal output
flabel metal3 s 1600 40368 2400 40488 0 FreeSans 480 0 0 0 io_west_out[9]
port 259 nsew signal output
flabel metal3 s 89200 12488 90000 12608 0 FreeSans 480 0 0 0 le_clk
port 260 nsew signal input
flabel metal3 s 89200 13168 90000 13288 0 FreeSans 480 0 0 0 le_en
port 261 nsew signal input
flabel metal3 s 89200 14528 90000 14648 0 FreeSans 480 0 0 0 le_nrst
port 262 nsew signal input
flabel metal2 s 40902 88000 40958 88800 0 FreeSans 224 90 0 0 nrst
port 263 nsew signal input
flabel metal4 s 3356 3376 3676 89104 0 FreeSans 1920 90 0 0 vccd1
port 264 nsew power bidirectional
flabel metal5 s 3356 3376 90116 3696 0 FreeSans 2560 0 0 0 vccd1
port 264 nsew power bidirectional
flabel metal5 s 3356 88784 90116 89104 0 FreeSans 2560 0 0 0 vccd1
port 264 nsew power bidirectional
flabel metal4 s 89796 3376 90116 89104 0 FreeSans 1920 90 0 0 vccd1
port 264 nsew power bidirectional
flabel metal4 s 17716 2716 18036 10187 0 FreeSans 1920 90 0 0 vccd1
port 264 nsew power bidirectional
flabel metal4 s 17716 81029 18036 89764 0 FreeSans 1920 90 0 0 vccd1
port 264 nsew power bidirectional
flabel metal4 s 36116 2716 36436 10187 0 FreeSans 1920 90 0 0 vccd1
port 264 nsew power bidirectional
flabel metal4 s 36116 81029 36436 89764 0 FreeSans 1920 90 0 0 vccd1
port 264 nsew power bidirectional
flabel metal4 s 54516 2716 54836 10187 0 FreeSans 1920 90 0 0 vccd1
port 264 nsew power bidirectional
flabel metal4 s 54516 81029 54836 89764 0 FreeSans 1920 90 0 0 vccd1
port 264 nsew power bidirectional
flabel metal4 s 72916 2716 73236 10187 0 FreeSans 1920 90 0 0 vccd1
port 264 nsew power bidirectional
flabel metal4 s 72916 81029 73236 89764 0 FreeSans 1920 90 0 0 vccd1
port 264 nsew power bidirectional
flabel metal5 s 2696 17736 90776 18056 0 FreeSans 2560 0 0 0 vccd1
port 264 nsew power bidirectional
flabel metal5 s 2696 36136 90776 36456 0 FreeSans 2560 0 0 0 vccd1
port 264 nsew power bidirectional
flabel metal5 s 2696 54536 90776 54856 0 FreeSans 2560 0 0 0 vccd1
port 264 nsew power bidirectional
flabel metal5 s 2696 72936 90776 73256 0 FreeSans 2560 0 0 0 vccd1
port 264 nsew power bidirectional
flabel metal4 s 5948 7024 6268 84912 0 FreeSans 1920 90 0 0 vccd1
port 264 nsew power bidirectional
flabel metal4 s 86540 7024 86860 84912 0 FreeSans 1920 90 0 0 vccd1
port 264 nsew power bidirectional
flabel metal4 s 2696 2716 3016 89764 0 FreeSans 1920 90 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal5 s 2696 2716 90776 3036 0 FreeSans 2560 0 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal5 s 2696 89444 90776 89764 0 FreeSans 2560 0 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal4 s 90456 2716 90776 89764 0 FreeSans 1920 90 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal4 s 18376 2716 18696 10187 0 FreeSans 1920 90 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal4 s 18376 81029 18696 89764 0 FreeSans 1920 90 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal4 s 36776 2716 37096 10187 0 FreeSans 1920 90 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal4 s 36776 81029 37096 89764 0 FreeSans 1920 90 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal4 s 55176 2716 55496 10187 0 FreeSans 1920 90 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal4 s 55176 81029 55496 89764 0 FreeSans 1920 90 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal4 s 73576 2716 73896 10187 0 FreeSans 1920 90 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal4 s 73576 81029 73896 89764 0 FreeSans 1920 90 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal5 s 2696 18396 90776 18716 0 FreeSans 2560 0 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal5 s 2696 36796 90776 37116 0 FreeSans 2560 0 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal5 s 2696 55196 90776 55516 0 FreeSans 2560 0 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal5 s 2696 73596 90776 73916 0 FreeSans 2560 0 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal4 s 6684 7024 7004 84912 0 FreeSans 1920 90 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal4 s 87276 7024 87596 84912 0 FreeSans 1920 90 0 0 vssd1
port 265 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 1600 1600 90000 88800
<< end >>
