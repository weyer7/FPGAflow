* NGSPICE file created from top.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

.subckt top VGND VPWR clk keypad_i[0] keypad_i[10] keypad_i[11] keypad_i[12] keypad_i[13]
+ keypad_i[1] keypad_i[2] keypad_i[3] keypad_i[4] keypad_i[5] keypad_i[6] keypad_i[7]
+ keypad_i[8] keypad_i[9] n_rst pwm
XTAP_TAPCELL_ROW_17_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0985_ clknet_4_0_0_clk _0048_ net47 VGND VGND VPWR VPWR waveshape.seq_div.dividend\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0770_ net81 _0323_ _0326_ VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__a21oi_1
XFILLER_5_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0968_ clknet_4_13_0_clk net73 net59 VGND VGND VPWR VPWR pwm_counter.active_sample\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_34_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_12_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_12_0_clk sky130_fd_sc_hd__clkbuf_8
X_0899_ _0404_ _0427_ _0414_ VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__o21bai_1
XTAP_TAPCELL_ROW_25_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0822_ _0115_ _0190_ VGND VGND VPWR VPWR _0366_ sky130_fd_sc_hd__and2_1
X_0753_ net78 pwm_counter.active_sample\[0\] _0197_ VGND VGND VPWR VPWR _0028_ sky130_fd_sc_hd__mux2_1
X_0684_ net147 _0278_ _0279_ _0284_ _0282_ VGND VGND VPWR VPWR waveshape.shaper.n_sample\[2\]
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_39_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Left_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1021_ clknet_4_11_0_clk net10 net54 VGND VGND VPWR VPWR keypad.keypad_reg\[5\] sky130_fd_sc_hd__dfrtp_1
X_0805_ _0163_ _0184_ VGND VGND VPWR VPWR _0353_ sky130_fd_sc_hd__nor2_1
X_0667_ _0271_ net121 VGND VGND VPWR VPWR pwm_counter.n_count\[5\] sky130_fd_sc_hd__nor2_1
X_0598_ count\[13\] _0100_ _0109_ count\[12\] VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__a22o_1
X_0736_ net45 waveshape.seq_div.dividend\[15\] net29 count\[8\] net19 VGND VGND VPWR
+ VPWR _0314_ sky130_fd_sc_hd__a221o_1
XFILLER_44_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold41 waveshape.seq_div.state\[1\] VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 freq_div.keycode\[3\] VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 waveshape.seq_div.dividend\[24\] VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__dlygate4sd3_1
Xhold30 waveshape.seq_div.dividend\[12\] VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 waveshape.scaled_count\[3\] VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0452_ sample_rate.count\[5\] sample_rate.count\[4\] _0091_ VGND VGND VPWR VPWR _0092_
+ sky130_fd_sc_hd__and3_1
XFILLER_6_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0521_ waveshape.seq_div.dividend\[28\] _0122_ _0148_ _0146_ VGND VGND VPWR VPWR
+ _0160_ sky130_fd_sc_hd__a31o_1
XFILLER_13_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1004_ clknet_4_13_0_clk pwm_counter.n_count\[2\] net59 VGND VGND VPWR VPWR pwm_counter.count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_34_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0719_ net45 waveshape.scaled_count\[6\] net23 VGND VGND VPWR VPWR _0306_ sky130_fd_sc_hd__and3_1
XFILLER_25_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0435_ pwm_counter.count\[6\] VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__inv_2
X_0504_ _0131_ _0142_ VGND VGND VPWR VPWR _0143_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_17_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_37_Left_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0984_ clknet_4_0_0_clk _0047_ net47 VGND VGND VPWR VPWR waveshape.seq_div.dividend\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0967_ clknet_4_13_0_clk net77 net61 VGND VGND VPWR VPWR pwm_counter.active_sample\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_34_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0898_ keypad.keypad_reg\[4\] keypad.keypad_reg\[5\] keypad.keypad_reg\[6\] keypad.keypad_reg\[7\]
+ VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__or4b_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0821_ net133 net26 _0362_ _0365_ VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__a22o_1
X_0752_ net145 net25 net21 VGND VGND VPWR VPWR _0027_ sky130_fd_sc_hd__o21a_1
XFILLER_43_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0683_ waveshape.scaled_count\[7\] waveshape.scaled_count\[1\] VGND VGND VPWR VPWR
+ _0284_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_24_Left_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_4_11_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_11_0_clk sky130_fd_sc_hd__clkbuf_8
X_1020_ clknet_4_11_0_clk net9 net53 VGND VGND VPWR VPWR keypad.keypad_reg\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0804_ waveshape.seq_div.dividend\[31\] net24 _0351_ _0352_ VGND VGND VPWR VPWR _0048_
+ sky130_fd_sc_hd__o22a_1
X_0735_ net103 net22 _0313_ VGND VGND VPWR VPWR _0018_ sky130_fd_sc_hd__o21a_1
X_0666_ pwm_counter.count\[4\] _0270_ net120 VGND VGND VPWR VPWR _0275_ sky130_fd_sc_hd__a21oi_1
X_0597_ count\[11\] _0165_ _0169_ count\[10\] VGND VGND VPWR VPWR _0232_ sky130_fd_sc_hd__a22o_1
Xhold42 _0036_ VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 waveshape.seq_div.dividend\[9\] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 waveshape.seq_div.dividend\[8\] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 waveshape.scaled_count\[6\] VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 waveshape.seq_div.dividend\[38\] VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 waveshape.scaled_count\[4\] VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_43_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0451_ sample_rate.count\[3\] _0090_ VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__and2_1
X_0520_ _0149_ _0153_ _0158_ VGND VGND VPWR VPWR _0159_ sky130_fd_sc_hd__nand3_1
X_1003_ clknet_4_13_0_clk pwm_counter.n_count\[1\] net61 VGND VGND VPWR VPWR pwm_counter.count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_19_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0718_ net140 net20 _0305_ VGND VGND VPWR VPWR _0009_ sky130_fd_sc_hd__a21o_1
X_0649_ _0091_ _0101_ VGND VGND VPWR VPWR _0266_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_11_Left_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0434_ pwm_counter.count\[7\] VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__inv_2
XFILLER_39_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_235 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0503_ _0134_ _0140_ _0141_ VGND VGND VPWR VPWR _0142_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_17_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0983_ clknet_4_0_0_clk _0046_ net46 VGND VGND VPWR VPWR waveshape.seq_div.dividend\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_6_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_131 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0966_ clknet_4_13_0_clk net84 net56 VGND VGND VPWR VPWR pwm_counter.active_sample\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_0897_ _0407_ _0419_ _0426_ _0214_ net33 VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__o32a_1
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0751_ net98 net23 _0321_ VGND VGND VPWR VPWR _0026_ sky130_fd_sc_hd__o21a_1
X_0820_ net40 waveshape.seq_div.dividend\[34\] _0364_ net39 VGND VGND VPWR VPWR _0365_
+ sky130_fd_sc_hd__a22o_1
XFILLER_36_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0682_ net149 _0278_ _0279_ _0283_ _0282_ VGND VGND VPWR VPWR waveshape.shaper.n_sample\[1\]
+ sky130_fd_sc_hd__a221o_1
XFILLER_49_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0949_ clknet_4_3_0_clk _0020_ net57 VGND VGND VPWR VPWR waveshape.seq_div.dividend\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_41_Left_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_55 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0665_ _0077_ _0270_ VGND VGND VPWR VPWR pwm_counter.n_count\[4\] sky130_fd_sc_hd__xnor2_1
X_0803_ net37 _0349_ _0350_ net27 VGND VGND VPWR VPWR _0352_ sky130_fd_sc_hd__a31o_1
X_0734_ net45 waveshape.seq_div.dividend\[14\] net29 count\[7\] net19 VGND VGND VPWR
+ VPWR _0313_ sky130_fd_sc_hd__a221o_1
X_0596_ _0227_ _0229_ _0230_ VGND VGND VPWR VPWR _0231_ sky130_fd_sc_hd__o21a_1
XFILLER_29_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold65 sample_rate.count\[4\] VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 sample_rate.count\[1\] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 _0032_ VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 waveshape.scaled_count\[0\] VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 waveshape.seq_div.state\[0\] VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 freq_div.keycode\[0\] VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 waveshape.seq_div.dividend\[11\] VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0450_ sample_rate.count\[1\] sample_rate.count\[0\] sample_rate.count\[2\] VGND
+ VGND VPWR VPWR _0090_ sky130_fd_sc_hd__and3_1
XFILLER_3_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1002_ clknet_4_15_0_clk pwm_counter.n_count\[0\] net59 VGND VGND VPWR VPWR pwm_counter.count\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_0648_ _0090_ _0101_ _0265_ VGND VGND VPWR VPWR sample_rate.n_count\[2\] sky130_fd_sc_hd__nor3_1
X_0717_ net45 waveshape.scaled_count\[5\] _0298_ VGND VGND VPWR VPWR _0305_ sky130_fd_sc_hd__and3_1
X_0579_ _0214_ VGND VGND VPWR VPWR keypad.n_modekey sky130_fd_sc_hd__inv_2
XFILLER_25_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_10_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_10_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0502_ waveshape.seq_div.dividend\[26\] _0130_ VGND VGND VPWR VPWR _0141_ sky130_fd_sc_hd__xor2_1
XFILLER_39_247 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0433_ waveshape.seq_div.dividend\[45\] VGND VGND VPWR VPWR _0073_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_17_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0982_ clknet_4_2_0_clk _0045_ net46 VGND VGND VPWR VPWR waveshape.seq_div.dividend\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_76 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_19_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0965_ clknet_4_13_0_clk net79 net56 VGND VGND VPWR VPWR pwm_counter.active_sample\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_0896_ keypad.keypad_reg\[3\] _0206_ _0415_ _0425_ VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_33_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_67 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0681_ waveshape.scaled_count\[0\] waveshape.scaled_count\[7\] VGND VGND VPWR VPWR
+ _0283_ sky130_fd_sc_hd__xor2_1
X_0750_ net40 waveshape.seq_div.dividend\[22\] net28 count\[15\] net21 VGND VGND VPWR
+ VPWR _0321_ sky130_fd_sc_hd__a221o_1
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_47_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0948_ clknet_4_9_0_clk _0019_ net55 VGND VGND VPWR VPWR waveshape.seq_div.dividend\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_22_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0879_ _0408_ _0410_ _0210_ VGND VGND VPWR VPWR _0411_ sky130_fd_sc_hd__o21a_1
XFILLER_18_67 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0802_ net40 waveshape.seq_div.dividend\[30\] VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__and2_1
X_0664_ _0270_ _0274_ VGND VGND VPWR VPWR pwm_counter.n_count\[3\] sky130_fd_sc_hd__nor2_1
X_0733_ net102 net22 _0312_ VGND VGND VPWR VPWR _0017_ sky130_fd_sc_hd__o21a_1
X_0595_ count\[10\] _0169_ _0225_ _0228_ VGND VGND VPWR VPWR _0230_ sky130_fd_sc_hd__o22a_1
Xhold22 sample_rate.n_count\[1\] VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__dlygate4sd3_1
Xhold11 pwm_counter.sample\[2\] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 pwm_counter.count\[5\] VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 pwm_counter.active_sample\[7\] VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 count\[4\] VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 waveshape.seq_div.dividend\[23\] VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 waveshape.scaled_count\[2\] VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1001_ clknet_4_5_0_clk _0064_ net50 VGND VGND VPWR VPWR waveshape.seq_div.dividend\[47\]
+ sky130_fd_sc_hd__dfrtp_1
X_0647_ sample_rate.count\[1\] sample_rate.count\[0\] net127 VGND VGND VPWR VPWR _0265_
+ sky130_fd_sc_hd__a21oi_1
X_0578_ keypad.keypad_reg\[12\] _0085_ _0211_ _0213_ VGND VGND VPWR VPWR _0214_ sky130_fd_sc_hd__or4_2
X_0716_ net132 net20 _0304_ VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__a21o_1
XFILLER_0_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0501_ waveshape.seq_div.dividend\[24\] _0137_ _0139_ VGND VGND VPWR VPWR _0140_
+ sky130_fd_sc_hd__o21ba_1
X_0432_ net37 VGND VGND VPWR VPWR _0072_ sky130_fd_sc_hd__inv_2
XFILLER_47_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0981_ clknet_4_2_0_clk _0044_ net46 VGND VGND VPWR VPWR waveshape.seq_div.dividend\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_88 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0964_ clknet_4_6_0_clk _0027_ net49 VGND VGND VPWR VPWR waveshape.scaled_count\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_0895_ _0408_ _0424_ _0210_ VGND VGND VPWR VPWR _0425_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_33_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0680_ net141 _0278_ _0282_ VGND VGND VPWR VPWR waveshape.shaper.n_sample\[0\] sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_47_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0947_ clknet_4_9_0_clk _0018_ net55 VGND VGND VPWR VPWR waveshape.seq_div.dividend\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_22_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0878_ _0402_ _0409_ VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__nor2_1
XFILLER_18_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload0 clknet_4_0_0_clk VGND VGND VPWR VPWR clkload0/Y sky130_fd_sc_hd__clkinv_2
XFILLER_46_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_28_Left_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0801_ _0157_ _0345_ _0153_ VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__o21ai_1
X_0663_ net125 _0269_ VGND VGND VPWR VPWR _0274_ sky130_fd_sc_hd__nor2_1
XFILLER_41_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0594_ count\[9\] _0176_ _0181_ count\[8\] VGND VGND VPWR VPWR _0229_ sky130_fd_sc_hd__a22o_1
X_0732_ net45 waveshape.seq_div.dividend\[13\] net29 count\[6\] net19 VGND VGND VPWR
+ VPWR _0312_ sky130_fd_sc_hd__a221o_1
XFILLER_37_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold56 _0275_ VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 waveshape.seq_div.n\[3\] VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 _0030_ VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 count\[7\] VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 waveshape.seq_div.dividend\[13\] VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold78 waveshape.seq_div.dividend\[30\] VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 waveshape.scaled_count\[5\] VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_41_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1000_ clknet_4_4_0_clk _0063_ net51 VGND VGND VPWR VPWR waveshape.seq_div.dividend\[46\]
+ sky130_fd_sc_hd__dfrtp_1
X_0715_ net44 waveshape.scaled_count\[4\] _0298_ VGND VGND VPWR VPWR _0304_ sky130_fd_sc_hd__and3_1
X_0646_ net86 sample_rate.count\[0\] _0264_ VGND VGND VPWR VPWR sample_rate.n_count\[1\]
+ sky130_fd_sc_hd__a21oi_1
X_0577_ keypad.keypad_reg\[8\] keypad.keypad_reg\[9\] keypad.keypad_reg\[11\] keypad.keypad_reg\[10\]
+ VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__or4_1
XFILLER_40_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0431_ net119 VGND VGND VPWR VPWR _0071_ sky130_fd_sc_hd__inv_2
X_0500_ waveshape.seq_div.dividend\[25\] _0133_ VGND VGND VPWR VPWR _0139_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Left_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0629_ _0253_ _0254_ VGND VGND VPWR VPWR oscill.n_count\[9\] sky130_fd_sc_hd__nor2_1
XFILLER_13_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0980_ clknet_4_2_0_clk _0043_ net46 VGND VGND VPWR VPWR waveshape.seq_div.dividend\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0894_ keypad.keypad_reg\[8\] keypad.keypad_reg\[9\] keypad.keypad_reg\[11\] _0403_
+ VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__and4bb_1
X_0963_ clknet_4_14_0_clk waveshape.shaper.n_sample\[7\] net58 VGND VGND VPWR VPWR
+ pwm_counter.sample\[7\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_2_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0877_ keypad.keypad_reg\[8\] keypad.keypad_reg\[9\] keypad.keypad_reg\[11\] keypad.keypad_reg\[10\]
+ VGND VGND VPWR VPWR _0409_ sky130_fd_sc_hd__or4b_1
XFILLER_9_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0946_ clknet_4_9_0_clk _0017_ net55 VGND VGND VPWR VPWR waveshape.seq_div.dividend\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload1 clknet_4_1_0_clk VGND VGND VPWR VPWR clkload1/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_3_Left_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0800_ _0153_ _0157_ _0345_ VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__or3_1
X_0731_ net99 net22 _0311_ VGND VGND VPWR VPWR _0016_ sky130_fd_sc_hd__o21a_1
X_0662_ _0269_ _0273_ VGND VGND VPWR VPWR pwm_counter.n_count\[2\] sky130_fd_sc_hd__nor2_1
XFILLER_34_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0593_ count\[8\] _0181_ VGND VGND VPWR VPWR _0228_ sky130_fd_sc_hd__nand2_1
XFILLER_37_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0929_ clknet_4_7_0_clk sample_rate.n_count\[4\] net50 VGND VGND VPWR VPWR sample_rate.count\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_20_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_45_Left_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold46 sample_rate.count\[3\] VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 _0039_ VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 pwm_counter.count\[2\] VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__dlygate4sd3_1
Xhold13 pwm_counter.sample\[0\] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 waveshape.seq_div.dividend\[35\] VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 waveshape.seq_div.dividend\[17\] VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold79 waveshape.seq_div.dividend\[42\] VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0645_ sample_rate.count\[1\] sample_rate.count\[0\] _0263_ VGND VGND VPWR VPWR _0264_
+ sky130_fd_sc_hd__o21ai_1
X_0714_ net129 net19 _0303_ VGND VGND VPWR VPWR _0007_ sky130_fd_sc_hd__a21o_1
X_0576_ keypad.keypad_reg\[8\] keypad.keypad_reg\[11\] VGND VGND VPWR VPWR _0212_
+ sky130_fd_sc_hd__nor2_1
XFILLER_15_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_139 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0430_ net34 VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__inv_2
XFILLER_47_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0628_ count\[9\] _0251_ net17 VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__o21ai_1
X_0559_ _0088_ _0196_ VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__nand2_4
XFILLER_26_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_32_Left_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0962_ clknet_4_14_0_clk waveshape.shaper.n_sample\[6\] net58 VGND VGND VPWR VPWR
+ pwm_counter.sample\[6\] sky130_fd_sc_hd__dfrtp_1
X_0893_ _0419_ _0421_ _0423_ _0214_ net35 VGND VGND VPWR VPWR _0066_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_2_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout60 net61 VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__clkbuf_2
XFILLER_49_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0876_ keypad.keypad_reg\[13\] _0213_ keypad.keypad_reg\[12\] VGND VGND VPWR VPWR
+ _0408_ sky130_fd_sc_hd__nor3b_1
XFILLER_9_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0945_ clknet_4_11_0_clk _0016_ net53 VGND VGND VPWR VPWR waveshape.seq_div.dividend\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_18_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload2 clknet_4_2_0_clk VGND VGND VPWR VPWR clkload2/Y sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_21_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0661_ pwm_counter.count\[1\] pwm_counter.count\[0\] net122 VGND VGND VPWR VPWR _0273_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_6_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0730_ net45 waveshape.seq_div.dividend\[12\] net29 count\[5\] net19 VGND VGND VPWR
+ VPWR _0311_ sky130_fd_sc_hd__a221o_1
X_0592_ _0223_ _0224_ _0226_ VGND VGND VPWR VPWR _0227_ sky130_fd_sc_hd__o21a_1
XFILLER_27_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0928_ clknet_4_7_0_clk sample_rate.n_count\[3\] net50 VGND VGND VPWR VPWR sample_rate.count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_0859_ _0073_ waveshape.seq_div.dividend\[44\] _0193_ VGND VGND VPWR VPWR _0394_
+ sky130_fd_sc_hd__or3_1
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold58 pwm_counter.count\[1\] VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__dlygate4sd3_1
Xhold14 _0028_ VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 waveshape.seq_div.dividend\[46\] VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 count\[10\] VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 waveshape.seq_div.dividend\[20\] VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 waveshape.seq_div.dividend\[19\] VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0644_ sample_rate.count\[0\] _0263_ VGND VGND VPWR VPWR sample_rate.n_count\[0\]
+ sky130_fd_sc_hd__and2b_1
X_0713_ net44 waveshape.scaled_count\[3\] net22 VGND VGND VPWR VPWR _0303_ sky130_fd_sc_hd__and3_1
X_0575_ _0208_ _0209_ VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__or2_1
XFILLER_33_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0558_ waveshape.seq_div.n\[1\] waveshape.seq_div.n\[0\] waveshape.seq_div.state\[1\]
+ VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__and3_1
X_0627_ count\[9\] _0251_ VGND VGND VPWR VPWR _0253_ sky130_fd_sc_hd__and2_1
X_0489_ _0127_ VGND VGND VPWR VPWR _0128_ sky130_fd_sc_hd__inv_2
XFILLER_26_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_28_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0961_ clknet_4_14_0_clk waveshape.shaper.n_sample\[5\] net59 VGND VGND VPWR VPWR
+ pwm_counter.sample\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_17_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0892_ _0210_ _0422_ keypad.n_modekey VGND VGND VPWR VPWR _0423_ sky130_fd_sc_hd__a21o_1
XFILLER_4_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_235 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout50 net51 VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__buf_2
XFILLER_13_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout61 net62 VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__clkbuf_2
XFILLER_49_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0944_ clknet_4_11_0_clk _0015_ net53 VGND VGND VPWR VPWR waveshape.seq_div.dividend\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_0875_ keypad.keypad_reg\[4\] _0084_ _0406_ keypad.n_modekey VGND VGND VPWR VPWR
+ _0407_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_30_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload3 clknet_4_3_0_clk VGND VGND VPWR VPWR clkload3/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_21_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0660_ net123 pwm_counter.count\[0\] VGND VGND VPWR VPWR pwm_counter.n_count\[1\]
+ sky130_fd_sc_hd__xor2_1
XFILLER_10_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0591_ count\[7\] _0150_ _0181_ count\[8\] _0225_ VGND VGND VPWR VPWR _0226_ sky130_fd_sc_hd__o221a_1
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0927_ clknet_4_5_0_clk sample_rate.n_count\[2\] net50 VGND VGND VPWR VPWR sample_rate.count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_0858_ waveshape.seq_div.dividend\[44\] net26 _0362_ _0393_ VGND VGND VPWR VPWR _0061_
+ sky130_fd_sc_hd__a22o_1
X_0789_ waveshape.seq_div.dividend\[28\] _0122_ _0144_ VGND VGND VPWR VPWR _0340_
+ sky130_fd_sc_hd__a21bo_1
Xhold59 pwm_counter.count\[7\] VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 waveshape.seq_div.state\[2\] VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 waveshape.seq_div.dividend\[14\] VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 count\[1\] VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 waveshape.seq_div.dividend\[18\] VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0643_ _0092_ _0101_ VGND VGND VPWR VPWR _0263_ sky130_fd_sc_hd__nor2_1
X_0574_ _0208_ _0209_ VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__nor2_1
X_0712_ net139 net19 _0302_ VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__a21o_1
XFILLER_15_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput16 net16 VGND VGND VPWR VPWR pwm sky130_fd_sc_hd__buf_2
XFILLER_16_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0557_ net80 _0195_ net38 VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__a21o_1
X_0626_ _0251_ _0252_ net17 VGND VGND VPWR VPWR oscill.n_count\[8\] sky130_fd_sc_hd__and3b_1
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0488_ waveshape.seq_div.dividend\[27\] _0125_ VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_19_Left_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0609_ count\[0\] count\[1\] count\[2\] VGND VGND VPWR VPWR _0242_ sky130_fd_sc_hd__and3_1
XFILLER_43_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0960_ clknet_4_15_0_clk waveshape.shaper.n_sample\[4\] net59 VGND VGND VPWR VPWR
+ pwm_counter.sample\[4\] sky130_fd_sc_hd__dfrtp_1
X_0891_ keypad.keypad_reg\[9\] _0212_ _0403_ _0410_ VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__a31o_1
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_247 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout62 net15 VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__buf_2
Xfanout40 net43 VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__buf_2
Xfanout51 net62 VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_2
XFILLER_13_83 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0874_ keypad.keypad_reg\[6\] _0405_ VGND VGND VPWR VPWR _0406_ sky130_fd_sc_hd__and2b_1
Xclkload10 clknet_4_10_0_clk VGND VGND VPWR VPWR clkload10/X sky130_fd_sc_hd__clkbuf_8
X_0943_ clknet_4_11_0_clk _0014_ net53 VGND VGND VPWR VPWR waveshape.seq_div.dividend\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload4 clknet_4_4_0_clk VGND VGND VPWR VPWR clkload4/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_21_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0590_ count\[9\] _0176_ VGND VGND VPWR VPWR _0225_ sky130_fd_sc_hd__or2_1
XFILLER_1_64 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0926_ clknet_4_5_0_clk net87 net48 VGND VGND VPWR VPWR sample_rate.count\[1\] sky130_fd_sc_hd__dfrtp_1
X_0857_ net41 waveshape.seq_div.dividend\[43\] _0392_ net39 VGND VGND VPWR VPWR _0393_
+ sky130_fd_sc_hd__a22o_1
XFILLER_20_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold16 waveshape.seq_div.n\[4\] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__dlygate4sd3_1
X_0788_ waveshape.seq_div.dividend\[28\] _0339_ net24 VGND VGND VPWR VPWR _0045_ sky130_fd_sc_hd__mux2_1
Xhold38 waveshape.seq_div.dividend\[15\] VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 waveshape.seq_div.dividend\[16\] VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold49 waveshape.seq_div.n\[2\] VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_7_Left_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0711_ net45 waveshape.scaled_count\[2\] net22 VGND VGND VPWR VPWR _0302_ sky130_fd_sc_hd__and3_1
XFILLER_32_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0573_ keypad.keypad_reg\[4\] keypad.keypad_reg\[5\] keypad.keypad_reg\[6\] keypad.keypad_reg\[7\]
+ VGND VGND VPWR VPWR _0209_ sky130_fd_sc_hd__or4_1
X_0642_ _0237_ _0238_ _0262_ VGND VGND VPWR VPWR oscill.n_count\[14\] sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_49_Left_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0909_ clknet_4_12_0_clk oscill.n_count\[0\] net57 VGND VGND VPWR VPWR count\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_48_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0625_ count\[6\] count\[7\] _0246_ count\[8\] VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__a31o_1
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0556_ waveshape.seq_div.dividend\[47\] _0194_ VGND VGND VPWR VPWR _0195_ sky130_fd_sc_hd__nor2_1
X_0487_ waveshape.seq_div.dividend\[27\] _0125_ VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__nand2_1
XFILLER_38_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0608_ count\[0\] count\[1\] count\[2\] VGND VGND VPWR VPWR _0241_ sky130_fd_sc_hd__a21o_1
XFILLER_37_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0539_ waveshape.seq_div.dividend\[33\] _0176_ VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_36_Left_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0890_ _0416_ _0420_ _0415_ VGND VGND VPWR VPWR _0421_ sky130_fd_sc_hd__a21boi_1
XTAP_TAPCELL_ROW_2_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout30 freq_div.keycode\[3\] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_2
Xfanout52 net54 VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__clkbuf_4
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout41 net42 VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__buf_2
XFILLER_13_95 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload11 clknet_4_12_0_clk VGND VGND VPWR VPWR clkload11/Y sky130_fd_sc_hd__bufinv_16
X_0873_ keypad.keypad_reg\[7\] _0404_ VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__nor2_1
XFILLER_13_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0942_ clknet_4_9_0_clk _0013_ net53 VGND VGND VPWR VPWR waveshape.seq_div.dividend\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload5 clknet_4_5_0_clk VGND VGND VPWR VPWR clkload5/Y sky130_fd_sc_hd__clkinv_2
XTAP_TAPCELL_ROW_21_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_23_Left_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0925_ clknet_4_5_0_clk sample_rate.n_count\[0\] net48 VGND VGND VPWR VPWR sample_rate.count\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_0856_ waveshape.seq_div.dividend\[44\] _0193_ VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__xnor2_1
X_0787_ net37 _0144_ _0338_ net43 waveshape.seq_div.dividend\[27\] VGND VGND VPWR
+ VPWR _0339_ sky130_fd_sc_hd__a32o_1
Xhold17 _0040_ VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 waveshape.seq_div.dividend\[10\] VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 waveshape.seq_div.dividend\[21\] VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0641_ count\[14\] _0260_ VGND VGND VPWR VPWR _0262_ sky130_fd_sc_hd__xnor2_1
X_0710_ net131 net20 _0301_ VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__a21o_1
X_0572_ _0205_ _0207_ VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__or2_1
XFILLER_25_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0839_ waveshape.seq_div.dividend\[40\] _0191_ VGND VGND VPWR VPWR _0379_ sky130_fd_sc_hd__xnor2_1
X_0908_ clknet_4_14_0_clk state_machine.nextState\[2\] net58 VGND VGND VPWR VPWR mode\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_21_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0624_ count\[7\] count\[8\] _0248_ VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__and3_1
XFILLER_38_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0555_ waveshape.seq_div.dividend\[46\] waveshape.seq_div.dividend\[45\] waveshape.seq_div.dividend\[44\]
+ _0193_ VGND VGND VPWR VPWR _0194_ sky130_fd_sc_hd__or4_2
X_0486_ net31 net34 _0094_ _0124_ VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__a31o_1
XFILLER_38_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_8_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_10_Left_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0538_ waveshape.seq_div.dividend\[33\] _0176_ VGND VGND VPWR VPWR _0177_ sky130_fd_sc_hd__nor2_1
X_0607_ net105 net113 _0240_ VGND VGND VPWR VPWR oscill.n_count\[1\] sky130_fd_sc_hd__a21oi_1
XFILLER_37_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0469_ net30 net34 VGND VGND VPWR VPWR _0108_ sky130_fd_sc_hd__or2_2
XFILLER_26_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_36_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_216 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout31 freq_div.keycode\[3\] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__buf_1
Xfanout53 net54 VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_4
Xfanout20 net21 VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout42 net43 VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_2
XFILLER_49_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0941_ clknet_4_12_0_clk _0012_ net58 VGND VGND VPWR VPWR waveshape.seq_div.dividend\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload12 clknet_4_13_0_clk VGND VGND VPWR VPWR clkload12/X sky130_fd_sc_hd__clkbuf_4
X_0872_ _0208_ _0213_ _0402_ VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_30_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload6 clknet_4_6_0_clk VGND VGND VPWR VPWR clkload6/Y sky130_fd_sc_hd__clkinv_2
XFILLER_34_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0924_ clknet_4_1_0_clk net65 net47 VGND VGND VPWR VPWR count\[15\] sky130_fd_sc_hd__dfrtp_1
X_0855_ waveshape.seq_div.dividend\[43\] net26 _0362_ _0391_ VGND VGND VPWR VPWR _0060_
+ sky130_fd_sc_hd__a22o_1
X_0786_ _0127_ _0143_ _0123_ _0126_ VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__o211ai_1
Xhold18 pwm_counter.sample\[1\] VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 waveshape.seq_div.dividend\[22\] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_40_Left_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0571_ keypad.keypad_reg\[2\] keypad.keypad_reg\[3\] VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__or2_1
X_0640_ net17 _0260_ _0261_ VGND VGND VPWR VPWR oscill.n_count\[13\] sky130_fd_sc_hd__and3_1
XFILLER_18_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0907_ clknet_4_14_0_clk state_machine.nextState\[1\] net58 VGND VGND VPWR VPWR state_machine.fsmState\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_0769_ waveshape.seq_div.n\[3\] _0323_ net81 VGND VGND VPWR VPWR _0326_ sky130_fd_sc_hd__a21oi_1
X_0838_ waveshape.seq_div.dividend\[39\] net26 _0362_ _0378_ VGND VGND VPWR VPWR _0056_
+ sky130_fd_sc_hd__a22o_1
XFILLER_24_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0623_ net110 _0248_ _0250_ VGND VGND VPWR VPWR oscill.n_count\[7\] sky130_fd_sc_hd__a21oi_1
X_0554_ _0117_ _0190_ _0192_ _0113_ VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__a211o_1
XFILLER_38_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0485_ net32 _0119_ _0120_ net31 VGND VGND VPWR VPWR _0124_ sky130_fd_sc_hd__a31oi_1
XFILLER_42_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0537_ _0174_ _0175_ VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__and2_1
X_0606_ count\[0\] count\[1\] net17 VGND VGND VPWR VPWR _0240_ sky130_fd_sc_hd__o21ai_1
X_0468_ freq_div.keycode\[0\] net35 net33 VGND VGND VPWR VPWR _0107_ sky130_fd_sc_hd__o21a_1
XFILLER_26_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_36_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout21 _0299_ VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__buf_2
Xfanout43 waveshape.seq_div.state\[3\] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_2
Xfanout32 net33 VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__clkbuf_2
Xfanout54 net55 VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__buf_2
XFILLER_22_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0940_ clknet_4_12_0_clk _0011_ net57 VGND VGND VPWR VPWR waveshape.seq_div.dividend\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload13 clknet_4_14_0_clk VGND VGND VPWR VPWR clkload13/Y sky130_fd_sc_hd__clkinv_2
X_0871_ keypad.keypad_reg\[10\] _0402_ VGND VGND VPWR VPWR _0403_ sky130_fd_sc_hd__nor2_1
XFILLER_9_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_30_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload7 clknet_4_7_0_clk VGND VGND VPWR VPWR clkload7/X sky130_fd_sc_hd__clkbuf_4
XFILLER_46_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0923_ clknet_4_3_0_clk oscill.n_count\[14\] net46 VGND VGND VPWR VPWR count\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_0854_ net39 _0389_ _0390_ net41 waveshape.seq_div.dividend\[42\] VGND VGND VPWR
+ VPWR _0391_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_49_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0785_ net137 _0337_ net24 VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__mux2_1
Xhold19 _0029_ VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_27_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0570_ keypad.keypad_reg\[2\] _0205_ VGND VGND VPWR VPWR _0206_ sky130_fd_sc_hd__nor2_1
XFILLER_2_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0906_ clknet_4_14_0_clk state_machine.nextState\[0\] net58 VGND VGND VPWR VPWR state_machine.fsmState\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_0837_ _0376_ _0377_ net41 waveshape.seq_div.dividend\[38\] VGND VGND VPWR VPWR _0378_
+ sky130_fd_sc_hd__a2bb2o_1
X_0768_ net88 _0323_ _0325_ VGND VGND VPWR VPWR _0039_ sky130_fd_sc_hd__a21oi_1
X_0699_ _0291_ _0292_ _0293_ VGND VGND VPWR VPWR _0294_ sky130_fd_sc_hd__or3_1
XFILLER_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0484_ waveshape.seq_div.dividend\[28\] _0122_ VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__xnor2_1
X_0622_ count\[7\] _0248_ _0239_ VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__o21ai_1
X_0553_ waveshape.seq_div.dividend\[42\] waveshape.seq_div.dividend\[43\] waveshape.seq_div.dividend\[41\]
+ waveshape.seq_div.dividend\[40\] VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__or4_1
XFILLER_30_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0536_ net30 _0093_ _0107_ _0118_ VGND VGND VPWR VPWR _0175_ sky130_fd_sc_hd__or4_1
X_0605_ net105 net17 VGND VGND VPWR VPWR oscill.n_count\[0\] sky130_fd_sc_hd__nand2_1
X_0467_ _0105_ VGND VGND VPWR VPWR _0106_ sky130_fd_sc_hd__inv_2
X_1019_ clknet_4_11_0_clk net8 net53 VGND VGND VPWR VPWR keypad.keypad_reg\[3\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_36_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_95 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0519_ waveshape.seq_div.dividend\[30\] _0156_ VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_1_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout44 net45 VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__buf_2
Xfanout55 net62 VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_4
Xfanout33 freq_div.keycode\[2\] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_2
Xfanout22 net23 VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__buf_2
XFILLER_22_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0870_ keypad.keypad_reg\[12\] keypad.keypad_reg\[13\] VGND VGND VPWR VPWR _0402_
+ sky130_fd_sc_hd__or2_1
XFILLER_9_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload14 clknet_4_15_0_clk VGND VGND VPWR VPWR clkload14/X sky130_fd_sc_hd__clkbuf_4
X_0999_ clknet_4_5_0_clk _0062_ net51 VGND VGND VPWR VPWR waveshape.seq_div.dividend\[45\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload8 clknet_4_8_0_clk VGND VGND VPWR VPWR clkload8/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_24_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0922_ clknet_4_3_0_clk oscill.n_count\[13\] net49 VGND VGND VPWR VPWR count\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_0853_ waveshape.seq_div.dividend\[43\] net18 VGND VGND VPWR VPWR _0390_ sky130_fd_sc_hd__or2_1
X_0784_ net37 _0335_ _0336_ net43 waveshape.seq_div.dividend\[26\] VGND VGND VPWR
+ VPWR _0337_ sky130_fd_sc_hd__a32o_1
Xinput1 keypad_i[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
XFILLER_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_27_Left_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0767_ waveshape.seq_div.n\[3\] _0323_ _0197_ VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__o21ai_1
X_0905_ clknet_4_7_0_clk _0000_ net49 VGND VGND VPWR VPWR waveshape.seq_div.state\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_0836_ waveshape.seq_div.dividend\[39\] _0106_ _0374_ _0072_ VGND VGND VPWR VPWR
+ _0377_ sky130_fd_sc_hd__a31o_1
XFILLER_0_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0698_ net8 net7 net10 net9 VGND VGND VPWR VPWR _0293_ sky130_fd_sc_hd__or4_1
XFILLER_21_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0621_ _0248_ _0249_ VGND VGND VPWR VPWR oscill.n_count\[6\] sky130_fd_sc_hd__nor2_1
X_0483_ _0069_ _0119_ _0120_ _0121_ VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__a31o_2
XFILLER_23_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0552_ _0117_ _0190_ _0113_ VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__a21o_1
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0819_ _0168_ _0363_ VGND VGND VPWR VPWR _0364_ sky130_fd_sc_hd__xnor2_1
XFILLER_29_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0604_ _0237_ _0238_ VGND VGND VPWR VPWR _0239_ sky130_fd_sc_hd__and2_1
X_0535_ net31 _0107_ _0119_ _0094_ VGND VGND VPWR VPWR _0174_ sky130_fd_sc_hd__a2bb2o_1
X_0466_ waveshape.seq_div.dividend\[38\] _0098_ VGND VGND VPWR VPWR _0105_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_36_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_14_Left_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1018_ clknet_4_11_0_clk net7 net53 VGND VGND VPWR VPWR keypad.keypad_reg\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_17_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0518_ waveshape.seq_div.dividend\[30\] _0156_ VGND VGND VPWR VPWR _0157_ sky130_fd_sc_hd__and2_1
X_0449_ waveshape.seq_div.n\[1\] waveshape.seq_div.n\[0\] _0088_ VGND VGND VPWR VPWR
+ _0089_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_1_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout56 net61 VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__clkbuf_4
Xfanout45 waveshape.seq_div.state\[3\] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__buf_2
Xfanout34 net35 VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__buf_2
XFILLER_22_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout23 _0298_ VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__buf_2
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0998_ clknet_4_5_0_clk _0061_ net48 VGND VGND VPWR VPWR waveshape.seq_div.dividend\[44\]
+ sky130_fd_sc_hd__dfrtp_2
Xclkload9 clknet_4_9_0_clk VGND VGND VPWR VPWR clkload9/X sky130_fd_sc_hd__clkbuf_8
X_0924__65 VGND VGND VPWR VPWR _0924__65/HI net65 sky130_fd_sc_hd__conb_1
XFILLER_10_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0921_ clknet_4_3_0_clk oscill.n_count\[12\] net49 VGND VGND VPWR VPWR count\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_0783_ _0143_ _0334_ VGND VGND VPWR VPWR _0336_ sky130_fd_sc_hd__or2_1
X_0852_ waveshape.seq_div.dividend\[43\] net18 VGND VGND VPWR VPWR _0389_ sky130_fd_sc_hd__nand2_1
XFILLER_5_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput2 keypad_i[10] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_2_Left_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0904_ clknet_4_6_0_clk _0003_ net56 VGND VGND VPWR VPWR waveshape.seq_div.state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_0766_ _0323_ _0324_ VGND VGND VPWR VPWR _0038_ sky130_fd_sc_hd__nor2_1
X_0697_ net12 net11 net14 net13 VGND VGND VPWR VPWR _0292_ sky130_fd_sc_hd__or4_1
X_0835_ _0106_ _0374_ waveshape.seq_div.dividend\[39\] VGND VGND VPWR VPWR _0376_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_24_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_44_Left_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0551_ _0163_ _0185_ _0189_ VGND VGND VPWR VPWR _0190_ sky130_fd_sc_hd__o21ai_2
X_0620_ count\[6\] _0246_ _0239_ VGND VGND VPWR VPWR _0249_ sky130_fd_sc_hd__o21ai_1
X_0482_ net32 net31 _0120_ VGND VGND VPWR VPWR _0121_ sky130_fd_sc_hd__mux2_1
XFILLER_16_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0818_ _0172_ _0359_ _0170_ VGND VGND VPWR VPWR _0363_ sky130_fd_sc_hd__a21oi_1
X_0749_ net94 net23 _0320_ VGND VGND VPWR VPWR _0025_ sky130_fd_sc_hd__o21a_1
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0534_ _0168_ _0172_ VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__nand2_1
X_0603_ count\[14\] _0098_ _0233_ _0234_ count\[15\] VGND VGND VPWR VPWR _0238_ sky130_fd_sc_hd__a221oi_1
X_0465_ net106 _0089_ _0104_ VGND VGND VPWR VPWR _0003_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_36_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1017_ clknet_4_11_0_clk net6 net53 VGND VGND VPWR VPWR keypad.keypad_reg\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_27_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_31_Left_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0517_ _0155_ _0107_ net30 VGND VGND VPWR VPWR _0156_ sky130_fd_sc_hd__mux2_2
X_0448_ waveshape.seq_div.n\[3\] waveshape.seq_div.n\[4\] waveshape.seq_div.n\[2\]
+ VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_1_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout35 freq_div.keycode\[1\] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_2
Xfanout24 _0297_ VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_4
Xfanout46 net47 VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_4
XFILLER_22_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout57 net61 VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_4
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0997_ clknet_4_4_0_clk _0060_ net48 VGND VGND VPWR VPWR waveshape.seq_div.dividend\[43\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_46_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0920_ clknet_4_3_0_clk oscill.n_count\[11\] net46 VGND VGND VPWR VPWR count\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_0782_ _0143_ _0334_ VGND VGND VPWR VPWR _0335_ sky130_fd_sc_hd__nand2_1
X_0851_ net144 net25 _0387_ _0388_ VGND VGND VPWR VPWR _0059_ sky130_fd_sc_hd__o22a_1
XFILLER_46_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput3 keypad_i[11] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0903_ clknet_4_4_0_clk net42 net49 VGND VGND VPWR VPWR waveshape.seq_div.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_0834_ net118 net27 _0362_ _0375_ VGND VGND VPWR VPWR _0055_ sky130_fd_sc_hd__a22o_1
X_0765_ net114 _0196_ VGND VGND VPWR VPWR _0324_ sky130_fd_sc_hd__nor2_1
X_0696_ net3 net2 net5 net4 VGND VGND VPWR VPWR _0291_ sky130_fd_sc_hd__or4_1
XFILLER_24_167 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0550_ _0173_ _0177_ _0187_ _0188_ _0166_ VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__o311a_1
X_0481_ net36 net35 VGND VGND VPWR VPWR _0120_ sky130_fd_sc_hd__nand2b_2
XFILLER_21_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0817_ _0071_ _0103_ net28 VGND VGND VPWR VPWR _0362_ sky130_fd_sc_hd__o21ba_2
XFILLER_21_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0748_ net40 waveshape.seq_div.dividend\[21\] net28 count\[14\] net21 VGND VGND VPWR
+ VPWR _0320_ sky130_fd_sc_hd__a221o_1
X_0679_ state_machine.fsmState\[1\] _0087_ waveshape.scaled_count\[7\] VGND VGND VPWR
+ VPWR _0282_ sky130_fd_sc_hd__and3_2
XFILLER_29_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0464_ waveshape.seq_div.state\[0\] _0103_ VGND VGND VPWR VPWR _0104_ sky130_fd_sc_hd__and2_1
X_0533_ _0170_ _0171_ VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__nor2_1
X_0602_ _0231_ _0232_ _0236_ VGND VGND VPWR VPWR _0237_ sky130_fd_sc_hd__o21ai_1
X_1016_ clknet_4_11_0_clk net1 net53 VGND VGND VPWR VPWR keypad.keypad_reg\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_27_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0516_ _0099_ _0154_ _0093_ VGND VGND VPWR VPWR _0155_ sky130_fd_sc_hd__a21o_1
X_0447_ mode\[1\] VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_1_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout36 freq_div.keycode\[0\] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__buf_2
Xfanout47 net62 VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_4
XFILLER_22_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_24_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout58 net60 VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__clkbuf_4
Xfanout25 _0297_ VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__buf_2
XFILLER_1_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0996_ clknet_4_4_0_clk _0059_ net48 VGND VGND VPWR VPWR waveshape.seq_div.dividend\[42\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_6_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0850_ net41 waveshape.seq_div.dividend\[41\] net26 VGND VGND VPWR VPWR _0388_ sky130_fd_sc_hd__a21o_1
X_0781_ _0126_ _0128_ VGND VGND VPWR VPWR _0334_ sky130_fd_sc_hd__nand2_1
XFILLER_39_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput4 keypad_i[12] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
X_0979_ clknet_4_0_0_clk _0042_ net46 VGND VGND VPWR VPWR waveshape.seq_div.dividend\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_35_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0902_ clknet_4_7_0_clk _0002_ net49 VGND VGND VPWR VPWR waveshape.seq_div.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_0833_ net38 _0373_ _0374_ net41 waveshape.seq_div.dividend\[37\] VGND VGND VPWR
+ VPWR _0375_ sky130_fd_sc_hd__a32o_1
X_0764_ waveshape.seq_div.n\[2\] _0196_ VGND VGND VPWR VPWR _0323_ sky130_fd_sc_hd__and2_1
X_0695_ state_machine.fsmState\[1\] mode\[1\] _0289_ _0290_ VGND VGND VPWR VPWR waveshape.shaper.n_sample\[7\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_24_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0480_ net34 net36 VGND VGND VPWR VPWR _0119_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_16_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0816_ net126 _0361_ net25 VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__mux2_1
X_0747_ net104 net23 _0319_ VGND VGND VPWR VPWR _0024_ sky130_fd_sc_hd__o21a_1
X_0678_ state_machine.fsmState\[1\] mode\[1\] _0280_ VGND VGND VPWR VPWR state_machine.nextState\[2\]
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_7_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0601_ count\[11\] _0165_ _0234_ _0235_ VGND VGND VPWR VPWR _0236_ sky130_fd_sc_hd__o211a_1
X_0532_ waveshape.seq_div.dividend\[34\] _0169_ VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__nor2_1
XFILLER_21_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0463_ _0101_ _0102_ VGND VGND VPWR VPWR _0103_ sky130_fd_sc_hd__nor2_1
X_1015_ clknet_4_11_0_clk keypad.n_modekey net53 VGND VGND VPWR VPWR keypad.modekey
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_34_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_18_Left_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0515_ net32 net34 net36 VGND VGND VPWR VPWR _0154_ sky130_fd_sc_hd__o21a_1
X_0446_ state_machine.fsmState\[1\] VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__inv_2
Xfanout37 net39 VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_24_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout26 net27 VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_4
Xfanout59 net60 VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__clkbuf_4
Xfanout48 net51 VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_4
XFILLER_1_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0995_ clknet_4_4_0_clk _0058_ net48 VGND VGND VPWR VPWR waveshape.seq_div.dividend\[41\]
+ sky130_fd_sc_hd__dfrtp_1
X_0429_ net33 VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__inv_2
XFILLER_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0780_ waveshape.seq_div.dividend\[26\] _0333_ net24 VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__mux2_1
Xinput5 keypad_i[13] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0978_ clknet_4_0_0_clk _0041_ net46 VGND VGND VPWR VPWR waveshape.seq_div.dividend\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_19_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0763_ _0196_ net116 VGND VGND VPWR VPWR _0037_ sky130_fd_sc_hd__nor2_1
X_0832_ waveshape.seq_div.dividend\[37\] _0100_ _0110_ _0366_ _0114_ VGND VGND VPWR
+ VPWR _0374_ sky130_fd_sc_hd__o221ai_4
X_0901_ clknet_4_6_0_clk _0001_ net49 VGND VGND VPWR VPWR waveshape.seq_div.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_0694_ _0086_ waveshape.scaled_count\[6\] waveshape.scaled_count\[7\] VGND VGND VPWR
+ VPWR _0290_ sky130_fd_sc_hd__a21o_1
XFILLER_24_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_6_Left_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_9_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_9_0_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_16_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0815_ net40 waveshape.seq_div.dividend\[33\] _0360_ net39 VGND VGND VPWR VPWR _0361_
+ sky130_fd_sc_hd__a22o_1
X_0746_ net42 waveshape.seq_div.dividend\[20\] net28 count\[13\] net21 VGND VGND VPWR
+ VPWR _0319_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_48_Left_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0677_ state_machine.fsmState\[1\] _0087_ _0277_ VGND VGND VPWR VPWR state_machine.nextState\[1\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0531_ waveshape.seq_div.dividend\[34\] _0169_ VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__and2_1
X_0600_ count\[12\] _0109_ _0233_ VGND VGND VPWR VPWR _0235_ sky130_fd_sc_hd__o21ba_1
XFILLER_14_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0462_ _0098_ _0100_ _0092_ VGND VGND VPWR VPWR _0102_ sky130_fd_sc_hd__a21bo_1
XFILLER_34_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1014_ clknet_4_10_0_clk _0068_ net52 VGND VGND VPWR VPWR freq_div.keycode\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_26_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0729_ net95 net22 _0310_ VGND VGND VPWR VPWR _0015_ sky130_fd_sc_hd__o21a_1
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0514_ _0151_ _0152_ VGND VGND VPWR VPWR _0153_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_49_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0445_ keypad.keypad_reg\[13\] VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__inv_2
Xfanout38 net39 VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__buf_2
XFILLER_13_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout49 net51 VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_24_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout27 _0296_ VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__buf_2
XFILLER_49_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_35_Left_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0994_ clknet_4_1_0_clk _0057_ net48 VGND VGND VPWR VPWR waveshape.seq_div.dividend\[40\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_10_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput6 keypad_i[1] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_1
X_0977_ clknet_4_7_0_clk net82 net56 VGND VGND VPWR VPWR waveshape.seq_div.n\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0900_ _0423_ _0425_ _0428_ _0214_ net117 VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__o32a_1
XFILLER_18_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0762_ waveshape.seq_div.n\[0\] waveshape.seq_div.state\[1\] net115 VGND VGND VPWR
+ VPWR _0322_ sky130_fd_sc_hd__a21oi_1
X_0831_ _0116_ _0366_ _0112_ _0114_ VGND VGND VPWR VPWR _0373_ sky130_fd_sc_hd__a211o_1
X_0693_ _0086_ waveshape.scaled_count\[7\] waveshape.scaled_count\[6\] VGND VGND VPWR
+ VPWR _0289_ sky130_fd_sc_hd__nand3_1
XFILLER_44_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_22_Left_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0814_ _0172_ _0359_ VGND VGND VPWR VPWR _0360_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_16_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0745_ net90 net23 _0318_ VGND VGND VPWR VPWR _0023_ sky130_fd_sc_hd__o21a_1
X_0676_ _0278_ _0281_ _0280_ VGND VGND VPWR VPWR state_machine.nextState\[0\] sky130_fd_sc_hd__o21a_1
XFILLER_12_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_188 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0530_ net30 _0155_ _0095_ _0154_ VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_11_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0461_ sample_rate.count\[7\] sample_rate.count\[6\] VGND VGND VPWR VPWR _0101_ sky130_fd_sc_hd__or2_2
X_1013_ clknet_4_8_0_clk _0067_ net52 VGND VGND VPWR VPWR freq_div.keycode\[2\] sky130_fd_sc_hd__dfrtp_1
X_0659_ net124 pwm_counter.count\[6\] _0271_ _0081_ VGND VGND VPWR VPWR pwm_counter.n_count\[0\]
+ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0728_ net45 waveshape.seq_div.dividend\[11\] net29 count\[4\] net19 VGND VGND VPWR
+ VPWR _0310_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_4_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_8_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_8_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0513_ waveshape.seq_div.dividend\[31\] _0150_ VGND VGND VPWR VPWR _0152_ sky130_fd_sc_hd__or2_1
X_0444_ keypad.keypad_reg\[5\] VGND VGND VPWR VPWR _0084_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_49_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout39 waveshape.seq_div.state\[4\] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__buf_2
XFILLER_13_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout17 _0239_ VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__buf_2
Xfanout28 _0295_ VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__buf_2
XFILLER_48_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0993_ clknet_4_4_0_clk _0056_ net48 VGND VGND VPWR VPWR waveshape.seq_div.dividend\[39\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_216 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput7 keypad_i[2] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_1
X_0976_ clknet_4_7_0_clk net89 net50 VGND VGND VPWR VPWR waveshape.seq_div.n\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_19_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0830_ waveshape.seq_div.dividend\[37\] net26 _0362_ _0372_ VGND VGND VPWR VPWR _0054_
+ sky130_fd_sc_hd__a22o_1
XFILLER_25_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0761_ waveshape.seq_div.n\[0\] net106 VGND VGND VPWR VPWR _0036_ sky130_fd_sc_hd__xor2_1
X_0692_ waveshape.scaled_count\[6\] _0278_ _0279_ _0288_ _0282_ VGND VGND VPWR VPWR
+ waveshape.shaper.n_sample\[6\] sky130_fd_sc_hd__a221o_1
XFILLER_49_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0959_ clknet_4_13_0_clk waveshape.shaper.n_sample\[3\] net56 VGND VGND VPWR VPWR
+ pwm_counter.sample\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_138 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0813_ _0186_ _0353_ _0177_ VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__o21ba_1
XFILLER_14_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput10 keypad_i[5] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_1
X_0744_ net44 waveshape.seq_div.dividend\[19\] net28 count\[12\] net21 VGND VGND VPWR
+ VPWR _0318_ sky130_fd_sc_hd__a221o_1
X_0675_ state_machine.fsmState\[1\] mode\[1\] keypad.modekey VGND VGND VPWR VPWR _0281_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_29_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0460_ net33 net35 net31 VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__a21bo_4
X_1012_ clknet_4_8_0_clk _0066_ net52 VGND VGND VPWR VPWR freq_div.keycode\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0727_ net97 net22 _0309_ VGND VGND VPWR VPWR _0014_ sky130_fd_sc_hd__o21a_1
X_0658_ pwm_counter.count\[6\] _0271_ VGND VGND VPWR VPWR _0272_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_4_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0589_ count\[7\] _0150_ _0156_ count\[6\] VGND VGND VPWR VPWR _0224_ sky130_fd_sc_hd__a22o_1
XFILLER_27_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0512_ waveshape.seq_div.dividend\[31\] _0150_ VGND VGND VPWR VPWR _0151_ sky130_fd_sc_hd__nand2_1
X_0443_ keypad.keypad_reg\[4\] VGND VGND VPWR VPWR _0083_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_49_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout29 _0295_ VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__buf_2
XFILLER_13_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0992_ clknet_4_4_0_clk _0055_ net49 VGND VGND VPWR VPWR waveshape.seq_div.dividend\[38\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_7_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_7_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_5_95 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput8 keypad_i[3] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_1
X_0975_ clknet_4_7_0_clk _0038_ net56 VGND VGND VPWR VPWR waveshape.seq_div.n\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_40_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0760_ net68 pwm_counter.active_sample\[7\] _0197_ VGND VGND VPWR VPWR _0035_ sky130_fd_sc_hd__mux2_1
X_0691_ waveshape.scaled_count\[7\] waveshape.scaled_count\[5\] VGND VGND VPWR VPWR
+ _0288_ sky130_fd_sc_hd__xor2_1
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0958_ clknet_4_13_0_clk waveshape.shaper.n_sample\[2\] net56 VGND VGND VPWR VPWR
+ pwm_counter.sample\[2\] sky130_fd_sc_hd__dfrtp_1
X_0889_ _0207_ keypad.keypad_reg\[0\] keypad.keypad_reg\[1\] VGND VGND VPWR VPWR _0420_
+ sky130_fd_sc_hd__or3b_1
XFILLER_15_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput11 keypad_i[6] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_1
X_0812_ net138 _0358_ net24 VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__mux2_1
X_0743_ net101 net23 _0317_ VGND VGND VPWR VPWR _0022_ sky130_fd_sc_hd__o21a_1
X_0674_ state_machine.fsmState\[0\] keypad.modekey VGND VGND VPWR VPWR _0280_ sky130_fd_sc_hd__or2_1
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1011_ clknet_4_10_0_clk _0065_ net52 VGND VGND VPWR VPWR freq_div.keycode\[0\] sky130_fd_sc_hd__dfrtp_1
X_0726_ net45 waveshape.seq_div.dividend\[10\] net29 count\[3\] net19 VGND VGND VPWR
+ VPWR _0309_ sky130_fd_sc_hd__a221o_1
X_0657_ pwm_counter.count\[5\] pwm_counter.count\[4\] _0270_ VGND VGND VPWR VPWR _0271_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_4_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0588_ count\[5\] _0145_ _0156_ count\[6\] _0222_ VGND VGND VPWR VPWR _0223_ sky130_fd_sc_hd__o221a_1
XFILLER_27_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0511_ _0096_ _0118_ _0108_ VGND VGND VPWR VPWR _0150_ sky130_fd_sc_hd__o21ai_2
XFILLER_12_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0442_ keypad.keypad_reg\[0\] VGND VGND VPWR VPWR _0082_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_49_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout19 _0299_ VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_32_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0709_ net44 waveshape.scaled_count\[1\] _0298_ VGND VGND VPWR VPWR _0301_ sky130_fd_sc_hd__and3_1
XFILLER_38_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0991_ clknet_4_1_0_clk _0054_ net47 VGND VGND VPWR VPWR waveshape.seq_div.dividend\[37\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_8_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_39_Left_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput9 keypad_i[4] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_1
X_0974_ clknet_4_7_0_clk _0037_ net50 VGND VGND VPWR VPWR waveshape.seq_div.n\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_6_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_6_0_clk sky130_fd_sc_hd__clkbuf_8
X_0690_ net148 _0278_ _0279_ _0287_ _0282_ VGND VGND VPWR VPWR waveshape.shaper.n_sample\[5\]
+ sky130_fd_sc_hd__a221o_1
XFILLER_2_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0957_ clknet_4_13_0_clk waveshape.shaper.n_sample\[1\] net56 VGND VGND VPWR VPWR
+ pwm_counter.sample\[1\] sky130_fd_sc_hd__dfrtp_1
X_0888_ _0083_ keypad.keypad_reg\[5\] _0406_ _0412_ VGND VGND VPWR VPWR _0419_ sky130_fd_sc_hd__a31o_1
XFILLER_46_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_92 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_26_Left_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput12 keypad_i[7] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_1
X_0811_ net40 waveshape.seq_div.dividend\[32\] _0357_ net37 VGND VGND VPWR VPWR _0358_
+ sky130_fd_sc_hd__a22o_1
X_0742_ net44 waveshape.seq_div.dividend\[18\] net28 count\[11\] net21 VGND VGND VPWR
+ VPWR _0317_ sky130_fd_sc_hd__a221o_1
X_0673_ state_machine.fsmState\[1\] _0087_ VGND VGND VPWR VPWR _0279_ sky130_fd_sc_hd__nor2_2
XFILLER_42_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_136 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1010_ clknet_4_11_0_clk pwm_counter.n_pwm net60 VGND VGND VPWR VPWR pwm1 sky130_fd_sc_hd__dfrtp_1
XFILLER_8_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0656_ pwm_counter.count\[3\] _0269_ VGND VGND VPWR VPWR _0270_ sky130_fd_sc_hd__and2_1
X_0725_ net93 net22 _0308_ VGND VGND VPWR VPWR _0013_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_4_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0587_ count\[5\] _0145_ _0215_ _0221_ VGND VGND VPWR VPWR _0222_ sky130_fd_sc_hd__a22o_1
XFILLER_27_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0510_ _0147_ _0148_ VGND VGND VPWR VPWR _0149_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_49_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0441_ pwm_counter.count\[0\] VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__inv_2
Xhold1 pwm_counter.sample\[5\] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Left_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0639_ count\[13\] _0258_ VGND VGND VPWR VPWR _0261_ sky130_fd_sc_hd__or2_1
X_0708_ net136 net21 _0300_ VGND VGND VPWR VPWR _0004_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0990_ clknet_4_1_0_clk _0053_ net47 VGND VGND VPWR VPWR waveshape.seq_div.dividend\[36\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_39_135 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0973_ clknet_4_7_0_clk net107 net56 VGND VGND VPWR VPWR waveshape.seq_div.n\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_40_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0956_ clknet_4_13_0_clk waveshape.shaper.n_sample\[0\] net56 VGND VGND VPWR VPWR
+ pwm_counter.sample\[0\] sky130_fd_sc_hd__dfrtp_1
X_0887_ _0407_ _0411_ _0418_ _0214_ net108 VGND VGND VPWR VPWR _0065_ sky130_fd_sc_hd__o32a_1
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Left_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput13 keypad_i[8] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_1
X_0810_ _0179_ _0356_ VGND VGND VPWR VPWR _0357_ sky130_fd_sc_hd__xnor2_1
X_0741_ net91 net23 _0316_ VGND VGND VPWR VPWR _0021_ sky130_fd_sc_hd__o21a_1
X_0672_ _0086_ _0087_ VGND VGND VPWR VPWR _0278_ sky130_fd_sc_hd__nor2_2
XFILLER_37_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0939_ clknet_4_14_0_clk _0010_ net58 VGND VGND VPWR VPWR waveshape.scaled_count\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_43_Left_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_5_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_5_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_43_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0655_ pwm_counter.count\[2\] pwm_counter.count\[1\] pwm_counter.count\[0\] VGND
+ VGND VPWR VPWR _0269_ sky130_fd_sc_hd__and3_1
X_0586_ _0218_ _0219_ _0220_ VGND VGND VPWR VPWR _0221_ sky130_fd_sc_hd__a21o_1
X_0724_ net44 waveshape.seq_div.dividend\[9\] net29 count\[2\] net19 VGND VGND VPWR
+ VPWR _0308_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_4_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0440_ pwm_counter.count\[1\] VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_49_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2 _0033_ VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0707_ net44 waveshape.scaled_count\[0\] net23 VGND VGND VPWR VPWR _0300_ sky130_fd_sc_hd__and3_1
X_0569_ keypad.keypad_reg\[0\] keypad.keypad_reg\[1\] VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__or2_1
X_0638_ count\[13\] _0258_ VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_23_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_30_Left_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0932__63 VGND VGND VPWR VPWR _0932__63/HI net63 sky130_fd_sc_hd__conb_1
XFILLER_39_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_95 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0972_ clknet_4_15_0_clk net69 net58 VGND VGND VPWR VPWR pwm_counter.active_sample\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_33_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0886_ _0415_ _0417_ _0412_ _0414_ VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__a211o_1
X_0955_ clknet_4_0_0_clk _0026_ net62 VGND VGND VPWR VPWR waveshape.seq_div.dividend\[23\]
+ sky130_fd_sc_hd__dfrtp_1
Xmax_cap18 _0385_ VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_1
XFILLER_23_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput14 keypad_i[9] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_1
XFILLER_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0740_ net44 waveshape.seq_div.dividend\[17\] net28 count\[10\] net21 VGND VGND VPWR
+ VPWR _0316_ sky130_fd_sc_hd__a221o_1
X_0671_ keypad.modekey state_machine.fsmState\[0\] VGND VGND VPWR VPWR _0277_ sky130_fd_sc_hd__and2b_1
XFILLER_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0869_ waveshape.seq_div.dividend\[47\] net27 _0362_ _0401_ VGND VGND VPWR VPWR _0064_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_15_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0938_ clknet_4_14_0_clk _0009_ net58 VGND VGND VPWR VPWR waveshape.scaled_count\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_38_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0723_ net96 net22 _0307_ VGND VGND VPWR VPWR _0012_ sky130_fd_sc_hd__o21a_1
X_0654_ _0263_ _0268_ VGND VGND VPWR VPWR sample_rate.n_count\[5\] sky130_fd_sc_hd__and2_1
X_0585_ count\[4\] _0122_ _0125_ count\[3\] VGND VGND VPWR VPWR _0220_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_49_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3 pwm_counter.sample\[7\] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_218 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_4_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_4_0_clk sky130_fd_sc_hd__clkbuf_8
X_0706_ _0072_ net25 VGND VGND VPWR VPWR _0299_ sky130_fd_sc_hd__nand2_1
XFILLER_38_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0568_ net142 _0074_ _0203_ _0204_ VGND VGND VPWR VPWR pwm_counter.n_pwm sky130_fd_sc_hd__a22o_1
X_0499_ waveshape.seq_div.dividend\[24\] _0137_ VGND VGND VPWR VPWR _0138_ sky130_fd_sc_hd__nor2_1
X_0637_ _0258_ _0259_ VGND VGND VPWR VPWR oscill.n_count\[12\] sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_0_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0971_ clknet_4_15_0_clk net71 net59 VGND VGND VPWR VPWR pwm_counter.active_sample\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_41_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0885_ _0082_ keypad.keypad_reg\[1\] _0207_ _0416_ VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__o31ai_1
X_0954_ clknet_4_3_0_clk _0025_ net62 VGND VGND VPWR VPWR waveshape.seq_div.dividend\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_46_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_143 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0670_ _0074_ _0272_ VGND VGND VPWR VPWR pwm_counter.n_count\[7\] sky130_fd_sc_hd__xnor2_1
Xinput15 n_rst VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_15_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0868_ net42 waveshape.seq_div.dividend\[46\] _0400_ net38 VGND VGND VPWR VPWR _0401_
+ sky130_fd_sc_hd__a22o_1
X_0799_ net143 net24 _0347_ _0348_ VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__o22a_1
X_0937_ clknet_4_12_0_clk _0008_ net58 VGND VGND VPWR VPWR waveshape.scaled_count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_38_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_29_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0653_ sample_rate.count\[3\] sample_rate.count\[4\] _0090_ sample_rate.count\[5\]
+ VGND VGND VPWR VPWR _0268_ sky130_fd_sc_hd__a31o_1
XFILLER_6_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0722_ net44 waveshape.seq_div.dividend\[8\] net29 count\[1\] net19 VGND VGND VPWR
+ VPWR _0307_ sky130_fd_sc_hd__a221o_1
XFILLER_40_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0584_ count\[3\] _0125_ _0130_ count\[2\] VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__o22a_1
XFILLER_33_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold4 _0035_ VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_49_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0636_ count\[12\] _0256_ net17 VGND VGND VPWR VPWR _0259_ sky130_fd_sc_hd__o21ai_1
X_0705_ net38 net26 VGND VGND VPWR VPWR _0298_ sky130_fd_sc_hd__nor2_1
X_0567_ pwm_counter.active_sample\[7\] _0074_ pwm_counter.active_sample\[6\] _0075_
+ VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__o22a_1
X_0498_ _0135_ _0136_ VGND VGND VPWR VPWR _0137_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_0_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Left_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0619_ count\[6\] _0246_ VGND VGND VPWR VPWR _0248_ sky130_fd_sc_hd__and2_1
XFILLER_14_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_3_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_3_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_44_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0970_ clknet_4_15_0_clk net67 net59 VGND VGND VPWR VPWR pwm_counter.active_sample\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0884_ keypad.keypad_reg\[3\] _0205_ keypad.keypad_reg\[2\] VGND VGND VPWR VPWR _0416_
+ sky130_fd_sc_hd__or3b_1
X_0953_ clknet_4_6_0_clk _0024_ net49 VGND VGND VPWR VPWR waveshape.seq_div.dividend\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_23_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0936_ clknet_4_12_0_clk _0007_ net57 VGND VGND VPWR VPWR waveshape.scaled_count\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_0867_ waveshape.seq_div.dividend\[47\] _0194_ VGND VGND VPWR VPWR _0400_ sky130_fd_sc_hd__xnor2_1
X_0798_ net40 waveshape.seq_div.dividend\[29\] net27 VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_38_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_5_Left_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_29_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0652_ net130 _0091_ _0267_ VGND VGND VPWR VPWR sample_rate.n_count\[4\] sky130_fd_sc_hd__o21a_1
XFILLER_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0583_ count\[2\] _0130_ _0216_ _0217_ VGND VGND VPWR VPWR _0218_ sky130_fd_sc_hd__a22o_1
X_0721_ count\[0\] _0104_ net29 net20 net85 VGND VGND VPWR VPWR _0011_ sky130_fd_sc_hd__a32o_1
XFILLER_33_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_47_Left_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0919_ clknet_4_2_0_clk oscill.n_count\[10\] net46 VGND VGND VPWR VPWR count\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_3_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5 pwm_counter.sample\[6\] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_49_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0566_ pwm_counter.active_sample\[6\] _0075_ pwm_counter.active_sample\[5\] _0076_
+ _0202_ VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__a221o_1
X_0635_ count\[12\] _0256_ VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__and2_1
X_0704_ waveshape.seq_div.state\[0\] net28 _0104_ VGND VGND VPWR VPWR _0297_ sky130_fd_sc_hd__o21bai_1
X_0497_ net32 _0119_ _0120_ _0095_ VGND VGND VPWR VPWR _0136_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_0_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0618_ _0246_ _0247_ _0239_ VGND VGND VPWR VPWR oscill.n_count\[5\] sky130_fd_sc_hd__and3b_1
X_0549_ _0167_ _0170_ VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_34_Left_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0952_ clknet_4_6_0_clk _0023_ net49 VGND VGND VPWR VPWR waveshape.seq_div.dividend\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_0883_ _0209_ _0213_ _0402_ VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__nor3_1
Xclkbuf_4_2_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_2_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_45_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0866_ net134 net26 _0362_ _0399_ VGND VGND VPWR VPWR _0063_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_15_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_21_Left_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0935_ clknet_4_12_0_clk _0006_ net57 VGND VGND VPWR VPWR waveshape.scaled_count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_0797_ _0345_ _0346_ net37 VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_38_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_29_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0720_ waveshape.scaled_count\[7\] net20 _0306_ VGND VGND VPWR VPWR _0010_ sky130_fd_sc_hd__a21o_1
X_0651_ sample_rate.count\[4\] _0091_ _0101_ VGND VGND VPWR VPWR _0267_ sky130_fd_sc_hd__a21oi_1
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0582_ count\[1\] _0133_ _0135_ _0136_ count\[0\] VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__a221o_1
XFILLER_10_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0918_ clknet_4_2_0_clk oscill.n_count\[9\] net46 VGND VGND VPWR VPWR count\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_0849_ _0385_ _0386_ net38 VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_3_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold6 _0034_ VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_15_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0703_ waveshape.seq_div.state\[0\] net28 _0104_ VGND VGND VPWR VPWR _0296_ sky130_fd_sc_hd__o21ba_1
X_0565_ pwm_counter.active_sample\[5\] _0076_ pwm_counter.active_sample\[4\] _0077_
+ _0201_ VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__o221a_1
X_0496_ _0069_ _0119_ _0120_ _0100_ VGND VGND VPWR VPWR _0135_ sky130_fd_sc_hd__a31o_1
X_0634_ _0256_ _0257_ net17 VGND VGND VPWR VPWR oscill.n_count\[11\] sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_0_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0479_ net34 net36 VGND VGND VPWR VPWR _0118_ sky130_fd_sc_hd__and2b_1
X_0548_ _0186_ VGND VGND VPWR VPWR _0187_ sky130_fd_sc_hd__inv_2
X_0617_ count\[3\] count\[4\] _0242_ count\[5\] VGND VGND VPWR VPWR _0247_ sky130_fd_sc_hd__a31o_1
XFILLER_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_143 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0882_ _0211_ _0413_ VGND VGND VPWR VPWR _0414_ sky130_fd_sc_hd__nor2_1
X_0951_ clknet_4_6_0_clk _0022_ net57 VGND VGND VPWR VPWR waveshape.seq_div.dividend\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0865_ net41 waveshape.seq_div.dividend\[45\] _0398_ VGND VGND VPWR VPWR _0399_ sky130_fd_sc_hd__a21o_1
X_0934_ clknet_4_12_0_clk _0005_ net57 VGND VGND VPWR VPWR waveshape.scaled_count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_0796_ _0146_ _0158_ _0344_ VGND VGND VPWR VPWR _0346_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_38_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0650_ net111 _0090_ _0266_ VGND VGND VPWR VPWR sample_rate.n_count\[3\] sky130_fd_sc_hd__o21a_1
XFILLER_6_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0581_ count\[1\] _0133_ VGND VGND VPWR VPWR _0216_ sky130_fd_sc_hd__or2_1
Xclkbuf_4_1_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_1_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_19_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0779_ net37 _0142_ _0332_ net43 waveshape.seq_div.dividend\[25\] VGND VGND VPWR
+ VPWR _0333_ sky130_fd_sc_hd__a32o_1
X_0917_ clknet_4_9_0_clk oscill.n_count\[8\] net55 VGND VGND VPWR VPWR count\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_0848_ waveshape.seq_div.dividend\[42\] _0381_ VGND VGND VPWR VPWR _0386_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_3_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold7 pwm_counter.sample\[3\] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__dlygate4sd3_1
X_0633_ count\[9\] count\[10\] _0251_ count\[11\] VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__a31o_1
X_0702_ net38 net42 VGND VGND VPWR VPWR _0295_ sky130_fd_sc_hd__nor2_1
X_0564_ pwm_counter.active_sample\[4\] _0077_ pwm_counter.active_sample\[3\] _0078_
+ _0200_ VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__a221o_1
X_0495_ waveshape.seq_div.dividend\[25\] _0133_ VGND VGND VPWR VPWR _0134_ sky130_fd_sc_hd__and2_1
XFILLER_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0616_ count\[4\] count\[5\] _0243_ VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__and3_1
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0547_ _0178_ _0182_ VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__or2_1
X_0478_ waveshape.seq_div.dividend\[39\] _0114_ _0115_ _0116_ VGND VGND VPWR VPWR
+ _0117_ sky130_fd_sc_hd__and4b_1
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0881_ keypad.keypad_reg\[9\] keypad.keypad_reg\[11\] _0403_ keypad.keypad_reg\[8\]
+ VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__or4bb_1
X_0950_ clknet_4_6_0_clk _0021_ net57 VGND VGND VPWR VPWR waveshape.seq_div.dividend\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_49_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0864_ _0194_ _0397_ _0072_ VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__a21oi_1
X_0795_ _0147_ _0344_ _0158_ VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__a21boi_1
X_0933_ clknet_4_6_0_clk _0004_ net57 VGND VGND VPWR VPWR waveshape.scaled_count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_3_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0580_ count\[4\] _0122_ VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__or2_1
X_0916_ clknet_4_9_0_clk oscill.n_count\[7\] net55 VGND VGND VPWR VPWR count\[7\]
+ sky130_fd_sc_hd__dfrtp_2
X_0778_ _0134_ _0140_ _0141_ VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__or3_1
X_0847_ waveshape.seq_div.dividend\[42\] waveshape.seq_div.dividend\[41\] waveshape.seq_div.dividend\[40\]
+ _0191_ VGND VGND VPWR VPWR _0385_ sky130_fd_sc_hd__nor4_1
XTAP_TAPCELL_ROW_3_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Left_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold8 _0031_ VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_15_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0563_ pwm_counter.active_sample\[3\] _0078_ pwm_counter.active_sample\[2\] _0079_
+ _0199_ VGND VGND VPWR VPWR _0200_ sky130_fd_sc_hd__o221a_1
X_0701_ waveshape.seq_div.dividend\[47\] _0194_ net80 VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__o21a_1
X_0632_ count\[10\] count\[11\] _0253_ VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__and3_1
X_0494_ _0093_ _0132_ _0108_ VGND VGND VPWR VPWR _0133_ sky130_fd_sc_hd__or3b_2
XFILLER_31_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_0_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_0_0_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_45_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0615_ net109 _0243_ _0245_ VGND VGND VPWR VPWR oscill.n_count\[4\] sky130_fd_sc_hd__a21oi_1
X_0546_ _0173_ _0177_ _0178_ _0184_ VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__or4_1
XFILLER_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0477_ waveshape.seq_div.dividend\[37\] _0100_ VGND VGND VPWR VPWR _0116_ sky130_fd_sc_hd__xor2_1
X_1029_ clknet_4_10_0_clk net5 net54 VGND VGND VPWR VPWR keypad.keypad_reg\[13\] sky130_fd_sc_hd__dfrtp_1
XFILLER_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0529_ _0166_ _0167_ VGND VGND VPWR VPWR _0168_ sky130_fd_sc_hd__and2_1
XFILLER_25_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_38_Left_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0880_ _0083_ _0084_ keypad.keypad_reg\[6\] _0405_ VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_18_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0932_ clknet_4_5_0_clk net63 net48 VGND VGND VPWR VPWR sample_rate.count\[7\] sky130_fd_sc_hd__dfrtp_1
X_0863_ waveshape.seq_div.dividend\[45\] waveshape.seq_div.dividend\[44\] _0193_ waveshape.seq_div.dividend\[46\]
+ VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__o31ai_1
X_0794_ _0148_ _0340_ VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__nand2_1
XFILLER_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_25_Left_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0915_ clknet_4_9_0_clk oscill.n_count\[6\] net55 VGND VGND VPWR VPWR count\[6\]
+ sky130_fd_sc_hd__dfrtp_2
X_0777_ _0331_ _0330_ net24 waveshape.seq_div.dividend\[25\] VGND VGND VPWR VPWR _0042_
+ sky130_fd_sc_hd__o2bb2a_1
X_0846_ waveshape.seq_div.dividend\[41\] net25 _0384_ VGND VGND VPWR VPWR _0058_ sky130_fd_sc_hd__o21a_1
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold9 pwm_counter.sample\[4\] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_3_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0700_ net6 net1 _0294_ pwm1 VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__o31a_1
X_0562_ pwm_counter.active_sample\[2\] _0079_ pwm_counter.active_sample\[1\] _0080_
+ _0198_ VGND VGND VPWR VPWR _0199_ sky130_fd_sc_hd__a221o_1
X_0631_ net112 _0253_ _0255_ VGND VGND VPWR VPWR oscill.n_count\[10\] sky130_fd_sc_hd__a21oi_1
X_0493_ net36 net32 net34 net30 VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_0_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0829_ net38 _0370_ _0371_ net41 waveshape.seq_div.dividend\[36\] VGND VGND VPWR
+ VPWR _0372_ sky130_fd_sc_hd__a32o_1
XFILLER_12_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0545_ _0182_ _0183_ VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__or2_1
X_0614_ count\[4\] _0243_ _0239_ VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__o21ai_1
X_0476_ waveshape.seq_div.dividend\[36\] _0109_ VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__xor2_1
X_1028_ clknet_4_10_0_clk net4 net54 VGND VGND VPWR VPWR keypad.keypad_reg\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_14_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_12_Left_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0459_ net32 net34 VGND VGND VPWR VPWR _0099_ sky130_fd_sc_hd__nand2_1
X_0528_ waveshape.seq_div.dividend\[35\] _0165_ VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__or2_1
XFILLER_25_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_90 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0931_ clknet_4_5_0_clk net64 net48 VGND VGND VPWR VPWR sample_rate.count\[6\] sky130_fd_sc_hd__dfrtp_1
X_0862_ waveshape.seq_div.dividend\[45\] net26 _0362_ _0396_ VGND VGND VPWR VPWR _0062_
+ sky130_fd_sc_hd__a22o_1
X_0793_ waveshape.seq_div.dividend\[29\] _0343_ net24 VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__mux2_1
XFILLER_22_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Left_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0914_ clknet_4_9_0_clk oscill.n_count\[5\] net55 VGND VGND VPWR VPWR count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_0845_ net42 waveshape.seq_div.dividend\[40\] _0383_ net38 net27 VGND VGND VPWR VPWR
+ _0384_ sky130_fd_sc_hd__a221o_1
X_0776_ net43 waveshape.seq_div.dividend\[24\] net27 VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__a21oi_1
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_42_Left_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0561_ pwm_counter.active_sample\[1\] _0080_ pwm_counter.active_sample\[0\] _0081_
+ VGND VGND VPWR VPWR _0198_ sky130_fd_sc_hd__o22a_1
X_0492_ waveshape.seq_div.dividend\[26\] _0130_ VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__nand2_1
X_0630_ count\[10\] _0253_ net17 VGND VGND VPWR VPWR _0255_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_0_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0759_ net70 pwm_counter.active_sample\[6\] _0197_ VGND VGND VPWR VPWR _0034_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_31_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0828_ _0116_ _0369_ VGND VGND VPWR VPWR _0371_ sky130_fd_sc_hd__or2_1
XFILLER_28_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0613_ _0243_ _0244_ net17 VGND VGND VPWR VPWR oscill.n_count\[3\] sky130_fd_sc_hd__and3b_1
X_0544_ waveshape.seq_div.dividend\[32\] _0181_ VGND VGND VPWR VPWR _0183_ sky130_fd_sc_hd__nor2_1
X_0475_ _0106_ _0111_ VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__and2_1
XFILLER_38_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1027_ clknet_4_10_0_clk net3 net54 VGND VGND VPWR VPWR keypad.keypad_reg\[11\] sky130_fd_sc_hd__dfrtp_1
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_59 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0458_ _0070_ _0093_ net30 VGND VGND VPWR VPWR _0098_ sky130_fd_sc_hd__a21o_1
X_0527_ waveshape.seq_div.dividend\[35\] _0165_ VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__nand2_1
XFILLER_26_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0930_ clknet_4_7_0_clk sample_rate.n_count\[5\] net50 VGND VGND VPWR VPWR sample_rate.count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_0861_ net39 _0394_ _0395_ net41 waveshape.seq_div.dividend\[44\] VGND VGND VPWR
+ VPWR _0396_ sky130_fd_sc_hd__a32o_1
X_0792_ net37 _0341_ _0342_ net40 waveshape.seq_div.dividend\[28\] VGND VGND VPWR
+ VPWR _0343_ sky130_fd_sc_hd__a32o_1
XFILLER_9_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0775_ _0072_ _0140_ _0329_ VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__or3_1
X_0913_ clknet_4_8_0_clk oscill.n_count\[4\] net52 VGND VGND VPWR VPWR count\[4\]
+ sky130_fd_sc_hd__dfrtp_2
X_0844_ _0381_ _0382_ VGND VGND VPWR VPWR _0383_ sky130_fd_sc_hd__nand2_1
XFILLER_33_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0560_ _0071_ _0103_ _0197_ VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__o21ai_1
X_0491_ _0096_ _0129_ _0108_ VGND VGND VPWR VPWR _0130_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0758_ net66 pwm_counter.active_sample\[5\] _0197_ VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__mux2_1
X_0827_ _0116_ _0369_ VGND VGND VPWR VPWR _0370_ sky130_fd_sc_hd__nand2_1
X_0689_ waveshape.scaled_count\[7\] waveshape.scaled_count\[4\] VGND VGND VPWR VPWR
+ _0287_ sky130_fd_sc_hd__xor2_1
XFILLER_12_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0612_ count\[3\] _0242_ VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__or2_1
XFILLER_38_112 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0543_ waveshape.seq_div.dividend\[32\] _0181_ VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__and2_1
X_0474_ _0111_ _0112_ waveshape.seq_div.dividend\[39\] _0105_ VGND VGND VPWR VPWR
+ _0113_ sky130_fd_sc_hd__a211o_1
XFILLER_38_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1026_ clknet_4_10_0_clk net2 net54 VGND VGND VPWR VPWR keypad.keypad_reg\[10\] sky130_fd_sc_hd__dfrtp_1
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold80 waveshape.scaled_count\[0\] VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__dlygate4sd3_1
X_0526_ net34 _0094_ _0098_ _0164_ VGND VGND VPWR VPWR _0165_ sky130_fd_sc_hd__a22o_1
X_0457_ net32 net34 VGND VGND VPWR VPWR _0097_ sky130_fd_sc_hd__nor2_1
X_1009_ clknet_4_15_0_clk pwm_counter.n_count\[7\] net60 VGND VGND VPWR VPWR pwm_counter.count\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0509_ waveshape.seq_div.dividend\[29\] _0145_ VGND VGND VPWR VPWR _0148_ sky130_fd_sc_hd__or2_1
XFILLER_36_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0860_ waveshape.seq_div.dividend\[44\] _0193_ _0073_ VGND VGND VPWR VPWR _0395_
+ sky130_fd_sc_hd__o21ai_1
X_0791_ _0149_ _0340_ VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__nand2_1
XFILLER_9_133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0989_ clknet_4_1_0_clk _0052_ net47 VGND VGND VPWR VPWR waveshape.seq_div.dividend\[35\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_47_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0912_ clknet_4_10_0_clk oscill.n_count\[3\] net52 VGND VGND VPWR VPWR count\[3\]
+ sky130_fd_sc_hd__dfrtp_2
X_0774_ _0138_ _0139_ VGND VGND VPWR VPWR _0329_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_11_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0843_ waveshape.seq_div.dividend\[40\] _0191_ waveshape.seq_div.dividend\[41\] VGND
+ VGND VPWR VPWR _0382_ sky130_fd_sc_hd__o21ai_1
XFILLER_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_29_Left_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0490_ _0069_ _0120_ _0107_ VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__a21oi_1
XFILLER_2_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0757_ net74 pwm_counter.active_sample\[4\] _0197_ VGND VGND VPWR VPWR _0032_ sky130_fd_sc_hd__mux2_1
X_0688_ net146 _0278_ _0279_ _0286_ _0282_ VGND VGND VPWR VPWR waveshape.shaper.n_sample\[4\]
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0826_ waveshape.seq_div.dividend\[36\] _0109_ _0366_ VGND VGND VPWR VPWR _0369_
+ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_39_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_15_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_15_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_44_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0542_ net30 _0129_ _0180_ VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__a21oi_2
X_0611_ count\[3\] _0242_ VGND VGND VPWR VPWR _0243_ sky130_fd_sc_hd__and2_1
XFILLER_38_124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0473_ waveshape.seq_div.dividend\[37\] _0100_ _0110_ VGND VGND VPWR VPWR _0112_
+ sky130_fd_sc_hd__o21a_1
X_1025_ clknet_4_10_0_clk net14 net52 VGND VGND VPWR VPWR keypad.keypad_reg\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_14_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0809_ _0182_ _0353_ VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__nor2_1
XFILLER_39_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold81 waveshape.scaled_count\[4\] VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__dlygate4sd3_1
Xhold70 waveshape.seq_div.dividend\[32\] VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0456_ net30 net32 VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__and2b_1
XFILLER_6_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0525_ net36 _0069_ _0070_ net30 VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__o211ai_1
XPHY_EDGE_ROW_16_Left_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1008_ clknet_4_15_0_clk pwm_counter.n_count\[6\] net60 VGND VGND VPWR VPWR pwm_counter.count\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0439_ pwm_counter.count\[2\] VGND VGND VPWR VPWR _0079_ sky130_fd_sc_hd__inv_2
X_0508_ waveshape.seq_div.dividend\[29\] _0145_ VGND VGND VPWR VPWR _0147_ sky130_fd_sc_hd__nand2_1
XFILLER_39_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0790_ _0149_ _0340_ VGND VGND VPWR VPWR _0341_ sky130_fd_sc_hd__or2_1
XFILLER_9_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0988_ clknet_4_1_0_clk _0051_ net47 VGND VGND VPWR VPWR waveshape.seq_div.dividend\[34\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_22_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0911_ clknet_4_8_0_clk oscill.n_count\[2\] net55 VGND VGND VPWR VPWR count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_0842_ waveshape.seq_div.dividend\[41\] waveshape.seq_div.dividend\[40\] _0191_ VGND
+ VGND VPWR VPWR _0381_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_11_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0773_ net24 _0327_ _0328_ net128 VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_34_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_4_Left_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0825_ waveshape.seq_div.dividend\[36\] _0368_ net25 VGND VGND VPWR VPWR _0053_ sky130_fd_sc_hd__mux2_1
X_0756_ net72 pwm_counter.active_sample\[3\] _0197_ VGND VGND VPWR VPWR _0031_ sky130_fd_sc_hd__mux2_1
X_0687_ waveshape.scaled_count\[7\] waveshape.scaled_count\[3\] VGND VGND VPWR VPWR
+ _0286_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_46_Left_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0541_ net32 _0070_ _0095_ VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__a21oi_1
XFILLER_7_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0610_ _0242_ net17 _0241_ VGND VGND VPWR VPWR oscill.n_count\[2\] sky130_fd_sc_hd__and3b_1
X_0472_ waveshape.seq_div.dividend\[38\] _0098_ VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__or2_1
XFILLER_38_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1024_ clknet_4_10_0_clk net13 net52 VGND VGND VPWR VPWR keypad.keypad_reg\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_15_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0808_ net135 _0355_ net24 VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__mux2_1
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0739_ net100 net23 _0315_ VGND VGND VPWR VPWR _0020_ sky130_fd_sc_hd__o21a_1
XFILLER_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold60 pwm_counter.count\[3\] VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 waveshape.scaled_count\[1\] VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 waveshape.scaled_count\[2\] VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_14_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_14_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_6_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0524_ _0144_ _0159_ _0162_ VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__o21a_1
X_0455_ net36 net33 net31 VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__o21bai_1
X_1007_ clknet_4_15_0_clk pwm_counter.n_count\[5\] net60 VGND VGND VPWR VPWR pwm_counter.count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_33_Left_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0438_ pwm_counter.count\[3\] VGND VGND VPWR VPWR _0078_ sky130_fd_sc_hd__inv_2
X_0507_ waveshape.seq_div.dividend\[29\] _0145_ VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__and2_1
XFILLER_22_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0987_ clknet_4_0_0_clk _0050_ net47 VGND VGND VPWR VPWR waveshape.seq_div.dividend\[33\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_6_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0772_ net37 _0137_ net27 VGND VGND VPWR VPWR _0328_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_11_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0910_ clknet_4_9_0_clk oscill.n_count\[1\] net57 VGND VGND VPWR VPWR count\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0841_ waveshape.seq_div.dividend\[40\] net25 _0380_ VGND VGND VPWR VPWR _0057_ sky130_fd_sc_hd__o21a_1
XFILLER_45_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_20_Left_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0755_ net76 pwm_counter.active_sample\[2\] _0197_ VGND VGND VPWR VPWR _0030_ sky130_fd_sc_hd__mux2_1
X_0824_ _0366_ _0367_ net41 waveshape.seq_div.dividend\[35\] VGND VGND VPWR VPWR _0368_
+ sky130_fd_sc_hd__a2bb2o_1
X_0686_ waveshape.scaled_count\[3\] _0278_ _0279_ _0285_ _0282_ VGND VGND VPWR VPWR
+ waveshape.shaper.n_sample\[3\] sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_39_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0540_ _0177_ _0178_ VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__nor2_1
X_0471_ waveshape.seq_div.dividend\[37\] _0100_ _0109_ waveshape.seq_div.dividend\[36\]
+ VGND VGND VPWR VPWR _0110_ sky130_fd_sc_hd__a22o_1
X_0931__64 VGND VGND VPWR VPWR _0931__64/HI net64 sky130_fd_sc_hd__conb_1
X_1023_ clknet_4_8_0_clk net12 net52 VGND VGND VPWR VPWR keypad.keypad_reg\[7\] sky130_fd_sc_hd__dfrtp_1
X_0807_ _0353_ _0354_ net40 waveshape.seq_div.dividend\[31\] VGND VGND VPWR VPWR _0355_
+ sky130_fd_sc_hd__a2bb2o_1
X_0738_ net44 waveshape.seq_div.dividend\[16\] net28 count\[9\] net21 VGND VGND VPWR
+ VPWR _0315_ sky130_fd_sc_hd__a221o_1
X_0669_ _0272_ _0276_ VGND VGND VPWR VPWR pwm_counter.n_count\[6\] sky130_fd_sc_hd__nor2_1
XFILLER_39_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold50 waveshape.seq_div.n\[1\] VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 waveshape.seq_div.dividend\[27\] VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 waveshape.seq_div.dividend\[34\] VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 waveshape.scaled_count\[5\] VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0523_ _0152_ _0157_ _0161_ VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__a21oi_1
X_0454_ net36 net33 VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__or2_1
X_1006_ clknet_4_15_0_clk pwm_counter.n_count\[4\] net59 VGND VGND VPWR VPWR pwm_counter.count\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_34_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0506_ net30 _0093_ _0118_ _0100_ _0097_ VGND VGND VPWR VPWR _0145_ sky130_fd_sc_hd__o32a_2
X_0437_ pwm_counter.count\[4\] VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__inv_2
XFILLER_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_13_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_13_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_62 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0986_ clknet_4_0_0_clk _0049_ net47 VGND VGND VPWR VPWR waveshape.seq_div.dividend\[32\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_6_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0771_ net40 waveshape.seq_div.dividend\[23\] _0138_ net37 VGND VGND VPWR VPWR _0327_
+ sky130_fd_sc_hd__a22o_1
X_0840_ net41 waveshape.seq_div.dividend\[39\] _0379_ net38 net26 VGND VGND VPWR VPWR
+ _0380_ sky130_fd_sc_hd__a221o_1
XFILLER_38_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0969_ clknet_4_15_0_clk net75 net59 VGND VGND VPWR VPWR pwm_counter.active_sample\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_3_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_48_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0754_ net83 pwm_counter.active_sample\[1\] _0197_ VGND VGND VPWR VPWR _0029_ sky130_fd_sc_hd__mux2_1
X_0823_ _0115_ _0190_ net38 VGND VGND VPWR VPWR _0367_ sky130_fd_sc_hd__o21ai_1
X_0685_ waveshape.scaled_count\[7\] waveshape.scaled_count\[2\] VGND VGND VPWR VPWR
+ _0285_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_39_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0470_ net36 _0108_ _0107_ VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__o21bai_4
XFILLER_38_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1022_ clknet_4_8_0_clk net11 net52 VGND VGND VPWR VPWR keypad.keypad_reg\[6\] sky130_fd_sc_hd__dfrtp_1
X_0668_ pwm_counter.count\[6\] _0271_ VGND VGND VPWR VPWR _0276_ sky130_fd_sc_hd__nor2_1
X_0806_ _0163_ _0184_ _0072_ VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__a21o_1
X_0737_ net92 net22 _0314_ VGND VGND VPWR VPWR _0019_ sky130_fd_sc_hd__o21a_1
X_0599_ count\[14\] _0098_ _0100_ count\[13\] VGND VGND VPWR VPWR _0234_ sky130_fd_sc_hd__o22a_1
XFILLER_20_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold40 count\[0\] VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 sample_rate.count\[2\] VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 _0322_ VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 waveshape.scaled_count\[1\] VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 waveshape.seq_div.dividend\[33\] VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0522_ _0153_ _0158_ _0160_ _0150_ waveshape.seq_div.dividend\[31\] VGND VGND VPWR
+ VPWR _0161_ sky130_fd_sc_hd__a32o_1
X_0453_ net36 net32 VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__nor2_1
XFILLER_20_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1005_ clknet_4_15_0_clk pwm_counter.n_count\[3\] net59 VGND VGND VPWR VPWR pwm_counter.count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_34_163 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0436_ pwm_counter.count\[5\] VGND VGND VPWR VPWR _0076_ sky130_fd_sc_hd__inv_2
X_0505_ _0126_ _0131_ _0142_ _0127_ _0123_ VGND VGND VPWR VPWR _0144_ sky130_fd_sc_hd__a311o_1
.ends

